-- File created by Bench2VHDL
-- Name: s1196b
-- File: bench/s1196b.bench
-- Timestamp: 2019-05-21T22:08:28.767691
--
-- Original File
-- =============
--	#  file :s1196.v
--	# //# 14 inputs 
--	# //# 14 outputs 
--	# //# 18 d-type flipflops 
--	# //# 141 inverters 
--	# //# 388 gates (118 ands + 119 nands + 101 ors + 50 nors) 
--	#  module :s1196
--	# 
--	# inputs
--	INPUT(G0)
--	INPUT(G1)
--	INPUT(G2)
--	INPUT(G3)
--	INPUT(G4)
--	INPUT(G5)
--	INPUT(G6)
--	INPUT(G7)
--	INPUT(G8)
--	INPUT(G9)
--	INPUT(G10)
--	INPUT(G11)
--	INPUT(G12)
--	INPUT(G13)
--	# 
--	# outputs
--	OUTPUT(G546)
--	OUTPUT(G539)
--	OUTPUT(G550)
--	OUTPUT(G551)
--	OUTPUT(G552)
--	OUTPUT(G547)
--	OUTPUT(G548)
--	OUTPUT(G549)
--	OUTPUT(G530)
--	OUTPUT(G45)
--	OUTPUT(G542)
--	OUTPUT(G532)
--	OUTPUT(G535)
--	OUTPUT(G537)
--	#
--	#      out =   type (input(s)...      )  # verilog node 
--	#
--	G29 = DFF( G502)
--	G30 = DFF( G503)
--	G31 = DFF( G504)
--	G32 = DFF( G505)
--	G33 = DFF( G506)
--	G34 = DFF( G507)
--	G35 = DFF( G508)
--	G36 = DFF( G509)
--	G37 = DFF( G510)
--	G38 = DFF( G511)
--	G39 = DFF( G512)
--	G40 = DFF( G513)
--	G41 = DFF( G514)
--	G42 = DFF( G515)
--	G43 = DFF( G516)
--	G44 = DFF( G517)
--	G45 = DFF( G518)
--	G46 = DFF( G519)
--	G520 = NOT( G0)
--	G521 = NOT( G1)
--	G522 = NOT( G2)
--	G524 = NOT( G3)
--	II156 = NOT( G4)
--	G334 = NOT( II156)
--	G527 = NOT( G4)
--	G528 = NOT( G5)
--	G529 = NOT( G6)
--	G531 = NOT( G7)
--	G533 = NOT( G8)
--	G536 = NOT( G9)
--	G538 = NOT( G10)
--	G540 = NOT( G11)
--	G541 = NOT( G12)
--	G543 = NOT( G13)
--	G476 = NOT( G30)
--	G484 = NOT( G30)
--	G125 = NOT( G40)
--	G140 = NOT( G33)
--	G546 = NOT( G41)
--	G132 = NOT( G42)
--	G70 = NOT( G43)
--	G67 = NOT( G44)
--	G99 = NOT( G29)
--	G475 = NOT( G57)
--	G59 = NOT( G58)
--	G228 = NOT( G524)
--	G272 = NOT( G271)
--	G98 = NOT( G97)
--	G135 = NOT( G134)
--	II218 = NOT( G528)
--	G333 = NOT( II218)
--	G55 = NOT( G54)
--	G165 = NOT( G529)
--	G72 = NOT( G71)
--	G236 = NOT( G274)
--	G275 = NOT( G274)
--	II249 = NOT( G538)
--	G370 = NOT( II249)
--	G75 = NOT( G74)
--	G490 = NOT( G190)
--	G482 = NOT( G241)
--	G153 = NOT( G522)
--	G192 = NOT( G193)
--	G123 = NOT( G122)
--	II272 = NOT( G209)
--	G458 = NOT( II272)
--	II276 = NOT( G238)
--	G332 = NOT( II276)
--	II280 = NOT( G272)
--	G309 = NOT( II280)
--	II287 = NOT( G135)
--	G347 = NOT( II287)
--	G498 = NOT( G195)
--	G78 = NOT( G77)
--	II295 = NOT( G198)
--	G459 = NOT( II295)
--	G199 = NOT( G200)
--	G90 = NOT( G89)
--	G221 = NOT( G222)
--	G223 = NOT( G224)
--	II316 = NOT( G239)
--	G369 = NOT( II316)
--	G234 = NOT( G235)
--	II327 = NOT( G135)
--	G435 = NOT( II327)
--	II330 = NOT( G236)
--	G441 = NOT( II330)
--	G50 = NOT( G49)
--	G130 = NOT( G9)
--	G501 = NOT( G156)
--	G477 = NOT( G276)
--	G485 = NOT( G276)
--	II352 = NOT( G77)
--	G299 = NOT( II352)
--	G497 = NOT( G205)
--	II371 = NOT( G1)
--	G335 = NOT( II371)
--	II374 = NOT( G520)
--	G456 = NOT( II374)
--	G87 = NOT( G86)
--	II386 = NOT( G199)
--	G414 = NOT( II386)
--	G486 = NOT( G68)
--	G231 = NOT( G232)
--	G160 = NOT( G161)
--	G265 = NOT( G50)
--	G64 = NOT( G63)
--	G180 = NOT( G181)
--	G107 = NOT( G456)
--	G207 = NOT( G208)
--	G167 = NOT( G168)
--	G124 = NOT( G206)
--	G203 = NOT( G204)
--	G489 = NOT( G273)
--	G495 = NOT( G273)
--	G177 = NOT( G357)
--	G212 = NOT( G213)
--	II493 = NOT( G218)
--	G404 = NOT( II493)
--	II502 = NOT( G124)
--	G468 = NOT( II502)
--	G173 = NOT( G495)
--	G487 = NOT( G534)
--	II529 = NOT( G468)
--	G149 = NOT( II529)
--	II536 = NOT( G79)
--	G446 = NOT( II536)
--	G494 = NOT( G173)
--	G500 = NOT( G173)
--	G214 = NOT( G215)
--	G492 = NOT( G62)
--	G483 = NOT( G182)
--	G282 = NOT( G281)
--	II573 = NOT( G176)
--	G403 = NOT( II573)
--	II576 = NOT( G175)
--	G447 = NOT( II576)
--	G479 = NOT( G194)
--	G491 = NOT( G194)
--	G554 = NOT( G553)
--	G170 = NOT( G171)
--	G172 = NOT( G171)
--	G525 = NOT( G526)
--	G493 = NOT( G544)
--	G545 = NOT( G544)
--	G488 = NOT( G172)
--	G499 = NOT( G280)
--	II624 = NOT( G120)
--	G303 = NOT( II624)
--	G480 = NOT( G179)
--	II631 = NOT( G188)
--	G336 = NOT( II631)
--	G496 = NOT( G188)
--	G174 = NOT( G496)
--	II662 = NOT( G174)
--	G405 = NOT( II662)
--	G478 = NOT( G279)
--	II692 = NOT( G145)
--	G432 = NOT( II692)
--	G359 = AND( G6, G31)
--	G469 = AND( G163, G3)
--	G461 = AND( G529, G531)
--	G431 = AND( G524, G67)
--	G362 = AND( G129, G77)
--	G81 = AND( G288, G240)
--	G348 = AND( G97, G55)
--	G352 = AND( G8, G135, G37, G164)
--	G511 = AND( G163, G164)
--	G379 = AND( G9, G211)
--	G385 = AND( G529, G7, G49)
--	G376 = AND( G533, G75)
--	G387 = AND( G6, G274, G75)
--	G462 = AND( G192, G538)
--	G436 = AND( G123, G77)
--	G363 = AND( G77, G205)
--	G410 = AND( G1, G205)
--	G399 = AND( G520, G1)
--	G437 = AND( G66, G229)
--	G307 = AND( G6, G104)
--	G306 = AND( G524, G78)
--	G283 = AND( G122, G219)
--	G339 = AND( G533, G199, G209)
--	G472 = AND( G136, G9, G190)
--	G351 = AND( G524, G169, G221, G234)
--	G440 = AND( G38, G234)
--	G382 = AND( G9, G100, G34)
--	G386 = AND( G536, G85)
--	G321 = AND( G90, G50)
--	G378 = AND( G89, G50)
--	G471 = AND( G191, G103, G112)
--	G377 = AND( G90, G56)
--	G358 = AND( G7, G83)
--	G400 = AND( G0, G277)
--	G308 = AND( G5, G151)
--	G411 = AND( G48, G59)
--	G413 = AND( G197, G201)
--	G434 = AND( G165, G231)
--	G373 = AND( G34, G160)
--	G357 = AND( G265, G232)
--	G444 = AND( G64, G78, G211)
--	G361 = AND( G6, G202)
--	G346 = AND( G2, G82)
--	G457 = AND( G4, G107)
--	G364 = AND( G2, G109)
--	G445 = AND( G53, G225)
--	G412 = AND( G3, G207)
--	G371 = AND( G161, G168, G267)
--	G353 = AND( G11, G92, G163)
--	G388 = AND( G11, G114)
--	G473 = AND( G11, G143)
--	G331 = AND( G213, G257)
--	G429 = AND( G51, G225)
--	G380 = AND( G6, G93)
--	G360 = AND( G8, G106)
--	G338 = AND( G202, G203)
--	G337 = AND( G270, G167)
--	G340 = AND( G8, G270)
--	G322 = AND( G522, G105, G196)
--	G330 = AND( G248, G249)
--	G430 = AND( G177, G196)
--	G344 = AND( G111, G189, G195)
--	G428 = AND( G212, G227)
--	G349 = AND( G6, G108)
--	G460 = AND( G2, G81, G115)
--	G463 = AND( G521, G148)
--	G393 = AND( G127, G34)
--	G470 = AND( G528, G149)
--	G341 = AND( G531, G118)
--	G342 = AND( G73, G197)
--	G324 = AND( G522, G183)
--	G323 = AND( G2, G144)
--	G354 = AND( G0, G214)
--	G312 = AND( G180, G182)
--	G315 = AND( G250, G251)
--	G474 = AND( G242, G77)
--	G343 = AND( G2, G528, G147)
--	G304 = AND( G52, G158)
--	G398 = AND( G94, G156, G158)
--	G365 = AND( G282, G137, G156)
--	G417 = AND( G13, G282, G70)
--	G290 = AND( G117, G135, G157)
--	G327 = AND( G4, G39, G157)
--	G367 = AND( G126, G157)
--	G397 = AND( G101, G98, G157)
--	G451 = AND( G541, G554, G187)
--	G406 = AND( G87, G172)
--	G418 = AND( G524, G60, G172)
--	G453 = AND( G545, G186)
--	G289 = AND( G2, G119, G156)
--	G311 = AND( G0, G178, G179)
--	G402 = AND( G154, G183)
--	G433 = AND( G91, G154)
--	G449 = AND( G88, G154)
--	G452 = AND( G526, G184)
--	G329 = AND( G150, G156)
--	G291 = AND( G138, G155)
--	G328 = AND( G5, G102, G155)
--	G366 = AND( G125, G155)
--	G372 = AND( G116, G275, G155)
--	G383 = AND( G131, G155)
--	G392 = AND( G132, G155)
--	G396 = AND( G76, G272, G155)
--	G401 = AND( G2, G110, G155)
--	G422 = AND( G0, G80, G155)
--	G415 = AND( G146, G142, G165)
--	G425 = AND( G146, G176)
--	G438 = AND( G8, G146, G133)
--	G424 = AND( G78, G174, G177)
--	G439 = AND( G174, G175)
--	G317 = AND( G159, G245)
--	G426 = AND( G37, G162, G38)
--	G443 = AND( G47, G162)
--	G416 = AND( G61, G167)
--	G427 = AND( G541, G95, G165)
--	G442 = AND( G541, G121)
--	G423 = AND( G541, G128)
--	G448 = AND( G139, G153)
--	G419 = OR( G3, G5)
--	G193 = OR( G6, G30)
--	G394 = OR( G5, G58)
--	G407 = OR( G6, G117)
--	G314 = OR( G527, G57)
--	G395 = OR( G4, G134)
--	G288 = OR( G1, G528)
--	G302 = OR( G4, G529)
--	G224 = OR( G533, G31)
--	G355 = OR( G11, G116)
--	G316 = OR( G531, G536)
--	G350 = OR( G6, G536)
--	G368 = OR( G533, G536)
--	G381 = OR( G7, G71)
--	G384 = OR( G529, G71)
--	G389 = OR( G9, G274)
--	G374 = OR( G536, G538)
--	G286 = OR( G9, G540)
--	G293 = OR( G7, G540)
--	G375 = OR( G10, G540)
--	G356 = OR( G6, G476)
--	G313 = OR( G521, G475)
--	G420 = OR( G522, G59)
--	G421 = OR( G521, G2, G228)
--	G320 = OR( G76, G272)
--	G310 = OR( G522, G135)
--	G408 = OR( G529, G77)
--	G305 = OR( G524, G55)
--	G409 = OR( G528, G55)
--	G296 = OR( G89, G484)
--	G325 = OR( G7, G536, G222)
--	G464 = OR( G72, G536)
--	G391 = OR( G74, G220)
--	G292 = OR( G538, G75)
--	G345 = OR( G529, G226)
--	G465 = OR( G524, G210)
--	G454 = OR( G122, G77)
--	G269 = OR( G362, G529)
--	G287 = OR( G522, G81)
--	G318 = OR( G6, G8, G232)
--	G326 = OR( G533, G232)
--	G390 = OR( G89, G50)
--	G298 = OR( G5, G497)
--	G300 = OR( G87, G97)
--	G261 = OR( G283, G528)
--	G301 = OR( G122, G486)
--	G92 = OR( G351, G352)
--	G47 = OR( G440, G441)
--	G114 = OR( G385, G386)
--	G297 = OR( G64, G274)
--	G93 = OR( G376, G377, G378)
--	G106 = OR( G358, G359)
--	G110 = OR( G399, G400)
--	G455 = OR( G78, G206)
--	G152 = OR( G306, G307, G308)
--	G60 = OR( G413, G414)
--	G133 = OR( G434, G435)
--	G105 = OR( G321, G273)
--	G108 = OR( G346, G347)
--	G115 = OR( G457, G458, G459)
--	G126 = OR( G363, G364)
--	G79 = OR( G444, G445)
--	G319 = OR( G529, G489)
--	G131 = OR( G379, G380)
--	G118 = OR( G337, G338)
--	G73 = OR( G339, G340)
--	G91 = OR( G430, G431)
--	G137 = OR( G348, G349)
--	G242 = OR( G469, G470)
--	G147 = OR( G341, G342)
--	G284 = OR( G528, G272, G281)
--	G294 = OR( G1, G117, G281)
--	G553 = OR( G322, G323, G324)
--	G141 = OR( G353, G354)
--	G142 = OR( G403, G404)
--	G88 = OR( G446, G447)
--	G544 = OR( G343, G344)
--	G285 = OR( G5, G479)
--	G295 = OR( G122, G491)
--	G450 = OR( G12, G171)
--	G150 = OR( G303, G304)
--	G146 = OR( G336, G170)
--	G539 = OR( G451, G452, G453)
--	G244 = OR( G371, G159)
--	G550 = OR( G289, G290, G291, G485)
--	G551 = OR( G327, G328, G329)
--	G552 = OR( G365, G366, G367)
--	G547 = OR( G382, G383)
--	G548 = OR( G392, G393)
--	G549 = OR( G396, G397, G398, G477)
--	G530 = OR( G401, G402)
--	G61 = OR( G405, G406)
--	G95 = OR( G424, G425)
--	G121 = OR( G438, G439)
--	G279 = OR( G317, G166)
--	G128 = OR( G415, G416, G417, G418)
--	G145 = OR( G426, G427)
--	G139 = OR( G442, G443)
--	G532 = OR( G422, G423)
--	G535 = OR( G432, G433)
--	G537 = OR( G448, G449)
--	G57 = NAND( G0, G2)
--	G58 = NAND( G1, G3)
--	G76 = NAND( G0, G3)
--	G101 = NAND( G3, G4)
--	G117 = NAND( G2, G4)
--	G271 = NAND( G1, G4)
--	G97 = NAND( G2, G5)
--	G134 = NAND( G3, G5)
--	G54 = NAND( G4, G6)
--	G116 = NAND( G6, G9)
--	G71 = NAND( G8, G10)
--	G274 = NAND( G7, G10)
--	G74 = NAND( G9, G11)
--	G112 = NAND( G8, G31)
--	G245 = NAND( G8, G34)
--	G122 = NAND( G522, G3)
--	G238 = NAND( G2, G524)
--	G129 = NAND( G527, G5)
--	G240 = NAND( G4, G134)
--	G252 = NAND( G3, G11, G35, G216)
--	G77 = NAND( G4, G528)
--	G103 = NAND( G529, G7, G30)
--	G200 = NAND( G527, G529)
--	G248 = NAND( G529, G36)
--	G89 = NAND( G531, G8)
--	G222 = NAND( G533, G10)
--	G239 = NAND( G7, G533)
--	G235 = NAND( G6, G536)
--	G220 = NAND( G7, G71)
--	G49 = NAND( G9, G538)
--	G251 = NAND( G543, G32)
--	G276 = NAND( G3, G543, G140)
--	G263 = NAND( G0, G99)
--	G226 = NAND( G527, G59)
--	G210 = NAND( G520, G272)
--	G66 = NAND( G129, G101)
--	G233 = NAND( G522, G135)
--	G104 = NAND( G122, G238, G240)
--	G86 = NAND( G55, G3)
--	G219 = NAND( G524, G55)
--	G68 = NAND( G302, G528)
--	G232 = NAND( G536, G164)
--	G136 = NAND( G222, G224)
--	G510 = NAND( G350, G235)
--	G161 = NAND( G316, G72)
--	G100 = NAND( G381, G220)
--	G85 = NAND( G384, G239)
--	G243 = NAND( G368, G275, G34)
--	G63 = NAND( G75, G8)
--	G237 = NAND( G10, G75, G201)
--	G503 = NAND( G286, G538)
--	G56 = NAND( G374, G375)
--	G83 = NAND( G355, G356)
--	G96 = NAND( G313, G314)
--	G278 = NAND( G332, G333)
--	G255 = NAND( G309, G2, G529)
--	G69 = NAND( G419, G420, G233)
--	G512 = NAND( G310, G233)
--	G181 = NAND( G2, G78)
--	G277 = NAND( G394, G395, G81)
--	G151 = NAND( G305, G200)
--	G48 = NAND( G407, G408, G409)
--	G264 = NAND( G227, G241)
--	G208 = NAND( G68, G229)
--	G168 = NAND( G75, G221)
--	G84 = NAND( G369, G370)
--	G258 = NAND( G464, G103, G223)
--	G166 = NAND( G7, G50)
--	G259 = NAND( G130, G225)
--	G504 = NAND( G292, G293)
--	G217 = NAND( G50, G230)
--	G257 = NAND( G538, G230)
--	G260 = NAND( G528, G529, G191)
--	G266 = NAND( G524, G96)
--	G262 = NAND( G527, G278)
--	G138 = NAND( G465, G263)
--	G256 = NAND( G4, G69)
--	G82 = NAND( G334, G335)
--	G109 = NAND( G269, G219)
--	G206 = NAND( G287, G524)
--	G204 = NAND( G521, G87)
--	G53 = NAND( G264, G237)
--	G273 = NAND( G325, G326)
--	G267 = NAND( G536, G84)
--	G113 = NAND( G389, G390)
--	G143 = NAND( G258, G193, G259)
--	G213 = NAND( G64, G275)
--	G51 = NAND( G260, G237)
--	G102 = NAND( G320, G266, G210)
--	G52 = NAND( G298, G299, G219)
--	G80 = NAND( G421, G226, G256)
--	G270 = NAND( G345, G204)
--	G94 = NAND( G261, G181, G262)
--	G505 = NAND( G300, G301, G181)
--	G249 = NAND( G11, G273, G201)
--	G268 = NAND( G11, G113)
--	G111 = NAND( G213, G217)
--	G534 = NAND( G296, G297, G166)
--	G253 = NAND( G87, G218)
--	G148 = NAND( G454, G455, G0)
--	G254 = NAND( G1, G152)
--	G127 = NAND( G391, G268)
--	G215 = NAND( G135, G55, G212)
--	G62 = NAND( G534, G32)
--	G523 = NAND( G254, G255, G208)
--	G508 = NAND( G318, G319)
--	G144 = NAND( G215, G252, G253)
--	G250 = NAND( G13, G523)
--	G281 = NAND( G523, G534)
--	G171 = NAND( G553, G187)
--	G526 = NAND( G1, G2, G141)
--	G280 = NAND( G46, G247)
--	G246 = NAND( G544, G186)
--	G119 = NAND( G284, G285)
--	G120 = NAND( G294, G295)
--	G185 = NAND( G525, G184)
--	G159 = NAND( G6, G155)
--	G518 = NAND( G450, G185, G246)
--	G542 = NAND( G243, G244, G279)
--	G163 = NOR( G0, G4)
--	G216 = NOR( G4, G5)
--	G169 = NOR( G5, G7)
--	G225 = NOR( G7, G8)
--	G190 = NOR( G7, G11)
--	G241 = NOR( G10, G11)
--	G198 = NOR( G520, G3)
--	G178 = NOR( G521, G4)
--	G229 = NOR( G1, G522)
--	G209 = NOR( G1, G524)
--	G195 = NOR( G521, G134)
--	G189 = NOR( G522, G54)
--	G201 = NOR( G528, G54)
--	G164 = NOR( G531, G10)
--	G211 = NOR( G6, G274)
--	G156 = NOR( G12, G543)
--	G205 = NOR( G529, G122)
--	G227 = NOR( G5, G200)
--	G230 = NOR( G8, G490)
--	G191 = NOR( G9, G482)
--	G196 = NOR( G5, G540, G86)
--	G197 = NOR( G540, G232)
--	G202 = NOR( G10, G63)
--	G502 = NOR( G436, G437)
--	G218 = NOR( G528, G217)
--	G516 = NOR( G410, G411, G412)
--	G515 = NOR( G387, G388)
--	G509 = NOR( G331, G5)
--	G513 = NOR( G360, G361)
--	G183 = NOR( G330, G3)
--	G517 = NOR( G428, G429)
--	G182 = NOR( G12, G62)
--	G519 = NOR( G460, G461, G462, G463)
--	G176 = NOR( G4, G494)
--	G175 = NOR( G86, G500)
--	G187 = NOR( G13, G492)
--	G158 = NOR( G521, G281)
--	G194 = NOR( G281, G271)
--	G157 = NOR( G13, G483)
--	G507 = NOR( G315, G12, G487)
--	G186 = NOR( G282, G501)
--	G247 = NOR( G471, G472, G473, G474)
--	G179 = NOR( G541, G280)
--	G188 = NOR( G543, G493)
--	G154 = NOR( G12, G488)
--	G184 = NOR( G541, G13, G499)
--	G506 = NOR( G311, G312)
--	G155 = NOR( G13, G480)
--	G162 = NOR( G185, G498)
--	G514 = NOR( G372, G373, G478)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s1196b is
	port (
		CLK: in std_logic;
		G0: in std_logic;
		G1: in std_logic;
		G2: in std_logic;
		G3: in std_logic;
		G4: in std_logic;
		G5: in std_logic;
		G6: in std_logic;
		G7: in std_logic;
		G8: in std_logic;
		G9: in std_logic;
		G10: in std_logic;
		G11: in std_logic;
		G12: in std_logic;
		G13: in std_logic;
		G45: out std_logic;
		G530: out std_logic;
		G532: out std_logic;
		G535: out std_logic;
		G537: out std_logic;
		G539: out std_logic;
		G542: out std_logic;
		G546: out std_logic;
		G547: out std_logic;
		G548: out std_logic;
		G549: out std_logic;
		G550: out std_logic;
		G551: out std_logic;
		G552: out std_logic
	);
end entity;

architecture RTL of s1196b is
	attribute dont_touch: boolean;

	signal G29: std_logic; attribute dont_touch of G29: signal is true;
	signal G30: std_logic; attribute dont_touch of G30: signal is true;
	signal G31: std_logic; attribute dont_touch of G31: signal is true;
	signal G32: std_logic; attribute dont_touch of G32: signal is true;
	signal G33: std_logic; attribute dont_touch of G33: signal is true;
	signal G34: std_logic; attribute dont_touch of G34: signal is true;
	signal G35: std_logic; attribute dont_touch of G35: signal is true;
	signal G36: std_logic; attribute dont_touch of G36: signal is true;
	signal G37: std_logic; attribute dont_touch of G37: signal is true;
	signal G38: std_logic; attribute dont_touch of G38: signal is true;
	signal G39: std_logic; attribute dont_touch of G39: signal is true;
	signal G40: std_logic; attribute dont_touch of G40: signal is true;
	signal G41: std_logic; attribute dont_touch of G41: signal is true;
	signal G42: std_logic; attribute dont_touch of G42: signal is true;
	signal G43: std_logic; attribute dont_touch of G43: signal is true;
	signal G44: std_logic; attribute dont_touch of G44: signal is true;
	signal G46: std_logic; attribute dont_touch of G46: signal is true;
	signal G47: std_logic; attribute dont_touch of G47: signal is true;
	signal G48: std_logic; attribute dont_touch of G48: signal is true;
	signal G49: std_logic; attribute dont_touch of G49: signal is true;
	signal G50: std_logic; attribute dont_touch of G50: signal is true;
	signal G51: std_logic; attribute dont_touch of G51: signal is true;
	signal G52: std_logic; attribute dont_touch of G52: signal is true;
	signal G53: std_logic; attribute dont_touch of G53: signal is true;
	signal G54: std_logic; attribute dont_touch of G54: signal is true;
	signal G55: std_logic; attribute dont_touch of G55: signal is true;
	signal G56: std_logic; attribute dont_touch of G56: signal is true;
	signal G57: std_logic; attribute dont_touch of G57: signal is true;
	signal G58: std_logic; attribute dont_touch of G58: signal is true;
	signal G59: std_logic; attribute dont_touch of G59: signal is true;
	signal G60: std_logic; attribute dont_touch of G60: signal is true;
	signal G61: std_logic; attribute dont_touch of G61: signal is true;
	signal G62: std_logic; attribute dont_touch of G62: signal is true;
	signal G63: std_logic; attribute dont_touch of G63: signal is true;
	signal G64: std_logic; attribute dont_touch of G64: signal is true;
	signal G66: std_logic; attribute dont_touch of G66: signal is true;
	signal G67: std_logic; attribute dont_touch of G67: signal is true;
	signal G68: std_logic; attribute dont_touch of G68: signal is true;
	signal G69: std_logic; attribute dont_touch of G69: signal is true;
	signal G70: std_logic; attribute dont_touch of G70: signal is true;
	signal G71: std_logic; attribute dont_touch of G71: signal is true;
	signal G72: std_logic; attribute dont_touch of G72: signal is true;
	signal G73: std_logic; attribute dont_touch of G73: signal is true;
	signal G74: std_logic; attribute dont_touch of G74: signal is true;
	signal G75: std_logic; attribute dont_touch of G75: signal is true;
	signal G76: std_logic; attribute dont_touch of G76: signal is true;
	signal G77: std_logic; attribute dont_touch of G77: signal is true;
	signal G78: std_logic; attribute dont_touch of G78: signal is true;
	signal G79: std_logic; attribute dont_touch of G79: signal is true;
	signal G80: std_logic; attribute dont_touch of G80: signal is true;
	signal G81: std_logic; attribute dont_touch of G81: signal is true;
	signal G82: std_logic; attribute dont_touch of G82: signal is true;
	signal G83: std_logic; attribute dont_touch of G83: signal is true;
	signal G84: std_logic; attribute dont_touch of G84: signal is true;
	signal G85: std_logic; attribute dont_touch of G85: signal is true;
	signal G86: std_logic; attribute dont_touch of G86: signal is true;
	signal G87: std_logic; attribute dont_touch of G87: signal is true;
	signal G88: std_logic; attribute dont_touch of G88: signal is true;
	signal G89: std_logic; attribute dont_touch of G89: signal is true;
	signal G90: std_logic; attribute dont_touch of G90: signal is true;
	signal G91: std_logic; attribute dont_touch of G91: signal is true;
	signal G92: std_logic; attribute dont_touch of G92: signal is true;
	signal G93: std_logic; attribute dont_touch of G93: signal is true;
	signal G94: std_logic; attribute dont_touch of G94: signal is true;
	signal G95: std_logic; attribute dont_touch of G95: signal is true;
	signal G96: std_logic; attribute dont_touch of G96: signal is true;
	signal G97: std_logic; attribute dont_touch of G97: signal is true;
	signal G98: std_logic; attribute dont_touch of G98: signal is true;
	signal G99: std_logic; attribute dont_touch of G99: signal is true;
	signal G100: std_logic; attribute dont_touch of G100: signal is true;
	signal G101: std_logic; attribute dont_touch of G101: signal is true;
	signal G102: std_logic; attribute dont_touch of G102: signal is true;
	signal G103: std_logic; attribute dont_touch of G103: signal is true;
	signal G104: std_logic; attribute dont_touch of G104: signal is true;
	signal G105: std_logic; attribute dont_touch of G105: signal is true;
	signal G106: std_logic; attribute dont_touch of G106: signal is true;
	signal G107: std_logic; attribute dont_touch of G107: signal is true;
	signal G108: std_logic; attribute dont_touch of G108: signal is true;
	signal G109: std_logic; attribute dont_touch of G109: signal is true;
	signal G110: std_logic; attribute dont_touch of G110: signal is true;
	signal G111: std_logic; attribute dont_touch of G111: signal is true;
	signal G112: std_logic; attribute dont_touch of G112: signal is true;
	signal G113: std_logic; attribute dont_touch of G113: signal is true;
	signal G114: std_logic; attribute dont_touch of G114: signal is true;
	signal G115: std_logic; attribute dont_touch of G115: signal is true;
	signal G116: std_logic; attribute dont_touch of G116: signal is true;
	signal G117: std_logic; attribute dont_touch of G117: signal is true;
	signal G118: std_logic; attribute dont_touch of G118: signal is true;
	signal G119: std_logic; attribute dont_touch of G119: signal is true;
	signal G120: std_logic; attribute dont_touch of G120: signal is true;
	signal G121: std_logic; attribute dont_touch of G121: signal is true;
	signal G122: std_logic; attribute dont_touch of G122: signal is true;
	signal G123: std_logic; attribute dont_touch of G123: signal is true;
	signal G124: std_logic; attribute dont_touch of G124: signal is true;
	signal G125: std_logic; attribute dont_touch of G125: signal is true;
	signal G126: std_logic; attribute dont_touch of G126: signal is true;
	signal G127: std_logic; attribute dont_touch of G127: signal is true;
	signal G128: std_logic; attribute dont_touch of G128: signal is true;
	signal G129: std_logic; attribute dont_touch of G129: signal is true;
	signal G130: std_logic; attribute dont_touch of G130: signal is true;
	signal G131: std_logic; attribute dont_touch of G131: signal is true;
	signal G132: std_logic; attribute dont_touch of G132: signal is true;
	signal G133: std_logic; attribute dont_touch of G133: signal is true;
	signal G134: std_logic; attribute dont_touch of G134: signal is true;
	signal G135: std_logic; attribute dont_touch of G135: signal is true;
	signal G136: std_logic; attribute dont_touch of G136: signal is true;
	signal G137: std_logic; attribute dont_touch of G137: signal is true;
	signal G138: std_logic; attribute dont_touch of G138: signal is true;
	signal G139: std_logic; attribute dont_touch of G139: signal is true;
	signal G140: std_logic; attribute dont_touch of G140: signal is true;
	signal G141: std_logic; attribute dont_touch of G141: signal is true;
	signal G142: std_logic; attribute dont_touch of G142: signal is true;
	signal G143: std_logic; attribute dont_touch of G143: signal is true;
	signal G144: std_logic; attribute dont_touch of G144: signal is true;
	signal G145: std_logic; attribute dont_touch of G145: signal is true;
	signal G146: std_logic; attribute dont_touch of G146: signal is true;
	signal G147: std_logic; attribute dont_touch of G147: signal is true;
	signal G148: std_logic; attribute dont_touch of G148: signal is true;
	signal G149: std_logic; attribute dont_touch of G149: signal is true;
	signal G150: std_logic; attribute dont_touch of G150: signal is true;
	signal G151: std_logic; attribute dont_touch of G151: signal is true;
	signal G152: std_logic; attribute dont_touch of G152: signal is true;
	signal G153: std_logic; attribute dont_touch of G153: signal is true;
	signal G154: std_logic; attribute dont_touch of G154: signal is true;
	signal G155: std_logic; attribute dont_touch of G155: signal is true;
	signal G156: std_logic; attribute dont_touch of G156: signal is true;
	signal G157: std_logic; attribute dont_touch of G157: signal is true;
	signal G158: std_logic; attribute dont_touch of G158: signal is true;
	signal G159: std_logic; attribute dont_touch of G159: signal is true;
	signal G160: std_logic; attribute dont_touch of G160: signal is true;
	signal G161: std_logic; attribute dont_touch of G161: signal is true;
	signal G162: std_logic; attribute dont_touch of G162: signal is true;
	signal G163: std_logic; attribute dont_touch of G163: signal is true;
	signal G164: std_logic; attribute dont_touch of G164: signal is true;
	signal G165: std_logic; attribute dont_touch of G165: signal is true;
	signal G166: std_logic; attribute dont_touch of G166: signal is true;
	signal G167: std_logic; attribute dont_touch of G167: signal is true;
	signal G168: std_logic; attribute dont_touch of G168: signal is true;
	signal G169: std_logic; attribute dont_touch of G169: signal is true;
	signal G170: std_logic; attribute dont_touch of G170: signal is true;
	signal G171: std_logic; attribute dont_touch of G171: signal is true;
	signal G172: std_logic; attribute dont_touch of G172: signal is true;
	signal G173: std_logic; attribute dont_touch of G173: signal is true;
	signal G174: std_logic; attribute dont_touch of G174: signal is true;
	signal G175: std_logic; attribute dont_touch of G175: signal is true;
	signal G176: std_logic; attribute dont_touch of G176: signal is true;
	signal G177: std_logic; attribute dont_touch of G177: signal is true;
	signal G178: std_logic; attribute dont_touch of G178: signal is true;
	signal G179: std_logic; attribute dont_touch of G179: signal is true;
	signal G180: std_logic; attribute dont_touch of G180: signal is true;
	signal G181: std_logic; attribute dont_touch of G181: signal is true;
	signal G182: std_logic; attribute dont_touch of G182: signal is true;
	signal G183: std_logic; attribute dont_touch of G183: signal is true;
	signal G184: std_logic; attribute dont_touch of G184: signal is true;
	signal G185: std_logic; attribute dont_touch of G185: signal is true;
	signal G186: std_logic; attribute dont_touch of G186: signal is true;
	signal G187: std_logic; attribute dont_touch of G187: signal is true;
	signal G188: std_logic; attribute dont_touch of G188: signal is true;
	signal G189: std_logic; attribute dont_touch of G189: signal is true;
	signal G190: std_logic; attribute dont_touch of G190: signal is true;
	signal G191: std_logic; attribute dont_touch of G191: signal is true;
	signal G192: std_logic; attribute dont_touch of G192: signal is true;
	signal G193: std_logic; attribute dont_touch of G193: signal is true;
	signal G194: std_logic; attribute dont_touch of G194: signal is true;
	signal G195: std_logic; attribute dont_touch of G195: signal is true;
	signal G196: std_logic; attribute dont_touch of G196: signal is true;
	signal G197: std_logic; attribute dont_touch of G197: signal is true;
	signal G198: std_logic; attribute dont_touch of G198: signal is true;
	signal G199: std_logic; attribute dont_touch of G199: signal is true;
	signal G200: std_logic; attribute dont_touch of G200: signal is true;
	signal G201: std_logic; attribute dont_touch of G201: signal is true;
	signal G202: std_logic; attribute dont_touch of G202: signal is true;
	signal G203: std_logic; attribute dont_touch of G203: signal is true;
	signal G204: std_logic; attribute dont_touch of G204: signal is true;
	signal G205: std_logic; attribute dont_touch of G205: signal is true;
	signal G206: std_logic; attribute dont_touch of G206: signal is true;
	signal G207: std_logic; attribute dont_touch of G207: signal is true;
	signal G208: std_logic; attribute dont_touch of G208: signal is true;
	signal G209: std_logic; attribute dont_touch of G209: signal is true;
	signal G210: std_logic; attribute dont_touch of G210: signal is true;
	signal G211: std_logic; attribute dont_touch of G211: signal is true;
	signal G212: std_logic; attribute dont_touch of G212: signal is true;
	signal G213: std_logic; attribute dont_touch of G213: signal is true;
	signal G214: std_logic; attribute dont_touch of G214: signal is true;
	signal G215: std_logic; attribute dont_touch of G215: signal is true;
	signal G216: std_logic; attribute dont_touch of G216: signal is true;
	signal G217: std_logic; attribute dont_touch of G217: signal is true;
	signal G218: std_logic; attribute dont_touch of G218: signal is true;
	signal G219: std_logic; attribute dont_touch of G219: signal is true;
	signal G220: std_logic; attribute dont_touch of G220: signal is true;
	signal G221: std_logic; attribute dont_touch of G221: signal is true;
	signal G222: std_logic; attribute dont_touch of G222: signal is true;
	signal G223: std_logic; attribute dont_touch of G223: signal is true;
	signal G224: std_logic; attribute dont_touch of G224: signal is true;
	signal G225: std_logic; attribute dont_touch of G225: signal is true;
	signal G226: std_logic; attribute dont_touch of G226: signal is true;
	signal G227: std_logic; attribute dont_touch of G227: signal is true;
	signal G228: std_logic; attribute dont_touch of G228: signal is true;
	signal G229: std_logic; attribute dont_touch of G229: signal is true;
	signal G230: std_logic; attribute dont_touch of G230: signal is true;
	signal G231: std_logic; attribute dont_touch of G231: signal is true;
	signal G232: std_logic; attribute dont_touch of G232: signal is true;
	signal G233: std_logic; attribute dont_touch of G233: signal is true;
	signal G234: std_logic; attribute dont_touch of G234: signal is true;
	signal G235: std_logic; attribute dont_touch of G235: signal is true;
	signal G236: std_logic; attribute dont_touch of G236: signal is true;
	signal G237: std_logic; attribute dont_touch of G237: signal is true;
	signal G238: std_logic; attribute dont_touch of G238: signal is true;
	signal G239: std_logic; attribute dont_touch of G239: signal is true;
	signal G240: std_logic; attribute dont_touch of G240: signal is true;
	signal G241: std_logic; attribute dont_touch of G241: signal is true;
	signal G242: std_logic; attribute dont_touch of G242: signal is true;
	signal G243: std_logic; attribute dont_touch of G243: signal is true;
	signal G244: std_logic; attribute dont_touch of G244: signal is true;
	signal G245: std_logic; attribute dont_touch of G245: signal is true;
	signal G246: std_logic; attribute dont_touch of G246: signal is true;
	signal G247: std_logic; attribute dont_touch of G247: signal is true;
	signal G248: std_logic; attribute dont_touch of G248: signal is true;
	signal G249: std_logic; attribute dont_touch of G249: signal is true;
	signal G250: std_logic; attribute dont_touch of G250: signal is true;
	signal G251: std_logic; attribute dont_touch of G251: signal is true;
	signal G252: std_logic; attribute dont_touch of G252: signal is true;
	signal G253: std_logic; attribute dont_touch of G253: signal is true;
	signal G254: std_logic; attribute dont_touch of G254: signal is true;
	signal G255: std_logic; attribute dont_touch of G255: signal is true;
	signal G256: std_logic; attribute dont_touch of G256: signal is true;
	signal G257: std_logic; attribute dont_touch of G257: signal is true;
	signal G258: std_logic; attribute dont_touch of G258: signal is true;
	signal G259: std_logic; attribute dont_touch of G259: signal is true;
	signal G260: std_logic; attribute dont_touch of G260: signal is true;
	signal G261: std_logic; attribute dont_touch of G261: signal is true;
	signal G262: std_logic; attribute dont_touch of G262: signal is true;
	signal G263: std_logic; attribute dont_touch of G263: signal is true;
	signal G264: std_logic; attribute dont_touch of G264: signal is true;
	signal G265: std_logic; attribute dont_touch of G265: signal is true;
	signal G266: std_logic; attribute dont_touch of G266: signal is true;
	signal G267: std_logic; attribute dont_touch of G267: signal is true;
	signal G268: std_logic; attribute dont_touch of G268: signal is true;
	signal G269: std_logic; attribute dont_touch of G269: signal is true;
	signal G270: std_logic; attribute dont_touch of G270: signal is true;
	signal G271: std_logic; attribute dont_touch of G271: signal is true;
	signal G272: std_logic; attribute dont_touch of G272: signal is true;
	signal G273: std_logic; attribute dont_touch of G273: signal is true;
	signal G274: std_logic; attribute dont_touch of G274: signal is true;
	signal G275: std_logic; attribute dont_touch of G275: signal is true;
	signal G276: std_logic; attribute dont_touch of G276: signal is true;
	signal G277: std_logic; attribute dont_touch of G277: signal is true;
	signal G278: std_logic; attribute dont_touch of G278: signal is true;
	signal G279: std_logic; attribute dont_touch of G279: signal is true;
	signal G280: std_logic; attribute dont_touch of G280: signal is true;
	signal G281: std_logic; attribute dont_touch of G281: signal is true;
	signal G282: std_logic; attribute dont_touch of G282: signal is true;
	signal G283: std_logic; attribute dont_touch of G283: signal is true;
	signal G284: std_logic; attribute dont_touch of G284: signal is true;
	signal G285: std_logic; attribute dont_touch of G285: signal is true;
	signal G286: std_logic; attribute dont_touch of G286: signal is true;
	signal G287: std_logic; attribute dont_touch of G287: signal is true;
	signal G288: std_logic; attribute dont_touch of G288: signal is true;
	signal G289: std_logic; attribute dont_touch of G289: signal is true;
	signal G290: std_logic; attribute dont_touch of G290: signal is true;
	signal G291: std_logic; attribute dont_touch of G291: signal is true;
	signal G292: std_logic; attribute dont_touch of G292: signal is true;
	signal G293: std_logic; attribute dont_touch of G293: signal is true;
	signal G294: std_logic; attribute dont_touch of G294: signal is true;
	signal G295: std_logic; attribute dont_touch of G295: signal is true;
	signal G296: std_logic; attribute dont_touch of G296: signal is true;
	signal G297: std_logic; attribute dont_touch of G297: signal is true;
	signal G298: std_logic; attribute dont_touch of G298: signal is true;
	signal G299: std_logic; attribute dont_touch of G299: signal is true;
	signal G300: std_logic; attribute dont_touch of G300: signal is true;
	signal G301: std_logic; attribute dont_touch of G301: signal is true;
	signal G302: std_logic; attribute dont_touch of G302: signal is true;
	signal G303: std_logic; attribute dont_touch of G303: signal is true;
	signal G304: std_logic; attribute dont_touch of G304: signal is true;
	signal G305: std_logic; attribute dont_touch of G305: signal is true;
	signal G306: std_logic; attribute dont_touch of G306: signal is true;
	signal G307: std_logic; attribute dont_touch of G307: signal is true;
	signal G308: std_logic; attribute dont_touch of G308: signal is true;
	signal G309: std_logic; attribute dont_touch of G309: signal is true;
	signal G310: std_logic; attribute dont_touch of G310: signal is true;
	signal G311: std_logic; attribute dont_touch of G311: signal is true;
	signal G312: std_logic; attribute dont_touch of G312: signal is true;
	signal G313: std_logic; attribute dont_touch of G313: signal is true;
	signal G314: std_logic; attribute dont_touch of G314: signal is true;
	signal G315: std_logic; attribute dont_touch of G315: signal is true;
	signal G316: std_logic; attribute dont_touch of G316: signal is true;
	signal G317: std_logic; attribute dont_touch of G317: signal is true;
	signal G318: std_logic; attribute dont_touch of G318: signal is true;
	signal G319: std_logic; attribute dont_touch of G319: signal is true;
	signal G320: std_logic; attribute dont_touch of G320: signal is true;
	signal G321: std_logic; attribute dont_touch of G321: signal is true;
	signal G322: std_logic; attribute dont_touch of G322: signal is true;
	signal G323: std_logic; attribute dont_touch of G323: signal is true;
	signal G324: std_logic; attribute dont_touch of G324: signal is true;
	signal G325: std_logic; attribute dont_touch of G325: signal is true;
	signal G326: std_logic; attribute dont_touch of G326: signal is true;
	signal G327: std_logic; attribute dont_touch of G327: signal is true;
	signal G328: std_logic; attribute dont_touch of G328: signal is true;
	signal G329: std_logic; attribute dont_touch of G329: signal is true;
	signal G330: std_logic; attribute dont_touch of G330: signal is true;
	signal G331: std_logic; attribute dont_touch of G331: signal is true;
	signal G332: std_logic; attribute dont_touch of G332: signal is true;
	signal G333: std_logic; attribute dont_touch of G333: signal is true;
	signal G334: std_logic; attribute dont_touch of G334: signal is true;
	signal G335: std_logic; attribute dont_touch of G335: signal is true;
	signal G336: std_logic; attribute dont_touch of G336: signal is true;
	signal G337: std_logic; attribute dont_touch of G337: signal is true;
	signal G338: std_logic; attribute dont_touch of G338: signal is true;
	signal G339: std_logic; attribute dont_touch of G339: signal is true;
	signal G340: std_logic; attribute dont_touch of G340: signal is true;
	signal G341: std_logic; attribute dont_touch of G341: signal is true;
	signal G342: std_logic; attribute dont_touch of G342: signal is true;
	signal G343: std_logic; attribute dont_touch of G343: signal is true;
	signal G344: std_logic; attribute dont_touch of G344: signal is true;
	signal G345: std_logic; attribute dont_touch of G345: signal is true;
	signal G346: std_logic; attribute dont_touch of G346: signal is true;
	signal G347: std_logic; attribute dont_touch of G347: signal is true;
	signal G348: std_logic; attribute dont_touch of G348: signal is true;
	signal G349: std_logic; attribute dont_touch of G349: signal is true;
	signal G350: std_logic; attribute dont_touch of G350: signal is true;
	signal G351: std_logic; attribute dont_touch of G351: signal is true;
	signal G352: std_logic; attribute dont_touch of G352: signal is true;
	signal G353: std_logic; attribute dont_touch of G353: signal is true;
	signal G354: std_logic; attribute dont_touch of G354: signal is true;
	signal G355: std_logic; attribute dont_touch of G355: signal is true;
	signal G356: std_logic; attribute dont_touch of G356: signal is true;
	signal G357: std_logic; attribute dont_touch of G357: signal is true;
	signal G358: std_logic; attribute dont_touch of G358: signal is true;
	signal G359: std_logic; attribute dont_touch of G359: signal is true;
	signal G360: std_logic; attribute dont_touch of G360: signal is true;
	signal G361: std_logic; attribute dont_touch of G361: signal is true;
	signal G362: std_logic; attribute dont_touch of G362: signal is true;
	signal G363: std_logic; attribute dont_touch of G363: signal is true;
	signal G364: std_logic; attribute dont_touch of G364: signal is true;
	signal G365: std_logic; attribute dont_touch of G365: signal is true;
	signal G366: std_logic; attribute dont_touch of G366: signal is true;
	signal G367: std_logic; attribute dont_touch of G367: signal is true;
	signal G368: std_logic; attribute dont_touch of G368: signal is true;
	signal G369: std_logic; attribute dont_touch of G369: signal is true;
	signal G370: std_logic; attribute dont_touch of G370: signal is true;
	signal G371: std_logic; attribute dont_touch of G371: signal is true;
	signal G372: std_logic; attribute dont_touch of G372: signal is true;
	signal G373: std_logic; attribute dont_touch of G373: signal is true;
	signal G374: std_logic; attribute dont_touch of G374: signal is true;
	signal G375: std_logic; attribute dont_touch of G375: signal is true;
	signal G376: std_logic; attribute dont_touch of G376: signal is true;
	signal G377: std_logic; attribute dont_touch of G377: signal is true;
	signal G378: std_logic; attribute dont_touch of G378: signal is true;
	signal G379: std_logic; attribute dont_touch of G379: signal is true;
	signal G380: std_logic; attribute dont_touch of G380: signal is true;
	signal G381: std_logic; attribute dont_touch of G381: signal is true;
	signal G382: std_logic; attribute dont_touch of G382: signal is true;
	signal G383: std_logic; attribute dont_touch of G383: signal is true;
	signal G384: std_logic; attribute dont_touch of G384: signal is true;
	signal G385: std_logic; attribute dont_touch of G385: signal is true;
	signal G386: std_logic; attribute dont_touch of G386: signal is true;
	signal G387: std_logic; attribute dont_touch of G387: signal is true;
	signal G388: std_logic; attribute dont_touch of G388: signal is true;
	signal G389: std_logic; attribute dont_touch of G389: signal is true;
	signal G390: std_logic; attribute dont_touch of G390: signal is true;
	signal G391: std_logic; attribute dont_touch of G391: signal is true;
	signal G392: std_logic; attribute dont_touch of G392: signal is true;
	signal G393: std_logic; attribute dont_touch of G393: signal is true;
	signal G394: std_logic; attribute dont_touch of G394: signal is true;
	signal G395: std_logic; attribute dont_touch of G395: signal is true;
	signal G396: std_logic; attribute dont_touch of G396: signal is true;
	signal G397: std_logic; attribute dont_touch of G397: signal is true;
	signal G398: std_logic; attribute dont_touch of G398: signal is true;
	signal G399: std_logic; attribute dont_touch of G399: signal is true;
	signal G400: std_logic; attribute dont_touch of G400: signal is true;
	signal G401: std_logic; attribute dont_touch of G401: signal is true;
	signal G402: std_logic; attribute dont_touch of G402: signal is true;
	signal G403: std_logic; attribute dont_touch of G403: signal is true;
	signal G404: std_logic; attribute dont_touch of G404: signal is true;
	signal G405: std_logic; attribute dont_touch of G405: signal is true;
	signal G406: std_logic; attribute dont_touch of G406: signal is true;
	signal G407: std_logic; attribute dont_touch of G407: signal is true;
	signal G408: std_logic; attribute dont_touch of G408: signal is true;
	signal G409: std_logic; attribute dont_touch of G409: signal is true;
	signal G410: std_logic; attribute dont_touch of G410: signal is true;
	signal G411: std_logic; attribute dont_touch of G411: signal is true;
	signal G412: std_logic; attribute dont_touch of G412: signal is true;
	signal G413: std_logic; attribute dont_touch of G413: signal is true;
	signal G414: std_logic; attribute dont_touch of G414: signal is true;
	signal G415: std_logic; attribute dont_touch of G415: signal is true;
	signal G416: std_logic; attribute dont_touch of G416: signal is true;
	signal G417: std_logic; attribute dont_touch of G417: signal is true;
	signal G418: std_logic; attribute dont_touch of G418: signal is true;
	signal G419: std_logic; attribute dont_touch of G419: signal is true;
	signal G420: std_logic; attribute dont_touch of G420: signal is true;
	signal G421: std_logic; attribute dont_touch of G421: signal is true;
	signal G422: std_logic; attribute dont_touch of G422: signal is true;
	signal G423: std_logic; attribute dont_touch of G423: signal is true;
	signal G424: std_logic; attribute dont_touch of G424: signal is true;
	signal G425: std_logic; attribute dont_touch of G425: signal is true;
	signal G426: std_logic; attribute dont_touch of G426: signal is true;
	signal G427: std_logic; attribute dont_touch of G427: signal is true;
	signal G428: std_logic; attribute dont_touch of G428: signal is true;
	signal G429: std_logic; attribute dont_touch of G429: signal is true;
	signal G430: std_logic; attribute dont_touch of G430: signal is true;
	signal G431: std_logic; attribute dont_touch of G431: signal is true;
	signal G432: std_logic; attribute dont_touch of G432: signal is true;
	signal G433: std_logic; attribute dont_touch of G433: signal is true;
	signal G434: std_logic; attribute dont_touch of G434: signal is true;
	signal G435: std_logic; attribute dont_touch of G435: signal is true;
	signal G436: std_logic; attribute dont_touch of G436: signal is true;
	signal G437: std_logic; attribute dont_touch of G437: signal is true;
	signal G438: std_logic; attribute dont_touch of G438: signal is true;
	signal G439: std_logic; attribute dont_touch of G439: signal is true;
	signal G440: std_logic; attribute dont_touch of G440: signal is true;
	signal G441: std_logic; attribute dont_touch of G441: signal is true;
	signal G442: std_logic; attribute dont_touch of G442: signal is true;
	signal G443: std_logic; attribute dont_touch of G443: signal is true;
	signal G444: std_logic; attribute dont_touch of G444: signal is true;
	signal G445: std_logic; attribute dont_touch of G445: signal is true;
	signal G446: std_logic; attribute dont_touch of G446: signal is true;
	signal G447: std_logic; attribute dont_touch of G447: signal is true;
	signal G448: std_logic; attribute dont_touch of G448: signal is true;
	signal G449: std_logic; attribute dont_touch of G449: signal is true;
	signal G450: std_logic; attribute dont_touch of G450: signal is true;
	signal G451: std_logic; attribute dont_touch of G451: signal is true;
	signal G452: std_logic; attribute dont_touch of G452: signal is true;
	signal G453: std_logic; attribute dont_touch of G453: signal is true;
	signal G454: std_logic; attribute dont_touch of G454: signal is true;
	signal G455: std_logic; attribute dont_touch of G455: signal is true;
	signal G456: std_logic; attribute dont_touch of G456: signal is true;
	signal G457: std_logic; attribute dont_touch of G457: signal is true;
	signal G458: std_logic; attribute dont_touch of G458: signal is true;
	signal G459: std_logic; attribute dont_touch of G459: signal is true;
	signal G460: std_logic; attribute dont_touch of G460: signal is true;
	signal G461: std_logic; attribute dont_touch of G461: signal is true;
	signal G462: std_logic; attribute dont_touch of G462: signal is true;
	signal G463: std_logic; attribute dont_touch of G463: signal is true;
	signal G464: std_logic; attribute dont_touch of G464: signal is true;
	signal G465: std_logic; attribute dont_touch of G465: signal is true;
	signal G468: std_logic; attribute dont_touch of G468: signal is true;
	signal G469: std_logic; attribute dont_touch of G469: signal is true;
	signal G470: std_logic; attribute dont_touch of G470: signal is true;
	signal G471: std_logic; attribute dont_touch of G471: signal is true;
	signal G472: std_logic; attribute dont_touch of G472: signal is true;
	signal G473: std_logic; attribute dont_touch of G473: signal is true;
	signal G474: std_logic; attribute dont_touch of G474: signal is true;
	signal G475: std_logic; attribute dont_touch of G475: signal is true;
	signal G476: std_logic; attribute dont_touch of G476: signal is true;
	signal G477: std_logic; attribute dont_touch of G477: signal is true;
	signal G478: std_logic; attribute dont_touch of G478: signal is true;
	signal G479: std_logic; attribute dont_touch of G479: signal is true;
	signal G480: std_logic; attribute dont_touch of G480: signal is true;
	signal G482: std_logic; attribute dont_touch of G482: signal is true;
	signal G483: std_logic; attribute dont_touch of G483: signal is true;
	signal G484: std_logic; attribute dont_touch of G484: signal is true;
	signal G485: std_logic; attribute dont_touch of G485: signal is true;
	signal G486: std_logic; attribute dont_touch of G486: signal is true;
	signal G487: std_logic; attribute dont_touch of G487: signal is true;
	signal G488: std_logic; attribute dont_touch of G488: signal is true;
	signal G489: std_logic; attribute dont_touch of G489: signal is true;
	signal G490: std_logic; attribute dont_touch of G490: signal is true;
	signal G491: std_logic; attribute dont_touch of G491: signal is true;
	signal G492: std_logic; attribute dont_touch of G492: signal is true;
	signal G493: std_logic; attribute dont_touch of G493: signal is true;
	signal G494: std_logic; attribute dont_touch of G494: signal is true;
	signal G495: std_logic; attribute dont_touch of G495: signal is true;
	signal G496: std_logic; attribute dont_touch of G496: signal is true;
	signal G497: std_logic; attribute dont_touch of G497: signal is true;
	signal G498: std_logic; attribute dont_touch of G498: signal is true;
	signal G499: std_logic; attribute dont_touch of G499: signal is true;
	signal G500: std_logic; attribute dont_touch of G500: signal is true;
	signal G501: std_logic; attribute dont_touch of G501: signal is true;
	signal G502: std_logic; attribute dont_touch of G502: signal is true;
	signal G503: std_logic; attribute dont_touch of G503: signal is true;
	signal G504: std_logic; attribute dont_touch of G504: signal is true;
	signal G505: std_logic; attribute dont_touch of G505: signal is true;
	signal G506: std_logic; attribute dont_touch of G506: signal is true;
	signal G507: std_logic; attribute dont_touch of G507: signal is true;
	signal G508: std_logic; attribute dont_touch of G508: signal is true;
	signal G509: std_logic; attribute dont_touch of G509: signal is true;
	signal G510: std_logic; attribute dont_touch of G510: signal is true;
	signal G511: std_logic; attribute dont_touch of G511: signal is true;
	signal G512: std_logic; attribute dont_touch of G512: signal is true;
	signal G513: std_logic; attribute dont_touch of G513: signal is true;
	signal G514: std_logic; attribute dont_touch of G514: signal is true;
	signal G515: std_logic; attribute dont_touch of G515: signal is true;
	signal G516: std_logic; attribute dont_touch of G516: signal is true;
	signal G517: std_logic; attribute dont_touch of G517: signal is true;
	signal G518: std_logic; attribute dont_touch of G518: signal is true;
	signal G519: std_logic; attribute dont_touch of G519: signal is true;
	signal G520: std_logic; attribute dont_touch of G520: signal is true;
	signal G521: std_logic; attribute dont_touch of G521: signal is true;
	signal G522: std_logic; attribute dont_touch of G522: signal is true;
	signal G523: std_logic; attribute dont_touch of G523: signal is true;
	signal G524: std_logic; attribute dont_touch of G524: signal is true;
	signal G525: std_logic; attribute dont_touch of G525: signal is true;
	signal G526: std_logic; attribute dont_touch of G526: signal is true;
	signal G527: std_logic; attribute dont_touch of G527: signal is true;
	signal G528: std_logic; attribute dont_touch of G528: signal is true;
	signal G529: std_logic; attribute dont_touch of G529: signal is true;
	signal G531: std_logic; attribute dont_touch of G531: signal is true;
	signal G533: std_logic; attribute dont_touch of G533: signal is true;
	signal G534: std_logic; attribute dont_touch of G534: signal is true;
	signal G536: std_logic; attribute dont_touch of G536: signal is true;
	signal G538: std_logic; attribute dont_touch of G538: signal is true;
	signal G540: std_logic; attribute dont_touch of G540: signal is true;
	signal G541: std_logic; attribute dont_touch of G541: signal is true;
	signal G543: std_logic; attribute dont_touch of G543: signal is true;
	signal G544: std_logic; attribute dont_touch of G544: signal is true;
	signal G545: std_logic; attribute dont_touch of G545: signal is true;
	signal G553: std_logic; attribute dont_touch of G553: signal is true;
	signal G554: std_logic; attribute dont_touch of G554: signal is true;
	signal II156: std_logic; attribute dont_touch of II156: signal is true;
	signal II218: std_logic; attribute dont_touch of II218: signal is true;
	signal II249: std_logic; attribute dont_touch of II249: signal is true;
	signal II272: std_logic; attribute dont_touch of II272: signal is true;
	signal II276: std_logic; attribute dont_touch of II276: signal is true;
	signal II280: std_logic; attribute dont_touch of II280: signal is true;
	signal II287: std_logic; attribute dont_touch of II287: signal is true;
	signal II295: std_logic; attribute dont_touch of II295: signal is true;
	signal II316: std_logic; attribute dont_touch of II316: signal is true;
	signal II327: std_logic; attribute dont_touch of II327: signal is true;
	signal II330: std_logic; attribute dont_touch of II330: signal is true;
	signal II352: std_logic; attribute dont_touch of II352: signal is true;
	signal II371: std_logic; attribute dont_touch of II371: signal is true;
	signal II374: std_logic; attribute dont_touch of II374: signal is true;
	signal II386: std_logic; attribute dont_touch of II386: signal is true;
	signal II493: std_logic; attribute dont_touch of II493: signal is true;
	signal II502: std_logic; attribute dont_touch of II502: signal is true;
	signal II529: std_logic; attribute dont_touch of II529: signal is true;
	signal II536: std_logic; attribute dont_touch of II536: signal is true;
	signal II573: std_logic; attribute dont_touch of II573: signal is true;
	signal II576: std_logic; attribute dont_touch of II576: signal is true;
	signal II624: std_logic; attribute dont_touch of II624: signal is true;
	signal II631: std_logic; attribute dont_touch of II631: signal is true;
	signal II662: std_logic; attribute dont_touch of II662: signal is true;
	signal II692: std_logic; attribute dont_touch of II692: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			G29<=G502;
			G30<=G503;
			G31<=G504;
			G32<=G505;
			G33<=G506;
			G34<=G507;
			G35<=G508;
			G36<=G509;
			G37<=G510;
			G38<=G511;
			G39<=G512;
			G40<=G513;
			G41<=G514;
			G42<=G515;
			G43<=G516;
			G44<=G517;
			G45<=G518;
			G46<=G519;
		end if;
	end process;
	G50<= not G49;
	G55<= not G54;
	G59<= not G58;
	G64<= not G63;
	G67<= not G44;
	G70<= not G43;
	G72<= not G71;
	G75<= not G74;
	G78<= not G77;
	G87<= not G86;
	G90<= not G89;
	G98<= not G97;
	G99<= not G29;
	G107<= not G456;
	G123<= not G122;
	G124<= not G206;
	G125<= not G40;
	G130<= not G9;
	G132<= not G42;
	G135<= not G134;
	G140<= not G33;
	G149<= not II529;
	G153<= not G522;
	G160<= not G161;
	G165<= not G529;
	G167<= not G168;
	G170<= not G171;
	G172<= not G171;
	G173<= not G495;
	G174<= not G496;
	G177<= not G357;
	G180<= not G181;
	G192<= not G193;
	G199<= not G200;
	G203<= not G204;
	G207<= not G208;
	G212<= not G213;
	G214<= not G215;
	G221<= not G222;
	G223<= not G224;
	G228<= not G524;
	G231<= not G232;
	G234<= not G235;
	G236<= not G274;
	G265<= not G50;
	G272<= not G271;
	G275<= not G274;
	G282<= not G281;
	G299<= not II352;
	G303<= not II624;
	G309<= not II280;
	G332<= not II276;
	G333<= not II218;
	G334<= not II156;
	G335<= not II371;
	G336<= not II631;
	G347<= not II287;
	G369<= not II316;
	G370<= not II249;
	G403<= not II573;
	G404<= not II493;
	G405<= not II662;
	G414<= not II386;
	G432<= not II692;
	G435<= not II327;
	G441<= not II330;
	G446<= not II536;
	G447<= not II576;
	G456<= not II374;
	G458<= not II272;
	G459<= not II295;
	G468<= not II502;
	G475<= not G57;
	G476<= not G30;
	G477<= not G276;
	G478<= not G279;
	G479<= not G194;
	G480<= not G179;
	G482<= not G241;
	G483<= not G182;
	G484<= not G30;
	G485<= not G276;
	G486<= not G68;
	G487<= not G534;
	G488<= not G172;
	G489<= not G273;
	G490<= not G190;
	G491<= not G194;
	G492<= not G62;
	G493<= not G544;
	G494<= not G173;
	G495<= not G273;
	G496<= not G188;
	G497<= not G205;
	G498<= not G195;
	G499<= not G280;
	G500<= not G173;
	G501<= not G156;
	G520<= not G0;
	G521<= not G1;
	G522<= not G2;
	G524<= not G3;
	G525<= not G526;
	G527<= not G4;
	G528<= not G5;
	G529<= not G6;
	G531<= not G7;
	G533<= not G8;
	G536<= not G9;
	G538<= not G10;
	G540<= not G11;
	G541<= not G12;
	G543<= not G13;
	G545<= not G544;
	G546<= not G41;
	G554<= not G553;
	II156<= not G4;
	II218<= not G528;
	II249<= not G538;
	II272<= not G209;
	II276<= not G238;
	II280<= not G272;
	II287<= not G135;
	II295<= not G198;
	II316<= not G239;
	II327<= not G135;
	II330<= not G236;
	II352<= not G77;
	II371<= not G1;
	II374<= not G520;
	II386<= not G199;
	II493<= not G218;
	II502<= not G124;
	II529<= not G468;
	II536<= not G79;
	II573<= not G176;
	II576<= not G175;
	II624<= not G120;
	II631<= not G188;
	II662<= not G174;
	II692<= not G145;
	G81<=G288 and G240;
	G283<=G122 and G219;
	G289<=G2 and G119 and G156;
	G290<=G117 and G135 and G157;
	G291<=G138 and G155;
	G304<=G52 and G158;
	G306<=G524 and G78;
	G307<=G6 and G104;
	G308<=G5 and G151;
	G311<=G0 and G178 and G179;
	G312<=G180 and G182;
	G315<=G250 and G251;
	G317<=G159 and G245;
	G321<=G90 and G50;
	G322<=G522 and G105 and G196;
	G323<=G2 and G144;
	G324<=G522 and G183;
	G327<=G4 and G39 and G157;
	G328<=G5 and G102 and G155;
	G329<=G150 and G156;
	G330<=G248 and G249;
	G331<=G213 and G257;
	G337<=G270 and G167;
	G338<=G202 and G203;
	G339<=G533 and G199 and G209;
	G340<=G8 and G270;
	G341<=G531 and G118;
	G342<=G73 and G197;
	G343<=G2 and G528 and G147;
	G344<=G111 and G189 and G195;
	G346<=G2 and G82;
	G348<=G97 and G55;
	G349<=G6 and G108;
	G351<=G524 and G169 and G221 and G234;
	G352<=G8 and G135 and G37 and G164;
	G353<=G11 and G92 and G163;
	G354<=G0 and G214;
	G357<=G265 and G232;
	G358<=G7 and G83;
	G359<=G6 and G31;
	G360<=G8 and G106;
	G361<=G6 and G202;
	G362<=G129 and G77;
	G363<=G77 and G205;
	G364<=G2 and G109;
	G365<=G282 and G137 and G156;
	G366<=G125 and G155;
	G367<=G126 and G157;
	G371<=G161 and G168 and G267;
	G372<=G116 and G275 and G155;
	G373<=G34 and G160;
	G376<=G533 and G75;
	G377<=G90 and G56;
	G378<=G89 and G50;
	G379<=G9 and G211;
	G380<=G6 and G93;
	G382<=G9 and G100 and G34;
	G383<=G131 and G155;
	G385<=G529 and G7 and G49;
	G386<=G536 and G85;
	G387<=G6 and G274 and G75;
	G388<=G11 and G114;
	G392<=G132 and G155;
	G393<=G127 and G34;
	G396<=G76 and G272 and G155;
	G397<=G101 and G98 and G157;
	G398<=G94 and G156 and G158;
	G399<=G520 and G1;
	G400<=G0 and G277;
	G401<=G2 and G110 and G155;
	G402<=G154 and G183;
	G406<=G87 and G172;
	G410<=G1 and G205;
	G411<=G48 and G59;
	G412<=G3 and G207;
	G413<=G197 and G201;
	G415<=G146 and G142 and G165;
	G416<=G61 and G167;
	G417<=G13 and G282 and G70;
	G418<=G524 and G60 and G172;
	G422<=G0 and G80 and G155;
	G423<=G541 and G128;
	G424<=G78 and G174 and G177;
	G425<=G146 and G176;
	G426<=G37 and G162 and G38;
	G427<=G541 and G95 and G165;
	G428<=G212 and G227;
	G429<=G51 and G225;
	G430<=G177 and G196;
	G431<=G524 and G67;
	G433<=G91 and G154;
	G434<=G165 and G231;
	G436<=G123 and G77;
	G437<=G66 and G229;
	G438<=G8 and G146 and G133;
	G439<=G174 and G175;
	G440<=G38 and G234;
	G442<=G541 and G121;
	G443<=G47 and G162;
	G444<=G64 and G78 and G211;
	G445<=G53 and G225;
	G448<=G139 and G153;
	G449<=G88 and G154;
	G451<=G541 and G554 and G187;
	G452<=G526 and G184;
	G453<=G545 and G186;
	G457<=G4 and G107;
	G460<=G2 and G81 and G115;
	G461<=G529 and G531;
	G462<=G192 and G538;
	G463<=G521 and G148;
	G469<=G163 and G3;
	G470<=G528 and G149;
	G471<=G191 and G103 and G112;
	G472<=G136 and G9 and G190;
	G473<=G11 and G143;
	G474<=G242 and G77;
	G511<=G163 and G164;
	G48<= not (G407 and G408 and G409);
	G49<= not (G9 and G538);
	G51<= not (G260 and G237);
	G52<= not (G298 and G299 and G219);
	G53<= not (G264 and G237);
	G54<= not (G4 and G6);
	G56<= not (G374 and G375);
	G57<= not (G0 and G2);
	G58<= not (G1 and G3);
	G62<= not (G534 and G32);
	G63<= not (G75 and G8);
	G66<= not (G129 and G101);
	G68<= not (G302 and G528);
	G69<= not (G419 and G420 and G233);
	G71<= not (G8 and G10);
	G74<= not (G9 and G11);
	G76<= not (G0 and G3);
	G77<= not (G4 and G528);
	G80<= not (G421 and G226 and G256);
	G82<= not (G334 and G335);
	G83<= not (G355 and G356);
	G84<= not (G369 and G370);
	G85<= not (G384 and G239);
	G86<= not (G55 and G3);
	G89<= not (G531 and G8);
	G94<= not (G261 and G181 and G262);
	G96<= not (G313 and G314);
	G97<= not (G2 and G5);
	G100<= not (G381 and G220);
	G101<= not (G3 and G4);
	G102<= not (G320 and G266 and G210);
	G103<= not (G529 and G7 and G30);
	G104<= not (G122 and G238 and G240);
	G109<= not (G269 and G219);
	G111<= not (G213 and G217);
	G112<= not (G8 and G31);
	G113<= not (G389 and G390);
	G116<= not (G6 and G9);
	G117<= not (G2 and G4);
	G119<= not (G284 and G285);
	G120<= not (G294 and G295);
	G122<= not (G522 and G3);
	G127<= not (G391 and G268);
	G129<= not (G527 and G5);
	G134<= not (G3 and G5);
	G136<= not (G222 and G224);
	G138<= not (G465 and G263);
	G143<= not (G258 and G193 and G259);
	G144<= not (G215 and G252 and G253);
	G148<= not (G454 and G455 and G0);
	G151<= not (G305 and G200);
	G159<= not (G6 and G155);
	G161<= not (G316 and G72);
	G166<= not (G7 and G50);
	G168<= not (G75 and G221);
	G171<= not (G553 and G187);
	G181<= not (G2 and G78);
	G185<= not (G525 and G184);
	G200<= not (G527 and G529);
	G204<= not (G521 and G87);
	G206<= not (G287 and G524);
	G208<= not (G68 and G229);
	G210<= not (G520 and G272);
	G213<= not (G64 and G275);
	G215<= not (G135 and G55 and G212);
	G217<= not (G50 and G230);
	G219<= not (G524 and G55);
	G220<= not (G7 and G71);
	G222<= not (G533 and G10);
	G226<= not (G527 and G59);
	G232<= not (G536 and G164);
	G233<= not (G522 and G135);
	G235<= not (G6 and G536);
	G237<= not (G10 and G75 and G201);
	G238<= not (G2 and G524);
	G239<= not (G7 and G533);
	G240<= not (G4 and G134);
	G243<= not (G368 and G275 and G34);
	G245<= not (G8 and G34);
	G246<= not (G544 and G186);
	G248<= not (G529 and G36);
	G249<= not (G11 and G273 and G201);
	G250<= not (G13 and G523);
	G251<= not (G543 and G32);
	G252<= not (G3 and G11 and G35 and G216);
	G253<= not (G87 and G218);
	G254<= not (G1 and G152);
	G255<= not (G309 and G2 and G529);
	G256<= not (G4 and G69);
	G257<= not (G538 and G230);
	G258<= not (G464 and G103 and G223);
	G259<= not (G130 and G225);
	G260<= not (G528 and G529 and G191);
	G262<= not (G527 and G278);
	G263<= not (G0 and G99);
	G264<= not (G227 and G241);
	G266<= not (G524 and G96);
	G267<= not (G536 and G84);
	G268<= not (G11 and G113);
	G270<= not (G345 and G204);
	G271<= not (G1 and G4);
	G273<= not (G325 and G326);
	G274<= not (G7 and G10);
	G276<= not (G3 and G543 and G140);
	G277<= not (G394 and G395 and G81);
	G278<= not (G332 and G333);
	G280<= not (G46 and G247);
	G281<= not (G523 and G534);
	G503<= not (G286 and G538);
	G504<= not (G292 and G293);
	G505<= not (G300 and G301 and G181);
	G508<= not (G318 and G319);
	G510<= not (G350 and G235);
	G512<= not (G310 and G233);
	G518<= not (G450 and G185 and G246);
	G523<= not (G254 and G255 and G208);
	G526<= not (G1 and G2 and G141);
	G534<= not (G296 and G297 and G166);
	G542<= not (G243 and G244 and G279);
	G47<=G440 or G441;
	G60<=G413 or G414;
	G61<=G405 or G406;
	G73<=G339 or G340;
	G79<=G444 or G445;
	G88<=G446 or G447;
	G91<=G430 or G431;
	G92<=G351 or G352;
	G93<=G376 or G377 or G378;
	G95<=G424 or G425;
	G105<=G321 or G273;
	G106<=G358 or G359;
	G108<=G346 or G347;
	G110<=G399 or G400;
	G114<=G385 or G386;
	G115<=G457 or G458 or G459;
	G118<=G337 or G338;
	G121<=G438 or G439;
	G126<=G363 or G364;
	G128<=G415 or G416 or G417 or G418;
	G131<=G379 or G380;
	G133<=G434 or G435;
	G137<=G348 or G349;
	G139<=G442 or G443;
	G141<=G353 or G354;
	G142<=G403 or G404;
	G145<=G426 or G427;
	G146<=G336 or G170;
	G147<=G341 or G342;
	G150<=G303 or G304;
	G152<=G306 or G307 or G308;
	G193<=G6 or G30;
	G224<=G533 or G31;
	G242<=G469 or G470;
	G244<=G371 or G159;
	G261<=G283 or G528;
	G269<=G362 or G529;
	G279<=G317 or G166;
	G284<=G528 or G272 or G281;
	G285<=G5 or G479;
	G286<=G9 or G540;
	G287<=G522 or G81;
	G288<=G1 or G528;
	G292<=G538 or G75;
	G293<=G7 or G540;
	G294<=G1 or G117 or G281;
	G295<=G122 or G491;
	G296<=G89 or G484;
	G297<=G64 or G274;
	G298<=G5 or G497;
	G300<=G87 or G97;
	G301<=G122 or G486;
	G302<=G4 or G529;
	G305<=G524 or G55;
	G310<=G522 or G135;
	G313<=G521 or G475;
	G314<=G527 or G57;
	G316<=G531 or G536;
	G318<=G6 or G8 or G232;
	G319<=G529 or G489;
	G320<=G76 or G272;
	G325<=G7 or G536 or G222;
	G326<=G533 or G232;
	G345<=G529 or G226;
	G350<=G6 or G536;
	G355<=G11 or G116;
	G356<=G6 or G476;
	G368<=G533 or G536;
	G374<=G536 or G538;
	G375<=G10 or G540;
	G381<=G7 or G71;
	G384<=G529 or G71;
	G389<=G9 or G274;
	G390<=G89 or G50;
	G391<=G74 or G220;
	G394<=G5 or G58;
	G395<=G4 or G134;
	G407<=G6 or G117;
	G408<=G529 or G77;
	G409<=G528 or G55;
	G419<=G3 or G5;
	G420<=G522 or G59;
	G421<=G521 or G2 or G228;
	G450<=G12 or G171;
	G454<=G122 or G77;
	G455<=G78 or G206;
	G464<=G72 or G536;
	G465<=G524 or G210;
	G530<=G401 or G402;
	G532<=G422 or G423;
	G535<=G432 or G433;
	G537<=G448 or G449;
	G539<=G451 or G452 or G453;
	G544<=G343 or G344;
	G547<=G382 or G383;
	G548<=G392 or G393;
	G549<=G396 or G397 or G398 or G477;
	G550<=G289 or G290 or G291 or G485;
	G551<=G327 or G328 or G329;
	G552<=G365 or G366 or G367;
	G553<=G322 or G323 or G324;
	G154<= not (G12 or G488);
	G155<= not (G13 or G480);
	G156<= not (G12 or G543);
	G157<= not (G13 or G483);
	G158<= not (G521 or G281);
	G162<= not (G185 or G498);
	G163<= not (G0 or G4);
	G164<= not (G531 or G10);
	G169<= not (G5 or G7);
	G175<= not (G86 or G500);
	G176<= not (G4 or G494);
	G178<= not (G521 or G4);
	G179<= not (G541 or G280);
	G182<= not (G12 or G62);
	G183<= not (G330 or G3);
	G184<= not (G541 or G13 or G499);
	G186<= not (G282 or G501);
	G187<= not (G13 or G492);
	G188<= not (G543 or G493);
	G189<= not (G522 or G54);
	G190<= not (G7 or G11);
	G191<= not (G9 or G482);
	G194<= not (G281 or G271);
	G195<= not (G521 or G134);
	G196<= not (G5 or G540 or G86);
	G197<= not (G540 or G232);
	G198<= not (G520 or G3);
	G201<= not (G528 or G54);
	G202<= not (G10 or G63);
	G205<= not (G529 or G122);
	G209<= not (G1 or G524);
	G211<= not (G6 or G274);
	G216<= not (G4 or G5);
	G218<= not (G528 or G217);
	G225<= not (G7 or G8);
	G227<= not (G5 or G200);
	G229<= not (G1 or G522);
	G230<= not (G8 or G490);
	G241<= not (G10 or G11);
	G247<= not (G471 or G472 or G473 or G474);
	G502<= not (G436 or G437);
	G506<= not (G311 or G312);
	G507<= not (G315 or G12 or G487);
	G509<= not (G331 or G5);
	G513<= not (G360 or G361);
	G514<= not (G372 or G373 or G478);
	G515<= not (G387 or G388);
	G516<= not (G410 or G411 or G412);
	G517<= not (G428 or G429);
	G519<= not (G460 or G461 or G462 or G463);
end RTL;
