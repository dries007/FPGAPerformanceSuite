-- File created by Bench2VHDL
-- Name: s5378
-- File: bench/s5378.bench
-- Timestamp: 2019-05-21T22:08:29.612803
--
-- Original File
-- =============
--	# s5378
--	# 35 inputs
--	# 49 outputs
--	# 179 D-type flipflops
--	# 1775 inverters
--	# 1004 gates (0 ANDs + 0 NANDs + 239 ORs + 765 NORs)
--	
--	INPUT(n3065gat)
--	INPUT(n3066gat)
--	INPUT(n3067gat)
--	INPUT(n3068gat)
--	INPUT(n3069gat)
--	INPUT(n3070gat)
--	INPUT(n3071gat)
--	INPUT(n3072gat)
--	INPUT(n3073gat)
--	INPUT(n3074gat)
--	INPUT(n3075gat)
--	INPUT(n3076gat)
--	INPUT(n3077gat)
--	INPUT(n3078gat)
--	INPUT(n3079gat)
--	INPUT(n3080gat)
--	INPUT(n3081gat)
--	INPUT(n3082gat)
--	INPUT(n3083gat)
--	INPUT(n3084gat)
--	INPUT(n3085gat)
--	INPUT(n3086gat)
--	INPUT(n3087gat)
--	INPUT(n3088gat)
--	INPUT(n3089gat)
--	INPUT(n3090gat)
--	INPUT(n3091gat)
--	INPUT(n3092gat)
--	INPUT(n3093gat)
--	INPUT(n3094gat)
--	INPUT(n3095gat)
--	INPUT(n3097gat)
--	INPUT(n3098gat)
--	INPUT(n3099gat)
--	INPUT(n3100gat)
--	
--	OUTPUT(n3104gat)
--	OUTPUT(n3105gat)
--	OUTPUT(n3106gat)
--	OUTPUT(n3107gat)
--	OUTPUT(n3108gat)
--	OUTPUT(n3109gat)
--	OUTPUT(n3110gat)
--	OUTPUT(n3111gat)
--	OUTPUT(n3112gat)
--	OUTPUT(n3113gat)
--	OUTPUT(n3114gat)
--	OUTPUT(n3115gat)
--	OUTPUT(n3116gat)
--	OUTPUT(n3117gat)
--	OUTPUT(n3118gat)
--	OUTPUT(n3119gat)
--	OUTPUT(n3120gat)
--	OUTPUT(n3121gat)
--	OUTPUT(n3122gat)
--	OUTPUT(n3123gat)
--	OUTPUT(n3124gat)
--	OUTPUT(n3125gat)
--	OUTPUT(n3126gat)
--	OUTPUT(n3127gat)
--	OUTPUT(n3128gat)
--	OUTPUT(n3129gat)
--	OUTPUT(n3130gat)
--	OUTPUT(n3131gat)
--	OUTPUT(n3132gat)
--	OUTPUT(n3133gat)
--	OUTPUT(n3134gat)
--	OUTPUT(n3135gat)
--	OUTPUT(n3136gat)
--	OUTPUT(n3137gat)
--	OUTPUT(n3138gat)
--	OUTPUT(n3139gat)
--	OUTPUT(n3140gat)
--	OUTPUT(n3141gat)
--	OUTPUT(n3142gat)
--	OUTPUT(n3143gat)
--	OUTPUT(n3144gat)
--	OUTPUT(n3145gat)
--	OUTPUT(n3146gat)
--	OUTPUT(n3147gat)
--	OUTPUT(n3148gat)
--	OUTPUT(n3149gat)
--	OUTPUT(n3150gat)
--	OUTPUT(n3151gat)
--	OUTPUT(n3152gat)
--	
--	n673gat = DFF(n2897gat)
--	n398gat = DFF(n2782gat)
--	n402gat = DFF(n2790gat)
--	n919gat = DFF(n2670gat)
--	n846gat = DFF(n2793gat)
--	n394gat = DFF(n2782gat)
--	n703gat = DFF(n2790gat)
--	n722gat = DFF(n2670gat)
--	n726gat = DFF(n2793gat)
--	n2510gat = DFF(n748gat)
--	n271gat = DFF(n2732gat)
--	n160gat = DFF(n2776gat)
--	n337gat = DFF(n2735gat)
--	n842gat = DFF(n2673gat)
--	n341gat = DFF(n2779gat)
--	n2522gat = DFF(n43gat)
--	n2472gat = DFF(n1620gat)
--	n2319gat = DFF(n2470gat)
--	n1821gat = DFF(n1827gat)
--	n1825gat = DFF(n1827gat)
--	n2029gat = DFF(n1816gat)
--	n1829gat = DFF(n2027gat)
--	n283gat = DFF(n2732gat)
--	n165gat = DFF(n2776gat)
--	n279gat = DFF(n2735gat)
--	n1026gat = DFF(n2673gat)
--	n275gat = DFF(n2779gat)
--	n2476gat = DFF(n55gat)
--	n1068gat = DFF(n2914gat)
--	n957gat = DFF(n2928gat)
--	n861gat = DFF(n2927gat)
--	n1294gat = DFF(n2896gat)
--	n1241gat = DFF(n2922gat)
--	n1298gat = DFF(n2897gat)
--	n865gat = DFF(n2894gat)
--	n1080gat = DFF(n2921gat)
--	n1148gat = DFF(n2895gat)
--	n2468gat = DFF(n933gat)
--	n618gat = DFF(n2790gat)
--	n491gat = DFF(n2782gat)
--	n622gat = DFF(n2793gat)
--	n626gat = DFF(n2670gat)
--	n834gat = DFF(n3064gat)
--	n707gat = DFF(n3055gat)
--	n838gat = DFF(n3063gat)
--	n830gat = DFF(n3062gat)
--	n614gat = DFF(n3056gat)
--	n2526gat = DFF(n504gat)
--	n680gat = DFF(n2913gat)
--	n816gat = DFF(n2920gat)
--	n580gat = DFF(n2905gat)
--	n824gat = DFF(n3057gat)
--	n820gat = DFF(n3059gat)
--	n883gat = DFF(n3058gat)
--	n584gat = DFF(n2898gat)
--	n684gat = DFF(n3060gat)
--	n699gat = DFF(n3061gat)
--	n2464gat = DFF(n567gat)
--	n2399gat = DFF(n3048gat)
--	n2343gat = DFF(n3049gat)
--	n2203gat = DFF(n3051gat)
--	n2562gat = DFF(n3047gat)
--	n2207gat = DFF(n3050gat)
--	n2626gat = DFF(n3040gat)
--	n2490gat = DFF(n3044gat)
--	n2622gat = DFF(n3042gat)
--	n2630gat = DFF(n3037gat)
--	n2543gat = DFF(n3041gat)
--	n2102gat = DFF(n1606gat)
--	n1880gat = DFF(n3052gat)
--	n1763gat = DFF(n1610gat)
--	n2155gat = DFF(n1858gat)
--	n1035gat = DFF(n2918gat)
--	n1121gat = DFF(n2952gat)
--	n1072gat = DFF(n2919gat)
--	n1282gat = DFF(n2910gat)
--	n1226gat = DFF(n2907gat)
--	n931gat = DFF(n2911gat)
--	n1135gat = DFF(n2912gat)
--	n1045gat = DFF(n2909gat)
--	n1197gat = DFF(n2908gat)
--	n2518gat = DFF(n2971gat)
--	n667gat = DFF(n2904gat)
--	n659gat = DFF(n2891gat)
--	n553gat = DFF(n2903gat)
--	n777gat = DFF(n2915gat)
--	n561gat = DFF(n2901gat)
--	n366gat = DFF(n2890gat)
--	n322gat = DFF(n2888gat)
--	n318gat = DFF(n2887gat)
--	n314gat = DFF(n2886gat)
--	n2599gat = DFF(n3010gat)
--	n2588gat = DFF(n3016gat)
--	n2640gat = DFF(n3054gat)
--	n2658gat = DFF(n2579gat)
--	n2495gat = DFF(n3036gat)
--	n2390gat = DFF(n3034gat)
--	n2270gat = DFF(n3031gat)
--	n2339gat = DFF(n3035gat)
--	n2502gat = DFF(n2646gat)
--	n2634gat = DFF(n3053gat)
--	n2506gat = DFF(n2613gat)
--	n1834gat = DFF(n1625gat)
--	n1767gat = DFF(n1626gat)
--	n2084gat = DFF(n1603gat)
--	n2143gat = DFF(n2541gat)
--	n2061gat = DFF(n2557gat)
--	n2139gat = DFF(n2487gat)
--	n1899gat = DFF(n2532gat)
--	n1850gat = DFF(n2628gat)
--	n2403gat = DFF(n2397gat)
--	n2394gat = DFF(n2341gat)
--	n2440gat = DFF(n2560gat)
--	n2407gat = DFF(n2205gat)
--	n2347gat = DFF(n2201gat)
--	n1389gat = DFF(n1793gat)
--	n2021gat = DFF(n1781gat)
--	n1394gat = DFF(n1516gat)
--	n1496gat = DFF(n1392gat)
--	n2091gat = DFF(n1685gat)
--	n1332gat = DFF(n1565gat)
--	n1740gat = DFF(n1330gat)
--	n2179gat = DFF(n1945gat)
--	n2190gat = DFF(n2268gat)
--	n2135gat = DFF(n2337gat)
--	n2262gat = DFF(n2388gat)
--	n2182gat = DFF(n1836gat)
--	n1433gat = DFF(n2983gat)
--	n1316gat = DFF(n1431gat)
--	n1363gat = DFF(n1314gat)
--	n1312gat = DFF(n1361gat)
--	n1775gat = DFF(n1696gat)
--	n1871gat = DFF(n2009gat)
--	n2592gat = DFF(n1773gat)
--	n1508gat = DFF(n1636gat)
--	n1678gat = DFF(n1712gat)
--	n2309gat = DFF(n3000gat)
--	n2450gat = DFF(n2307gat)
--	n2446gat = DFF(n2661gat)
--	n2095gat = DFF(n827gat)
--	n2176gat = DFF(n2093gat)
--	n2169gat = DFF(n2174gat)
--	n2454gat = DFF(n2163gat)
--	n2040gat = DFF(n1777gat)
--	n2044gat = DFF(n2015gat)
--	n2037gat = DFF(n2042gat)
--	n2025gat = DFF(n2017gat)
--	n2099gat = DFF(n2023gat)
--	n2266gat = DFF(n2493gat)
--	n2033gat = DFF(n2035gat)
--	n2110gat = DFF(n2031gat)
--	n2125gat = DFF(n2108gat)
--	n2121gat = DFF(n2123gat)
--	n2117gat = DFF(n2119gat)
--	n1975gat = DFF(n2632gat)
--	n2644gat = DFF(n2638gat)
--	n156gat = DFF(n612gat)
--	n152gat = DFF(n705gat)
--	n331gat = DFF(n822gat)
--	n388gat = DFF(n881gat)
--	n463gat = DFF(n818gat)
--	n327gat = DFF(n682gat)
--	n384gat = DFF(n697gat)
--	n256gat = DFF(n836gat)
--	n470gat = DFF(n828gat)
--	n148gat = DFF(n832gat)
--	n2458gat = DFF(n2590gat)
--	n2514gat = DFF(n2456gat)
--	n1771gat = DFF(n1613gat)
--	n1336gat = DFF(n1391gat)
--	n1748gat = DFF(n1927gat)
--	n1675gat = DFF(n1713gat)
--	n1807gat = DFF(n1717gat)
--	n1340gat = DFF(n1567gat)
--	n1456gat = DFF(n1564gat)
--	n1525gat = DFF(n1632gat)
--	n1462gat = DFF(n1915gat)
--	n1596gat = DFF(n1800gat)
--	n1588gat = DFF(n1593gat)
--	
--	I1 = NOT(n3088gat)
--	n2717gat = NOT(I1)
--	n2715gat = NOT(n2717gat)
--	I5 = NOT(n3087gat)
--	n2725gat = NOT(I5)
--	n2723gat = NOT(n2725gat)
--	n296gat = NOT(n421gat)
--	I11 = NOT(n3093gat)
--	n2768gat = NOT(I11)
--	I14 = NOT(n2768gat)
--	n2767gat = NOT(I14)
--	n373gat = NOT(n2767gat)
--	I18 = NOT(n3072gat)
--	n2671gat = NOT(I18)
--	n2669gat = NOT(n2671gat)
--	I23 = NOT(n3081gat)
--	n2845gat = NOT(I23)
--	n2844gat = NOT(n2845gat)
--	I27 = NOT(n3095gat)
--	n2668gat = NOT(I27)
--	I30 = NOT(n2668gat)
--	n2667gat = NOT(I30)
--	n856gat = NOT(n2667gat)
--	I44 = NOT(n673gat)
--	n672gat = NOT(I44)
--	I47 = NOT(n3069gat)
--	n2783gat = NOT(I47)
--	I50 = NOT(n2783gat)
--	n2782gat = NOT(I50)
--	n396gat = NOT(n398gat)
--	I62 = NOT(n3070gat)
--	n2791gat = NOT(I62)
--	I65 = NOT(n2791gat)
--	n2790gat = NOT(I65)
--	I76 = NOT(n402gat)
--	n401gat = NOT(I76)
--	n1645gat = NOT(n1499gat)
--	I81 = NOT(n2671gat)
--	n2670gat = NOT(I81)
--	I92 = NOT(n919gat)
--	n918gat = NOT(I92)
--	n1553gat = NOT(n1616gat)
--	I97 = NOT(n3071gat)
--	n2794gat = NOT(I97)
--	I100 = NOT(n2794gat)
--	n2793gat = NOT(I100)
--	I111 = NOT(n846gat)
--	n845gat = NOT(I111)
--	n1559gat = NOT(n1614gat)
--	n1643gat = NOT(n1641gat)
--	n1651gat = NOT(n1642gat)
--	n1562gat = NOT(n1556gat)
--	n1560gat = NOT(n1557gat)
--	n1640gat = NOT(n1639gat)
--	n1566gat = NOT(n1605gat)
--	n1554gat = NOT(n1555gat)
--	n1722gat = NOT(n1558gat)
--	n392gat = NOT(n394gat)
--	I149 = NOT(n703gat)
--	n702gat = NOT(I149)
--	n1319gat = NOT(n1256gat)
--	n720gat = NOT(n722gat)
--	I171 = NOT(n726gat)
--	n725gat = NOT(I171)
--	n1447gat = NOT(n1117gat)
--	n1627gat = NOT(n1618gat)
--	I178 = NOT(n722gat)
--	n721gat = NOT(I178)
--	n1380gat = NOT(n1114gat)
--	n1628gat = NOT(n1621gat)
--	n701gat = NOT(n703gat)
--	n1446gat = NOT(n1318gat)
--	n1705gat = NOT(n1619gat)
--	n1706gat = NOT(n1622gat)
--	I192 = NOT(n3083gat)
--	n2856gat = NOT(I192)
--	n2854gat = NOT(n2856gat)
--	I196 = NOT(n2854gat)
--	n1218gat = NOT(I196)
--	I199 = NOT(n3085gat)
--	n2861gat = NOT(I199)
--	n2859gat = NOT(n2861gat)
--	I203 = NOT(n2859gat)
--	n1219gat = NOT(I203)
--	I206 = NOT(n3084gat)
--	n2864gat = NOT(I206)
--	n2862gat = NOT(n2864gat)
--	I210 = NOT(n2862gat)
--	n1220gat = NOT(I210)
--	I214 = NOT(n2861gat)
--	n2860gat = NOT(I214)
--	I217 = NOT(n2860gat)
--	n1221gat = NOT(I217)
--	I220 = NOT(n2864gat)
--	n2863gat = NOT(I220)
--	I223 = NOT(n2863gat)
--	n1222gat = NOT(I223)
--	I227 = NOT(n2856gat)
--	n2855gat = NOT(I227)
--	I230 = NOT(n2855gat)
--	n1223gat = NOT(I230)
--	n640gat = NOT(n1213gat)
--	I237 = NOT(n640gat)
--	n753gat = NOT(I237)
--	I240 = NOT(n2717gat)
--	n2716gat = NOT(I240)
--	I243 = NOT(n3089gat)
--	n2869gat = NOT(I243)
--	n2867gat = NOT(n2869gat)
--	I248 = NOT(n2869gat)
--	n2868gat = NOT(I248)
--	I253 = NOT(n2906gat)
--	n754gat = NOT(I253)
--	I256 = NOT(n2725gat)
--	n2724gat = NOT(I256)
--	I259 = NOT(n3086gat)
--	n2728gat = NOT(I259)
--	n2726gat = NOT(n2728gat)
--	I264 = NOT(n2728gat)
--	n2727gat = NOT(I264)
--	n422gat = NOT(n2889gat)
--	I270 = NOT(n422gat)
--	n755gat = NOT(I270)
--	n747gat = NOT(n2906gat)
--	I275 = NOT(n747gat)
--	n756gat = NOT(I275)
--	I278 = NOT(n2889gat)
--	n757gat = NOT(I278)
--	I282 = NOT(n1213gat)
--	n758gat = NOT(I282)
--	n2508gat = NOT(n2510gat)
--	I297 = NOT(n3065gat)
--	n2733gat = NOT(I297)
--	I300 = NOT(n2733gat)
--	n2732gat = NOT(I300)
--	I311 = NOT(n271gat)
--	n270gat = NOT(I311)
--	I314 = NOT(n270gat)
--	n263gat = NOT(I314)
--	I317 = NOT(n3067gat)
--	n2777gat = NOT(I317)
--	I320 = NOT(n2777gat)
--	n2776gat = NOT(I320)
--	I331 = NOT(n160gat)
--	n159gat = NOT(I331)
--	I334 = NOT(n159gat)
--	n264gat = NOT(I334)
--	I337 = NOT(n3066gat)
--	n2736gat = NOT(I337)
--	I340 = NOT(n2736gat)
--	n2735gat = NOT(I340)
--	I351 = NOT(n337gat)
--	n336gat = NOT(I351)
--	I354 = NOT(n336gat)
--	n265gat = NOT(I354)
--	n158gat = NOT(n160gat)
--	I359 = NOT(n158gat)
--	n266gat = NOT(I359)
--	n335gat = NOT(n337gat)
--	I363 = NOT(n335gat)
--	n267gat = NOT(I363)
--	n269gat = NOT(n271gat)
--	I368 = NOT(n269gat)
--	n268gat = NOT(I368)
--	n41gat = NOT(n258gat)
--	I375 = NOT(n41gat)
--	n48gat = NOT(I375)
--	I378 = NOT(n725gat)
--	n1018gat = NOT(I378)
--	I381 = NOT(n3073gat)
--	n2674gat = NOT(I381)
--	I384 = NOT(n2674gat)
--	n2673gat = NOT(I384)
--	I395 = NOT(n842gat)
--	n841gat = NOT(I395)
--	I398 = NOT(n841gat)
--	n1019gat = NOT(I398)
--	I401 = NOT(n721gat)
--	n1020gat = NOT(I401)
--	n840gat = NOT(n842gat)
--	I406 = NOT(n840gat)
--	n1021gat = NOT(I406)
--	I409 = NOT(n720gat)
--	n1022gat = NOT(I409)
--	n724gat = NOT(n726gat)
--	I414 = NOT(n724gat)
--	n1023gat = NOT(I414)
--	I420 = NOT(n1013gat)
--	n49gat = NOT(I420)
--	I423 = NOT(n3068gat)
--	n2780gat = NOT(I423)
--	I426 = NOT(n2780gat)
--	n2779gat = NOT(I426)
--	I437 = NOT(n341gat)
--	n340gat = NOT(I437)
--	I440 = NOT(n340gat)
--	n480gat = NOT(I440)
--	I443 = NOT(n702gat)
--	n481gat = NOT(I443)
--	I446 = NOT(n394gat)
--	n393gat = NOT(I446)
--	I449 = NOT(n393gat)
--	n482gat = NOT(I449)
--	I453 = NOT(n701gat)
--	n483gat = NOT(I453)
--	I456 = NOT(n392gat)
--	n484gat = NOT(I456)
--	n339gat = NOT(n341gat)
--	I461 = NOT(n339gat)
--	n485gat = NOT(I461)
--	n42gat = NOT(n475gat)
--	I468 = NOT(n42gat)
--	n50gat = NOT(I468)
--	n162gat = NOT(n1013gat)
--	I473 = NOT(n162gat)
--	n51gat = NOT(I473)
--	I476 = NOT(n475gat)
--	n52gat = NOT(I476)
--	I480 = NOT(n258gat)
--	n53gat = NOT(I480)
--	n2520gat = NOT(n2522gat)
--	n1448gat = NOT(n1376gat)
--	n1701gat = NOT(n1617gat)
--	n1379gat = NOT(n1377gat)
--	n1615gat = NOT(n1624gat)
--	n1500gat = NOT(n1113gat)
--	n1503gat = NOT(n1501gat)
--	n1779gat = NOT(n1623gat)
--	I509 = NOT(n3099gat)
--	n2730gat = NOT(I509)
--	I512 = NOT(n2730gat)
--	n2729gat = NOT(I512)
--	n2470gat = NOT(n2472gat)
--	n2317gat = NOT(n2319gat)
--	n1819gat = NOT(n1821gat)
--	n1823gat = NOT(n1825gat)
--	n1816gat = NOT(n1817gat)
--	n2027gat = NOT(n2029gat)
--	I572 = NOT(n1829gat)
--	n1828gat = NOT(I572)
--	I576 = NOT(n3100gat)
--	n2851gat = NOT(I576)
--	I579 = NOT(n2851gat)
--	n2850gat = NOT(I579)
--	I583 = NOT(n2786gat)
--	n2785gat = NOT(I583)
--	n92gat = NOT(n2785gat)
--	n637gat = NOT(n529gat)
--	n293gat = NOT(n361gat)
--	I591 = NOT(n3094gat)
--	n2722gat = NOT(I591)
--	I594 = NOT(n2722gat)
--	n2721gat = NOT(I594)
--	n297gat = NOT(n2721gat)
--	I606 = NOT(n283gat)
--	n282gat = NOT(I606)
--	I609 = NOT(n282gat)
--	n172gat = NOT(I609)
--	I620 = NOT(n165gat)
--	n164gat = NOT(I620)
--	I623 = NOT(n164gat)
--	n173gat = NOT(I623)
--	I634 = NOT(n279gat)
--	n278gat = NOT(I634)
--	I637 = NOT(n278gat)
--	n174gat = NOT(I637)
--	n163gat = NOT(n165gat)
--	I642 = NOT(n163gat)
--	n175gat = NOT(I642)
--	n277gat = NOT(n279gat)
--	I646 = NOT(n277gat)
--	n176gat = NOT(I646)
--	n281gat = NOT(n283gat)
--	I651 = NOT(n281gat)
--	n177gat = NOT(I651)
--	n54gat = NOT(n167gat)
--	I658 = NOT(n54gat)
--	n60gat = NOT(I658)
--	I661 = NOT(n845gat)
--	n911gat = NOT(I661)
--	I672 = NOT(n1026gat)
--	n1025gat = NOT(I672)
--	I675 = NOT(n1025gat)
--	n912gat = NOT(I675)
--	I678 = NOT(n918gat)
--	n913gat = NOT(I678)
--	n1024gat = NOT(n1026gat)
--	I683 = NOT(n1024gat)
--	n914gat = NOT(I683)
--	n917gat = NOT(n919gat)
--	I687 = NOT(n917gat)
--	n915gat = NOT(I687)
--	n844gat = NOT(n846gat)
--	I692 = NOT(n844gat)
--	n916gat = NOT(I692)
--	I698 = NOT(n906gat)
--	n61gat = NOT(I698)
--	I709 = NOT(n275gat)
--	n274gat = NOT(I709)
--	I712 = NOT(n274gat)
--	n348gat = NOT(I712)
--	I715 = NOT(n401gat)
--	n349gat = NOT(I715)
--	I718 = NOT(n398gat)
--	n397gat = NOT(I718)
--	I721 = NOT(n397gat)
--	n350gat = NOT(I721)
--	n400gat = NOT(n402gat)
--	I726 = NOT(n400gat)
--	n351gat = NOT(I726)
--	I729 = NOT(n396gat)
--	n352gat = NOT(I729)
--	n273gat = NOT(n275gat)
--	I734 = NOT(n273gat)
--	n353gat = NOT(I734)
--	n178gat = NOT(n343gat)
--	I741 = NOT(n178gat)
--	n62gat = NOT(I741)
--	n66gat = NOT(n906gat)
--	I746 = NOT(n66gat)
--	n63gat = NOT(I746)
--	I749 = NOT(n343gat)
--	n64gat = NOT(I749)
--	I753 = NOT(n167gat)
--	n65gat = NOT(I753)
--	n2474gat = NOT(n2476gat)
--	I768 = NOT(n3090gat)
--	n2832gat = NOT(I768)
--	I771 = NOT(n2832gat)
--	n2831gat = NOT(I771)
--	n2731gat = NOT(n2733gat)
--	I776 = NOT(n3074gat)
--	n2719gat = NOT(I776)
--	n2718gat = NOT(n2719gat)
--	I790 = NOT(n1068gat)
--	n1067gat = NOT(I790)
--	I793 = NOT(n1067gat)
--	n949gat = NOT(I793)
--	I796 = NOT(n3076gat)
--	n2839gat = NOT(I796)
--	n2838gat = NOT(n2839gat)
--	n2775gat = NOT(n2777gat)
--	I812 = NOT(n957gat)
--	n956gat = NOT(I812)
--	I815 = NOT(n956gat)
--	n950gat = NOT(I815)
--	I818 = NOT(n3075gat)
--	n2712gat = NOT(I818)
--	n2711gat = NOT(n2712gat)
--	n2734gat = NOT(n2736gat)
--	I834 = NOT(n861gat)
--	n860gat = NOT(I834)
--	I837 = NOT(n860gat)
--	n951gat = NOT(I837)
--	n955gat = NOT(n957gat)
--	I842 = NOT(n955gat)
--	n952gat = NOT(I842)
--	n859gat = NOT(n861gat)
--	I846 = NOT(n859gat)
--	n953gat = NOT(I846)
--	n1066gat = NOT(n1068gat)
--	I851 = NOT(n1066gat)
--	n954gat = NOT(I851)
--	n857gat = NOT(n944gat)
--	I858 = NOT(n857gat)
--	n938gat = NOT(I858)
--	n2792gat = NOT(n2794gat)
--	I863 = NOT(n3080gat)
--	n2847gat = NOT(I863)
--	n2846gat = NOT(n2847gat)
--	I877 = NOT(n1294gat)
--	n1293gat = NOT(I877)
--	I880 = NOT(n1293gat)
--	n1233gat = NOT(I880)
--	n2672gat = NOT(n2674gat)
--	I885 = NOT(n3082gat)
--	n2853gat = NOT(I885)
--	n2852gat = NOT(n2853gat)
--	I899 = NOT(n1241gat)
--	n1240gat = NOT(I899)
--	I902 = NOT(n1240gat)
--	n1234gat = NOT(I902)
--	I913 = NOT(n1298gat)
--	n1297gat = NOT(I913)
--	I916 = NOT(n1297gat)
--	n1235gat = NOT(I916)
--	n1239gat = NOT(n1241gat)
--	I921 = NOT(n1239gat)
--	n1236gat = NOT(I921)
--	n1296gat = NOT(n1298gat)
--	I925 = NOT(n1296gat)
--	n1237gat = NOT(I925)
--	n1292gat = NOT(n1294gat)
--	I930 = NOT(n1292gat)
--	n1238gat = NOT(I930)
--	I936 = NOT(n1228gat)
--	n939gat = NOT(I936)
--	n2778gat = NOT(n2780gat)
--	I941 = NOT(n3077gat)
--	n2837gat = NOT(I941)
--	n2836gat = NOT(n2837gat)
--	I955 = NOT(n865gat)
--	n864gat = NOT(I955)
--	I958 = NOT(n864gat)
--	n1055gat = NOT(I958)
--	n2789gat = NOT(n2791gat)
--	I963 = NOT(n3079gat)
--	n2841gat = NOT(I963)
--	n2840gat = NOT(n2841gat)
--	I977 = NOT(n1080gat)
--	n1079gat = NOT(I977)
--	I980 = NOT(n1079gat)
--	n1056gat = NOT(I980)
--	n2781gat = NOT(n2783gat)
--	I985 = NOT(n3078gat)
--	n2843gat = NOT(I985)
--	n2842gat = NOT(n2843gat)
--	I999 = NOT(n1148gat)
--	n1147gat = NOT(I999)
--	I1002 = NOT(n1147gat)
--	n1057gat = NOT(I1002)
--	n1078gat = NOT(n1080gat)
--	I1007 = NOT(n1078gat)
--	n1058gat = NOT(I1007)
--	n1146gat = NOT(n1148gat)
--	I1011 = NOT(n1146gat)
--	n1059gat = NOT(I1011)
--	n863gat = NOT(n865gat)
--	I1016 = NOT(n863gat)
--	n1060gat = NOT(I1016)
--	n928gat = NOT(n1050gat)
--	I1023 = NOT(n928gat)
--	n940gat = NOT(I1023)
--	n858gat = NOT(n1228gat)
--	I1028 = NOT(n858gat)
--	n941gat = NOT(I1028)
--	I1031 = NOT(n1050gat)
--	n942gat = NOT(I1031)
--	I1035 = NOT(n944gat)
--	n943gat = NOT(I1035)
--	n2466gat = NOT(n2468gat)
--	n2720gat = NOT(n2722gat)
--	n740gat = NOT(n2667gat)
--	n2784gat = NOT(n2786gat)
--	n743gat = NOT(n746gat)
--	n294gat = NOT(n360gat)
--	n374gat = NOT(n2767gat)
--	n616gat = NOT(n618gat)
--	I1067 = NOT(n616gat)
--	n501gat = NOT(I1067)
--	n489gat = NOT(n491gat)
--	I1079 = NOT(n489gat)
--	n502gat = NOT(I1079)
--	I1082 = NOT(n618gat)
--	n617gat = NOT(I1082)
--	I1085 = NOT(n617gat)
--	n499gat = NOT(I1085)
--	I1088 = NOT(n491gat)
--	n490gat = NOT(I1088)
--	I1091 = NOT(n490gat)
--	n500gat = NOT(I1091)
--	n620gat = NOT(n622gat)
--	I1103 = NOT(n620gat)
--	n738gat = NOT(I1103)
--	n624gat = NOT(n626gat)
--	I1115 = NOT(n624gat)
--	n737gat = NOT(I1115)
--	I1118 = NOT(n622gat)
--	n621gat = NOT(I1118)
--	I1121 = NOT(n621gat)
--	n733gat = NOT(I1121)
--	I1124 = NOT(n626gat)
--	n625gat = NOT(I1124)
--	I1127 = NOT(n625gat)
--	n735gat = NOT(I1127)
--	I1138 = NOT(n834gat)
--	n833gat = NOT(I1138)
--	I1141 = NOT(n833gat)
--	n714gat = NOT(I1141)
--	I1152 = NOT(n707gat)
--	n706gat = NOT(I1152)
--	I1155 = NOT(n706gat)
--	n715gat = NOT(I1155)
--	I1166 = NOT(n838gat)
--	n837gat = NOT(I1166)
--	I1169 = NOT(n837gat)
--	n716gat = NOT(I1169)
--	n705gat = NOT(n707gat)
--	I1174 = NOT(n705gat)
--	n717gat = NOT(I1174)
--	n836gat = NOT(n838gat)
--	I1178 = NOT(n836gat)
--	n718gat = NOT(I1178)
--	n832gat = NOT(n834gat)
--	I1183 = NOT(n832gat)
--	n719gat = NOT(I1183)
--	n515gat = NOT(n709gat)
--	I1190 = NOT(n515gat)
--	n509gat = NOT(I1190)
--	I1201 = NOT(n830gat)
--	n829gat = NOT(I1201)
--	I1204 = NOT(n829gat)
--	n734gat = NOT(I1204)
--	n828gat = NOT(n830gat)
--	I1209 = NOT(n828gat)
--	n736gat = NOT(I1209)
--	I1216 = NOT(n728gat)
--	n510gat = NOT(I1216)
--	I1227 = NOT(n614gat)
--	n613gat = NOT(I1227)
--	I1230 = NOT(n613gat)
--	n498gat = NOT(I1230)
--	n612gat = NOT(n614gat)
--	I1236 = NOT(n612gat)
--	n503gat = NOT(I1236)
--	n404gat = NOT(n493gat)
--	I1243 = NOT(n404gat)
--	n511gat = NOT(I1243)
--	n405gat = NOT(n728gat)
--	I1248 = NOT(n405gat)
--	n512gat = NOT(I1248)
--	I1251 = NOT(n493gat)
--	n513gat = NOT(I1251)
--	I1255 = NOT(n709gat)
--	n514gat = NOT(I1255)
--	n2524gat = NOT(n2526gat)
--	n17gat = NOT(n564gat)
--	n79gat = NOT(n86gat)
--	n219gat = NOT(n78gat)
--	n563gat = NOT(I1278)
--	n289gat = NOT(n563gat)
--	n179gat = NOT(n287gat)
--	n188gat = NOT(n288gat)
--	n72gat = NOT(n181gat)
--	n111gat = NOT(n182gat)
--	I1302 = NOT(n680gat)
--	n679gat = NOT(I1302)
--	I1305 = NOT(n679gat)
--	n808gat = NOT(I1305)
--	I1319 = NOT(n816gat)
--	n815gat = NOT(I1319)
--	I1322 = NOT(n815gat)
--	n809gat = NOT(I1322)
--	I1336 = NOT(n580gat)
--	n579gat = NOT(I1336)
--	I1339 = NOT(n579gat)
--	n810gat = NOT(I1339)
--	n814gat = NOT(n816gat)
--	I1344 = NOT(n814gat)
--	n811gat = NOT(I1344)
--	n578gat = NOT(n580gat)
--	I1348 = NOT(n578gat)
--	n812gat = NOT(I1348)
--	n678gat = NOT(n680gat)
--	I1353 = NOT(n678gat)
--	n813gat = NOT(I1353)
--	n677gat = NOT(n803gat)
--	I1360 = NOT(n677gat)
--	n572gat = NOT(I1360)
--	I1371 = NOT(n824gat)
--	n823gat = NOT(I1371)
--	I1374 = NOT(n823gat)
--	n591gat = NOT(I1374)
--	I1385 = NOT(n820gat)
--	n819gat = NOT(I1385)
--	I1388 = NOT(n819gat)
--	n592gat = NOT(I1388)
--	I1399 = NOT(n883gat)
--	n882gat = NOT(I1399)
--	I1402 = NOT(n882gat)
--	n593gat = NOT(I1402)
--	n818gat = NOT(n820gat)
--	I1407 = NOT(n818gat)
--	n594gat = NOT(I1407)
--	n881gat = NOT(n883gat)
--	I1411 = NOT(n881gat)
--	n595gat = NOT(I1411)
--	n822gat = NOT(n824gat)
--	I1416 = NOT(n822gat)
--	n596gat = NOT(I1416)
--	I1422 = NOT(n586gat)
--	n573gat = NOT(I1422)
--	I1436 = NOT(n584gat)
--	n583gat = NOT(I1436)
--	I1439 = NOT(n583gat)
--	n691gat = NOT(I1439)
--	I1450 = NOT(n684gat)
--	n683gat = NOT(I1450)
--	I1453 = NOT(n683gat)
--	n692gat = NOT(I1453)
--	I1464 = NOT(n699gat)
--	n698gat = NOT(I1464)
--	I1467 = NOT(n698gat)
--	n693gat = NOT(I1467)
--	n682gat = NOT(n684gat)
--	I1472 = NOT(n682gat)
--	n694gat = NOT(I1472)
--	n697gat = NOT(n699gat)
--	I1476 = NOT(n697gat)
--	n695gat = NOT(I1476)
--	n582gat = NOT(n584gat)
--	I1481 = NOT(n582gat)
--	n696gat = NOT(I1481)
--	n456gat = NOT(n686gat)
--	I1488 = NOT(n456gat)
--	n574gat = NOT(I1488)
--	n565gat = NOT(n586gat)
--	I1493 = NOT(n565gat)
--	n575gat = NOT(I1493)
--	I1496 = NOT(n686gat)
--	n576gat = NOT(I1496)
--	I1500 = NOT(n803gat)
--	n577gat = NOT(I1500)
--	n2462gat = NOT(n2464gat)
--	n2665gat = NOT(I1516)
--	n2596gat = NOT(n2665gat)
--	n189gat = NOT(n286gat)
--	n194gat = NOT(n187gat)
--	n21gat = NOT(n15gat)
--	I1538 = NOT(n2399gat)
--	n2398gat = NOT(I1538)
--	n2353gat = NOT(n2398gat)
--	I1550 = NOT(n2343gat)
--	n2342gat = NOT(I1550)
--	n2284gat = NOT(n2342gat)
--	n2201gat = NOT(n2203gat)
--	n2354gat = NOT(n2201gat)
--	n2560gat = NOT(n2562gat)
--	n2356gat = NOT(n2560gat)
--	n2205gat = NOT(n2207gat)
--	n2214gat = NOT(n2205gat)
--	n2286gat = NOT(I1585)
--	n2624gat = NOT(n2626gat)
--	I1606 = NOT(n2490gat)
--	n2489gat = NOT(I1606)
--	I1617 = NOT(n2622gat)
--	n2621gat = NOT(I1617)
--	n2533gat = NOT(n2534gat)
--	I1630 = NOT(n2630gat)
--	n2629gat = NOT(I1630)
--	n2486gat = NOT(n2629gat)
--	n2541gat = NOT(n2543gat)
--	n2429gat = NOT(n2541gat)
--	n2432gat = NOT(n2430gat)
--	I1655 = NOT(n2102gat)
--	n2101gat = NOT(I1655)
--	n1693gat = NOT(n2101gat)
--	I1667 = NOT(n1880gat)
--	n1879gat = NOT(I1667)
--	n1698gat = NOT(n1934gat)
--	n1543gat = NOT(n1606gat)
--	I1683 = NOT(n1763gat)
--	n1762gat = NOT(I1683)
--	n1673gat = NOT(n2989gat)
--	n1858gat = NOT(n1673gat)
--	I1698 = NOT(n2155gat)
--	n2154gat = NOT(I1698)
--	n2488gat = NOT(n2490gat)
--	I1703 = NOT(n2626gat)
--	n2625gat = NOT(I1703)
--	n2530gat = NOT(n2531gat)
--	I1708 = NOT(n2543gat)
--	n2542gat = NOT(I1708)
--	n2482gat = NOT(n2542gat)
--	n2426gat = NOT(n2480gat)
--	n2153gat = NOT(n2155gat)
--	n2341gat = NOT(n2343gat)
--	n2355gat = NOT(n2341gat)
--	I1719 = NOT(n2562gat)
--	n2561gat = NOT(I1719)
--	n2443gat = NOT(n2561gat)
--	n2289gat = NOT(I1724)
--	n2148gat = NOT(I1734)
--	n855gat = NOT(n2148gat)
--	n759gat = NOT(n855gat)
--	I1749 = NOT(n1035gat)
--	n1034gat = NOT(I1749)
--	I1752 = NOT(n1034gat)
--	n1189gat = NOT(I1752)
--	n1075gat = NOT(n855gat)
--	I1766 = NOT(n1121gat)
--	n1120gat = NOT(I1766)
--	I1769 = NOT(n1120gat)
--	n1190gat = NOT(I1769)
--	n760gat = NOT(n855gat)
--	I1783 = NOT(n1072gat)
--	n1071gat = NOT(I1783)
--	I1786 = NOT(n1071gat)
--	n1191gat = NOT(I1786)
--	n1119gat = NOT(n1121gat)
--	I1791 = NOT(n1119gat)
--	n1192gat = NOT(I1791)
--	n1070gat = NOT(n1072gat)
--	I1795 = NOT(n1070gat)
--	n1193gat = NOT(I1795)
--	n1033gat = NOT(n1035gat)
--	I1800 = NOT(n1033gat)
--	n1194gat = NOT(I1800)
--	n1183gat = NOT(n1184gat)
--	I1807 = NOT(n1183gat)
--	n1274gat = NOT(I1807)
--	n644gat = NOT(n855gat)
--	n1280gat = NOT(n1282gat)
--	n641gat = NOT(n855gat)
--	I1833 = NOT(n1226gat)
--	n1225gat = NOT(I1833)
--	I1837 = NOT(n1282gat)
--	n1281gat = NOT(I1837)
--	n1224gat = NOT(n1226gat)
--	I1843 = NOT(n2970gat)
--	n1275gat = NOT(I1843)
--	n761gat = NOT(n855gat)
--	I1857 = NOT(n931gat)
--	n930gat = NOT(I1857)
--	I1860 = NOT(n930gat)
--	n1206gat = NOT(I1860)
--	n762gat = NOT(n855gat)
--	I1874 = NOT(n1135gat)
--	n1134gat = NOT(I1874)
--	I1877 = NOT(n1134gat)
--	n1207gat = NOT(I1877)
--	n643gat = NOT(n855gat)
--	I1891 = NOT(n1045gat)
--	n1044gat = NOT(I1891)
--	I1894 = NOT(n1044gat)
--	n1208gat = NOT(I1894)
--	n1133gat = NOT(n1135gat)
--	I1899 = NOT(n1133gat)
--	n1209gat = NOT(I1899)
--	n1043gat = NOT(n1045gat)
--	I1903 = NOT(n1043gat)
--	n1210gat = NOT(I1903)
--	n929gat = NOT(n931gat)
--	I1908 = NOT(n929gat)
--	n1211gat = NOT(I1908)
--	n1268gat = NOT(n1201gat)
--	I1915 = NOT(n1268gat)
--	n1276gat = NOT(I1915)
--	n1329gat = NOT(n2970gat)
--	I1920 = NOT(n1329gat)
--	n1277gat = NOT(I1920)
--	I1923 = NOT(n1201gat)
--	n1278gat = NOT(I1923)
--	I1927 = NOT(n1184gat)
--	n1279gat = NOT(I1927)
--	n1284gat = NOT(n1269gat)
--	n642gat = NOT(n855gat)
--	n1195gat = NOT(n1197gat)
--	I1947 = NOT(n1197gat)
--	n1196gat = NOT(I1947)
--	n2516gat = NOT(n2518gat)
--	I1961 = NOT(n2516gat)
--	n3017gat = NOT(I1961)
--	n851gat = NOT(n853gat)
--	n1725gat = NOT(n2148gat)
--	n664gat = NOT(n1725gat)
--	n852gat = NOT(n854gat)
--	I1981 = NOT(n667gat)
--	n666gat = NOT(I1981)
--	n368gat = NOT(n1725gat)
--	I1996 = NOT(n659gat)
--	n658gat = NOT(I1996)
--	I1999 = NOT(n658gat)
--	n784gat = NOT(I1999)
--	n662gat = NOT(n1725gat)
--	I2014 = NOT(n553gat)
--	n552gat = NOT(I2014)
--	I2017 = NOT(n552gat)
--	n785gat = NOT(I2017)
--	n661gat = NOT(n1725gat)
--	I2032 = NOT(n777gat)
--	n776gat = NOT(I2032)
--	I2035 = NOT(n776gat)
--	n786gat = NOT(I2035)
--	n551gat = NOT(n553gat)
--	I2040 = NOT(n551gat)
--	n787gat = NOT(I2040)
--	n775gat = NOT(n777gat)
--	I2044 = NOT(n775gat)
--	n788gat = NOT(I2044)
--	n657gat = NOT(n659gat)
--	I2049 = NOT(n657gat)
--	n789gat = NOT(I2049)
--	n35gat = NOT(n779gat)
--	I2056 = NOT(n35gat)
--	n125gat = NOT(I2056)
--	n558gat = NOT(n1725gat)
--	n559gat = NOT(n561gat)
--	n371gat = NOT(n1725gat)
--	I2084 = NOT(n366gat)
--	n365gat = NOT(I2084)
--	I2088 = NOT(n561gat)
--	n560gat = NOT(I2088)
--	n364gat = NOT(n366gat)
--	I2094 = NOT(n2876gat)
--	n126gat = NOT(I2094)
--	n663gat = NOT(n1725gat)
--	I2109 = NOT(n322gat)
--	n321gat = NOT(I2109)
--	I2112 = NOT(n321gat)
--	n226gat = NOT(I2112)
--	n370gat = NOT(n1725gat)
--	I2127 = NOT(n318gat)
--	n317gat = NOT(I2127)
--	I2130 = NOT(n317gat)
--	n227gat = NOT(I2130)
--	n369gat = NOT(n1725gat)
--	I2145 = NOT(n314gat)
--	n313gat = NOT(I2145)
--	I2148 = NOT(n313gat)
--	n228gat = NOT(I2148)
--	n316gat = NOT(n318gat)
--	I2153 = NOT(n316gat)
--	n229gat = NOT(I2153)
--	n312gat = NOT(n314gat)
--	I2157 = NOT(n312gat)
--	n230gat = NOT(I2157)
--	n320gat = NOT(n322gat)
--	I2162 = NOT(n320gat)
--	n231gat = NOT(I2162)
--	n34gat = NOT(n221gat)
--	I2169 = NOT(n34gat)
--	n127gat = NOT(I2169)
--	n133gat = NOT(n2876gat)
--	I2174 = NOT(n133gat)
--	n128gat = NOT(I2174)
--	I2177 = NOT(n221gat)
--	n129gat = NOT(I2177)
--	I2181 = NOT(n779gat)
--	n130gat = NOT(I2181)
--	n665gat = NOT(n667gat)
--	n1601gat = NOT(n120gat)
--	n2597gat = NOT(n2599gat)
--	n2595gat = NOT(n2594gat)
--	n2586gat = NOT(n2588gat)
--	I2213 = NOT(n2342gat)
--	n2573gat = NOT(I2213)
--	n2638gat = NOT(n2640gat)
--	I2225 = NOT(n2638gat)
--	n2574gat = NOT(I2225)
--	I2228 = NOT(n2561gat)
--	n2575gat = NOT(I2228)
--	I2232 = NOT(n2640gat)
--	n2639gat = NOT(I2232)
--	I2235 = NOT(n2639gat)
--	n2576gat = NOT(I2235)
--	I2238 = NOT(n2560gat)
--	n2577gat = NOT(I2238)
--	I2242 = NOT(n2341gat)
--	n2578gat = NOT(I2242)
--	I2248 = NOT(n2568gat)
--	n2582gat = NOT(I2248)
--	I2251 = NOT(n2207gat)
--	n2206gat = NOT(I2251)
--	I2254 = NOT(n2206gat)
--	n2414gat = NOT(I2254)
--	I2257 = NOT(n2398gat)
--	n2415gat = NOT(I2257)
--	I2260 = NOT(n2203gat)
--	n2202gat = NOT(I2260)
--	I2263 = NOT(n2202gat)
--	n2416gat = NOT(I2263)
--	n2397gat = NOT(n2399gat)
--	I2268 = NOT(n2397gat)
--	n2417gat = NOT(I2268)
--	I2271 = NOT(n2201gat)
--	n2418gat = NOT(I2271)
--	I2275 = NOT(n2205gat)
--	n2419gat = NOT(I2275)
--	I2281 = NOT(n2409gat)
--	n2585gat = NOT(I2281)
--	n2656gat = NOT(n2658gat)
--	n2493gat = NOT(n2495gat)
--	n2388gat = NOT(n2390gat)
--	I2316 = NOT(n2390gat)
--	n2389gat = NOT(I2316)
--	I2319 = NOT(n2495gat)
--	n2494gat = NOT(I2319)
--	I2324 = NOT(n3014gat)
--	n2649gat = NOT(I2324)
--	n2268gat = NOT(n2270gat)
--	I2344 = NOT(n2339gat)
--	n2338gat = NOT(I2344)
--	n2337gat = NOT(n2339gat)
--	I2349 = NOT(n2270gat)
--	n2269gat = NOT(I2349)
--	I2354 = NOT(n2880gat)
--	n2652gat = NOT(I2354)
--	n2500gat = NOT(n2502gat)
--	n2620gat = NOT(n2622gat)
--	n2612gat = NOT(n2620gat)
--	I2372 = NOT(n2612gat)
--	n2606gat = NOT(I2372)
--	n2532gat = NOT(n2625gat)
--	I2376 = NOT(n2532gat)
--	n2607gat = NOT(I2376)
--	n2540gat = NOT(n2488gat)
--	I2380 = NOT(n2540gat)
--	n2608gat = NOT(I2380)
--	n2536gat = NOT(n2624gat)
--	I2385 = NOT(n2536gat)
--	n2609gat = NOT(I2385)
--	n2487gat = NOT(n2489gat)
--	I2389 = NOT(n2487gat)
--	n2610gat = NOT(I2389)
--	n2557gat = NOT(n2621gat)
--	I2394 = NOT(n2557gat)
--	n2611gat = NOT(I2394)
--	I2400 = NOT(n2601gat)
--	n2616gat = NOT(I2400)
--	I2403 = NOT(n2629gat)
--	n2550gat = NOT(I2403)
--	I2414 = NOT(n2634gat)
--	n2633gat = NOT(I2414)
--	I2417 = NOT(n2633gat)
--	n2551gat = NOT(I2417)
--	I2420 = NOT(n2542gat)
--	n2552gat = NOT(I2420)
--	n2632gat = NOT(n2634gat)
--	I2425 = NOT(n2632gat)
--	n2553gat = NOT(I2425)
--	I2428 = NOT(n2541gat)
--	n2554gat = NOT(I2428)
--	n2628gat = NOT(n2630gat)
--	I2433 = NOT(n2628gat)
--	n2555gat = NOT(I2433)
--	I2439 = NOT(n2545gat)
--	n2619gat = NOT(I2439)
--	n2504gat = NOT(n2506gat)
--	n2660gat = NOT(n2655gat)
--	n1528gat = NOT(n2293gat)
--	n1523gat = NOT(n2219gat)
--	n1592gat = NOT(n1529gat)
--	n2666gat = NOT(n1704gat)
--	n2422gat = NOT(n3013gat)
--	n2290gat = NOT(n2202gat)
--	n2081gat = NOT(n2218gat)
--	n2285gat = NOT(n2397gat)
--	n2359gat = NOT(n2358gat)
--	n1414gat = NOT(n1415gat)
--	n566gat = NOT(n364gat)
--	n1480gat = NOT(n2292gat)
--	n1301gat = NOT(n1416gat)
--	n1150gat = NOT(n312gat)
--	n873gat = NOT(n316gat)
--	n2011gat = NOT(n2306gat)
--	n1478gat = NOT(n1481gat)
--	n875gat = NOT(n559gat)
--	n1410gat = NOT(n2357gat)
--	n876gat = NOT(n1347gat)
--	n1160gat = NOT(n1484gat)
--	n1084gat = NOT(n657gat)
--	n983gat = NOT(n320gat)
--	n1482gat = NOT(n2363gat)
--	n1157gat = NOT(n1483gat)
--	n985gat = NOT(n775gat)
--	n1530gat = NOT(n2364gat)
--	n1307gat = NOT(n1308gat)
--	n1085gat = NOT(n551gat)
--	n1479gat = NOT(n2291gat)
--	n1348gat = NOT(n1349gat)
--	n2217gat = NOT(n2206gat)
--	n1591gat = NOT(n2223gat)
--	n1437gat = NOT(n1438gat)
--	n1832gat = NOT(n1834gat)
--	n1765gat = NOT(n1767gat)
--	n1878gat = NOT(n1880gat)
--	n1442gat = NOT(n1831gat)
--	n1444gat = NOT(n1442gat)
--	n1378gat = NOT(n2975gat)
--	n1322gat = NOT(n2974gat)
--	n1439gat = NOT(n1486gat)
--	n1370gat = NOT(n1426gat)
--	n1369gat = NOT(n2966gat)
--	n1366gat = NOT(n1365gat)
--	n1374gat = NOT(n2979gat)
--	n2162gat = NOT(n2220gat)
--	n1450gat = NOT(n1423gat)
--	n1427gat = NOT(n1608gat)
--	n1603gat = NOT(n1831gat)
--	n2082gat = NOT(n2084gat)
--	n1449gat = NOT(n1494gat)
--	n1590gat = NOT(n1603gat)
--	n1248gat = NOT(n2954gat)
--	n1418gat = NOT(n1417gat)
--	n1306gat = NOT(n2964gat)
--	n1353gat = NOT(n1419gat)
--	n1247gat = NOT(n2958gat)
--	n1355gat = NOT(n1422gat)
--	n1300gat = NOT(n2963gat)
--	n1487gat = NOT(n1485gat)
--	n1164gat = NOT(n2953gat)
--	n1356gat = NOT(n1354gat)
--	n1436gat = NOT(n1435gat)
--	n1106gat = NOT(n2949gat)
--	n1425gat = NOT(n1421gat)
--	n1105gat = NOT(n2934gat)
--	n1424gat = NOT(n1420gat)
--	n1309gat = NOT(n2959gat)
--	I2672 = NOT(n2143gat)
--	n2142gat = NOT(I2672)
--	n1788gat = NOT(n2142gat)
--	I2684 = NOT(n2061gat)
--	n2060gat = NOT(I2684)
--	n1786gat = NOT(n2060gat)
--	I2696 = NOT(n2139gat)
--	n2138gat = NOT(I2696)
--	n1839gat = NOT(n2138gat)
--	n1897gat = NOT(n1899gat)
--	n1884gat = NOT(n1897gat)
--	n1848gat = NOT(n1850gat)
--	n1783gat = NOT(n1848gat)
--	n1548gat = NOT(I2721)
--	n1719gat = NOT(n1548gat)
--	n2137gat = NOT(n2139gat)
--	n1633gat = NOT(n2137gat)
--	n2059gat = NOT(n2061gat)
--	n1785gat = NOT(n2059gat)
--	I2731 = NOT(n1850gat)
--	n1849gat = NOT(I2731)
--	n1784gat = NOT(n1849gat)
--	n1716gat = NOT(I2736)
--	n1635gat = NOT(n1716gat)
--	n2401gat = NOT(n2403gat)
--	n1989gat = NOT(n2401gat)
--	n2392gat = NOT(n2394gat)
--	n1918gat = NOT(n2392gat)
--	I2771 = NOT(n2440gat)
--	n2439gat = NOT(I2771)
--	n1986gat = NOT(n2439gat)
--	n1866gat = NOT(n1865gat)
--	I2785 = NOT(n2407gat)
--	n2406gat = NOT(I2785)
--	n2216gat = NOT(n2406gat)
--	n2345gat = NOT(n2347gat)
--	n1988gat = NOT(n2345gat)
--	n1735gat = NOT(n1861gat)
--	n1387gat = NOT(n1389gat)
--	n1694gat = NOT(I2813)
--	n1777gat = NOT(n1694gat)
--	n1781gat = NOT(n1780gat)
--	n2019gat = NOT(n2021gat)
--	n1549gat = NOT(I2832)
--	n1551gat = NOT(n1549gat)
--	I2837 = NOT(n2347gat)
--	n2346gat = NOT(I2837)
--	n2152gat = NOT(n2346gat)
--	n2405gat = NOT(n2407gat)
--	n2351gat = NOT(n2405gat)
--	I2843 = NOT(n2403gat)
--	n2402gat = NOT(I2843)
--	n2212gat = NOT(n2402gat)
--	I2847 = NOT(n2394gat)
--	n2393gat = NOT(I2847)
--	n1991gat = NOT(n2393gat)
--	n1665gat = NOT(n1666gat)
--	n1517gat = NOT(n1578gat)
--	n1392gat = NOT(n1394gat)
--	I2873 = NOT(n1496gat)
--	n1495gat = NOT(I2873)
--	n1685gat = NOT(n1604gat)
--	I2885 = NOT(n2091gat)
--	n2090gat = NOT(I2885)
--	n1550gat = NOT(I2890)
--	n1552gat = NOT(n1550gat)
--	n1330gat = NOT(n1332gat)
--	n1738gat = NOT(n1740gat)
--	I2915 = NOT(n1740gat)
--	n1739gat = NOT(I2915)
--	n1925gat = NOT(n1920gat)
--	n1917gat = NOT(n1921gat)
--	n2141gat = NOT(n2143gat)
--	n1787gat = NOT(n2141gat)
--	n1717gat = NOT(I2926)
--	n1859gat = NOT(n1717gat)
--	n1922gat = NOT(n1798gat)
--	n1713gat = NOT(I2935)
--	n1743gat = NOT(n1713gat)
--	n1923gat = NOT(n1864gat)
--	n1945gat = NOT(n1690gat)
--	I2953 = NOT(n2179gat)
--	n2178gat = NOT(I2953)
--	n1661gat = NOT(n1660gat)
--	n1572gat = NOT(n1576gat)
--	n2438gat = NOT(n2440gat)
--	n2283gat = NOT(n2438gat)
--	n1520gat = NOT(n1582gat)
--	n1580gat = NOT(n1577gat)
--	n1990gat = NOT(n2988gat)
--	I2978 = NOT(n2190gat)
--	n2189gat = NOT(I2978)
--	I2989 = NOT(n2135gat)
--	n2134gat = NOT(I2989)
--	I3000 = NOT(n2262gat)
--	n2261gat = NOT(I3000)
--	n2128gat = NOT(n2129gat)
--	n1836gat = NOT(n1695gat)
--	I3016 = NOT(n2182gat)
--	n2181gat = NOT(I3016)
--	n1431gat = NOT(n1433gat)
--	n1314gat = NOT(n1316gat)
--	n1361gat = NOT(n1363gat)
--	I3056 = NOT(n1312gat)
--	n1311gat = NOT(I3056)
--	n1707gat = NOT(n1626gat)
--	n1773gat = NOT(n1775gat)
--	n1659gat = NOT(n2987gat)
--	n1515gat = NOT(n1521gat)
--	n1736gat = NOT(n1737gat)
--	n1658gat = NOT(n2216gat)
--	n1724gat = NOT(n1732gat)
--	n1662gat = NOT(n1663gat)
--	n1656gat = NOT(n1655gat)
--	n1670gat = NOT(n1667gat)
--	n1569gat = NOT(n1570gat)
--	n1568gat = NOT(n1575gat)
--	n1727gat = NOT(n1728gat)
--	n1797gat = NOT(n1801gat)
--	n1730gat = NOT(n1731gat)
--	n1561gat = NOT(n1571gat)
--	n1668gat = NOT(n1734gat)
--	n1742gat = NOT(n2216gat)
--	n1671gat = NOT(n1669gat)
--	n1652gat = NOT(n1657gat)
--	n1648gat = NOT(n1729gat)
--	n1790gat = NOT(n1726gat)
--	n2004gat = NOT(n1929gat)
--	n1869gat = NOT(n1871gat)
--	I3143 = NOT(n2592gat)
--	n2591gat = NOT(I3143)
--	n1584gat = NOT(n2989gat)
--	n1714gat = NOT(I3149)
--	n1718gat = NOT(n1714gat)
--	I3163 = NOT(n1508gat)
--	n1507gat = NOT(I3163)
--	n1396gat = NOT(n1401gat)
--	I3168 = NOT(n1394gat)
--	n1393gat = NOT(I3168)
--	n1409gat = NOT(n1476gat)
--	I3174 = NOT(n1899gat)
--	n1898gat = NOT(I3174)
--	n1838gat = NOT(n1898gat)
--	n1712gat = NOT(I3179)
--	I3191 = NOT(n1678gat)
--	n1677gat = NOT(I3191)
--	n2000gat = NOT(n1412gat)
--	n2001gat = NOT(n1412gat)
--	n1999gat = NOT(n2001gat)
--	n2307gat = NOT(n2309gat)
--	I3211 = NOT(n2663gat)
--	n3018gat = NOT(I3211)
--	n2448gat = NOT(n2450gat)
--	n2661gat = NOT(n2662gat)
--	n2444gat = NOT(n2446gat)
--	I3235 = NOT(n2238gat)
--	n3019gat = NOT(I3235)
--	n1310gat = NOT(n1312gat)
--	n199gat = NOT(n87gat)
--	n195gat = NOT(n184gat)
--	n827gat = NOT(n204gat)
--	n2093gat = NOT(n2095gat)
--	n2174gat = NOT(n2176gat)
--	I3273 = NOT(n2169gat)
--	n2168gat = NOT(I3273)
--	n2452gat = NOT(n2454gat)
--	n1691gat = NOT(n2452gat)
--	I3287 = NOT(n1691gat)
--	n3020gat = NOT(I3287)
--	I3290 = NOT(n1691gat)
--	n3021gat = NOT(I3290)
--	I3293 = NOT(n1691gat)
--	n3022gat = NOT(I3293)
--	n1699gat = NOT(n2452gat)
--	I3297 = NOT(n1699gat)
--	n3023gat = NOT(I3297)
--	I3300 = NOT(n1699gat)
--	n3024gat = NOT(I3300)
--	I3303 = NOT(n1691gat)
--	n3025gat = NOT(I3303)
--	I3306 = NOT(n1699gat)
--	n3026gat = NOT(I3306)
--	I3309 = NOT(n1699gat)
--	n3027gat = NOT(I3309)
--	I3312 = NOT(n1699gat)
--	n3028gat = NOT(I3312)
--	I3315 = NOT(n1869gat)
--	n3029gat = NOT(I3315)
--	I3318 = NOT(n1869gat)
--	n3030gat = NOT(I3318)
--	n2260gat = NOT(n2262gat)
--	n2257gat = NOT(n2189gat)
--	n2188gat = NOT(n2190gat)
--	n2187gat = NOT(n3004gat)
--	I3336 = NOT(n2040gat)
--	n2039gat = NOT(I3336)
--	I3339 = NOT(n1775gat)
--	n1774gat = NOT(I3339)
--	I3342 = NOT(n1316gat)
--	n1315gat = NOT(I3342)
--	n2042gat = NOT(n2044gat)
--	n2035gat = NOT(n2037gat)
--	n2023gat = NOT(n2025gat)
--	n2097gat = NOT(n2099gat)
--	n1855gat = NOT(n2014gat)
--	I3387 = NOT(n2194gat)
--	n3031gat = NOT(I3387)
--	I3390 = NOT(n2261gat)
--	n3032gat = NOT(I3390)
--	n2256gat = NOT(n3032gat)
--	I3394 = NOT(n2260gat)
--	n3033gat = NOT(I3394)
--	n2251gat = NOT(n3033gat)
--	n2184gat = NOT(n3003gat)
--	I3401 = NOT(n2192gat)
--	n3034gat = NOT(I3401)
--	n2133gat = NOT(n2135gat)
--	n2131gat = NOT(n2185gat)
--	n2049gat = NOT(n3001gat)
--	I3412 = NOT(n2057gat)
--	n3035gat = NOT(I3412)
--	n2253gat = NOT(n2189gat)
--	n2252gat = NOT(n2260gat)
--	n2248gat = NOT(n3006gat)
--	n2264gat = NOT(n2266gat)
--	I3429 = NOT(n2266gat)
--	n2265gat = NOT(I3429)
--	n2492gat = NOT(n2329gat)
--	I3436 = NOT(n2492gat)
--	n3036gat = NOT(I3436)
--	n1709gat = NOT(n1849gat)
--	n1845gat = NOT(n2141gat)
--	n1891gat = NOT(n2059gat)
--	n1963gat = NOT(n2137gat)
--	n1886gat = NOT(n1897gat)
--	n1968gat = NOT(n1958gat)
--	n1629gat = NOT(n1895gat)
--	n1631gat = NOT(n1848gat)
--	n1711gat = NOT(n2990gat)
--	n2200gat = NOT(n2078gat)
--	n2437gat = NOT(n2195gat)
--	I3457 = NOT(n2556gat)
--	n3037gat = NOT(I3457)
--	n1956gat = NOT(n1898gat)
--	I3461 = NOT(n1956gat)
--	n3038gat = NOT(I3461)
--	n1954gat = NOT(n3038gat)
--	I3465 = NOT(n1886gat)
--	n3039gat = NOT(I3465)
--	n1888gat = NOT(n3039gat)
--	n2048gat = NOT(n2994gat)
--	I3472 = NOT(n2539gat)
--	n3040gat = NOT(I3472)
--	n1969gat = NOT(n2142gat)
--	n1893gat = NOT(n2060gat)
--	n1892gat = NOT(n2993gat)
--	I3483 = NOT(n2436gat)
--	n3041gat = NOT(I3483)
--	n2056gat = NOT(n2998gat)
--	I3491 = NOT(n2387gat)
--	n3042gat = NOT(I3491)
--	I3494 = NOT(n1963gat)
--	n3043gat = NOT(I3494)
--	n1960gat = NOT(n3043gat)
--	n1887gat = NOT(n2138gat)
--	n1961gat = NOT(n2996gat)
--	I3504 = NOT(n2330gat)
--	n3044gat = NOT(I3504)
--	n2199gat = NOT(n2147gat)
--	I3509 = NOT(n2438gat)
--	n3045gat = NOT(I3509)
--	n2332gat = NOT(n3045gat)
--	I3513 = NOT(n2439gat)
--	n3046gat = NOT(I3513)
--	n2259gat = NOT(n3046gat)
--	n2328gat = NOT(n3008gat)
--	I3520 = NOT(n2498gat)
--	n3047gat = NOT(I3520)
--	n2151gat = NOT(n2193gat)
--	n2209gat = NOT(n3005gat)
--	I3530 = NOT(n2396gat)
--	n3048gat = NOT(I3530)
--	n2052gat = NOT(n2393gat)
--	n2058gat = NOT(n2997gat)
--	I3539 = NOT(n2198gat)
--	n3049gat = NOT(I3539)
--	n2349gat = NOT(n2215gat)
--	n2281gat = NOT(n3009gat)
--	I3549 = NOT(n2197gat)
--	n3050gat = NOT(I3549)
--	n2146gat = NOT(n3002gat)
--	I3558 = NOT(n2196gat)
--	n3051gat = NOT(I3558)
--	n2031gat = NOT(n2033gat)
--	n2108gat = NOT(n2110gat)
--	I3587 = NOT(n2125gat)
--	n2124gat = NOT(I3587)
--	n2123gat = NOT(n2125gat)
--	n2119gat = NOT(n2121gat)
--	n2115gat = NOT(n2117gat)
--	I3610 = NOT(n1882gat)
--	n3052gat = NOT(I3610)
--	I3621 = NOT(n1975gat)
--	n1974gat = NOT(I3621)
--	n1955gat = NOT(n1956gat)
--	n1970gat = NOT(n1896gat)
--	n1973gat = NOT(n1975gat)
--	n2558gat = NOT(n2559gat)
--	I3635 = NOT(n2558gat)
--	n3053gat = NOT(I3635)
--	I3646 = NOT(n2644gat)
--	n2643gat = NOT(I3646)
--	n2333gat = NOT(n2438gat)
--	n2564gat = NOT(n2352gat)
--	n2642gat = NOT(n2644gat)
--	n2636gat = NOT(n2637gat)
--	I3660 = NOT(n2636gat)
--	n3054gat = NOT(I3660)
--	n88gat = NOT(n84gat)
--	n375gat = NOT(n110gat)
--	I3677 = NOT(n156gat)
--	n155gat = NOT(I3677)
--	n253gat = NOT(n1702gat)
--	n150gat = NOT(n152gat)
--	I3691 = NOT(n152gat)
--	n151gat = NOT(I3691)
--	n243gat = NOT(n1702gat)
--	n233gat = NOT(n243gat)
--	n154gat = NOT(n156gat)
--	n800gat = NOT(n2874gat)
--	I3703 = NOT(n2917gat)
--	n3055gat = NOT(I3703)
--	n235gat = NOT(n2878gat)
--	I3713 = NOT(n2892gat)
--	n3056gat = NOT(I3713)
--	n372gat = NOT(n212gat)
--	n329gat = NOT(n331gat)
--	I3736 = NOT(n388gat)
--	n387gat = NOT(I3736)
--	n334gat = NOT(n1700gat)
--	n386gat = NOT(n388gat)
--	I3742 = NOT(n331gat)
--	n330gat = NOT(I3742)
--	n1430gat = NOT(n1700gat)
--	n1490gat = NOT(n1430gat)
--	n452gat = NOT(n2885gat)
--	I3754 = NOT(n2900gat)
--	n3057gat = NOT(I3754)
--	n333gat = NOT(n2883gat)
--	I3765 = NOT(n2929gat)
--	n3058gat = NOT(I3765)
--	I3777 = NOT(n463gat)
--	n462gat = NOT(I3777)
--	n325gat = NOT(n327gat)
--	n457gat = NOT(n2884gat)
--	n461gat = NOT(n463gat)
--	n458gat = NOT(n2902gat)
--	I3801 = NOT(n2925gat)
--	n3059gat = NOT(I3801)
--	n144gat = NOT(n247gat)
--	I3808 = NOT(n327gat)
--	n326gat = NOT(I3808)
--	n878gat = NOT(n2879gat)
--	I3817 = NOT(n2916gat)
--	n3060gat = NOT(I3817)
--	n382gat = NOT(n384gat)
--	I3831 = NOT(n384gat)
--	n383gat = NOT(I3831)
--	n134gat = NOT(n2875gat)
--	I3841 = NOT(n2899gat)
--	n3061gat = NOT(I3841)
--	n254gat = NOT(n256gat)
--	n252gat = NOT(n2877gat)
--	n468gat = NOT(n470gat)
--	I3867 = NOT(n470gat)
--	n469gat = NOT(I3867)
--	n381gat = NOT(n2893gat)
--	I3876 = NOT(n2926gat)
--	n3062gat = NOT(I3876)
--	n241gat = NOT(n140gat)
--	I3882 = NOT(n256gat)
--	n255gat = NOT(I3882)
--	n802gat = NOT(n2882gat)
--	I3891 = NOT(n2924gat)
--	n3063gat = NOT(I3891)
--	n146gat = NOT(n148gat)
--	I3904 = NOT(n148gat)
--	n147gat = NOT(I3904)
--	n380gat = NOT(n2881gat)
--	I3914 = NOT(n2923gat)
--	n3064gat = NOT(I3914)
--	n69gat = NOT(n68gat)
--	n1885gat = NOT(n2048gat)
--	I3923 = NOT(n2710gat)
--	n2707gat = NOT(I3923)
--	n16gat = NOT(n564gat)
--	n295gat = NOT(n357gat)
--	n11gat = NOT(n12gat)
--	n1889gat = NOT(n1961gat)
--	I3935 = NOT(n2704gat)
--	n2700gat = NOT(I3935)
--	n2051gat = NOT(n2056gat)
--	I3941 = NOT(n2684gat)
--	n2680gat = NOT(I3941)
--	n1350gat = NOT(n1831gat)
--	I3945 = NOT(n1350gat)
--	n2696gat = NOT(I3945)
--	I3948 = NOT(n2696gat)
--	n2692gat = NOT(I3948)
--	I3951 = NOT(n2448gat)
--	n2683gat = NOT(I3951)
--	I3954 = NOT(n2683gat)
--	n2679gat = NOT(I3954)
--	I3957 = NOT(n2450gat)
--	n2449gat = NOT(I3957)
--	n1754gat = NOT(n2449gat)
--	I3962 = NOT(n2830gat)
--	n2827gat = NOT(I3962)
--	n2590gat = NOT(n2592gat)
--	n2456gat = NOT(n2458gat)
--	n2512gat = NOT(n2514gat)
--	n1544gat = NOT(n1625gat)
--	n1769gat = NOT(n1771gat)
--	n1683gat = NOT(n1756gat)
--	n2167gat = NOT(n2169gat)
--	n2013gat = NOT(I4000)
--	n1791gat = NOT(n2013gat)
--	n2691gat = NOT(n2695gat)
--	n1518gat = NOT(n1694gat)
--	n2699gat = NOT(n2703gat)
--	n2159gat = NOT(n1412gat)
--	n2478gat = NOT(n2579gat)
--	I4014 = NOT(n2744gat)
--	n2740gat = NOT(I4014)
--	n2158gat = NOT(n1412gat)
--	n2186gat = NOT(n2613gat)
--	I4020 = NOT(n2800gat)
--	n2797gat = NOT(I4020)
--	n2288gat = NOT(I4024)
--	n1513gat = NOT(n2288gat)
--	n2537gat = NOT(n2538gat)
--	n2442gat = NOT(n2483gat)
--	n1334gat = NOT(n1336gat)
--	I4055 = NOT(n1748gat)
--	n1747gat = NOT(I4055)
--	I4067 = NOT(n1675gat)
--	n1674gat = NOT(I4067)
--	n1403gat = NOT(n1402gat)
--	I4081 = NOT(n1807gat)
--	n1806gat = NOT(I4081)
--	n1634gat = NOT(n1712gat)
--	n1338gat = NOT(n1340gat)
--	I4105 = NOT(n1456gat)
--	n1455gat = NOT(I4105)
--	I4108 = NOT(n1340gat)
--	n1339gat = NOT(I4108)
--	n1505gat = NOT(n2980gat)
--	I4117 = NOT(n1505gat)
--	n2758gat = NOT(I4117)
--	n2755gat = NOT(n2758gat)
--	n1546gat = NOT(n2980gat)
--	I4122 = NOT(n1546gat)
--	n2752gat = NOT(I4122)
--	n2748gat = NOT(n2752gat)
--	n2012gat = NOT(n2016gat)
--	n2002gat = NOT(n2008gat)
--	I4129 = NOT(n3097gat)
--	n2858gat = NOT(I4129)
--	n2857gat = NOT(n2858gat)
--	I4135 = NOT(n3098gat)
--	n2766gat = NOT(I4135)
--	I4138 = NOT(n2766gat)
--	n2765gat = NOT(I4138)
--	n1684gat = NOT(n1759gat)
--	n1632gat = NOT(I4145)
--	I4157 = NOT(n1525gat)
--	n1524gat = NOT(I4157)
--	n1862gat = NOT(n1863gat)
--	n1919gat = NOT(n1860gat)
--	n1460gat = NOT(n1462gat)
--	I4185 = NOT(n1596gat)
--	n1595gat = NOT(I4185)
--	n1454gat = NOT(n1469gat)
--	n1468gat = NOT(n1519gat)
--	I4194 = NOT(n1462gat)
--	n1461gat = NOT(I4194)
--	n1477gat = NOT(n2984gat)
--	n1594gat = NOT(n1596gat)
--	I4212 = NOT(n1588gat)
--	n1587gat = NOT(I4212)
--	n1681gat = NOT(I4217)
--	I4222 = NOT(n1761gat)
--	n2751gat = NOT(I4222)
--	n2747gat = NOT(n2751gat)
--	I4227 = NOT(n1760gat)
--	n2743gat = NOT(I4227)
--	n2739gat = NOT(n2743gat)
--	n1978gat = NOT(n2286gat)
--	I4233 = NOT(n1721gat)
--	n2808gat = NOT(I4233)
--	I4236 = NOT(n2808gat)
--	n2804gat = NOT(I4236)
--	n517gat = NOT(n518gat)
--	n417gat = NOT(n418gat)
--	n413gat = NOT(n411gat)
--	n412gat = NOT(n522gat)
--	n406gat = NOT(n516gat)
--	n407gat = NOT(n355gat)
--	n290gat = NOT(n525gat)
--	n527gat = NOT(n356gat)
--	n416gat = NOT(n415gat)
--	n528gat = NOT(n521gat)
--	n358gat = NOT(n532gat)
--	n639gat = NOT(n523gat)
--	n1111gat = NOT(n635gat)
--	n524gat = NOT(n414gat)
--	n1112gat = NOT(n630gat)
--	n741gat = NOT(n629gat)
--	n633gat = NOT(n634gat)
--	n926gat = NOT(n632gat)
--	n670gat = NOT(n636gat)
--	n1123gat = NOT(n632gat)
--	n1007gat = NOT(n635gat)
--	n1006gat = NOT(n630gat)
--	I4309 = NOT(n2941gat)
--	n2814gat = NOT(I4309)
--	I4312 = NOT(n2814gat)
--	n2811gat = NOT(I4312)
--	n1002gat = NOT(n2946gat)
--	I4329 = NOT(n2950gat)
--	n2813gat = NOT(I4329)
--	I4332 = NOT(n2813gat)
--	n2810gat = NOT(I4332)
--	n888gat = NOT(n2933gat)
--	I4349 = NOT(n2935gat)
--	n2818gat = NOT(I4349)
--	I4352 = NOT(n2818gat)
--	n2816gat = NOT(I4352)
--	n898gat = NOT(n2940gat)
--	I4369 = NOT(n2937gat)
--	n2817gat = NOT(I4369)
--	I4372 = NOT(n2817gat)
--	n2815gat = NOT(I4372)
--	n1179gat = NOT(n2947gat)
--	I4389 = NOT(n2956gat)
--	n2824gat = NOT(I4389)
--	I4392 = NOT(n2824gat)
--	n2821gat = NOT(I4392)
--	n897gat = NOT(n2939gat)
--	I4409 = NOT(n2938gat)
--	n2823gat = NOT(I4409)
--	I4412 = NOT(n2823gat)
--	n2820gat = NOT(I4412)
--	n894gat = NOT(n2932gat)
--	I4429 = NOT(n2936gat)
--	n2829gat = NOT(I4429)
--	I4432 = NOT(n2829gat)
--	n2826gat = NOT(I4432)
--	n1180gat = NOT(n2948gat)
--	I4449 = NOT(n2955gat)
--	n2828gat = NOT(I4449)
--	I4452 = NOT(n2828gat)
--	n2825gat = NOT(I4452)
--	n671gat = NOT(n673gat)
--	n628gat = NOT(n631gat)
--	n976gat = NOT(n628gat)
--	I4475 = NOT(n2951gat)
--	n2807gat = NOT(I4475)
--	I4478 = NOT(n2807gat)
--	n2803gat = NOT(I4478)
--	n2127gat = NOT(n2389gat)
--	I4482 = NOT(n2127gat)
--	n2682gat = NOT(I4482)
--	I4485 = NOT(n2682gat)
--	n2678gat = NOT(I4485)
--	n2046gat = NOT(n2269gat)
--	I4489 = NOT(n2046gat)
--	n2681gat = NOT(I4489)
--	I4492 = NOT(n2681gat)
--	n2677gat = NOT(I4492)
--	n1708gat = NOT(n2338gat)
--	I4496 = NOT(n1708gat)
--	n2688gat = NOT(I4496)
--	I4499 = NOT(n2688gat)
--	n2686gat = NOT(I4499)
--	n455gat = NOT(n291gat)
--	n2237gat = NOT(n2646gat)
--	I4506 = NOT(n2764gat)
--	n2763gat = NOT(I4506)
--	n1782gat = NOT(n2971gat)
--	I4512 = NOT(n2762gat)
--	n2760gat = NOT(I4512)
--	n2325gat = NOT(n3010gat)
--	I4518 = NOT(n2761gat)
--	n2759gat = NOT(I4518)
--	n2245gat = NOT(n504gat)
--	I4524 = NOT(n2757gat)
--	n2754gat = NOT(I4524)
--	n2244gat = NOT(n567gat)
--	I4530 = NOT(n2756gat)
--	n2753gat = NOT(I4530)
--	n2243gat = NOT(n55gat)
--	I4536 = NOT(n2750gat)
--	n2746gat = NOT(I4536)
--	n2246gat = NOT(n933gat)
--	I4542 = NOT(n2749gat)
--	n2745gat = NOT(I4542)
--	n2384gat = NOT(n43gat)
--	I4548 = NOT(n2742gat)
--	n2738gat = NOT(I4548)
--	n2385gat = NOT(n748gat)
--	I4554 = NOT(n2741gat)
--	n2737gat = NOT(I4554)
--	n1286gat = NOT(n1269gat)
--	I4558 = NOT(n1286gat)
--	n2687gat = NOT(I4558)
--	n2685gat = NOT(n2687gat)
--	n1328gat = NOT(n1224gat)
--	n1381gat = NOT(n1328gat)
--	n1384gat = NOT(n2184gat)
--	I4566 = NOT(n2694gat)
--	n2690gat = NOT(I4566)
--	n1382gat = NOT(n1280gat)
--	n1451gat = NOT(n1382gat)
--	n1453gat = NOT(n2187gat)
--	I4573 = NOT(n2693gat)
--	n2689gat = NOT(I4573)
--	n927gat = NOT(n1133gat)
--	n925gat = NOT(n927gat)
--	n1452gat = NOT(n2049gat)
--	I4580 = NOT(n2702gat)
--	n2698gat = NOT(I4580)
--	n923gat = NOT(n1043gat)
--	n921gat = NOT(n923gat)
--	n1890gat = NOT(n2328gat)
--	I4587 = NOT(n2701gat)
--	n2697gat = NOT(I4587)
--	n850gat = NOT(n929gat)
--	n739gat = NOT(n850gat)
--	n1841gat = NOT(n2058gat)
--	I4594 = NOT(n2709gat)
--	n2706gat = NOT(I4594)
--	n922gat = NOT(n1119gat)
--	n848gat = NOT(n922gat)
--	n2047gat = NOT(n2209gat)
--	I4601 = NOT(n2708gat)
--	n2705gat = NOT(I4601)
--	n924gat = NOT(n1070gat)
--	n849gat = NOT(n924gat)
--	n2050gat = NOT(n2146gat)
--	I4608 = NOT(n2799gat)
--	n2796gat = NOT(I4608)
--	n1118gat = NOT(n1033gat)
--	n1032gat = NOT(n1118gat)
--	n2054gat = NOT(n2281gat)
--	I4615 = NOT(n2798gat)
--	n2795gat = NOT(I4615)
--	I4620 = NOT(n1745gat)
--	n2806gat = NOT(I4620)
--	I4623 = NOT(n2806gat)
--	n2802gat = NOT(I4623)
--	I4626 = NOT(n1871gat)
--	n1870gat = NOT(I4626)
--	n1086gat = NOT(n1870gat)
--	I4630 = NOT(n1086gat)
--	n2805gat = NOT(I4630)
--	I4633 = NOT(n2805gat)
--	n2801gat = NOT(I4633)
--	n67gat = NOT(n85gat)
--	n71gat = NOT(n180gat)
--	n1840gat = NOT(n1892gat)
--	I4642 = NOT(n2812gat)
--	n2809gat = NOT(I4642)
--	n76gat = NOT(n82gat)
--	n14gat = NOT(n186gat)
--	n1842gat = NOT(n1711gat)
--	I4651 = NOT(n2822gat)
--	n2819gat = NOT(I4651)
--	I4654 = NOT(n2819gat)
--	n3104gat = NOT(I4654)
--	I4657 = NOT(n2809gat)
--	n3105gat = NOT(I4657)
--	I4660 = NOT(n2801gat)
--	n3106gat = NOT(I4660)
--	I4663 = NOT(n2802gat)
--	n3107gat = NOT(I4663)
--	I4666 = NOT(n2795gat)
--	n3108gat = NOT(I4666)
--	I4669 = NOT(n2796gat)
--	n3109gat = NOT(I4669)
--	I4672 = NOT(n2705gat)
--	n3110gat = NOT(I4672)
--	I4675 = NOT(n2706gat)
--	n3111gat = NOT(I4675)
--	I4678 = NOT(n2697gat)
--	n3112gat = NOT(I4678)
--	I4681 = NOT(n2698gat)
--	n3113gat = NOT(I4681)
--	I4684 = NOT(n2689gat)
--	n3114gat = NOT(I4684)
--	I4687 = NOT(n2690gat)
--	n3115gat = NOT(I4687)
--	I4690 = NOT(n2685gat)
--	n3116gat = NOT(I4690)
--	I4693 = NOT(n2737gat)
--	n3117gat = NOT(I4693)
--	I4696 = NOT(n2738gat)
--	n3118gat = NOT(I4696)
--	I4699 = NOT(n2745gat)
--	n3119gat = NOT(I4699)
--	I4702 = NOT(n2746gat)
--	n3120gat = NOT(I4702)
--	I4705 = NOT(n2753gat)
--	n3121gat = NOT(I4705)
--	I4708 = NOT(n2754gat)
--	n3122gat = NOT(I4708)
--	I4711 = NOT(n2759gat)
--	n3123gat = NOT(I4711)
--	I4714 = NOT(n2760gat)
--	n3124gat = NOT(I4714)
--	I4717 = NOT(n2763gat)
--	n3125gat = NOT(I4717)
--	I4720 = NOT(n2686gat)
--	n3126gat = NOT(I4720)
--	I4723 = NOT(n2677gat)
--	n3127gat = NOT(I4723)
--	I4726 = NOT(n2678gat)
--	n3128gat = NOT(I4726)
--	I4729 = NOT(n2803gat)
--	n3129gat = NOT(I4729)
--	I4732 = NOT(n2825gat)
--	n3130gat = NOT(I4732)
--	I4735 = NOT(n2826gat)
--	n3131gat = NOT(I4735)
--	I4738 = NOT(n2820gat)
--	n3132gat = NOT(I4738)
--	I4741 = NOT(n2821gat)
--	n3133gat = NOT(I4741)
--	I4744 = NOT(n2815gat)
--	n3134gat = NOT(I4744)
--	I4747 = NOT(n2816gat)
--	n3135gat = NOT(I4747)
--	I4750 = NOT(n2810gat)
--	n3136gat = NOT(I4750)
--	I4753 = NOT(n2811gat)
--	n3137gat = NOT(I4753)
--	I4756 = NOT(n2804gat)
--	n3138gat = NOT(I4756)
--	I4759 = NOT(n2739gat)
--	n3139gat = NOT(I4759)
--	I4762 = NOT(n2747gat)
--	n3140gat = NOT(I4762)
--	I4765 = NOT(n2748gat)
--	n3141gat = NOT(I4765)
--	I4768 = NOT(n2755gat)
--	n3142gat = NOT(I4768)
--	I4771 = NOT(n2797gat)
--	n3143gat = NOT(I4771)
--	I4774 = NOT(n2740gat)
--	n3144gat = NOT(I4774)
--	I4777 = NOT(n2699gat)
--	n3145gat = NOT(I4777)
--	I4780 = NOT(n2691gat)
--	n3146gat = NOT(I4780)
--	I4783 = NOT(n2827gat)
--	n3147gat = NOT(I4783)
--	I4786 = NOT(n2679gat)
--	n3148gat = NOT(I4786)
--	I4789 = NOT(n2692gat)
--	n3149gat = NOT(I4789)
--	I4792 = NOT(n2680gat)
--	n3150gat = NOT(I4792)
--	I4795 = NOT(n2700gat)
--	n3151gat = NOT(I4795)
--	I4798 = NOT(n2707gat)
--	n3152gat = NOT(I4798)
--	
--	n2897gat = OR(n648gat, n442gat)
--	n1213gat = OR(n1214gat, n1215gat, n1216gat, n1217gat)
--	n2906gat = OR(n745gat, n638gat)
--	n2889gat = OR(n423gat, n362gat)
--	n748gat = OR(n749gat, n750gat, n751gat, n752gat)
--	n258gat = OR(n259gat, n260gat, n261gat, n262gat)
--	n1013gat = OR(n1014gat, n1015gat, n1016gat, n1017gat)
--	n475gat = OR(n476gat, n477gat, n478gat, n479gat)
--	n43gat = OR(n44gat, n45gat, n46gat, n47gat)
--	n2786gat = OR(n3091gat, n3092gat)
--	n167gat = OR(n168gat, n169gat, n170gat, n171gat)
--	n906gat = OR(n907gat, n908gat, n909gat, n910gat)
--	n343gat = OR(n344gat, n345gat, n346gat, n347gat)
--	n55gat = OR(n56gat, n57gat, n58gat, n59gat)
--	n2914gat = OR(n768gat, n655gat)
--	n2928gat = OR(n963gat, n868gat)
--	n2927gat = OR(n962gat, n959gat)
--	n944gat = OR(n945gat, n946gat, n947gat, n948gat)
--	n2896gat = OR(n647gat, n441gat)
--	n2922gat = OR(n967gat, n792gat)
--	n1228gat = OR(n1229gat, n1230gat, n1231gat, n1232gat)
--	n2894gat = OR(n443gat, n439gat)
--	n2921gat = OR(n966gat, n790gat)
--	n2895gat = OR(n444gat, n440gat)
--	n1050gat = OR(n1051gat, n1052gat, n1053gat, n1054gat)
--	n933gat = OR(n934gat, n935gat, n936gat, n937gat)
--	n709gat = OR(n710gat, n711gat, n712gat, n713gat)
--	n728gat = OR(n729gat, n730gat, n731gat, n732gat)
--	n493gat = OR(n494gat, n495gat, n496gat, n497gat)
--	n504gat = OR(n505gat, n506gat, n507gat, n508gat)
--	I1277 = OR(n2860gat, n2855gat, n2863gat)
--	I1278 = OR(n740gat, n3030gat, I1277)
--	n2913gat = OR(n767gat, n653gat)
--	n2920gat = OR(n867gat, n771gat)
--	n2905gat = OR(n964gat, n961gat)
--	n803gat = OR(n804gat, n805gat, n806gat, n807gat)
--	n586gat = OR(n587gat, n588gat, n589gat, n590gat)
--	n2898gat = OR(n447gat, n445gat)
--	n686gat = OR(n687gat, n688gat, n689gat, n690gat)
--	n567gat = OR(n568gat, n569gat, n570gat, n571gat)
--	I1515 = OR(n2474gat, n2524gat, n2831gat)
--	I1516 = OR(n2466gat, n2462gat, I1515)
--	I1584 = OR(n2353gat, n2284gat, n2354gat)
--	I1585 = OR(n2356gat, n2214gat, I1584)
--	n2989gat = OR(n1693gat, n1692gat)
--	I1723 = OR(n2354gat, n2353gat, n2214gat)
--	I1724 = OR(n2355gat, n2443gat, I1723)
--	I1733 = OR(n2286gat, n2428gat, n2289gat)
--	I1734 = OR(n1604gat, n2214gat, I1733)
--	n2918gat = OR(n769gat, n759gat)
--	n2952gat = OR(n1076gat, n1075gat)
--	n2919gat = OR(n766gat, n760gat)
--	n1184gat = OR(n1185gat, n1186gat, n1187gat, n1188gat)
--	n2910gat = OR(n645gat, n644gat)
--	n2907gat = OR(n646gat, n641gat)
--	n2970gat = OR(n1383gat, n1327gat)
--	n2911gat = OR(n761gat, n651gat)
--	n2912gat = OR(n762gat, n652gat)
--	n2909gat = OR(n765gat, n643gat)
--	n1201gat = OR(n1202gat, n1203gat, n1204gat, n1205gat)
--	n1269gat = OR(n1270gat, n1271gat, n1272gat, n1273gat)
--	n2908gat = OR(n763gat, n642gat)
--	n2971gat = OR(n1287gat, n1285gat)
--	n2904gat = OR(n793gat, n664gat, n556gat)
--	n2891gat = OR(n795gat, n656gat, n368gat)
--	n2903gat = OR(n794gat, n773gat, n662gat)
--	n2915gat = OR(n965gat, n960gat, n661gat)
--	n779gat = OR(n780gat, n781gat, n782gat, n783gat)
--	n2901gat = OR(n558gat, n555gat, n450gat)
--	n2890gat = OR(n654gat, n557gat, n371gat)
--	n2876gat = OR(n874gat, n132gat)
--	n2888gat = OR(n663gat, n649gat, n449gat)
--	n2887gat = OR(n791gat, n650gat, n370gat)
--	n2886gat = OR(n774gat, n764gat, n369gat)
--	n221gat = OR(n222gat, n223gat, n224gat, n225gat)
--	n120gat = OR(n121gat, n122gat, n123gat, n124gat)
--	n3010gat = OR(n2460gat, n2423gat)
--	n3016gat = OR(n2596gat, n2595gat)
--	n2568gat = OR(n2569gat, n2570gat, n2571gat, n2572gat)
--	n2409gat = OR(n2410gat, n2411gat, n2412gat, n2413gat)
--	n2579gat = OR(n2580gat, n2581gat)
--	n3014gat = OR(n2567gat, n2499gat)
--	n2880gat = OR(n299gat, n207gat)
--	n2646gat = OR(n2647gat, n2648gat)
--	n2601gat = OR(n2602gat, n2603gat, n2604gat, n2605gat)
--	n2545gat = OR(n2546gat, n2547gat, n2548gat, n2549gat)
--	n2613gat = OR(n2614gat, n2615gat)
--	n3013gat = OR(n2461gat, n2421gat)
--	n2930gat = OR(n1153gat, n1151gat, n982gat, n877gat)
--	n2957gat = OR(n1159gat, n1158gat, n1156gat, n1155gat)
--	n2975gat = OR(n1443gat, n1325gat)
--	n2974gat = OR(n1321gat, n1320gat)
--	n2966gat = OR(n1368gat, n1258gat)
--	n2979gat = OR(n1373gat, n1372gat)
--	n2978gat = OR(n1441gat, n1440gat, n1371gat, n1367gat)
--	n2982gat = OR(n1504gat, n1502gat)
--	n2954gat = OR(n1250gat, n1103gat)
--	n2964gat = OR(n1304gat, n1249gat)
--	n2958gat = OR(n1246gat, n1161gat)
--	n2963gat = OR(n1291gat, n1245gat)
--	n2973gat = OR(n1352gat, n1351gat, n1303gat, n1302gat)
--	n2953gat = OR(n1163gat, n1102gat)
--	n2949gat = OR(n1101gat, n996gat)
--	n2934gat = OR(n1104gat, n887gat)
--	n2959gat = OR(n1305gat, n1162gat)
--	n2977gat = OR(n1360gat, n1359gat, n1358gat, n1357gat)
--	I2720 = OR(n1788gat, n1786gat, n1839gat)
--	I2721 = OR(n1884gat, n1783gat, I2720)
--	I2735 = OR(n1788gat, n1884gat, n1633gat)
--	I2736 = OR(n1785gat, n1784gat, I2735)
--	I2812 = OR(n1703gat, n1704gat, n1778gat)
--	I2813 = OR(n1609gat, n1702gat, n1700gat, I2812)
--	I2831 = OR(n1839gat, n1786gat, n1788gat)
--	I2832 = OR(n1884gat, n1784gat, I2831)
--	I2889 = OR(n1784gat, n1633gat, n1884gat)
--	I2890 = OR(n1788gat, n1786gat, I2889)
--	I2925 = OR(n1784gat, n1785gat, n1633gat)
--	I2926 = OR(n1884gat, n1787gat, I2925)
--	I2934 = OR(n1784gat, n1839gat, n1788gat)
--	I2935 = OR(n1785gat, n1884gat, I2934)
--	n2988gat = OR(n1733gat, n1581gat)
--	n2983gat = OR(n2079gat, n2073gat)
--	n2987gat = OR(n1574gat, n1573gat)
--	n2992gat = OR(n1723gat, n1647gat, n1646gat)
--	n2986gat = OR(n1650gat, n1649gat, n1563gat)
--	n2991gat = OR(n1654gat, n1653gat, n1644gat)
--	I3148 = OR(n1839gat, n1884gat, n1784gat)
--	I3149 = OR(n1786gat, n1787gat, I3148)
--	I3178 = OR(n1838gat, n1785gat, n1788gat)
--	I3179 = OR(n1839gat, n1784gat, I3178)
--	n2981gat = OR(n1413gat, n1408gat, n1407gat)
--	n3000gat = OR(n2000gat, n1999gat)
--	n3004gat = OR(n2258gat, n2257gat, n2255gat)
--	n3003gat = OR(n2256gat, n2251gat)
--	n3001gat = OR(n2132gat, n2130gat)
--	n3006gat = OR(n2253gat, n2252gat)
--	n3007gat = OR(n2250gat, n2249gat)
--	n2990gat = OR(n1710gat, n1630gat)
--	n2994gat = OR(n1954gat, n1888gat)
--	n2993gat = OR(n1894gat, n1847gat, n1846gat)
--	n2998gat = OR(n2055gat, n1967gat)
--	n2996gat = OR(n1960gat, n1959gat, n1957gat)
--	n3008gat = OR(n2332gat, n2259gat)
--	n3005gat = OR(n2211gat, n2210gat)
--	n2997gat = OR(n2053gat, n2052gat, n1964gat)
--	n3009gat = OR(n2350gat, n2282gat)
--	n3002gat = OR(n2213gat, n2150gat, n2149gat)
--	n2995gat = OR(n1962gat, n1955gat)
--	n2999gat = OR(n1972gat, n1971gat)
--	n3011gat = OR(n2333gat, n2331gat)
--	n3015gat = OR(n2566gat, n2565gat)
--	n2874gat = OR(n141gat, n38gat, n37gat)
--	n2917gat = OR(n1074gat, n872gat)
--	n2878gat = OR(n234gat, n137gat)
--	n2892gat = OR(n378gat, n377gat)
--	n2885gat = OR(n250gat, n249gat, n248gat)
--	n2900gat = OR(n869gat, n453gat, n448gat)
--	n2883gat = OR(n251gat, n244gat)
--	n2929gat = OR(n974gat, n973gat, n870gat)
--	n2884gat = OR(n246gat, n245gat)
--	n2902gat = OR(n460gat, n459gat)
--	n2925gat = OR(n975gat, n972gat, n969gat)
--	n2879gat = OR(n145gat, n143gat)
--	n2916gat = OR(n971gat, n970gat, n968gat)
--	n2875gat = OR(n142gat, n40gat, n39gat)
--	n2899gat = OR(n772gat, n451gat, n446gat)
--	n2877gat = OR(n139gat, n136gat)
--	n2893gat = OR(n391gat, n390gat)
--	n2926gat = OR(n1083gat, n1077gat)
--	n2882gat = OR(n242gat, n240gat)
--	n2924gat = OR(n871gat, n797gat)
--	n2881gat = OR(n324gat, n238gat, n237gat)
--	n2923gat = OR(n1082gat, n796gat)
--	n2710gat = OR(n69gat, n1885gat)
--	n2704gat = OR(n11gat, n1889gat)
--	n2684gat = OR(n1599gat, n2051gat)
--	n2830gat = OR(n2444gat, n1754gat)
--	I3999 = OR(n2167gat, n2031gat, n2174gat)
--	I4000 = OR(n2108gat, n2093gat, n2035gat, I3999)
--	n2695gat = OR(n1586gat, n1791gat)
--	n2703gat = OR(n1755gat, n1518gat)
--	n2744gat = OR(n2159gat, n2478gat)
--	n2800gat = OR(n2158gat, n2186gat)
--	I4023 = OR(n2443gat, n2290gat, n2214gat)
--	I4024 = OR(n2353gat, n2284gat, I4023)
--	n2980gat = OR(n1470gat, n1400gat, n1399gat, n1398gat)
--	I4144 = OR(n1633gat, n1838gat, n1786gat)
--	I4145 = OR(n1788gat, n1784gat, I4144)
--	n2984gat = OR(n1467gat, n1466gat)
--	n2985gat = OR(n1686gat, n1533gat, n1532gat, n1531gat)
--	I4216 = OR(n1427gat, n1595gat, n1677gat)
--	I4217 = OR(n1392gat, n2989gat, I4216)
--	n2931gat = OR(n1100gat, n994gat, n989gat, n880gat)
--	n2943gat = OR(n1012gat, n905gat)
--	n2941gat = OR(n1003gat, n902gat)
--	n2946gat = OR(n1099gat, n998gat, n995gat, n980gat)
--	n2960gat = OR(n1175gat, n1174gat)
--	n2950gat = OR(n1001gat, n999gat)
--	n2969gat = OR(n1323gat, n1264gat)
--	n2933gat = OR(n981gat, n890gat, n889gat, n886gat)
--	n2935gat = OR(n892gat, n891gat)
--	n2942gat = OR(n904gat, n903gat)
--	n2940gat = OR(n1152gat, n1092gat, n997gat, n993gat)
--	n2937gat = OR(n900gat, n895gat)
--	n2947gat = OR(n1094gat, n1093gat, n988gat, n984gat)
--	n2965gat = OR(n1267gat, n1257gat)
--	n2956gat = OR(n1178gat, n1116gat)
--	n2961gat = OR(n1375gat, n1324gat)
--	n2939gat = OR(n1091gat, n1088gat, n992gat, n987gat)
--	n2938gat = OR(n899gat, n896gat)
--	n2967gat = OR(n1262gat, n1260gat)
--	n2932gat = OR(n1098gat, n1090gat, n986gat, n885gat)
--	n2936gat = OR(n901gat, n893gat)
--	n2948gat = OR(n1097gat, n1089gat, n1087gat, n991gat)
--	n2968gat = OR(n1326gat, n1261gat)
--	n2955gat = OR(n1177gat, n1115gat)
--	n2944gat = OR(n977gat, n976gat)
--	n2945gat = OR(n1096gat, n1095gat, n990gat, n979gat)
--	n2962gat = OR(n1176gat, n1173gat)
--	n2951gat = OR(n1004gat, n1000gat)
--	n2764gat = OR(n1029gat, n2237gat)
--	n2762gat = OR(n1028gat, n1782gat)
--	n2761gat = OR(n1031gat, n2325gat)
--	n2757gat = OR(n1030gat, n2245gat)
--	n2756gat = OR(n1011gat, n2244gat)
--	n2750gat = OR(n1181gat, n2243gat)
--	n2749gat = OR(n1010gat, n2246gat)
--	n2742gat = OR(n1005gat, n2384gat)
--	n2741gat = OR(n1182gat, n2385gat)
--	n2694gat = OR(n1381gat, n1384gat)
--	n2693gat = OR(n1451gat, n1453gat)
--	n2702gat = OR(n925gat, n1452gat)
--	n2701gat = OR(n921gat, n1890gat)
--	n2709gat = OR(n739gat, n1841gat)
--	n2708gat = OR(n848gat, n2047gat)
--	n2799gat = OR(n849gat, n2050gat)
--	n2798gat = OR(n1032gat, n2054gat)
--	n2812gat = OR(n73gat, n70gat, n1840gat)
--	n2822gat = OR(n77gat, n13gat, n1842gat)
--	
--	n421gat = NOR(n2715gat, n2723gat)
--	n648gat = NOR(n373gat, n2669gat)
--	n442gat = NOR(n2844gat, n856gat)
--	n1499gat = NOR(n396gat, n401gat)
--	n1616gat = NOR(n918gat, n396gat)
--	n1614gat = NOR(n396gat, n845gat)
--	n1641gat = NOR(n1645gat, n1553gat, n1559gat)
--	n1642gat = NOR(n1559gat, n1616gat, n1645gat)
--	n1556gat = NOR(n1614gat, n1645gat, n1616gat)
--	n1557gat = NOR(n1553gat, n1645gat, n1614gat)
--	n1639gat = NOR(n1499gat, n1559gat, n1553gat)
--	n1605gat = NOR(n1614gat, n1616gat, n1499gat, n396gat)
--	n1555gat = NOR(n1616gat, n1559gat, n1499gat)
--	n1558gat = NOR(n1614gat, n1553gat, n1499gat)
--	n1256gat = NOR(n392gat, n702gat)
--	n1117gat = NOR(n720gat, n725gat)
--	n1618gat = NOR(n1319gat, n1447gat)
--	n1114gat = NOR(n725gat, n721gat)
--	n1621gat = NOR(n1319gat, n1380gat)
--	n1318gat = NOR(n392gat, n701gat)
--	n1619gat = NOR(n1447gat, n1446gat)
--	n1622gat = NOR(n1380gat, n1446gat)
--	n1214gat = NOR(n1218gat, n1219gat, n1220gat)
--	n1215gat = NOR(n1218gat, n1221gat, n1222gat)
--	n1216gat = NOR(n1223gat, n1219gat, n1222gat)
--	n1217gat = NOR(n1223gat, n1221gat, n1220gat)
--	n745gat = NOR(n2716gat, n2867gat)
--	n638gat = NOR(n2715gat, n2868gat)
--	n423gat = NOR(n2724gat, n2726gat)
--	n362gat = NOR(n2723gat, n2727gat)
--	n749gat = NOR(n753gat, n754gat, n755gat)
--	n750gat = NOR(n753gat, n756gat, n757gat)
--	n751gat = NOR(n758gat, n754gat, n757gat)
--	n752gat = NOR(n758gat, n756gat, n755gat)
--	n259gat = NOR(n263gat, n264gat, n265gat)
--	n260gat = NOR(n263gat, n266gat, n267gat)
--	n261gat = NOR(n268gat, n264gat, n267gat)
--	n262gat = NOR(n268gat, n266gat, n265gat)
--	n1014gat = NOR(n1018gat, n1019gat, n1020gat)
--	n1015gat = NOR(n1018gat, n1021gat, n1022gat)
--	n1016gat = NOR(n1023gat, n1019gat, n1022gat)
--	n1017gat = NOR(n1023gat, n1021gat, n1020gat)
--	n476gat = NOR(n480gat, n481gat, n482gat)
--	n477gat = NOR(n480gat, n483gat, n484gat)
--	n478gat = NOR(n485gat, n481gat, n484gat)
--	n479gat = NOR(n485gat, n483gat, n482gat)
--	n44gat = NOR(n48gat, n49gat, n50gat)
--	n45gat = NOR(n48gat, n51gat, n52gat)
--	n46gat = NOR(n53gat, n49gat, n52gat)
--	n47gat = NOR(n53gat, n51gat, n50gat)
--	n1376gat = NOR(n724gat, n720gat)
--	n1617gat = NOR(n1319gat, n1448gat)
--	n1377gat = NOR(n724gat, n721gat)
--	n1624gat = NOR(n1319gat, n1379gat)
--	n1113gat = NOR(n393gat, n701gat)
--	n1501gat = NOR(n1448gat, n1500gat)
--	n1623gat = NOR(n1379gat, n1446gat)
--	n1620gat = NOR(n1448gat, n1446gat)
--	n1827gat = NOR(n2729gat, n2317gat)
--	n1817gat = NOR(n1819gat, n1823gat)
--	n1935gat = NOR(n1816gat, n1828gat)
--	n529gat = NOR(n2724gat, n2715gat)
--	n361gat = NOR(n2859gat, n2726gat)
--	n168gat = NOR(n172gat, n173gat, n174gat)
--	n169gat = NOR(n172gat, n175gat, n176gat)
--	n170gat = NOR(n177gat, n173gat, n176gat)
--	n171gat = NOR(n177gat, n175gat, n174gat)
--	n907gat = NOR(n911gat, n912gat, n913gat)
--	n908gat = NOR(n911gat, n914gat, n915gat)
--	n909gat = NOR(n916gat, n912gat, n915gat)
--	n910gat = NOR(n916gat, n914gat, n913gat)
--	n344gat = NOR(n348gat, n349gat, n350gat)
--	n345gat = NOR(n348gat, n351gat, n352gat)
--	n346gat = NOR(n353gat, n349gat, n352gat)
--	n347gat = NOR(n353gat, n351gat, n350gat)
--	n56gat = NOR(n60gat, n61gat, n62gat)
--	n57gat = NOR(n60gat, n63gat, n64gat)
--	n58gat = NOR(n65gat, n61gat, n64gat)
--	n59gat = NOR(n65gat, n63gat, n62gat)
--	n768gat = NOR(n373gat, n2731gat)
--	n655gat = NOR(n856gat, n2718gat)
--	n963gat = NOR(n856gat, n2838gat)
--	n868gat = NOR(n2775gat, n373gat)
--	n962gat = NOR(n856gat, n2711gat)
--	n959gat = NOR(n373gat, n2734gat)
--	n945gat = NOR(n949gat, n950gat, n951gat)
--	n946gat = NOR(n949gat, n952gat, n953gat)
--	n947gat = NOR(n954gat, n950gat, n953gat)
--	n948gat = NOR(n954gat, n952gat, n951gat)
--	n647gat = NOR(n2792gat, n373gat)
--	n441gat = NOR(n856gat, n2846gat)
--	n967gat = NOR(n373gat, n2672gat)
--	n792gat = NOR(n2852gat, n856gat)
--	n1229gat = NOR(n1233gat, n1234gat, n1235gat)
--	n1230gat = NOR(n1233gat, n1236gat, n1237gat)
--	n1231gat = NOR(n1238gat, n1234gat, n1237gat)
--	n1232gat = NOR(n1238gat, n1236gat, n1235gat)
--	n443gat = NOR(n2778gat, n373gat)
--	n439gat = NOR(n856gat, n2836gat)
--	n966gat = NOR(n2789gat, n373gat)
--	n790gat = NOR(n856gat, n2840gat)
--	n444gat = NOR(n373gat, n2781gat)
--	n440gat = NOR(n856gat, n2842gat)
--	n1051gat = NOR(n1055gat, n1056gat, n1057gat)
--	n1052gat = NOR(n1055gat, n1058gat, n1059gat)
--	n1053gat = NOR(n1060gat, n1056gat, n1059gat)
--	n1054gat = NOR(n1060gat, n1058gat, n1057gat)
--	n934gat = NOR(n938gat, n939gat, n940gat)
--	n935gat = NOR(n938gat, n941gat, n942gat)
--	n936gat = NOR(n943gat, n939gat, n942gat)
--	n937gat = NOR(n943gat, n941gat, n940gat)
--	n746gat = NOR(n2716gat, n2723gat)
--	n360gat = NOR(n2859gat, n2727gat)
--	n710gat = NOR(n714gat, n715gat, n716gat)
--	n711gat = NOR(n714gat, n717gat, n718gat)
--	n712gat = NOR(n719gat, n715gat, n718gat)
--	n713gat = NOR(n719gat, n717gat, n716gat)
--	n729gat = NOR(n733gat, n734gat, n735gat)
--	n730gat = NOR(n733gat, n736gat, n737gat)
--	n731gat = NOR(n738gat, n734gat, n737gat)
--	n732gat = NOR(n738gat, n736gat, n735gat)
--	n494gat = NOR(n498gat, n499gat, n500gat)
--	n495gat = NOR(n498gat, n501gat, n502gat)
--	n496gat = NOR(n503gat, n499gat, n502gat)
--	n497gat = NOR(n503gat, n501gat, n500gat)
--	n505gat = NOR(n509gat, n510gat, n511gat)
--	n506gat = NOR(n509gat, n512gat, n513gat)
--	n507gat = NOR(n514gat, n510gat, n513gat)
--	n508gat = NOR(n514gat, n512gat, n511gat)
--	n564gat = NOR(n3029gat, n2863gat, n2855gat, n374gat)
--	n86gat = NOR(n743gat, n294gat, n17gat)
--	n78gat = NOR(n2784gat, n79gat)
--	n767gat = NOR(n219gat, n2731gat)
--	n286gat = NOR(n289gat, n2723gat)
--	n287gat = NOR(n289gat, n2715gat)
--	n288gat = NOR(n289gat, n2726gat)
--	n181gat = NOR(n286gat, n179gat, n188gat)
--	n182gat = NOR(n72gat, n2720gat)
--	n653gat = NOR(n2718gat, n111gat)
--	n867gat = NOR(n219gat, n2775gat)
--	n771gat = NOR(n2838gat, n111gat)
--	n964gat = NOR(n111gat, n2711gat)
--	n961gat = NOR(n219gat, n2734gat)
--	n804gat = NOR(n808gat, n809gat, n810gat)
--	n805gat = NOR(n808gat, n811gat, n812gat)
--	n806gat = NOR(n813gat, n809gat, n812gat)
--	n807gat = NOR(n813gat, n811gat, n810gat)
--	n587gat = NOR(n591gat, n592gat, n593gat)
--	n588gat = NOR(n591gat, n594gat, n595gat)
--	n589gat = NOR(n596gat, n592gat, n595gat)
--	n590gat = NOR(n596gat, n594gat, n593gat)
--	n447gat = NOR(n2836gat, n111gat)
--	n445gat = NOR(n2778gat, n219gat)
--	n687gat = NOR(n691gat, n692gat, n693gat)
--	n688gat = NOR(n691gat, n694gat, n695gat)
--	n689gat = NOR(n696gat, n692gat, n695gat)
--	n690gat = NOR(n696gat, n694gat, n693gat)
--	n568gat = NOR(n572gat, n573gat, n574gat)
--	n569gat = NOR(n572gat, n575gat, n576gat)
--	n570gat = NOR(n577gat, n573gat, n576gat)
--	n571gat = NOR(n577gat, n575gat, n574gat)
--	n187gat = NOR(n189gat, n287gat, n188gat)
--	n197gat = NOR(n194gat, n297gat)
--	n15gat = NOR(n637gat, n17gat, n293gat)
--	n22gat = NOR(n92gat, n21gat)
--	n93gat = NOR(n197gat, n22gat)
--	n769gat = NOR(n93gat, n2731gat)
--	n2534gat = NOR(n2624gat, n2489gat, n2621gat)
--	n2430gat = NOR(n2533gat, n2486gat, n2429gat)
--	n1606gat = NOR(n3020gat, n270gat)
--	n2239gat = NOR(n2850gat, n3019gat)
--	n1934gat = NOR(n2470gat, n1935gat, n2239gat)
--	n1610gat = NOR(n1698gat, n1543gat)
--	n1692gat = NOR(n1879gat, n1762gat)
--	n2433gat = NOR(n2432gat, n2154gat)
--	n2531gat = NOR(n2488gat, n2625gat, n2621gat)
--	n2480gat = NOR(n2530gat, n2482gat, n2486gat)
--	n2427gat = NOR(n2426gat, n2153gat)
--	n2428gat = NOR(n2433gat, n2427gat)
--	n1778gat = NOR(n3026gat, n1779gat)
--	n1609gat = NOR(n1503gat, n3025gat)
--	n1702gat = NOR(n3024gat, n1615gat)
--	n1700gat = NOR(n1701gat, n3023gat)
--	n1604gat = NOR(n1778gat, n1609gat, n1702gat, n1700gat)
--	n1076gat = NOR(n93gat, n2775gat)
--	n766gat = NOR(n93gat, n2734gat)
--	n1185gat = NOR(n1189gat, n1190gat, n1191gat)
--	n1186gat = NOR(n1189gat, n1192gat, n1193gat)
--	n1187gat = NOR(n1194gat, n1190gat, n1193gat)
--	n1188gat = NOR(n1194gat, n1192gat, n1191gat)
--	n645gat = NOR(n2792gat, n93gat)
--	n646gat = NOR(n93gat, n2669gat)
--	n1383gat = NOR(n1280gat, n1225gat)
--	n1327gat = NOR(n1281gat, n1224gat)
--	n651gat = NOR(n93gat, n2778gat)
--	n652gat = NOR(n2789gat, n93gat)
--	n765gat = NOR(n2781gat, n93gat)
--	n1202gat = NOR(n1206gat, n1207gat, n1208gat)
--	n1203gat = NOR(n1206gat, n1209gat, n1210gat)
--	n1204gat = NOR(n1211gat, n1207gat, n1210gat)
--	n1205gat = NOR(n1211gat, n1209gat, n1208gat)
--	n1270gat = NOR(n1274gat, n1275gat, n1276gat)
--	n1271gat = NOR(n1274gat, n1277gat, n1278gat)
--	n1272gat = NOR(n1279gat, n1275gat, n1278gat)
--	n1273gat = NOR(n1279gat, n1277gat, n1276gat)
--	n763gat = NOR(n2672gat, n93gat)
--	n1287gat = NOR(n1284gat, n1195gat)
--	n1285gat = NOR(n1196gat, n1269gat)
--	n853gat = NOR(n740gat, n2148gat)
--	n793gat = NOR(n2852gat, n851gat)
--	n854gat = NOR(n2148gat, n374gat)
--	n556gat = NOR(n2672gat, n852gat)
--	n795gat = NOR(n2731gat, n852gat)
--	n656gat = NOR(n851gat, n2718gat)
--	n794gat = NOR(n852gat, n2775gat)
--	n773gat = NOR(n851gat, n2838gat)
--	n965gat = NOR(n2711gat, n851gat)
--	n960gat = NOR(n2734gat, n852gat)
--	n780gat = NOR(n784gat, n785gat, n786gat)
--	n781gat = NOR(n784gat, n787gat, n788gat)
--	n782gat = NOR(n789gat, n785gat, n788gat)
--	n783gat = NOR(n789gat, n787gat, n786gat)
--	n555gat = NOR(n852gat, n2792gat)
--	n450gat = NOR(n851gat, n2846gat)
--	n654gat = NOR(n851gat, n2844gat)
--	n557gat = NOR(n2669gat, n852gat)
--	n874gat = NOR(n559gat, n365gat)
--	n132gat = NOR(n560gat, n364gat)
--	n649gat = NOR(n2778gat, n852gat)
--	n449gat = NOR(n2836gat, n851gat)
--	n791gat = NOR(n851gat, n2840gat)
--	n650gat = NOR(n852gat, n2789gat)
--	n774gat = NOR(n2842gat, n851gat)
--	n764gat = NOR(n852gat, n2781gat)
--	n222gat = NOR(n226gat, n227gat, n228gat)
--	n223gat = NOR(n226gat, n229gat, n230gat)
--	n224gat = NOR(n231gat, n227gat, n230gat)
--	n225gat = NOR(n231gat, n229gat, n228gat)
--	n121gat = NOR(n125gat, n126gat, n127gat)
--	n122gat = NOR(n125gat, n128gat, n129gat)
--	n123gat = NOR(n130gat, n126gat, n129gat)
--	n124gat = NOR(n130gat, n128gat, n127gat)
--	n2460gat = NOR(n666gat, n120gat)
--	n2423gat = NOR(n665gat, n1601gat)
--	n2594gat = NOR(n3017gat, n2520gat, n2597gat)
--	n2569gat = NOR(n2573gat, n2574gat, n2575gat)
--	n2570gat = NOR(n2573gat, n2576gat, n2577gat)
--	n2571gat = NOR(n2578gat, n2574gat, n2577gat)
--	n2572gat = NOR(n2578gat, n2576gat, n2575gat)
--	n2410gat = NOR(n2414gat, n2415gat, n2416gat)
--	n2411gat = NOR(n2414gat, n2417gat, n2418gat)
--	n2412gat = NOR(n2419gat, n2415gat, n2418gat)
--	n2413gat = NOR(n2419gat, n2417gat, n2416gat)
--	n2583gat = NOR(n2582gat, n2585gat)
--	n2580gat = NOR(n2582gat, n2583gat)
--	n2581gat = NOR(n2583gat, n2585gat)
--	n2567gat = NOR(n2493gat, n2388gat)
--	n2499gat = NOR(n2389gat, n2494gat)
--	n299gat = NOR(n2268gat, n2338gat)
--	n207gat = NOR(n2337gat, n2269gat)
--	n2650gat = NOR(n2649gat, n2652gat)
--	n2647gat = NOR(n2649gat, n2650gat)
--	n2648gat = NOR(n2650gat, n2652gat)
--	n2602gat = NOR(n2606gat, n2607gat, n2608gat)
--	n2603gat = NOR(n2606gat, n2609gat, n2610gat)
--	n2604gat = NOR(n2611gat, n2607gat, n2610gat)
--	n2605gat = NOR(n2611gat, n2609gat, n2608gat)
--	n2546gat = NOR(n2550gat, n2551gat, n2552gat)
--	n2547gat = NOR(n2550gat, n2553gat, n2554gat)
--	n2548gat = NOR(n2555gat, n2551gat, n2554gat)
--	n2549gat = NOR(n2555gat, n2553gat, n2552gat)
--	n2617gat = NOR(n2616gat, n2619gat)
--	n2614gat = NOR(n2616gat, n2617gat)
--	n2615gat = NOR(n2617gat, n2619gat)
--	n2655gat = NOR(n2508gat, n2656gat, n2500gat, n2504gat)
--	n2293gat = NOR(n2353gat, n2284gat, n2443gat)
--	n2219gat = NOR(n2354gat, n2214gat)
--	n1529gat = NOR(n1528gat, n1523gat)
--	n1704gat = NOR(n3027gat, n1706gat)
--	n2461gat = NOR(n120gat, n2666gat)
--	n2421gat = NOR(n1601gat, n1704gat)
--	n1598gat = NOR(n1592gat, n2422gat)
--	n2218gat = NOR(n2214gat, n2290gat)
--	n2358gat = NOR(n2285gat, n2356gat, n2355gat)
--	n1415gat = NOR(n2081gat, n2359gat)
--	n1153gat = NOR(n1414gat, n566gat)
--	n2292gat = NOR(n2443gat, n2284gat, n2285gat)
--	n1416gat = NOR(n2081gat, n1480gat)
--	n1151gat = NOR(n1301gat, n1150gat)
--	n2306gat = NOR(n2356gat, n2284gat, n2285gat)
--	n1481gat = NOR(n2081gat, n2011gat)
--	n982gat = NOR(n873gat, n1478gat)
--	n2357gat = NOR(n2285gat, n2355gat, n2443gat)
--	n1347gat = NOR(n2081gat, n1410gat)
--	n877gat = NOR(n875gat, n876gat)
--	n1484gat = NOR(n2081gat, n1528gat)
--	n1159gat = NOR(n1160gat, n1084gat)
--	n2363gat = NOR(n2353gat, n2356gat, n2355gat)
--	n1483gat = NOR(n2081gat, n1482gat)
--	n1158gat = NOR(n983gat, n1157gat)
--	n2364gat = NOR(n2353gat, n2284gat, n2356gat)
--	n1308gat = NOR(n2081gat, n1530gat)
--	n1156gat = NOR(n985gat, n1307gat)
--	n2291gat = NOR(n2353gat, n2355gat, n2443gat)
--	n1349gat = NOR(n1479gat, n2081gat)
--	n1155gat = NOR(n1085gat, n1348gat)
--	n1154gat = NOR(n1598gat, n2930gat, n2957gat)
--	n1703gat = NOR(n1705gat, n3028gat)
--	n1608gat = NOR(n1704gat, n1703gat)
--	n1411gat = NOR(n1154gat, n1608gat)
--	n2223gat = NOR(n2354gat, n2217gat)
--	n1438gat = NOR(n1591gat, n1480gat)
--	n1625gat = NOR(n3021gat, n1628gat)
--	n1626gat = NOR(n1627gat, n3022gat)
--	n1831gat = NOR(n1832gat, n1765gat, n1878gat)
--	n1443gat = NOR(n1442gat, n706gat)
--	n1325gat = NOR(n1444gat, n164gat)
--	n1441gat = NOR(n1437gat, n1378gat)
--	n1321gat = NOR(n1442gat, n837gat)
--	n1320gat = NOR(n1444gat, n278gat)
--	n1486gat = NOR(n1482gat, n1591gat)
--	n1440gat = NOR(n1322gat, n1439gat)
--	n1426gat = NOR(n2011gat, n1591gat)
--	n1368gat = NOR(n1442gat, n613gat)
--	n1258gat = NOR(n274gat, n1444gat)
--	n1371gat = NOR(n1370gat, n1369gat)
--	n1365gat = NOR(n1479gat, n1591gat)
--	n1373gat = NOR(n833gat, n1442gat)
--	n1372gat = NOR(n282gat, n1444gat)
--	n1367gat = NOR(n1366gat, n1374gat)
--	n2220gat = NOR(n2290gat, n2217gat)
--	n1423gat = NOR(n2162gat, n1530gat)
--	n1498gat = NOR(n1609gat, n1427gat)
--	n1504gat = NOR(n1450gat, n1498gat)
--	n1607gat = NOR(n2082gat, n1609gat)
--	n1494gat = NOR(n1528gat, n2162gat)
--	n1502gat = NOR(n1607gat, n1449gat)
--	n1250gat = NOR(n1603gat, n815gat)
--	n1103gat = NOR(n956gat, n1590gat)
--	n1417gat = NOR(n2162gat, n1480gat)
--	n1352gat = NOR(n1248gat, n1418gat)
--	n1304gat = NOR(n1590gat, n1067gat)
--	n1249gat = NOR(n679gat, n1603gat)
--	n1419gat = NOR(n2162gat, n1479gat)
--	n1351gat = NOR(n1306gat, n1353gat)
--	n1246gat = NOR(n864gat, n1590gat)
--	n1161gat = NOR(n583gat, n1603gat)
--	n1422gat = NOR(n2011gat, n2162gat)
--	n1303gat = NOR(n1247gat, n1355gat)
--	n1291gat = NOR(n1603gat, n579gat)
--	n1245gat = NOR(n1590gat, n860gat)
--	n1485gat = NOR(n1482gat, n2162gat)
--	n1302gat = NOR(n1300gat, n1487gat)
--	n1163gat = NOR(n882gat, n1603gat)
--	n1102gat = NOR(n1297gat, n1590gat)
--	n1354gat = NOR(n1591gat, n1530gat)
--	n1360gat = NOR(n1164gat, n1356gat)
--	n1435gat = NOR(n1591gat, n1528gat)
--	n1101gat = NOR(n1590gat, n1293gat)
--	n996gat = NOR(n1603gat, n823gat)
--	n1359gat = NOR(n1436gat, n1106gat)
--	n1421gat = NOR(n2162gat, n2359gat)
--	n1104gat = NOR(n1079gat, n1590gat)
--	n887gat = NOR(n1603gat, n683gat)
--	n1358gat = NOR(n1425gat, n1105gat)
--	n1420gat = NOR(n1410gat, n2162gat)
--	n1305gat = NOR(n1147gat, n1590gat)
--	n1162gat = NOR(n698gat, n1603gat)
--	n1357gat = NOR(n1424gat, n1309gat)
--	n1428gat = NOR(n2978gat, n2982gat, n2973gat, n2977gat)
--	n1794gat = NOR(n1673gat, n1719gat)
--	n1796gat = NOR(n1858gat, n1635gat)
--	n1792gat = NOR(n1794gat, n1796gat)
--	n1865gat = NOR(n1989gat, n1918gat, n1986gat)
--	n1861gat = NOR(n1866gat, n2216gat, n1988gat)
--	n1793gat = NOR(n1792gat, n1735gat)
--	n1406gat = NOR(n1428gat, n1387gat)
--	n1780gat = NOR(n1777gat, n1625gat, n1626gat)
--	n2016gat = NOR(n2019gat, n1878gat)
--	n2664gat = NOR(n2850gat, n3018gat)
--	n1666gat = NOR(n1986gat, n2212gat, n1991gat)
--	n1578gat = NOR(n2152gat, n2351gat, n1665gat)
--	n1516gat = NOR(n1551gat, n1517gat)
--	n1864gat = NOR(n1858gat, n1495gat, n2090gat)
--	n1565gat = NOR(n1735gat, n1552gat)
--	n1921gat = NOR(n1738gat, n1673gat)
--	n1798gat = NOR(n1739gat, n1673gat)
--	n1920gat = NOR(n1864gat, n1921gat, n1798gat)
--	n1926gat = NOR(n1925gat, n1635gat)
--	n1916gat = NOR(n1917gat, n1859gat)
--	n1994gat = NOR(n1719gat, n1922gat)
--	n1924gat = NOR(n1743gat, n1923gat)
--	n2078gat = NOR(n1926gat, n1916gat, n1994gat, n1924gat)
--	n1690gat = NOR(n1700gat, n1702gat)
--	n1660gat = NOR(n1918gat, n1986gat, n2212gat)
--	n1576gat = NOR(n2351gat, n1988gat, n1661gat)
--	n1733gat = NOR(n1673gat, n1572gat)
--	n1582gat = NOR(n2283gat, n1991gat, n2212gat)
--	n1577gat = NOR(n1520gat, n2351gat, n1988gat)
--	n1581gat = NOR(n1858gat, n1580gat)
--	n2129gat = NOR(n2189gat, n2134gat, n2261gat)
--	n2079gat = NOR(n2078gat, n2178gat, n1990gat, n2128gat)
--	n1695gat = NOR(n1609gat, n1778gat, n1704gat, n1703gat)
--	n2073gat = NOR(n2078gat, n1990gat, n2181gat)
--	n1696gat = NOR(n1707gat, n1698gat)
--	n1758gat = NOR(n1311gat, n1773gat)
--	n1574gat = NOR(n1719gat, n1673gat, n1444gat)
--	n1573gat = NOR(n1444gat, n1858gat, n1635gat)
--	n1521gat = NOR(n2283gat, n1991gat)
--	n1737gat = NOR(n2212gat, n2152gat)
--	n1732gat = NOR(n1515gat, n1736gat, n1658gat)
--	n1723gat = NOR(n1659gat, n1722gat, n1724gat)
--	n1663gat = NOR(n1986gat, n1918gat)
--	n1655gat = NOR(n1736gat, n1662gat, n1658gat)
--	n1647gat = NOR(n1656gat, n1659gat, n1554gat)
--	n1667gat = NOR(n1991gat, n1986gat)
--	n1570gat = NOR(n1736gat, n1658gat, n1670gat)
--	n1646gat = NOR(n1569gat, n1659gat, n1566gat)
--	n1575gat = NOR(n1918gat, n2283gat)
--	n1728gat = NOR(n1568gat, n1736gat, n1658gat)
--	n1650gat = NOR(n1727gat, n1659gat, n1640gat)
--	n1801gat = NOR(n2152gat, n1989gat)
--	n1731gat = NOR(n1658gat, n1515gat, n1797gat)
--	n1649gat = NOR(n1560gat, n1659gat, n1730gat)
--	n1571gat = NOR(n1670gat, n1658gat, n1797gat)
--	n1563gat = NOR(n1561gat, n1562gat, n1659gat)
--	n1734gat = NOR(n1988gat, n2212gat)
--	n1669gat = NOR(n1668gat, n1742gat, n1670gat)
--	n1654gat = NOR(n1671gat, n1659gat)
--	n1657gat = NOR(n1662gat, n1797gat, n1658gat)
--	n1653gat = NOR(n1651gat, n1652gat, n1659gat)
--	n1729gat = NOR(n1658gat, n1797gat, n1568gat)
--	n1644gat = NOR(n1643gat, n1648gat, n1659gat)
--	n1726gat = NOR(n2992gat, n2986gat, n2991gat)
--	n1929gat = NOR(n1758gat, n1790gat)
--	n2009gat = NOR(n2016gat, n2664gat, n2004gat)
--	n1413gat = NOR(n1869gat, n672gat, n2591gat)
--	n1636gat = NOR(n1584gat, n1718gat)
--	n1401gat = NOR(n1584gat, n1590gat)
--	n1408gat = NOR(n1507gat, n1396gat, n1393gat)
--	n1476gat = NOR(n1858gat, n1590gat)
--	n1407gat = NOR(n1393gat, n1409gat, n1677gat)
--	n1412gat = NOR(n1411gat, n1406gat, n2981gat)
--	n2663gat = NOR(n2586gat, n2660gat, n2307gat)
--	n2662gat = NOR(n2660gat, n2586gat)
--	n2238gat = NOR(n2448gat, n2444gat)
--	n87gat = NOR(n743gat, n17gat, n293gat)
--	n200gat = NOR(n199gat, n92gat)
--	n184gat = NOR(n189gat, n188gat, n179gat)
--	n196gat = NOR(n297gat, n195gat)
--	n204gat = NOR(n200gat, n196gat)
--	n2163gat = NOR(n1790gat, n1310gat, n2664gat, n2168gat)
--	n2258gat = NOR(n2260gat, n2189gat)
--	n2255gat = NOR(n2261gat, n2188gat)
--	n2015gat = NOR(n2039gat, n1774gat, n1315gat)
--	n2017gat = NOR(n1790gat, n2016gat)
--	n2018gat = NOR(n2016gat, n2097gat)
--	n2014gat = NOR(n2035gat, n2093gat, n2018gat, n2664gat)
--	n2194gat = NOR(n2187gat, n1855gat)
--	n2192gat = NOR(n2184gat, n1855gat)
--	n2185gat = NOR(n2261gat, n2189gat)
--	n2132gat = NOR(n2133gat, n2131gat)
--	n2130gat = NOR(n2134gat, n2185gat)
--	n2057gat = NOR(n2049gat, n1855gat)
--	n2250gat = NOR(n2248gat, n2264gat)
--	n2249gat = NOR(n2265gat, n3006gat)
--	n2329gat = NOR(n1855gat, n3007gat)
--	n1958gat = NOR(n1963gat, n1886gat)
--	n1895gat = NOR(n1845gat, n1891gat, n1968gat)
--	n1710gat = NOR(n1709gat, n1629gat)
--	n1630gat = NOR(n1895gat, n1631gat)
--	n2195gat = NOR(n2200gat, n1855gat)
--	n2556gat = NOR(n1711gat, n2437gat)
--	n2539gat = NOR(n2048gat, n2437gat)
--	n1894gat = NOR(n1968gat, n1891gat, n1969gat)
--	n1847gat = NOR(n1958gat, n1845gat)
--	n1846gat = NOR(n1845gat, n1893gat)
--	n2436gat = NOR(n2437gat, n1892gat)
--	n2055gat = NOR(n1891gat, n1958gat)
--	n1967gat = NOR(n1893gat, n1968gat)
--	n2387gat = NOR(n2056gat, n2437gat)
--	n1959gat = NOR(n1956gat, n1963gat)
--	n1957gat = NOR(n1886gat, n1887gat)
--	n2330gat = NOR(n2437gat, n1961gat)
--	n2147gat = NOR(n2988gat, n1855gat)
--	n2498gat = NOR(n2199gat, n2328gat)
--	n2193gat = NOR(n2393gat, n2439gat)
--	n2211gat = NOR(n2193gat, n2402gat)
--	n2210gat = NOR(n2401gat, n2151gat)
--	n2396gat = NOR(n2199gat, n2209gat)
--	n2053gat = NOR(n2393gat, n2438gat)
--	n1964gat = NOR(n2392gat, n2439gat)
--	n2198gat = NOR(n2199gat, n2058gat)
--	n2215gat = NOR(n2346gat, n2151gat, n2402gat)
--	n2350gat = NOR(n2405gat, n2349gat)
--	n2282gat = NOR(n2406gat, n2215gat)
--	n2197gat = NOR(n2199gat, n2281gat)
--	n2213gat = NOR(n2402gat, n2151gat, n2345gat)
--	n2150gat = NOR(n2401gat, n2346gat)
--	n2149gat = NOR(n2193gat, n2346gat)
--	n2196gat = NOR(n2199gat, n2146gat)
--	n1882gat = NOR(n2124gat, n2115gat, n2239gat)
--	n1962gat = NOR(n1963gat, n1893gat)
--	n1896gat = NOR(n2995gat, n1895gat)
--	n1972gat = NOR(n1974gat, n1970gat)
--	n1971gat = NOR(n1896gat, n1973gat)
--	n2559gat = NOR(n2999gat, n2437gat)
--	n2331gat = NOR(n2393gat, n2401gat)
--	n2352gat = NOR(n3011gat, n2215gat)
--	n2566gat = NOR(n2643gat, n2564gat)
--	n2565gat = NOR(n2352gat, n2642gat)
--	n2637gat = NOR(n3015gat, n2199gat)
--	n84gat = NOR(n296gat, n17gat, n294gat)
--	n89gat = NOR(n88gat, n2784gat)
--	n110gat = NOR(n182gat, n89gat)
--	n1074gat = NOR(n2775gat, n110gat)
--	n141gat = NOR(n155gat, n253gat, n150gat)
--	n38gat = NOR(n151gat, n233gat)
--	n37gat = NOR(n151gat, n154gat)
--	n872gat = NOR(n375gat, n800gat)
--	n234gat = NOR(n155gat, n233gat)
--	n137gat = NOR(n154gat, n253gat)
--	n378gat = NOR(n375gat, n235gat)
--	n377gat = NOR(n110gat, n2778gat)
--	n869gat = NOR(n219gat, n2792gat)
--	n212gat = NOR(n182gat, n78gat)
--	n250gat = NOR(n329gat, n387gat, n334gat)
--	n249gat = NOR(n386gat, n330gat)
--	n248gat = NOR(n330gat, n1490gat)
--	n453gat = NOR(n372gat, n452gat)
--	n448gat = NOR(n111gat, n2846gat)
--	n974gat = NOR(n2844gat, n111gat)
--	n251gat = NOR(n1490gat, n387gat)
--	n244gat = NOR(n334gat, n386gat)
--	n973gat = NOR(n372gat, n333gat)
--	n870gat = NOR(n2669gat, n219gat)
--	n975gat = NOR(n111gat, n2852gat)
--	n246gat = NOR(n330gat, n325gat, n334gat)
--	n245gat = NOR(n386gat, n334gat)
--	n460gat = NOR(n462gat, n2884gat)
--	n459gat = NOR(n457gat, n461gat)
--	n972gat = NOR(n372gat, n458gat)
--	n969gat = NOR(n219gat, n2672gat)
--	n971gat = NOR(n111gat, n2840gat)
--	n247gat = NOR(n334gat, n387gat, n330gat)
--	n145gat = NOR(n144gat, n325gat)
--	n143gat = NOR(n326gat, n247gat)
--	n970gat = NOR(n372gat, n878gat)
--	n968gat = NOR(n2789gat, n219gat)
--	n772gat = NOR(n111gat, n2842gat)
--	n142gat = NOR(n382gat, n326gat, n144gat)
--	n40gat = NOR(n325gat, n383gat)
--	n39gat = NOR(n383gat, n247gat)
--	n451gat = NOR(n134gat, n372gat)
--	n446gat = NOR(n219gat, n2781gat)
--	n139gat = NOR(n253gat, n151gat, n254gat)
--	n136gat = NOR(n253gat, n154gat)
--	n391gat = NOR(n252gat, n468gat)
--	n390gat = NOR(n469gat, n2877gat)
--	n1083gat = NOR(n381gat, n375gat)
--	n1077gat = NOR(n110gat, n2672gat)
--	n140gat = NOR(n151gat, n253gat, n155gat)
--	n242gat = NOR(n254gat, n241gat)
--	n240gat = NOR(n255gat, n140gat)
--	n871gat = NOR(n802gat, n375gat)
--	n797gat = NOR(n110gat, n2734gat)
--	n324gat = NOR(n255gat, n146gat, n241gat)
--	n238gat = NOR(n147gat, n254gat)
--	n237gat = NOR(n140gat, n147gat)
--	n1082gat = NOR(n375gat, n380gat)
--	n796gat = NOR(n2731gat, n110gat)
--	n85gat = NOR(n17gat, n294gat, n637gat)
--	n180gat = NOR(n286gat, n188gat, n287gat)
--	n68gat = NOR(n85gat, n180gat)
--	n186gat = NOR(n189gat, n287gat, n288gat)
--	n357gat = NOR(n2726gat, n2860gat)
--	n82gat = NOR(n16gat, n295gat, n637gat)
--	n12gat = NOR(n186gat, n82gat)
--	n1599gat = NOR(n1691gat, n336gat)
--	n1613gat = NOR(n1544gat, n1698gat)
--	n1756gat = NOR(n2512gat, n1769gat, n1773gat)
--	n1586gat = NOR(n1869gat, n1683gat)
--	n1755gat = NOR(n1769gat, n1773gat, n2512gat)
--	n2538gat = NOR(n2620gat, n2625gat, n2488gat)
--	n2483gat = NOR(n2537gat, n2482gat, n2486gat)
--	n1391gat = NOR(n1513gat, n2442gat)
--	n1471gat = NOR(n1334gat, n1858gat, n1604gat)
--	n1469gat = NOR(n1858gat, n1608gat)
--	n1472gat = NOR(n1476gat, n1471gat, n1469gat)
--	n1927gat = NOR(n1790gat, n1635gat)
--	n1470gat = NOR(n1472gat, n1747gat)
--	n1402gat = NOR(n1858gat, n1393gat, n1604gat)
--	n1400gat = NOR(n1674gat, n1403gat)
--	n1567gat = NOR(n1634gat, n1735gat)
--	n1399gat = NOR(n1806gat, n1338gat, n1584gat)
--	n1564gat = NOR(n1584gat, n1719gat, n1790gat, n1576gat)
--	n1600gat = NOR(n1685gat, n1427gat)
--	n1519gat = NOR(n1584gat, n1339gat, n1600gat)
--	n1397gat = NOR(n1519gat, n1401gat)
--	n1398gat = NOR(n1455gat, n1397gat)
--	n2008gat = NOR(n2012gat, n1774gat)
--	n2005gat = NOR(n2002gat, n2857gat)
--	n1818gat = NOR(n1823gat, n2005gat)
--	n1759gat = NOR(n1818gat, n1935gat, n2765gat)
--	n1686gat = NOR(n1774gat, n1869gat, n1684gat)
--	n1533gat = NOR(n1524gat, n1403gat)
--	n1863gat = NOR(n1991gat, n2283gat, n1989gat)
--	n1860gat = NOR(n1988gat, n2216gat, n1862gat)
--	n1915gat = NOR(n1859gat, n1919gat)
--	n1510gat = NOR(n1584gat, n1460gat)
--	n1800gat = NOR(n1635gat, n1919gat)
--	n1459gat = NOR(n1595gat, n1454gat)
--	n1458gat = NOR(n1510gat, n1459gat)
--	n1532gat = NOR(n1677gat, n1458gat)
--	n1467gat = NOR(n2289gat, n1468gat)
--	n1466gat = NOR(n1392gat, n1461gat, n1396gat)
--	n1531gat = NOR(n1507gat, n1477gat)
--	n1593gat = NOR(n1551gat, n1310gat)
--	n1602gat = NOR(n1594gat, n1587gat, n2989gat)
--	n1761gat = NOR(n2985gat, n1602gat, n1681gat)
--	n1760gat = NOR(n1681gat, n1602gat, n2985gat)
--	n1721gat = NOR(n2442gat, n1690gat, n1978gat)
--	n520gat = NOR(n374gat, n2862gat)
--	n519gat = NOR(n2854gat, n374gat)
--	n518gat = NOR(n520gat, n519gat)
--	n418gat = NOR(n374gat, n2723gat)
--	n411gat = NOR(n374gat, n2726gat)
--	n522gat = NOR(n374gat, n2859gat)
--	n516gat = NOR(n374gat, n2715gat)
--	n410gat = NOR(n417gat, n413gat, n412gat, n406gat)
--	n354gat = NOR(n411gat, n522gat)
--	n355gat = NOR(n517gat, n410gat, n354gat)
--	n408gat = NOR(n516gat, n407gat)
--	n526gat = NOR(n2859gat, n740gat)
--	n531gat = NOR(n740gat, n2854gat)
--	n530gat = NOR(n2862gat, n740gat)
--	n525gat = NOR(n526gat, n531gat, n530gat)
--	n356gat = NOR(n2726gat, n740gat)
--	n415gat = NOR(n2723gat, n740gat)
--	n521gat = NOR(n740gat, n2715gat)
--	n532gat = NOR(n527gat, n416gat, n528gat)
--	n359gat = NOR(n290gat, n358gat)
--	n420gat = NOR(n408gat, n359gat)
--	n523gat = NOR(n522gat, n356gat)
--	n634gat = NOR(n418gat, n521gat)
--	n414gat = NOR(n411gat, n415gat)
--	n635gat = NOR(n639gat, n634gat, n414gat)
--	n1100gat = NOR(n1297gat, n1111gat)
--	n630gat = NOR(n634gat, n523gat, n524gat)
--	n994gat = NOR(n1112gat, n882gat)
--	n629gat = NOR(n414gat, n634gat, n523gat)
--	n989gat = NOR(n721gat, n741gat)
--	n632gat = NOR(n414gat, n523gat, n633gat)
--	n880gat = NOR(n926gat, n566gat)
--	n636gat = NOR(n414gat, n633gat, n639gat)
--	n801gat = NOR(n672gat, n670gat)
--	n879gat = NOR(n2931gat, n801gat)
--	n1003gat = NOR(n420gat, n879gat)
--	n1255gat = NOR(n1123gat, n1225gat)
--	n1012gat = NOR(n1007gat, n918gat)
--	n905gat = NOR(n625gat, n1006gat)
--	n1009gat = NOR(n1255gat, n2943gat)
--	n409gat = NOR(n406gat, n407gat)
--	n292gat = NOR(n415gat, n356gat)
--	n291gat = NOR(n290gat, n292gat)
--	n419gat = NOR(n409gat, n291gat)
--	n902gat = NOR(n1009gat, n419gat)
--	n1099gat = NOR(n1111gat, n1293gat)
--	n998gat = NOR(n725gat, n741gat)
--	n995gat = NOR(n823gat, n1112gat)
--	n980gat = NOR(n875gat, n926gat)
--	n1001gat = NOR(n420gat, n1002gat)
--	n1175gat = NOR(n621gat, n1006gat)
--	n1174gat = NOR(n845gat, n1007gat)
--	n1243gat = NOR(n1281gat, n1123gat)
--	n1171gat = NOR(n2960gat, n1243gat)
--	n999gat = NOR(n419gat, n1171gat)
--	n1244gat = NOR(n1123gat, n1134gat)
--	n1323gat = NOR(n1007gat, n401gat)
--	n1264gat = NOR(n1006gat, n617gat)
--	n1265gat = NOR(n1244gat, n2969gat)
--	n892gat = NOR(n419gat, n1265gat)
--	n981gat = NOR(n926gat, n873gat)
--	n890gat = NOR(n741gat, n702gat)
--	n889gat = NOR(n1111gat, n1079gat)
--	n886gat = NOR(n683gat, n1112gat)
--	n891gat = NOR(n420gat, n888gat)
--	n904gat = NOR(n1006gat, n490gat)
--	n903gat = NOR(n1007gat, n397gat)
--	n1254gat = NOR(n1123gat, n1044gat)
--	n1008gat = NOR(n2942gat, n1254gat)
--	n900gat = NOR(n419gat, n1008gat)
--	n1152gat = NOR(n926gat, n1150gat)
--	n1092gat = NOR(n1147gat, n1111gat)
--	n997gat = NOR(n741gat, n393gat)
--	n993gat = NOR(n1112gat, n698gat)
--	n895gat = NOR(n420gat, n898gat)
--	n1094gat = NOR(n1112gat, n583gat)
--	n1093gat = NOR(n1111gat, n864gat)
--	n988gat = NOR(n340gat, n741gat)
--	n984gat = NOR(n926gat, n983gat)
--	n1178gat = NOR(n420gat, n1179gat)
--	n1267gat = NOR(n613gat, n1006gat)
--	n1257gat = NOR(n1007gat, n274gat)
--	n1253gat = NOR(n930gat, n1123gat)
--	n1266gat = NOR(n2965gat, n1253gat)
--	n1116gat = NOR(n419gat, n1266gat)
--	n1375gat = NOR(n1006gat, n706gat)
--	n1324gat = NOR(n164gat, n1007gat)
--	n1200gat = NOR(n1120gat, n1123gat)
--	n1172gat = NOR(n2961gat, n1200gat)
--	n899gat = NOR(n419gat, n1172gat)
--	n1091gat = NOR(n1111gat, n956gat)
--	n1088gat = NOR(n1085gat, n926gat)
--	n992gat = NOR(n815gat, n1112gat)
--	n987gat = NOR(n741gat, n159gat)
--	n896gat = NOR(n897gat, n420gat)
--	n1262gat = NOR(n837gat, n1006gat)
--	n1260gat = NOR(n1007gat, n278gat)
--	n1251gat = NOR(n1123gat, n1071gat)
--	n1259gat = NOR(n2967gat, n1251gat)
--	n901gat = NOR(n419gat, n1259gat)
--	n1098gat = NOR(n336gat, n741gat)
--	n1090gat = NOR(n1111gat, n860gat)
--	n986gat = NOR(n985gat, n926gat)
--	n885gat = NOR(n579gat, n1112gat)
--	n893gat = NOR(n894gat, n420gat)
--	n1097gat = NOR(n270gat, n741gat)
--	n1089gat = NOR(n1067gat, n1111gat)
--	n1087gat = NOR(n926gat, n1084gat)
--	n991gat = NOR(n1112gat, n679gat)
--	n1177gat = NOR(n1180gat, n420gat)
--	n1212gat = NOR(n1123gat, n1034gat)
--	n1326gat = NOR(n1007gat, n282gat)
--	n1261gat = NOR(n833gat, n1006gat)
--	n1263gat = NOR(n1212gat, n2968gat)
--	n1115gat = NOR(n1263gat, n419gat)
--	n977gat = NOR(n670gat, n671gat)
--	n631gat = NOR(n523gat, n633gat, n524gat)
--	n1096gat = NOR(n819gat, n1112gat)
--	n1095gat = NOR(n1240gat, n1111gat)
--	n990gat = NOR(n841gat, n741gat)
--	n979gat = NOR(n1601gat, n926gat)
--	n978gat = NOR(n2944gat, n2945gat)
--	n1004gat = NOR(n978gat, n420gat)
--	n1199gat = NOR(n1123gat, n1284gat)
--	n1176gat = NOR(n829gat, n1006gat)
--	n1173gat = NOR(n1007gat, n1025gat)
--	n1252gat = NOR(n1199gat, n2962gat)
--	n1000gat = NOR(n419gat, n1252gat)
--	n1029gat = NOR(n978gat, n455gat)
--	n1028gat = NOR(n455gat, n879gat)
--	n1031gat = NOR(n1002gat, n455gat)
--	n1030gat = NOR(n455gat, n888gat)
--	n1011gat = NOR(n455gat, n898gat)
--	n1181gat = NOR(n455gat, n1179gat)
--	n1010gat = NOR(n897gat, n455gat)
--	n1005gat = NOR(n894gat, n455gat)
--	n1182gat = NOR(n1180gat, n455gat)
--	n1757gat = NOR(n1773gat, n1769gat)
--	n1745gat = NOR(n1869gat, n1757gat)
--	n73gat = NOR(n67gat, n2784gat)
--	n70gat = NOR(n71gat, n2720gat)
--	n77gat = NOR(n76gat, n2784gat)
--	n13gat = NOR(n2720gat, n14gat)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s5378 is
	port (
		CLK: in std_logic;
		N3065GAT: in std_logic;
		N3066GAT: in std_logic;
		N3067GAT: in std_logic;
		N3068GAT: in std_logic;
		N3069GAT: in std_logic;
		N3070GAT: in std_logic;
		N3071GAT: in std_logic;
		N3072GAT: in std_logic;
		N3073GAT: in std_logic;
		N3074GAT: in std_logic;
		N3075GAT: in std_logic;
		N3076GAT: in std_logic;
		N3077GAT: in std_logic;
		N3078GAT: in std_logic;
		N3079GAT: in std_logic;
		N3080GAT: in std_logic;
		N3081GAT: in std_logic;
		N3082GAT: in std_logic;
		N3083GAT: in std_logic;
		N3084GAT: in std_logic;
		N3085GAT: in std_logic;
		N3086GAT: in std_logic;
		N3087GAT: in std_logic;
		N3088GAT: in std_logic;
		N3089GAT: in std_logic;
		N3090GAT: in std_logic;
		N3091GAT: in std_logic;
		N3092GAT: in std_logic;
		N3093GAT: in std_logic;
		N3094GAT: in std_logic;
		N3095GAT: in std_logic;
		N3097GAT: in std_logic;
		N3098GAT: in std_logic;
		N3099GAT: in std_logic;
		N3100GAT: in std_logic;
		N3104GAT: out std_logic;
		N3105GAT: out std_logic;
		N3106GAT: out std_logic;
		N3107GAT: out std_logic;
		N3108GAT: out std_logic;
		N3109GAT: out std_logic;
		N3110GAT: out std_logic;
		N3111GAT: out std_logic;
		N3112GAT: out std_logic;
		N3113GAT: out std_logic;
		N3114GAT: out std_logic;
		N3115GAT: out std_logic;
		N3116GAT: out std_logic;
		N3117GAT: out std_logic;
		N3118GAT: out std_logic;
		N3119GAT: out std_logic;
		N3120GAT: out std_logic;
		N3121GAT: out std_logic;
		N3122GAT: out std_logic;
		N3123GAT: out std_logic;
		N3124GAT: out std_logic;
		N3125GAT: out std_logic;
		N3126GAT: out std_logic;
		N3127GAT: out std_logic;
		N3128GAT: out std_logic;
		N3129GAT: out std_logic;
		N3130GAT: out std_logic;
		N3131GAT: out std_logic;
		N3132GAT: out std_logic;
		N3133GAT: out std_logic;
		N3134GAT: out std_logic;
		N3135GAT: out std_logic;
		N3136GAT: out std_logic;
		N3137GAT: out std_logic;
		N3138GAT: out std_logic;
		N3139GAT: out std_logic;
		N3140GAT: out std_logic;
		N3141GAT: out std_logic;
		N3142GAT: out std_logic;
		N3143GAT: out std_logic;
		N3144GAT: out std_logic;
		N3145GAT: out std_logic;
		N3146GAT: out std_logic;
		N3147GAT: out std_logic;
		N3148GAT: out std_logic;
		N3149GAT: out std_logic;
		N3150GAT: out std_logic;
		N3151GAT: out std_logic;
		N3152GAT: out std_logic
	);
end entity;

architecture RTL of s5378 is
	attribute dont_touch: boolean;

	signal I1: std_logic; attribute dont_touch of I1: signal is true;
	signal I5: std_logic; attribute dont_touch of I5: signal is true;
	signal I11: std_logic; attribute dont_touch of I11: signal is true;
	signal I14: std_logic; attribute dont_touch of I14: signal is true;
	signal I18: std_logic; attribute dont_touch of I18: signal is true;
	signal I23: std_logic; attribute dont_touch of I23: signal is true;
	signal I27: std_logic; attribute dont_touch of I27: signal is true;
	signal I30: std_logic; attribute dont_touch of I30: signal is true;
	signal I44: std_logic; attribute dont_touch of I44: signal is true;
	signal I47: std_logic; attribute dont_touch of I47: signal is true;
	signal I50: std_logic; attribute dont_touch of I50: signal is true;
	signal I62: std_logic; attribute dont_touch of I62: signal is true;
	signal I65: std_logic; attribute dont_touch of I65: signal is true;
	signal I76: std_logic; attribute dont_touch of I76: signal is true;
	signal I81: std_logic; attribute dont_touch of I81: signal is true;
	signal I92: std_logic; attribute dont_touch of I92: signal is true;
	signal I97: std_logic; attribute dont_touch of I97: signal is true;
	signal I100: std_logic; attribute dont_touch of I100: signal is true;
	signal I111: std_logic; attribute dont_touch of I111: signal is true;
	signal I149: std_logic; attribute dont_touch of I149: signal is true;
	signal I171: std_logic; attribute dont_touch of I171: signal is true;
	signal I178: std_logic; attribute dont_touch of I178: signal is true;
	signal I192: std_logic; attribute dont_touch of I192: signal is true;
	signal I196: std_logic; attribute dont_touch of I196: signal is true;
	signal I199: std_logic; attribute dont_touch of I199: signal is true;
	signal I203: std_logic; attribute dont_touch of I203: signal is true;
	signal I206: std_logic; attribute dont_touch of I206: signal is true;
	signal I210: std_logic; attribute dont_touch of I210: signal is true;
	signal I214: std_logic; attribute dont_touch of I214: signal is true;
	signal I217: std_logic; attribute dont_touch of I217: signal is true;
	signal I220: std_logic; attribute dont_touch of I220: signal is true;
	signal I223: std_logic; attribute dont_touch of I223: signal is true;
	signal I227: std_logic; attribute dont_touch of I227: signal is true;
	signal I230: std_logic; attribute dont_touch of I230: signal is true;
	signal I237: std_logic; attribute dont_touch of I237: signal is true;
	signal I240: std_logic; attribute dont_touch of I240: signal is true;
	signal I243: std_logic; attribute dont_touch of I243: signal is true;
	signal I248: std_logic; attribute dont_touch of I248: signal is true;
	signal I253: std_logic; attribute dont_touch of I253: signal is true;
	signal I256: std_logic; attribute dont_touch of I256: signal is true;
	signal I259: std_logic; attribute dont_touch of I259: signal is true;
	signal I264: std_logic; attribute dont_touch of I264: signal is true;
	signal I270: std_logic; attribute dont_touch of I270: signal is true;
	signal I275: std_logic; attribute dont_touch of I275: signal is true;
	signal I278: std_logic; attribute dont_touch of I278: signal is true;
	signal I282: std_logic; attribute dont_touch of I282: signal is true;
	signal I297: std_logic; attribute dont_touch of I297: signal is true;
	signal I300: std_logic; attribute dont_touch of I300: signal is true;
	signal I311: std_logic; attribute dont_touch of I311: signal is true;
	signal I314: std_logic; attribute dont_touch of I314: signal is true;
	signal I317: std_logic; attribute dont_touch of I317: signal is true;
	signal I320: std_logic; attribute dont_touch of I320: signal is true;
	signal I331: std_logic; attribute dont_touch of I331: signal is true;
	signal I334: std_logic; attribute dont_touch of I334: signal is true;
	signal I337: std_logic; attribute dont_touch of I337: signal is true;
	signal I340: std_logic; attribute dont_touch of I340: signal is true;
	signal I351: std_logic; attribute dont_touch of I351: signal is true;
	signal I354: std_logic; attribute dont_touch of I354: signal is true;
	signal I359: std_logic; attribute dont_touch of I359: signal is true;
	signal I363: std_logic; attribute dont_touch of I363: signal is true;
	signal I368: std_logic; attribute dont_touch of I368: signal is true;
	signal I375: std_logic; attribute dont_touch of I375: signal is true;
	signal I378: std_logic; attribute dont_touch of I378: signal is true;
	signal I381: std_logic; attribute dont_touch of I381: signal is true;
	signal I384: std_logic; attribute dont_touch of I384: signal is true;
	signal I395: std_logic; attribute dont_touch of I395: signal is true;
	signal I398: std_logic; attribute dont_touch of I398: signal is true;
	signal I401: std_logic; attribute dont_touch of I401: signal is true;
	signal I406: std_logic; attribute dont_touch of I406: signal is true;
	signal I409: std_logic; attribute dont_touch of I409: signal is true;
	signal I414: std_logic; attribute dont_touch of I414: signal is true;
	signal I420: std_logic; attribute dont_touch of I420: signal is true;
	signal I423: std_logic; attribute dont_touch of I423: signal is true;
	signal I426: std_logic; attribute dont_touch of I426: signal is true;
	signal I437: std_logic; attribute dont_touch of I437: signal is true;
	signal I440: std_logic; attribute dont_touch of I440: signal is true;
	signal I443: std_logic; attribute dont_touch of I443: signal is true;
	signal I446: std_logic; attribute dont_touch of I446: signal is true;
	signal I449: std_logic; attribute dont_touch of I449: signal is true;
	signal I453: std_logic; attribute dont_touch of I453: signal is true;
	signal I456: std_logic; attribute dont_touch of I456: signal is true;
	signal I461: std_logic; attribute dont_touch of I461: signal is true;
	signal I468: std_logic; attribute dont_touch of I468: signal is true;
	signal I473: std_logic; attribute dont_touch of I473: signal is true;
	signal I476: std_logic; attribute dont_touch of I476: signal is true;
	signal I480: std_logic; attribute dont_touch of I480: signal is true;
	signal I509: std_logic; attribute dont_touch of I509: signal is true;
	signal I512: std_logic; attribute dont_touch of I512: signal is true;
	signal I572: std_logic; attribute dont_touch of I572: signal is true;
	signal I576: std_logic; attribute dont_touch of I576: signal is true;
	signal I579: std_logic; attribute dont_touch of I579: signal is true;
	signal I583: std_logic; attribute dont_touch of I583: signal is true;
	signal I591: std_logic; attribute dont_touch of I591: signal is true;
	signal I594: std_logic; attribute dont_touch of I594: signal is true;
	signal I606: std_logic; attribute dont_touch of I606: signal is true;
	signal I609: std_logic; attribute dont_touch of I609: signal is true;
	signal I620: std_logic; attribute dont_touch of I620: signal is true;
	signal I623: std_logic; attribute dont_touch of I623: signal is true;
	signal I634: std_logic; attribute dont_touch of I634: signal is true;
	signal I637: std_logic; attribute dont_touch of I637: signal is true;
	signal I642: std_logic; attribute dont_touch of I642: signal is true;
	signal I646: std_logic; attribute dont_touch of I646: signal is true;
	signal I651: std_logic; attribute dont_touch of I651: signal is true;
	signal I658: std_logic; attribute dont_touch of I658: signal is true;
	signal I661: std_logic; attribute dont_touch of I661: signal is true;
	signal I672: std_logic; attribute dont_touch of I672: signal is true;
	signal I675: std_logic; attribute dont_touch of I675: signal is true;
	signal I678: std_logic; attribute dont_touch of I678: signal is true;
	signal I683: std_logic; attribute dont_touch of I683: signal is true;
	signal I687: std_logic; attribute dont_touch of I687: signal is true;
	signal I692: std_logic; attribute dont_touch of I692: signal is true;
	signal I698: std_logic; attribute dont_touch of I698: signal is true;
	signal I709: std_logic; attribute dont_touch of I709: signal is true;
	signal I712: std_logic; attribute dont_touch of I712: signal is true;
	signal I715: std_logic; attribute dont_touch of I715: signal is true;
	signal I718: std_logic; attribute dont_touch of I718: signal is true;
	signal I721: std_logic; attribute dont_touch of I721: signal is true;
	signal I726: std_logic; attribute dont_touch of I726: signal is true;
	signal I729: std_logic; attribute dont_touch of I729: signal is true;
	signal I734: std_logic; attribute dont_touch of I734: signal is true;
	signal I741: std_logic; attribute dont_touch of I741: signal is true;
	signal I746: std_logic; attribute dont_touch of I746: signal is true;
	signal I749: std_logic; attribute dont_touch of I749: signal is true;
	signal I753: std_logic; attribute dont_touch of I753: signal is true;
	signal I768: std_logic; attribute dont_touch of I768: signal is true;
	signal I771: std_logic; attribute dont_touch of I771: signal is true;
	signal I776: std_logic; attribute dont_touch of I776: signal is true;
	signal I790: std_logic; attribute dont_touch of I790: signal is true;
	signal I793: std_logic; attribute dont_touch of I793: signal is true;
	signal I796: std_logic; attribute dont_touch of I796: signal is true;
	signal I812: std_logic; attribute dont_touch of I812: signal is true;
	signal I815: std_logic; attribute dont_touch of I815: signal is true;
	signal I818: std_logic; attribute dont_touch of I818: signal is true;
	signal I834: std_logic; attribute dont_touch of I834: signal is true;
	signal I837: std_logic; attribute dont_touch of I837: signal is true;
	signal I842: std_logic; attribute dont_touch of I842: signal is true;
	signal I846: std_logic; attribute dont_touch of I846: signal is true;
	signal I851: std_logic; attribute dont_touch of I851: signal is true;
	signal I858: std_logic; attribute dont_touch of I858: signal is true;
	signal I863: std_logic; attribute dont_touch of I863: signal is true;
	signal I877: std_logic; attribute dont_touch of I877: signal is true;
	signal I880: std_logic; attribute dont_touch of I880: signal is true;
	signal I885: std_logic; attribute dont_touch of I885: signal is true;
	signal I899: std_logic; attribute dont_touch of I899: signal is true;
	signal I902: std_logic; attribute dont_touch of I902: signal is true;
	signal I913: std_logic; attribute dont_touch of I913: signal is true;
	signal I916: std_logic; attribute dont_touch of I916: signal is true;
	signal I921: std_logic; attribute dont_touch of I921: signal is true;
	signal I925: std_logic; attribute dont_touch of I925: signal is true;
	signal I930: std_logic; attribute dont_touch of I930: signal is true;
	signal I936: std_logic; attribute dont_touch of I936: signal is true;
	signal I941: std_logic; attribute dont_touch of I941: signal is true;
	signal I955: std_logic; attribute dont_touch of I955: signal is true;
	signal I958: std_logic; attribute dont_touch of I958: signal is true;
	signal I963: std_logic; attribute dont_touch of I963: signal is true;
	signal I977: std_logic; attribute dont_touch of I977: signal is true;
	signal I980: std_logic; attribute dont_touch of I980: signal is true;
	signal I985: std_logic; attribute dont_touch of I985: signal is true;
	signal I999: std_logic; attribute dont_touch of I999: signal is true;
	signal I1002: std_logic; attribute dont_touch of I1002: signal is true;
	signal I1007: std_logic; attribute dont_touch of I1007: signal is true;
	signal I1011: std_logic; attribute dont_touch of I1011: signal is true;
	signal I1016: std_logic; attribute dont_touch of I1016: signal is true;
	signal I1023: std_logic; attribute dont_touch of I1023: signal is true;
	signal I1028: std_logic; attribute dont_touch of I1028: signal is true;
	signal I1031: std_logic; attribute dont_touch of I1031: signal is true;
	signal I1035: std_logic; attribute dont_touch of I1035: signal is true;
	signal I1067: std_logic; attribute dont_touch of I1067: signal is true;
	signal I1079: std_logic; attribute dont_touch of I1079: signal is true;
	signal I1082: std_logic; attribute dont_touch of I1082: signal is true;
	signal I1085: std_logic; attribute dont_touch of I1085: signal is true;
	signal I1088: std_logic; attribute dont_touch of I1088: signal is true;
	signal I1091: std_logic; attribute dont_touch of I1091: signal is true;
	signal I1103: std_logic; attribute dont_touch of I1103: signal is true;
	signal I1115: std_logic; attribute dont_touch of I1115: signal is true;
	signal I1118: std_logic; attribute dont_touch of I1118: signal is true;
	signal I1121: std_logic; attribute dont_touch of I1121: signal is true;
	signal I1124: std_logic; attribute dont_touch of I1124: signal is true;
	signal I1127: std_logic; attribute dont_touch of I1127: signal is true;
	signal I1138: std_logic; attribute dont_touch of I1138: signal is true;
	signal I1141: std_logic; attribute dont_touch of I1141: signal is true;
	signal I1152: std_logic; attribute dont_touch of I1152: signal is true;
	signal I1155: std_logic; attribute dont_touch of I1155: signal is true;
	signal I1166: std_logic; attribute dont_touch of I1166: signal is true;
	signal I1169: std_logic; attribute dont_touch of I1169: signal is true;
	signal I1174: std_logic; attribute dont_touch of I1174: signal is true;
	signal I1178: std_logic; attribute dont_touch of I1178: signal is true;
	signal I1183: std_logic; attribute dont_touch of I1183: signal is true;
	signal I1190: std_logic; attribute dont_touch of I1190: signal is true;
	signal I1201: std_logic; attribute dont_touch of I1201: signal is true;
	signal I1204: std_logic; attribute dont_touch of I1204: signal is true;
	signal I1209: std_logic; attribute dont_touch of I1209: signal is true;
	signal I1216: std_logic; attribute dont_touch of I1216: signal is true;
	signal I1227: std_logic; attribute dont_touch of I1227: signal is true;
	signal I1230: std_logic; attribute dont_touch of I1230: signal is true;
	signal I1236: std_logic; attribute dont_touch of I1236: signal is true;
	signal I1243: std_logic; attribute dont_touch of I1243: signal is true;
	signal I1248: std_logic; attribute dont_touch of I1248: signal is true;
	signal I1251: std_logic; attribute dont_touch of I1251: signal is true;
	signal I1255: std_logic; attribute dont_touch of I1255: signal is true;
	signal I1277: std_logic; attribute dont_touch of I1277: signal is true;
	signal I1278: std_logic; attribute dont_touch of I1278: signal is true;
	signal I1302: std_logic; attribute dont_touch of I1302: signal is true;
	signal I1305: std_logic; attribute dont_touch of I1305: signal is true;
	signal I1319: std_logic; attribute dont_touch of I1319: signal is true;
	signal I1322: std_logic; attribute dont_touch of I1322: signal is true;
	signal I1336: std_logic; attribute dont_touch of I1336: signal is true;
	signal I1339: std_logic; attribute dont_touch of I1339: signal is true;
	signal I1344: std_logic; attribute dont_touch of I1344: signal is true;
	signal I1348: std_logic; attribute dont_touch of I1348: signal is true;
	signal I1353: std_logic; attribute dont_touch of I1353: signal is true;
	signal I1360: std_logic; attribute dont_touch of I1360: signal is true;
	signal I1371: std_logic; attribute dont_touch of I1371: signal is true;
	signal I1374: std_logic; attribute dont_touch of I1374: signal is true;
	signal I1385: std_logic; attribute dont_touch of I1385: signal is true;
	signal I1388: std_logic; attribute dont_touch of I1388: signal is true;
	signal I1399: std_logic; attribute dont_touch of I1399: signal is true;
	signal I1402: std_logic; attribute dont_touch of I1402: signal is true;
	signal I1407: std_logic; attribute dont_touch of I1407: signal is true;
	signal I1411: std_logic; attribute dont_touch of I1411: signal is true;
	signal I1416: std_logic; attribute dont_touch of I1416: signal is true;
	signal I1422: std_logic; attribute dont_touch of I1422: signal is true;
	signal I1436: std_logic; attribute dont_touch of I1436: signal is true;
	signal I1439: std_logic; attribute dont_touch of I1439: signal is true;
	signal I1450: std_logic; attribute dont_touch of I1450: signal is true;
	signal I1453: std_logic; attribute dont_touch of I1453: signal is true;
	signal I1464: std_logic; attribute dont_touch of I1464: signal is true;
	signal I1467: std_logic; attribute dont_touch of I1467: signal is true;
	signal I1472: std_logic; attribute dont_touch of I1472: signal is true;
	signal I1476: std_logic; attribute dont_touch of I1476: signal is true;
	signal I1481: std_logic; attribute dont_touch of I1481: signal is true;
	signal I1488: std_logic; attribute dont_touch of I1488: signal is true;
	signal I1493: std_logic; attribute dont_touch of I1493: signal is true;
	signal I1496: std_logic; attribute dont_touch of I1496: signal is true;
	signal I1500: std_logic; attribute dont_touch of I1500: signal is true;
	signal I1515: std_logic; attribute dont_touch of I1515: signal is true;
	signal I1516: std_logic; attribute dont_touch of I1516: signal is true;
	signal I1538: std_logic; attribute dont_touch of I1538: signal is true;
	signal I1550: std_logic; attribute dont_touch of I1550: signal is true;
	signal I1584: std_logic; attribute dont_touch of I1584: signal is true;
	signal I1585: std_logic; attribute dont_touch of I1585: signal is true;
	signal I1606: std_logic; attribute dont_touch of I1606: signal is true;
	signal I1617: std_logic; attribute dont_touch of I1617: signal is true;
	signal I1630: std_logic; attribute dont_touch of I1630: signal is true;
	signal I1655: std_logic; attribute dont_touch of I1655: signal is true;
	signal I1667: std_logic; attribute dont_touch of I1667: signal is true;
	signal I1683: std_logic; attribute dont_touch of I1683: signal is true;
	signal I1698: std_logic; attribute dont_touch of I1698: signal is true;
	signal I1703: std_logic; attribute dont_touch of I1703: signal is true;
	signal I1708: std_logic; attribute dont_touch of I1708: signal is true;
	signal I1719: std_logic; attribute dont_touch of I1719: signal is true;
	signal I1723: std_logic; attribute dont_touch of I1723: signal is true;
	signal I1724: std_logic; attribute dont_touch of I1724: signal is true;
	signal I1733: std_logic; attribute dont_touch of I1733: signal is true;
	signal I1734: std_logic; attribute dont_touch of I1734: signal is true;
	signal I1749: std_logic; attribute dont_touch of I1749: signal is true;
	signal I1752: std_logic; attribute dont_touch of I1752: signal is true;
	signal I1766: std_logic; attribute dont_touch of I1766: signal is true;
	signal I1769: std_logic; attribute dont_touch of I1769: signal is true;
	signal I1783: std_logic; attribute dont_touch of I1783: signal is true;
	signal I1786: std_logic; attribute dont_touch of I1786: signal is true;
	signal I1791: std_logic; attribute dont_touch of I1791: signal is true;
	signal I1795: std_logic; attribute dont_touch of I1795: signal is true;
	signal I1800: std_logic; attribute dont_touch of I1800: signal is true;
	signal I1807: std_logic; attribute dont_touch of I1807: signal is true;
	signal I1833: std_logic; attribute dont_touch of I1833: signal is true;
	signal I1837: std_logic; attribute dont_touch of I1837: signal is true;
	signal I1843: std_logic; attribute dont_touch of I1843: signal is true;
	signal I1857: std_logic; attribute dont_touch of I1857: signal is true;
	signal I1860: std_logic; attribute dont_touch of I1860: signal is true;
	signal I1874: std_logic; attribute dont_touch of I1874: signal is true;
	signal I1877: std_logic; attribute dont_touch of I1877: signal is true;
	signal I1891: std_logic; attribute dont_touch of I1891: signal is true;
	signal I1894: std_logic; attribute dont_touch of I1894: signal is true;
	signal I1899: std_logic; attribute dont_touch of I1899: signal is true;
	signal I1903: std_logic; attribute dont_touch of I1903: signal is true;
	signal I1908: std_logic; attribute dont_touch of I1908: signal is true;
	signal I1915: std_logic; attribute dont_touch of I1915: signal is true;
	signal I1920: std_logic; attribute dont_touch of I1920: signal is true;
	signal I1923: std_logic; attribute dont_touch of I1923: signal is true;
	signal I1927: std_logic; attribute dont_touch of I1927: signal is true;
	signal I1947: std_logic; attribute dont_touch of I1947: signal is true;
	signal I1961: std_logic; attribute dont_touch of I1961: signal is true;
	signal I1981: std_logic; attribute dont_touch of I1981: signal is true;
	signal I1996: std_logic; attribute dont_touch of I1996: signal is true;
	signal I1999: std_logic; attribute dont_touch of I1999: signal is true;
	signal I2014: std_logic; attribute dont_touch of I2014: signal is true;
	signal I2017: std_logic; attribute dont_touch of I2017: signal is true;
	signal I2032: std_logic; attribute dont_touch of I2032: signal is true;
	signal I2035: std_logic; attribute dont_touch of I2035: signal is true;
	signal I2040: std_logic; attribute dont_touch of I2040: signal is true;
	signal I2044: std_logic; attribute dont_touch of I2044: signal is true;
	signal I2049: std_logic; attribute dont_touch of I2049: signal is true;
	signal I2056: std_logic; attribute dont_touch of I2056: signal is true;
	signal I2084: std_logic; attribute dont_touch of I2084: signal is true;
	signal I2088: std_logic; attribute dont_touch of I2088: signal is true;
	signal I2094: std_logic; attribute dont_touch of I2094: signal is true;
	signal I2109: std_logic; attribute dont_touch of I2109: signal is true;
	signal I2112: std_logic; attribute dont_touch of I2112: signal is true;
	signal I2127: std_logic; attribute dont_touch of I2127: signal is true;
	signal I2130: std_logic; attribute dont_touch of I2130: signal is true;
	signal I2145: std_logic; attribute dont_touch of I2145: signal is true;
	signal I2148: std_logic; attribute dont_touch of I2148: signal is true;
	signal I2153: std_logic; attribute dont_touch of I2153: signal is true;
	signal I2157: std_logic; attribute dont_touch of I2157: signal is true;
	signal I2162: std_logic; attribute dont_touch of I2162: signal is true;
	signal I2169: std_logic; attribute dont_touch of I2169: signal is true;
	signal I2174: std_logic; attribute dont_touch of I2174: signal is true;
	signal I2177: std_logic; attribute dont_touch of I2177: signal is true;
	signal I2181: std_logic; attribute dont_touch of I2181: signal is true;
	signal I2213: std_logic; attribute dont_touch of I2213: signal is true;
	signal I2225: std_logic; attribute dont_touch of I2225: signal is true;
	signal I2228: std_logic; attribute dont_touch of I2228: signal is true;
	signal I2232: std_logic; attribute dont_touch of I2232: signal is true;
	signal I2235: std_logic; attribute dont_touch of I2235: signal is true;
	signal I2238: std_logic; attribute dont_touch of I2238: signal is true;
	signal I2242: std_logic; attribute dont_touch of I2242: signal is true;
	signal I2248: std_logic; attribute dont_touch of I2248: signal is true;
	signal I2251: std_logic; attribute dont_touch of I2251: signal is true;
	signal I2254: std_logic; attribute dont_touch of I2254: signal is true;
	signal I2257: std_logic; attribute dont_touch of I2257: signal is true;
	signal I2260: std_logic; attribute dont_touch of I2260: signal is true;
	signal I2263: std_logic; attribute dont_touch of I2263: signal is true;
	signal I2268: std_logic; attribute dont_touch of I2268: signal is true;
	signal I2271: std_logic; attribute dont_touch of I2271: signal is true;
	signal I2275: std_logic; attribute dont_touch of I2275: signal is true;
	signal I2281: std_logic; attribute dont_touch of I2281: signal is true;
	signal I2316: std_logic; attribute dont_touch of I2316: signal is true;
	signal I2319: std_logic; attribute dont_touch of I2319: signal is true;
	signal I2324: std_logic; attribute dont_touch of I2324: signal is true;
	signal I2344: std_logic; attribute dont_touch of I2344: signal is true;
	signal I2349: std_logic; attribute dont_touch of I2349: signal is true;
	signal I2354: std_logic; attribute dont_touch of I2354: signal is true;
	signal I2372: std_logic; attribute dont_touch of I2372: signal is true;
	signal I2376: std_logic; attribute dont_touch of I2376: signal is true;
	signal I2380: std_logic; attribute dont_touch of I2380: signal is true;
	signal I2385: std_logic; attribute dont_touch of I2385: signal is true;
	signal I2389: std_logic; attribute dont_touch of I2389: signal is true;
	signal I2394: std_logic; attribute dont_touch of I2394: signal is true;
	signal I2400: std_logic; attribute dont_touch of I2400: signal is true;
	signal I2403: std_logic; attribute dont_touch of I2403: signal is true;
	signal I2414: std_logic; attribute dont_touch of I2414: signal is true;
	signal I2417: std_logic; attribute dont_touch of I2417: signal is true;
	signal I2420: std_logic; attribute dont_touch of I2420: signal is true;
	signal I2425: std_logic; attribute dont_touch of I2425: signal is true;
	signal I2428: std_logic; attribute dont_touch of I2428: signal is true;
	signal I2433: std_logic; attribute dont_touch of I2433: signal is true;
	signal I2439: std_logic; attribute dont_touch of I2439: signal is true;
	signal I2672: std_logic; attribute dont_touch of I2672: signal is true;
	signal I2684: std_logic; attribute dont_touch of I2684: signal is true;
	signal I2696: std_logic; attribute dont_touch of I2696: signal is true;
	signal I2720: std_logic; attribute dont_touch of I2720: signal is true;
	signal I2721: std_logic; attribute dont_touch of I2721: signal is true;
	signal I2731: std_logic; attribute dont_touch of I2731: signal is true;
	signal I2735: std_logic; attribute dont_touch of I2735: signal is true;
	signal I2736: std_logic; attribute dont_touch of I2736: signal is true;
	signal I2771: std_logic; attribute dont_touch of I2771: signal is true;
	signal I2785: std_logic; attribute dont_touch of I2785: signal is true;
	signal I2812: std_logic; attribute dont_touch of I2812: signal is true;
	signal I2813: std_logic; attribute dont_touch of I2813: signal is true;
	signal I2831: std_logic; attribute dont_touch of I2831: signal is true;
	signal I2832: std_logic; attribute dont_touch of I2832: signal is true;
	signal I2837: std_logic; attribute dont_touch of I2837: signal is true;
	signal I2843: std_logic; attribute dont_touch of I2843: signal is true;
	signal I2847: std_logic; attribute dont_touch of I2847: signal is true;
	signal I2873: std_logic; attribute dont_touch of I2873: signal is true;
	signal I2885: std_logic; attribute dont_touch of I2885: signal is true;
	signal I2889: std_logic; attribute dont_touch of I2889: signal is true;
	signal I2890: std_logic; attribute dont_touch of I2890: signal is true;
	signal I2915: std_logic; attribute dont_touch of I2915: signal is true;
	signal I2925: std_logic; attribute dont_touch of I2925: signal is true;
	signal I2926: std_logic; attribute dont_touch of I2926: signal is true;
	signal I2934: std_logic; attribute dont_touch of I2934: signal is true;
	signal I2935: std_logic; attribute dont_touch of I2935: signal is true;
	signal I2953: std_logic; attribute dont_touch of I2953: signal is true;
	signal I2978: std_logic; attribute dont_touch of I2978: signal is true;
	signal I2989: std_logic; attribute dont_touch of I2989: signal is true;
	signal I3000: std_logic; attribute dont_touch of I3000: signal is true;
	signal I3016: std_logic; attribute dont_touch of I3016: signal is true;
	signal I3056: std_logic; attribute dont_touch of I3056: signal is true;
	signal I3143: std_logic; attribute dont_touch of I3143: signal is true;
	signal I3148: std_logic; attribute dont_touch of I3148: signal is true;
	signal I3149: std_logic; attribute dont_touch of I3149: signal is true;
	signal I3163: std_logic; attribute dont_touch of I3163: signal is true;
	signal I3168: std_logic; attribute dont_touch of I3168: signal is true;
	signal I3174: std_logic; attribute dont_touch of I3174: signal is true;
	signal I3178: std_logic; attribute dont_touch of I3178: signal is true;
	signal I3179: std_logic; attribute dont_touch of I3179: signal is true;
	signal I3191: std_logic; attribute dont_touch of I3191: signal is true;
	signal I3211: std_logic; attribute dont_touch of I3211: signal is true;
	signal I3235: std_logic; attribute dont_touch of I3235: signal is true;
	signal I3273: std_logic; attribute dont_touch of I3273: signal is true;
	signal I3287: std_logic; attribute dont_touch of I3287: signal is true;
	signal I3290: std_logic; attribute dont_touch of I3290: signal is true;
	signal I3293: std_logic; attribute dont_touch of I3293: signal is true;
	signal I3297: std_logic; attribute dont_touch of I3297: signal is true;
	signal I3300: std_logic; attribute dont_touch of I3300: signal is true;
	signal I3303: std_logic; attribute dont_touch of I3303: signal is true;
	signal I3306: std_logic; attribute dont_touch of I3306: signal is true;
	signal I3309: std_logic; attribute dont_touch of I3309: signal is true;
	signal I3312: std_logic; attribute dont_touch of I3312: signal is true;
	signal I3315: std_logic; attribute dont_touch of I3315: signal is true;
	signal I3318: std_logic; attribute dont_touch of I3318: signal is true;
	signal I3336: std_logic; attribute dont_touch of I3336: signal is true;
	signal I3339: std_logic; attribute dont_touch of I3339: signal is true;
	signal I3342: std_logic; attribute dont_touch of I3342: signal is true;
	signal I3387: std_logic; attribute dont_touch of I3387: signal is true;
	signal I3390: std_logic; attribute dont_touch of I3390: signal is true;
	signal I3394: std_logic; attribute dont_touch of I3394: signal is true;
	signal I3401: std_logic; attribute dont_touch of I3401: signal is true;
	signal I3412: std_logic; attribute dont_touch of I3412: signal is true;
	signal I3429: std_logic; attribute dont_touch of I3429: signal is true;
	signal I3436: std_logic; attribute dont_touch of I3436: signal is true;
	signal I3457: std_logic; attribute dont_touch of I3457: signal is true;
	signal I3461: std_logic; attribute dont_touch of I3461: signal is true;
	signal I3465: std_logic; attribute dont_touch of I3465: signal is true;
	signal I3472: std_logic; attribute dont_touch of I3472: signal is true;
	signal I3483: std_logic; attribute dont_touch of I3483: signal is true;
	signal I3491: std_logic; attribute dont_touch of I3491: signal is true;
	signal I3494: std_logic; attribute dont_touch of I3494: signal is true;
	signal I3504: std_logic; attribute dont_touch of I3504: signal is true;
	signal I3509: std_logic; attribute dont_touch of I3509: signal is true;
	signal I3513: std_logic; attribute dont_touch of I3513: signal is true;
	signal I3520: std_logic; attribute dont_touch of I3520: signal is true;
	signal I3530: std_logic; attribute dont_touch of I3530: signal is true;
	signal I3539: std_logic; attribute dont_touch of I3539: signal is true;
	signal I3549: std_logic; attribute dont_touch of I3549: signal is true;
	signal I3558: std_logic; attribute dont_touch of I3558: signal is true;
	signal I3587: std_logic; attribute dont_touch of I3587: signal is true;
	signal I3610: std_logic; attribute dont_touch of I3610: signal is true;
	signal I3621: std_logic; attribute dont_touch of I3621: signal is true;
	signal I3635: std_logic; attribute dont_touch of I3635: signal is true;
	signal I3646: std_logic; attribute dont_touch of I3646: signal is true;
	signal I3660: std_logic; attribute dont_touch of I3660: signal is true;
	signal I3677: std_logic; attribute dont_touch of I3677: signal is true;
	signal I3691: std_logic; attribute dont_touch of I3691: signal is true;
	signal I3703: std_logic; attribute dont_touch of I3703: signal is true;
	signal I3713: std_logic; attribute dont_touch of I3713: signal is true;
	signal I3736: std_logic; attribute dont_touch of I3736: signal is true;
	signal I3742: std_logic; attribute dont_touch of I3742: signal is true;
	signal I3754: std_logic; attribute dont_touch of I3754: signal is true;
	signal I3765: std_logic; attribute dont_touch of I3765: signal is true;
	signal I3777: std_logic; attribute dont_touch of I3777: signal is true;
	signal I3801: std_logic; attribute dont_touch of I3801: signal is true;
	signal I3808: std_logic; attribute dont_touch of I3808: signal is true;
	signal I3817: std_logic; attribute dont_touch of I3817: signal is true;
	signal I3831: std_logic; attribute dont_touch of I3831: signal is true;
	signal I3841: std_logic; attribute dont_touch of I3841: signal is true;
	signal I3867: std_logic; attribute dont_touch of I3867: signal is true;
	signal I3876: std_logic; attribute dont_touch of I3876: signal is true;
	signal I3882: std_logic; attribute dont_touch of I3882: signal is true;
	signal I3891: std_logic; attribute dont_touch of I3891: signal is true;
	signal I3904: std_logic; attribute dont_touch of I3904: signal is true;
	signal I3914: std_logic; attribute dont_touch of I3914: signal is true;
	signal I3923: std_logic; attribute dont_touch of I3923: signal is true;
	signal I3935: std_logic; attribute dont_touch of I3935: signal is true;
	signal I3941: std_logic; attribute dont_touch of I3941: signal is true;
	signal I3945: std_logic; attribute dont_touch of I3945: signal is true;
	signal I3948: std_logic; attribute dont_touch of I3948: signal is true;
	signal I3951: std_logic; attribute dont_touch of I3951: signal is true;
	signal I3954: std_logic; attribute dont_touch of I3954: signal is true;
	signal I3957: std_logic; attribute dont_touch of I3957: signal is true;
	signal I3962: std_logic; attribute dont_touch of I3962: signal is true;
	signal I3999: std_logic; attribute dont_touch of I3999: signal is true;
	signal I4000: std_logic; attribute dont_touch of I4000: signal is true;
	signal I4014: std_logic; attribute dont_touch of I4014: signal is true;
	signal I4020: std_logic; attribute dont_touch of I4020: signal is true;
	signal I4023: std_logic; attribute dont_touch of I4023: signal is true;
	signal I4024: std_logic; attribute dont_touch of I4024: signal is true;
	signal I4055: std_logic; attribute dont_touch of I4055: signal is true;
	signal I4067: std_logic; attribute dont_touch of I4067: signal is true;
	signal I4081: std_logic; attribute dont_touch of I4081: signal is true;
	signal I4105: std_logic; attribute dont_touch of I4105: signal is true;
	signal I4108: std_logic; attribute dont_touch of I4108: signal is true;
	signal I4117: std_logic; attribute dont_touch of I4117: signal is true;
	signal I4122: std_logic; attribute dont_touch of I4122: signal is true;
	signal I4129: std_logic; attribute dont_touch of I4129: signal is true;
	signal I4135: std_logic; attribute dont_touch of I4135: signal is true;
	signal I4138: std_logic; attribute dont_touch of I4138: signal is true;
	signal I4144: std_logic; attribute dont_touch of I4144: signal is true;
	signal I4145: std_logic; attribute dont_touch of I4145: signal is true;
	signal I4157: std_logic; attribute dont_touch of I4157: signal is true;
	signal I4185: std_logic; attribute dont_touch of I4185: signal is true;
	signal I4194: std_logic; attribute dont_touch of I4194: signal is true;
	signal I4212: std_logic; attribute dont_touch of I4212: signal is true;
	signal I4216: std_logic; attribute dont_touch of I4216: signal is true;
	signal I4217: std_logic; attribute dont_touch of I4217: signal is true;
	signal I4222: std_logic; attribute dont_touch of I4222: signal is true;
	signal I4227: std_logic; attribute dont_touch of I4227: signal is true;
	signal I4233: std_logic; attribute dont_touch of I4233: signal is true;
	signal I4236: std_logic; attribute dont_touch of I4236: signal is true;
	signal I4309: std_logic; attribute dont_touch of I4309: signal is true;
	signal I4312: std_logic; attribute dont_touch of I4312: signal is true;
	signal I4329: std_logic; attribute dont_touch of I4329: signal is true;
	signal I4332: std_logic; attribute dont_touch of I4332: signal is true;
	signal I4349: std_logic; attribute dont_touch of I4349: signal is true;
	signal I4352: std_logic; attribute dont_touch of I4352: signal is true;
	signal I4369: std_logic; attribute dont_touch of I4369: signal is true;
	signal I4372: std_logic; attribute dont_touch of I4372: signal is true;
	signal I4389: std_logic; attribute dont_touch of I4389: signal is true;
	signal I4392: std_logic; attribute dont_touch of I4392: signal is true;
	signal I4409: std_logic; attribute dont_touch of I4409: signal is true;
	signal I4412: std_logic; attribute dont_touch of I4412: signal is true;
	signal I4429: std_logic; attribute dont_touch of I4429: signal is true;
	signal I4432: std_logic; attribute dont_touch of I4432: signal is true;
	signal I4449: std_logic; attribute dont_touch of I4449: signal is true;
	signal I4452: std_logic; attribute dont_touch of I4452: signal is true;
	signal I4475: std_logic; attribute dont_touch of I4475: signal is true;
	signal I4478: std_logic; attribute dont_touch of I4478: signal is true;
	signal I4482: std_logic; attribute dont_touch of I4482: signal is true;
	signal I4485: std_logic; attribute dont_touch of I4485: signal is true;
	signal I4489: std_logic; attribute dont_touch of I4489: signal is true;
	signal I4492: std_logic; attribute dont_touch of I4492: signal is true;
	signal I4496: std_logic; attribute dont_touch of I4496: signal is true;
	signal I4499: std_logic; attribute dont_touch of I4499: signal is true;
	signal I4506: std_logic; attribute dont_touch of I4506: signal is true;
	signal I4512: std_logic; attribute dont_touch of I4512: signal is true;
	signal I4518: std_logic; attribute dont_touch of I4518: signal is true;
	signal I4524: std_logic; attribute dont_touch of I4524: signal is true;
	signal I4530: std_logic; attribute dont_touch of I4530: signal is true;
	signal I4536: std_logic; attribute dont_touch of I4536: signal is true;
	signal I4542: std_logic; attribute dont_touch of I4542: signal is true;
	signal I4548: std_logic; attribute dont_touch of I4548: signal is true;
	signal I4554: std_logic; attribute dont_touch of I4554: signal is true;
	signal I4558: std_logic; attribute dont_touch of I4558: signal is true;
	signal I4566: std_logic; attribute dont_touch of I4566: signal is true;
	signal I4573: std_logic; attribute dont_touch of I4573: signal is true;
	signal I4580: std_logic; attribute dont_touch of I4580: signal is true;
	signal I4587: std_logic; attribute dont_touch of I4587: signal is true;
	signal I4594: std_logic; attribute dont_touch of I4594: signal is true;
	signal I4601: std_logic; attribute dont_touch of I4601: signal is true;
	signal I4608: std_logic; attribute dont_touch of I4608: signal is true;
	signal I4615: std_logic; attribute dont_touch of I4615: signal is true;
	signal I4620: std_logic; attribute dont_touch of I4620: signal is true;
	signal I4623: std_logic; attribute dont_touch of I4623: signal is true;
	signal I4626: std_logic; attribute dont_touch of I4626: signal is true;
	signal I4630: std_logic; attribute dont_touch of I4630: signal is true;
	signal I4633: std_logic; attribute dont_touch of I4633: signal is true;
	signal I4642: std_logic; attribute dont_touch of I4642: signal is true;
	signal I4651: std_logic; attribute dont_touch of I4651: signal is true;
	signal I4654: std_logic; attribute dont_touch of I4654: signal is true;
	signal I4657: std_logic; attribute dont_touch of I4657: signal is true;
	signal I4660: std_logic; attribute dont_touch of I4660: signal is true;
	signal I4663: std_logic; attribute dont_touch of I4663: signal is true;
	signal I4666: std_logic; attribute dont_touch of I4666: signal is true;
	signal I4669: std_logic; attribute dont_touch of I4669: signal is true;
	signal I4672: std_logic; attribute dont_touch of I4672: signal is true;
	signal I4675: std_logic; attribute dont_touch of I4675: signal is true;
	signal I4678: std_logic; attribute dont_touch of I4678: signal is true;
	signal I4681: std_logic; attribute dont_touch of I4681: signal is true;
	signal I4684: std_logic; attribute dont_touch of I4684: signal is true;
	signal I4687: std_logic; attribute dont_touch of I4687: signal is true;
	signal I4690: std_logic; attribute dont_touch of I4690: signal is true;
	signal I4693: std_logic; attribute dont_touch of I4693: signal is true;
	signal I4696: std_logic; attribute dont_touch of I4696: signal is true;
	signal I4699: std_logic; attribute dont_touch of I4699: signal is true;
	signal I4702: std_logic; attribute dont_touch of I4702: signal is true;
	signal I4705: std_logic; attribute dont_touch of I4705: signal is true;
	signal I4708: std_logic; attribute dont_touch of I4708: signal is true;
	signal I4711: std_logic; attribute dont_touch of I4711: signal is true;
	signal I4714: std_logic; attribute dont_touch of I4714: signal is true;
	signal I4717: std_logic; attribute dont_touch of I4717: signal is true;
	signal I4720: std_logic; attribute dont_touch of I4720: signal is true;
	signal I4723: std_logic; attribute dont_touch of I4723: signal is true;
	signal I4726: std_logic; attribute dont_touch of I4726: signal is true;
	signal I4729: std_logic; attribute dont_touch of I4729: signal is true;
	signal I4732: std_logic; attribute dont_touch of I4732: signal is true;
	signal I4735: std_logic; attribute dont_touch of I4735: signal is true;
	signal I4738: std_logic; attribute dont_touch of I4738: signal is true;
	signal I4741: std_logic; attribute dont_touch of I4741: signal is true;
	signal I4744: std_logic; attribute dont_touch of I4744: signal is true;
	signal I4747: std_logic; attribute dont_touch of I4747: signal is true;
	signal I4750: std_logic; attribute dont_touch of I4750: signal is true;
	signal I4753: std_logic; attribute dont_touch of I4753: signal is true;
	signal I4756: std_logic; attribute dont_touch of I4756: signal is true;
	signal I4759: std_logic; attribute dont_touch of I4759: signal is true;
	signal I4762: std_logic; attribute dont_touch of I4762: signal is true;
	signal I4765: std_logic; attribute dont_touch of I4765: signal is true;
	signal I4768: std_logic; attribute dont_touch of I4768: signal is true;
	signal I4771: std_logic; attribute dont_touch of I4771: signal is true;
	signal I4774: std_logic; attribute dont_touch of I4774: signal is true;
	signal I4777: std_logic; attribute dont_touch of I4777: signal is true;
	signal I4780: std_logic; attribute dont_touch of I4780: signal is true;
	signal I4783: std_logic; attribute dont_touch of I4783: signal is true;
	signal I4786: std_logic; attribute dont_touch of I4786: signal is true;
	signal I4789: std_logic; attribute dont_touch of I4789: signal is true;
	signal I4792: std_logic; attribute dont_touch of I4792: signal is true;
	signal I4795: std_logic; attribute dont_touch of I4795: signal is true;
	signal I4798: std_logic; attribute dont_touch of I4798: signal is true;
	signal N11GAT: std_logic; attribute dont_touch of N11GAT: signal is true;
	signal N12GAT: std_logic; attribute dont_touch of N12GAT: signal is true;
	signal N13GAT: std_logic; attribute dont_touch of N13GAT: signal is true;
	signal N14GAT: std_logic; attribute dont_touch of N14GAT: signal is true;
	signal N15GAT: std_logic; attribute dont_touch of N15GAT: signal is true;
	signal N16GAT: std_logic; attribute dont_touch of N16GAT: signal is true;
	signal N17GAT: std_logic; attribute dont_touch of N17GAT: signal is true;
	signal N21GAT: std_logic; attribute dont_touch of N21GAT: signal is true;
	signal N22GAT: std_logic; attribute dont_touch of N22GAT: signal is true;
	signal N34GAT: std_logic; attribute dont_touch of N34GAT: signal is true;
	signal N35GAT: std_logic; attribute dont_touch of N35GAT: signal is true;
	signal N37GAT: std_logic; attribute dont_touch of N37GAT: signal is true;
	signal N38GAT: std_logic; attribute dont_touch of N38GAT: signal is true;
	signal N39GAT: std_logic; attribute dont_touch of N39GAT: signal is true;
	signal N40GAT: std_logic; attribute dont_touch of N40GAT: signal is true;
	signal N41GAT: std_logic; attribute dont_touch of N41GAT: signal is true;
	signal N42GAT: std_logic; attribute dont_touch of N42GAT: signal is true;
	signal N43GAT: std_logic; attribute dont_touch of N43GAT: signal is true;
	signal N44GAT: std_logic; attribute dont_touch of N44GAT: signal is true;
	signal N45GAT: std_logic; attribute dont_touch of N45GAT: signal is true;
	signal N46GAT: std_logic; attribute dont_touch of N46GAT: signal is true;
	signal N47GAT: std_logic; attribute dont_touch of N47GAT: signal is true;
	signal N48GAT: std_logic; attribute dont_touch of N48GAT: signal is true;
	signal N49GAT: std_logic; attribute dont_touch of N49GAT: signal is true;
	signal N50GAT: std_logic; attribute dont_touch of N50GAT: signal is true;
	signal N51GAT: std_logic; attribute dont_touch of N51GAT: signal is true;
	signal N52GAT: std_logic; attribute dont_touch of N52GAT: signal is true;
	signal N53GAT: std_logic; attribute dont_touch of N53GAT: signal is true;
	signal N54GAT: std_logic; attribute dont_touch of N54GAT: signal is true;
	signal N55GAT: std_logic; attribute dont_touch of N55GAT: signal is true;
	signal N56GAT: std_logic; attribute dont_touch of N56GAT: signal is true;
	signal N57GAT: std_logic; attribute dont_touch of N57GAT: signal is true;
	signal N58GAT: std_logic; attribute dont_touch of N58GAT: signal is true;
	signal N59GAT: std_logic; attribute dont_touch of N59GAT: signal is true;
	signal N60GAT: std_logic; attribute dont_touch of N60GAT: signal is true;
	signal N61GAT: std_logic; attribute dont_touch of N61GAT: signal is true;
	signal N62GAT: std_logic; attribute dont_touch of N62GAT: signal is true;
	signal N63GAT: std_logic; attribute dont_touch of N63GAT: signal is true;
	signal N64GAT: std_logic; attribute dont_touch of N64GAT: signal is true;
	signal N65GAT: std_logic; attribute dont_touch of N65GAT: signal is true;
	signal N66GAT: std_logic; attribute dont_touch of N66GAT: signal is true;
	signal N67GAT: std_logic; attribute dont_touch of N67GAT: signal is true;
	signal N68GAT: std_logic; attribute dont_touch of N68GAT: signal is true;
	signal N69GAT: std_logic; attribute dont_touch of N69GAT: signal is true;
	signal N70GAT: std_logic; attribute dont_touch of N70GAT: signal is true;
	signal N71GAT: std_logic; attribute dont_touch of N71GAT: signal is true;
	signal N72GAT: std_logic; attribute dont_touch of N72GAT: signal is true;
	signal N73GAT: std_logic; attribute dont_touch of N73GAT: signal is true;
	signal N76GAT: std_logic; attribute dont_touch of N76GAT: signal is true;
	signal N77GAT: std_logic; attribute dont_touch of N77GAT: signal is true;
	signal N78GAT: std_logic; attribute dont_touch of N78GAT: signal is true;
	signal N79GAT: std_logic; attribute dont_touch of N79GAT: signal is true;
	signal N82GAT: std_logic; attribute dont_touch of N82GAT: signal is true;
	signal N84GAT: std_logic; attribute dont_touch of N84GAT: signal is true;
	signal N85GAT: std_logic; attribute dont_touch of N85GAT: signal is true;
	signal N86GAT: std_logic; attribute dont_touch of N86GAT: signal is true;
	signal N87GAT: std_logic; attribute dont_touch of N87GAT: signal is true;
	signal N88GAT: std_logic; attribute dont_touch of N88GAT: signal is true;
	signal N89GAT: std_logic; attribute dont_touch of N89GAT: signal is true;
	signal N92GAT: std_logic; attribute dont_touch of N92GAT: signal is true;
	signal N93GAT: std_logic; attribute dont_touch of N93GAT: signal is true;
	signal N110GAT: std_logic; attribute dont_touch of N110GAT: signal is true;
	signal N111GAT: std_logic; attribute dont_touch of N111GAT: signal is true;
	signal N120GAT: std_logic; attribute dont_touch of N120GAT: signal is true;
	signal N121GAT: std_logic; attribute dont_touch of N121GAT: signal is true;
	signal N122GAT: std_logic; attribute dont_touch of N122GAT: signal is true;
	signal N123GAT: std_logic; attribute dont_touch of N123GAT: signal is true;
	signal N124GAT: std_logic; attribute dont_touch of N124GAT: signal is true;
	signal N125GAT: std_logic; attribute dont_touch of N125GAT: signal is true;
	signal N126GAT: std_logic; attribute dont_touch of N126GAT: signal is true;
	signal N127GAT: std_logic; attribute dont_touch of N127GAT: signal is true;
	signal N128GAT: std_logic; attribute dont_touch of N128GAT: signal is true;
	signal N129GAT: std_logic; attribute dont_touch of N129GAT: signal is true;
	signal N130GAT: std_logic; attribute dont_touch of N130GAT: signal is true;
	signal N132GAT: std_logic; attribute dont_touch of N132GAT: signal is true;
	signal N133GAT: std_logic; attribute dont_touch of N133GAT: signal is true;
	signal N134GAT: std_logic; attribute dont_touch of N134GAT: signal is true;
	signal N136GAT: std_logic; attribute dont_touch of N136GAT: signal is true;
	signal N137GAT: std_logic; attribute dont_touch of N137GAT: signal is true;
	signal N139GAT: std_logic; attribute dont_touch of N139GAT: signal is true;
	signal N140GAT: std_logic; attribute dont_touch of N140GAT: signal is true;
	signal N141GAT: std_logic; attribute dont_touch of N141GAT: signal is true;
	signal N142GAT: std_logic; attribute dont_touch of N142GAT: signal is true;
	signal N143GAT: std_logic; attribute dont_touch of N143GAT: signal is true;
	signal N144GAT: std_logic; attribute dont_touch of N144GAT: signal is true;
	signal N145GAT: std_logic; attribute dont_touch of N145GAT: signal is true;
	signal N146GAT: std_logic; attribute dont_touch of N146GAT: signal is true;
	signal N147GAT: std_logic; attribute dont_touch of N147GAT: signal is true;
	signal N148GAT: std_logic; attribute dont_touch of N148GAT: signal is true;
	signal N150GAT: std_logic; attribute dont_touch of N150GAT: signal is true;
	signal N151GAT: std_logic; attribute dont_touch of N151GAT: signal is true;
	signal N152GAT: std_logic; attribute dont_touch of N152GAT: signal is true;
	signal N154GAT: std_logic; attribute dont_touch of N154GAT: signal is true;
	signal N155GAT: std_logic; attribute dont_touch of N155GAT: signal is true;
	signal N156GAT: std_logic; attribute dont_touch of N156GAT: signal is true;
	signal N158GAT: std_logic; attribute dont_touch of N158GAT: signal is true;
	signal N159GAT: std_logic; attribute dont_touch of N159GAT: signal is true;
	signal N160GAT: std_logic; attribute dont_touch of N160GAT: signal is true;
	signal N162GAT: std_logic; attribute dont_touch of N162GAT: signal is true;
	signal N163GAT: std_logic; attribute dont_touch of N163GAT: signal is true;
	signal N164GAT: std_logic; attribute dont_touch of N164GAT: signal is true;
	signal N165GAT: std_logic; attribute dont_touch of N165GAT: signal is true;
	signal N167GAT: std_logic; attribute dont_touch of N167GAT: signal is true;
	signal N168GAT: std_logic; attribute dont_touch of N168GAT: signal is true;
	signal N169GAT: std_logic; attribute dont_touch of N169GAT: signal is true;
	signal N170GAT: std_logic; attribute dont_touch of N170GAT: signal is true;
	signal N171GAT: std_logic; attribute dont_touch of N171GAT: signal is true;
	signal N172GAT: std_logic; attribute dont_touch of N172GAT: signal is true;
	signal N173GAT: std_logic; attribute dont_touch of N173GAT: signal is true;
	signal N174GAT: std_logic; attribute dont_touch of N174GAT: signal is true;
	signal N175GAT: std_logic; attribute dont_touch of N175GAT: signal is true;
	signal N176GAT: std_logic; attribute dont_touch of N176GAT: signal is true;
	signal N177GAT: std_logic; attribute dont_touch of N177GAT: signal is true;
	signal N178GAT: std_logic; attribute dont_touch of N178GAT: signal is true;
	signal N179GAT: std_logic; attribute dont_touch of N179GAT: signal is true;
	signal N180GAT: std_logic; attribute dont_touch of N180GAT: signal is true;
	signal N181GAT: std_logic; attribute dont_touch of N181GAT: signal is true;
	signal N182GAT: std_logic; attribute dont_touch of N182GAT: signal is true;
	signal N184GAT: std_logic; attribute dont_touch of N184GAT: signal is true;
	signal N186GAT: std_logic; attribute dont_touch of N186GAT: signal is true;
	signal N187GAT: std_logic; attribute dont_touch of N187GAT: signal is true;
	signal N188GAT: std_logic; attribute dont_touch of N188GAT: signal is true;
	signal N189GAT: std_logic; attribute dont_touch of N189GAT: signal is true;
	signal N194GAT: std_logic; attribute dont_touch of N194GAT: signal is true;
	signal N195GAT: std_logic; attribute dont_touch of N195GAT: signal is true;
	signal N196GAT: std_logic; attribute dont_touch of N196GAT: signal is true;
	signal N197GAT: std_logic; attribute dont_touch of N197GAT: signal is true;
	signal N199GAT: std_logic; attribute dont_touch of N199GAT: signal is true;
	signal N200GAT: std_logic; attribute dont_touch of N200GAT: signal is true;
	signal N204GAT: std_logic; attribute dont_touch of N204GAT: signal is true;
	signal N207GAT: std_logic; attribute dont_touch of N207GAT: signal is true;
	signal N212GAT: std_logic; attribute dont_touch of N212GAT: signal is true;
	signal N219GAT: std_logic; attribute dont_touch of N219GAT: signal is true;
	signal N221GAT: std_logic; attribute dont_touch of N221GAT: signal is true;
	signal N222GAT: std_logic; attribute dont_touch of N222GAT: signal is true;
	signal N223GAT: std_logic; attribute dont_touch of N223GAT: signal is true;
	signal N224GAT: std_logic; attribute dont_touch of N224GAT: signal is true;
	signal N225GAT: std_logic; attribute dont_touch of N225GAT: signal is true;
	signal N226GAT: std_logic; attribute dont_touch of N226GAT: signal is true;
	signal N227GAT: std_logic; attribute dont_touch of N227GAT: signal is true;
	signal N228GAT: std_logic; attribute dont_touch of N228GAT: signal is true;
	signal N229GAT: std_logic; attribute dont_touch of N229GAT: signal is true;
	signal N230GAT: std_logic; attribute dont_touch of N230GAT: signal is true;
	signal N231GAT: std_logic; attribute dont_touch of N231GAT: signal is true;
	signal N233GAT: std_logic; attribute dont_touch of N233GAT: signal is true;
	signal N234GAT: std_logic; attribute dont_touch of N234GAT: signal is true;
	signal N235GAT: std_logic; attribute dont_touch of N235GAT: signal is true;
	signal N237GAT: std_logic; attribute dont_touch of N237GAT: signal is true;
	signal N238GAT: std_logic; attribute dont_touch of N238GAT: signal is true;
	signal N240GAT: std_logic; attribute dont_touch of N240GAT: signal is true;
	signal N241GAT: std_logic; attribute dont_touch of N241GAT: signal is true;
	signal N242GAT: std_logic; attribute dont_touch of N242GAT: signal is true;
	signal N243GAT: std_logic; attribute dont_touch of N243GAT: signal is true;
	signal N244GAT: std_logic; attribute dont_touch of N244GAT: signal is true;
	signal N245GAT: std_logic; attribute dont_touch of N245GAT: signal is true;
	signal N246GAT: std_logic; attribute dont_touch of N246GAT: signal is true;
	signal N247GAT: std_logic; attribute dont_touch of N247GAT: signal is true;
	signal N248GAT: std_logic; attribute dont_touch of N248GAT: signal is true;
	signal N249GAT: std_logic; attribute dont_touch of N249GAT: signal is true;
	signal N250GAT: std_logic; attribute dont_touch of N250GAT: signal is true;
	signal N251GAT: std_logic; attribute dont_touch of N251GAT: signal is true;
	signal N252GAT: std_logic; attribute dont_touch of N252GAT: signal is true;
	signal N253GAT: std_logic; attribute dont_touch of N253GAT: signal is true;
	signal N254GAT: std_logic; attribute dont_touch of N254GAT: signal is true;
	signal N255GAT: std_logic; attribute dont_touch of N255GAT: signal is true;
	signal N256GAT: std_logic; attribute dont_touch of N256GAT: signal is true;
	signal N258GAT: std_logic; attribute dont_touch of N258GAT: signal is true;
	signal N259GAT: std_logic; attribute dont_touch of N259GAT: signal is true;
	signal N260GAT: std_logic; attribute dont_touch of N260GAT: signal is true;
	signal N261GAT: std_logic; attribute dont_touch of N261GAT: signal is true;
	signal N262GAT: std_logic; attribute dont_touch of N262GAT: signal is true;
	signal N263GAT: std_logic; attribute dont_touch of N263GAT: signal is true;
	signal N264GAT: std_logic; attribute dont_touch of N264GAT: signal is true;
	signal N265GAT: std_logic; attribute dont_touch of N265GAT: signal is true;
	signal N266GAT: std_logic; attribute dont_touch of N266GAT: signal is true;
	signal N267GAT: std_logic; attribute dont_touch of N267GAT: signal is true;
	signal N268GAT: std_logic; attribute dont_touch of N268GAT: signal is true;
	signal N269GAT: std_logic; attribute dont_touch of N269GAT: signal is true;
	signal N270GAT: std_logic; attribute dont_touch of N270GAT: signal is true;
	signal N271GAT: std_logic; attribute dont_touch of N271GAT: signal is true;
	signal N273GAT: std_logic; attribute dont_touch of N273GAT: signal is true;
	signal N274GAT: std_logic; attribute dont_touch of N274GAT: signal is true;
	signal N275GAT: std_logic; attribute dont_touch of N275GAT: signal is true;
	signal N277GAT: std_logic; attribute dont_touch of N277GAT: signal is true;
	signal N278GAT: std_logic; attribute dont_touch of N278GAT: signal is true;
	signal N279GAT: std_logic; attribute dont_touch of N279GAT: signal is true;
	signal N281GAT: std_logic; attribute dont_touch of N281GAT: signal is true;
	signal N282GAT: std_logic; attribute dont_touch of N282GAT: signal is true;
	signal N283GAT: std_logic; attribute dont_touch of N283GAT: signal is true;
	signal N286GAT: std_logic; attribute dont_touch of N286GAT: signal is true;
	signal N287GAT: std_logic; attribute dont_touch of N287GAT: signal is true;
	signal N288GAT: std_logic; attribute dont_touch of N288GAT: signal is true;
	signal N289GAT: std_logic; attribute dont_touch of N289GAT: signal is true;
	signal N290GAT: std_logic; attribute dont_touch of N290GAT: signal is true;
	signal N291GAT: std_logic; attribute dont_touch of N291GAT: signal is true;
	signal N292GAT: std_logic; attribute dont_touch of N292GAT: signal is true;
	signal N293GAT: std_logic; attribute dont_touch of N293GAT: signal is true;
	signal N294GAT: std_logic; attribute dont_touch of N294GAT: signal is true;
	signal N295GAT: std_logic; attribute dont_touch of N295GAT: signal is true;
	signal N296GAT: std_logic; attribute dont_touch of N296GAT: signal is true;
	signal N297GAT: std_logic; attribute dont_touch of N297GAT: signal is true;
	signal N299GAT: std_logic; attribute dont_touch of N299GAT: signal is true;
	signal N312GAT: std_logic; attribute dont_touch of N312GAT: signal is true;
	signal N313GAT: std_logic; attribute dont_touch of N313GAT: signal is true;
	signal N314GAT: std_logic; attribute dont_touch of N314GAT: signal is true;
	signal N316GAT: std_logic; attribute dont_touch of N316GAT: signal is true;
	signal N317GAT: std_logic; attribute dont_touch of N317GAT: signal is true;
	signal N318GAT: std_logic; attribute dont_touch of N318GAT: signal is true;
	signal N320GAT: std_logic; attribute dont_touch of N320GAT: signal is true;
	signal N321GAT: std_logic; attribute dont_touch of N321GAT: signal is true;
	signal N322GAT: std_logic; attribute dont_touch of N322GAT: signal is true;
	signal N324GAT: std_logic; attribute dont_touch of N324GAT: signal is true;
	signal N325GAT: std_logic; attribute dont_touch of N325GAT: signal is true;
	signal N326GAT: std_logic; attribute dont_touch of N326GAT: signal is true;
	signal N327GAT: std_logic; attribute dont_touch of N327GAT: signal is true;
	signal N329GAT: std_logic; attribute dont_touch of N329GAT: signal is true;
	signal N330GAT: std_logic; attribute dont_touch of N330GAT: signal is true;
	signal N331GAT: std_logic; attribute dont_touch of N331GAT: signal is true;
	signal N333GAT: std_logic; attribute dont_touch of N333GAT: signal is true;
	signal N334GAT: std_logic; attribute dont_touch of N334GAT: signal is true;
	signal N335GAT: std_logic; attribute dont_touch of N335GAT: signal is true;
	signal N336GAT: std_logic; attribute dont_touch of N336GAT: signal is true;
	signal N337GAT: std_logic; attribute dont_touch of N337GAT: signal is true;
	signal N339GAT: std_logic; attribute dont_touch of N339GAT: signal is true;
	signal N340GAT: std_logic; attribute dont_touch of N340GAT: signal is true;
	signal N341GAT: std_logic; attribute dont_touch of N341GAT: signal is true;
	signal N343GAT: std_logic; attribute dont_touch of N343GAT: signal is true;
	signal N344GAT: std_logic; attribute dont_touch of N344GAT: signal is true;
	signal N345GAT: std_logic; attribute dont_touch of N345GAT: signal is true;
	signal N346GAT: std_logic; attribute dont_touch of N346GAT: signal is true;
	signal N347GAT: std_logic; attribute dont_touch of N347GAT: signal is true;
	signal N348GAT: std_logic; attribute dont_touch of N348GAT: signal is true;
	signal N349GAT: std_logic; attribute dont_touch of N349GAT: signal is true;
	signal N350GAT: std_logic; attribute dont_touch of N350GAT: signal is true;
	signal N351GAT: std_logic; attribute dont_touch of N351GAT: signal is true;
	signal N352GAT: std_logic; attribute dont_touch of N352GAT: signal is true;
	signal N353GAT: std_logic; attribute dont_touch of N353GAT: signal is true;
	signal N354GAT: std_logic; attribute dont_touch of N354GAT: signal is true;
	signal N355GAT: std_logic; attribute dont_touch of N355GAT: signal is true;
	signal N356GAT: std_logic; attribute dont_touch of N356GAT: signal is true;
	signal N357GAT: std_logic; attribute dont_touch of N357GAT: signal is true;
	signal N358GAT: std_logic; attribute dont_touch of N358GAT: signal is true;
	signal N359GAT: std_logic; attribute dont_touch of N359GAT: signal is true;
	signal N360GAT: std_logic; attribute dont_touch of N360GAT: signal is true;
	signal N361GAT: std_logic; attribute dont_touch of N361GAT: signal is true;
	signal N362GAT: std_logic; attribute dont_touch of N362GAT: signal is true;
	signal N364GAT: std_logic; attribute dont_touch of N364GAT: signal is true;
	signal N365GAT: std_logic; attribute dont_touch of N365GAT: signal is true;
	signal N366GAT: std_logic; attribute dont_touch of N366GAT: signal is true;
	signal N368GAT: std_logic; attribute dont_touch of N368GAT: signal is true;
	signal N369GAT: std_logic; attribute dont_touch of N369GAT: signal is true;
	signal N370GAT: std_logic; attribute dont_touch of N370GAT: signal is true;
	signal N371GAT: std_logic; attribute dont_touch of N371GAT: signal is true;
	signal N372GAT: std_logic; attribute dont_touch of N372GAT: signal is true;
	signal N373GAT: std_logic; attribute dont_touch of N373GAT: signal is true;
	signal N374GAT: std_logic; attribute dont_touch of N374GAT: signal is true;
	signal N375GAT: std_logic; attribute dont_touch of N375GAT: signal is true;
	signal N377GAT: std_logic; attribute dont_touch of N377GAT: signal is true;
	signal N378GAT: std_logic; attribute dont_touch of N378GAT: signal is true;
	signal N380GAT: std_logic; attribute dont_touch of N380GAT: signal is true;
	signal N381GAT: std_logic; attribute dont_touch of N381GAT: signal is true;
	signal N382GAT: std_logic; attribute dont_touch of N382GAT: signal is true;
	signal N383GAT: std_logic; attribute dont_touch of N383GAT: signal is true;
	signal N384GAT: std_logic; attribute dont_touch of N384GAT: signal is true;
	signal N386GAT: std_logic; attribute dont_touch of N386GAT: signal is true;
	signal N387GAT: std_logic; attribute dont_touch of N387GAT: signal is true;
	signal N388GAT: std_logic; attribute dont_touch of N388GAT: signal is true;
	signal N390GAT: std_logic; attribute dont_touch of N390GAT: signal is true;
	signal N391GAT: std_logic; attribute dont_touch of N391GAT: signal is true;
	signal N392GAT: std_logic; attribute dont_touch of N392GAT: signal is true;
	signal N393GAT: std_logic; attribute dont_touch of N393GAT: signal is true;
	signal N394GAT: std_logic; attribute dont_touch of N394GAT: signal is true;
	signal N396GAT: std_logic; attribute dont_touch of N396GAT: signal is true;
	signal N397GAT: std_logic; attribute dont_touch of N397GAT: signal is true;
	signal N398GAT: std_logic; attribute dont_touch of N398GAT: signal is true;
	signal N400GAT: std_logic; attribute dont_touch of N400GAT: signal is true;
	signal N401GAT: std_logic; attribute dont_touch of N401GAT: signal is true;
	signal N402GAT: std_logic; attribute dont_touch of N402GAT: signal is true;
	signal N404GAT: std_logic; attribute dont_touch of N404GAT: signal is true;
	signal N405GAT: std_logic; attribute dont_touch of N405GAT: signal is true;
	signal N406GAT: std_logic; attribute dont_touch of N406GAT: signal is true;
	signal N407GAT: std_logic; attribute dont_touch of N407GAT: signal is true;
	signal N408GAT: std_logic; attribute dont_touch of N408GAT: signal is true;
	signal N409GAT: std_logic; attribute dont_touch of N409GAT: signal is true;
	signal N410GAT: std_logic; attribute dont_touch of N410GAT: signal is true;
	signal N411GAT: std_logic; attribute dont_touch of N411GAT: signal is true;
	signal N412GAT: std_logic; attribute dont_touch of N412GAT: signal is true;
	signal N413GAT: std_logic; attribute dont_touch of N413GAT: signal is true;
	signal N414GAT: std_logic; attribute dont_touch of N414GAT: signal is true;
	signal N415GAT: std_logic; attribute dont_touch of N415GAT: signal is true;
	signal N416GAT: std_logic; attribute dont_touch of N416GAT: signal is true;
	signal N417GAT: std_logic; attribute dont_touch of N417GAT: signal is true;
	signal N418GAT: std_logic; attribute dont_touch of N418GAT: signal is true;
	signal N419GAT: std_logic; attribute dont_touch of N419GAT: signal is true;
	signal N420GAT: std_logic; attribute dont_touch of N420GAT: signal is true;
	signal N421GAT: std_logic; attribute dont_touch of N421GAT: signal is true;
	signal N422GAT: std_logic; attribute dont_touch of N422GAT: signal is true;
	signal N423GAT: std_logic; attribute dont_touch of N423GAT: signal is true;
	signal N439GAT: std_logic; attribute dont_touch of N439GAT: signal is true;
	signal N440GAT: std_logic; attribute dont_touch of N440GAT: signal is true;
	signal N441GAT: std_logic; attribute dont_touch of N441GAT: signal is true;
	signal N442GAT: std_logic; attribute dont_touch of N442GAT: signal is true;
	signal N443GAT: std_logic; attribute dont_touch of N443GAT: signal is true;
	signal N444GAT: std_logic; attribute dont_touch of N444GAT: signal is true;
	signal N445GAT: std_logic; attribute dont_touch of N445GAT: signal is true;
	signal N446GAT: std_logic; attribute dont_touch of N446GAT: signal is true;
	signal N447GAT: std_logic; attribute dont_touch of N447GAT: signal is true;
	signal N448GAT: std_logic; attribute dont_touch of N448GAT: signal is true;
	signal N449GAT: std_logic; attribute dont_touch of N449GAT: signal is true;
	signal N450GAT: std_logic; attribute dont_touch of N450GAT: signal is true;
	signal N451GAT: std_logic; attribute dont_touch of N451GAT: signal is true;
	signal N452GAT: std_logic; attribute dont_touch of N452GAT: signal is true;
	signal N453GAT: std_logic; attribute dont_touch of N453GAT: signal is true;
	signal N455GAT: std_logic; attribute dont_touch of N455GAT: signal is true;
	signal N456GAT: std_logic; attribute dont_touch of N456GAT: signal is true;
	signal N457GAT: std_logic; attribute dont_touch of N457GAT: signal is true;
	signal N458GAT: std_logic; attribute dont_touch of N458GAT: signal is true;
	signal N459GAT: std_logic; attribute dont_touch of N459GAT: signal is true;
	signal N460GAT: std_logic; attribute dont_touch of N460GAT: signal is true;
	signal N461GAT: std_logic; attribute dont_touch of N461GAT: signal is true;
	signal N462GAT: std_logic; attribute dont_touch of N462GAT: signal is true;
	signal N463GAT: std_logic; attribute dont_touch of N463GAT: signal is true;
	signal N468GAT: std_logic; attribute dont_touch of N468GAT: signal is true;
	signal N469GAT: std_logic; attribute dont_touch of N469GAT: signal is true;
	signal N470GAT: std_logic; attribute dont_touch of N470GAT: signal is true;
	signal N475GAT: std_logic; attribute dont_touch of N475GAT: signal is true;
	signal N476GAT: std_logic; attribute dont_touch of N476GAT: signal is true;
	signal N477GAT: std_logic; attribute dont_touch of N477GAT: signal is true;
	signal N478GAT: std_logic; attribute dont_touch of N478GAT: signal is true;
	signal N479GAT: std_logic; attribute dont_touch of N479GAT: signal is true;
	signal N480GAT: std_logic; attribute dont_touch of N480GAT: signal is true;
	signal N481GAT: std_logic; attribute dont_touch of N481GAT: signal is true;
	signal N482GAT: std_logic; attribute dont_touch of N482GAT: signal is true;
	signal N483GAT: std_logic; attribute dont_touch of N483GAT: signal is true;
	signal N484GAT: std_logic; attribute dont_touch of N484GAT: signal is true;
	signal N485GAT: std_logic; attribute dont_touch of N485GAT: signal is true;
	signal N489GAT: std_logic; attribute dont_touch of N489GAT: signal is true;
	signal N490GAT: std_logic; attribute dont_touch of N490GAT: signal is true;
	signal N491GAT: std_logic; attribute dont_touch of N491GAT: signal is true;
	signal N493GAT: std_logic; attribute dont_touch of N493GAT: signal is true;
	signal N494GAT: std_logic; attribute dont_touch of N494GAT: signal is true;
	signal N495GAT: std_logic; attribute dont_touch of N495GAT: signal is true;
	signal N496GAT: std_logic; attribute dont_touch of N496GAT: signal is true;
	signal N497GAT: std_logic; attribute dont_touch of N497GAT: signal is true;
	signal N498GAT: std_logic; attribute dont_touch of N498GAT: signal is true;
	signal N499GAT: std_logic; attribute dont_touch of N499GAT: signal is true;
	signal N500GAT: std_logic; attribute dont_touch of N500GAT: signal is true;
	signal N501GAT: std_logic; attribute dont_touch of N501GAT: signal is true;
	signal N502GAT: std_logic; attribute dont_touch of N502GAT: signal is true;
	signal N503GAT: std_logic; attribute dont_touch of N503GAT: signal is true;
	signal N504GAT: std_logic; attribute dont_touch of N504GAT: signal is true;
	signal N505GAT: std_logic; attribute dont_touch of N505GAT: signal is true;
	signal N506GAT: std_logic; attribute dont_touch of N506GAT: signal is true;
	signal N507GAT: std_logic; attribute dont_touch of N507GAT: signal is true;
	signal N508GAT: std_logic; attribute dont_touch of N508GAT: signal is true;
	signal N509GAT: std_logic; attribute dont_touch of N509GAT: signal is true;
	signal N510GAT: std_logic; attribute dont_touch of N510GAT: signal is true;
	signal N511GAT: std_logic; attribute dont_touch of N511GAT: signal is true;
	signal N512GAT: std_logic; attribute dont_touch of N512GAT: signal is true;
	signal N513GAT: std_logic; attribute dont_touch of N513GAT: signal is true;
	signal N514GAT: std_logic; attribute dont_touch of N514GAT: signal is true;
	signal N515GAT: std_logic; attribute dont_touch of N515GAT: signal is true;
	signal N516GAT: std_logic; attribute dont_touch of N516GAT: signal is true;
	signal N517GAT: std_logic; attribute dont_touch of N517GAT: signal is true;
	signal N518GAT: std_logic; attribute dont_touch of N518GAT: signal is true;
	signal N519GAT: std_logic; attribute dont_touch of N519GAT: signal is true;
	signal N520GAT: std_logic; attribute dont_touch of N520GAT: signal is true;
	signal N521GAT: std_logic; attribute dont_touch of N521GAT: signal is true;
	signal N522GAT: std_logic; attribute dont_touch of N522GAT: signal is true;
	signal N523GAT: std_logic; attribute dont_touch of N523GAT: signal is true;
	signal N524GAT: std_logic; attribute dont_touch of N524GAT: signal is true;
	signal N525GAT: std_logic; attribute dont_touch of N525GAT: signal is true;
	signal N526GAT: std_logic; attribute dont_touch of N526GAT: signal is true;
	signal N527GAT: std_logic; attribute dont_touch of N527GAT: signal is true;
	signal N528GAT: std_logic; attribute dont_touch of N528GAT: signal is true;
	signal N529GAT: std_logic; attribute dont_touch of N529GAT: signal is true;
	signal N530GAT: std_logic; attribute dont_touch of N530GAT: signal is true;
	signal N531GAT: std_logic; attribute dont_touch of N531GAT: signal is true;
	signal N532GAT: std_logic; attribute dont_touch of N532GAT: signal is true;
	signal N551GAT: std_logic; attribute dont_touch of N551GAT: signal is true;
	signal N552GAT: std_logic; attribute dont_touch of N552GAT: signal is true;
	signal N553GAT: std_logic; attribute dont_touch of N553GAT: signal is true;
	signal N555GAT: std_logic; attribute dont_touch of N555GAT: signal is true;
	signal N556GAT: std_logic; attribute dont_touch of N556GAT: signal is true;
	signal N557GAT: std_logic; attribute dont_touch of N557GAT: signal is true;
	signal N558GAT: std_logic; attribute dont_touch of N558GAT: signal is true;
	signal N559GAT: std_logic; attribute dont_touch of N559GAT: signal is true;
	signal N560GAT: std_logic; attribute dont_touch of N560GAT: signal is true;
	signal N561GAT: std_logic; attribute dont_touch of N561GAT: signal is true;
	signal N563GAT: std_logic; attribute dont_touch of N563GAT: signal is true;
	signal N564GAT: std_logic; attribute dont_touch of N564GAT: signal is true;
	signal N565GAT: std_logic; attribute dont_touch of N565GAT: signal is true;
	signal N566GAT: std_logic; attribute dont_touch of N566GAT: signal is true;
	signal N567GAT: std_logic; attribute dont_touch of N567GAT: signal is true;
	signal N568GAT: std_logic; attribute dont_touch of N568GAT: signal is true;
	signal N569GAT: std_logic; attribute dont_touch of N569GAT: signal is true;
	signal N570GAT: std_logic; attribute dont_touch of N570GAT: signal is true;
	signal N571GAT: std_logic; attribute dont_touch of N571GAT: signal is true;
	signal N572GAT: std_logic; attribute dont_touch of N572GAT: signal is true;
	signal N573GAT: std_logic; attribute dont_touch of N573GAT: signal is true;
	signal N574GAT: std_logic; attribute dont_touch of N574GAT: signal is true;
	signal N575GAT: std_logic; attribute dont_touch of N575GAT: signal is true;
	signal N576GAT: std_logic; attribute dont_touch of N576GAT: signal is true;
	signal N577GAT: std_logic; attribute dont_touch of N577GAT: signal is true;
	signal N578GAT: std_logic; attribute dont_touch of N578GAT: signal is true;
	signal N579GAT: std_logic; attribute dont_touch of N579GAT: signal is true;
	signal N580GAT: std_logic; attribute dont_touch of N580GAT: signal is true;
	signal N582GAT: std_logic; attribute dont_touch of N582GAT: signal is true;
	signal N583GAT: std_logic; attribute dont_touch of N583GAT: signal is true;
	signal N584GAT: std_logic; attribute dont_touch of N584GAT: signal is true;
	signal N586GAT: std_logic; attribute dont_touch of N586GAT: signal is true;
	signal N587GAT: std_logic; attribute dont_touch of N587GAT: signal is true;
	signal N588GAT: std_logic; attribute dont_touch of N588GAT: signal is true;
	signal N589GAT: std_logic; attribute dont_touch of N589GAT: signal is true;
	signal N590GAT: std_logic; attribute dont_touch of N590GAT: signal is true;
	signal N591GAT: std_logic; attribute dont_touch of N591GAT: signal is true;
	signal N592GAT: std_logic; attribute dont_touch of N592GAT: signal is true;
	signal N593GAT: std_logic; attribute dont_touch of N593GAT: signal is true;
	signal N594GAT: std_logic; attribute dont_touch of N594GAT: signal is true;
	signal N595GAT: std_logic; attribute dont_touch of N595GAT: signal is true;
	signal N596GAT: std_logic; attribute dont_touch of N596GAT: signal is true;
	signal N612GAT: std_logic; attribute dont_touch of N612GAT: signal is true;
	signal N613GAT: std_logic; attribute dont_touch of N613GAT: signal is true;
	signal N614GAT: std_logic; attribute dont_touch of N614GAT: signal is true;
	signal N616GAT: std_logic; attribute dont_touch of N616GAT: signal is true;
	signal N617GAT: std_logic; attribute dont_touch of N617GAT: signal is true;
	signal N618GAT: std_logic; attribute dont_touch of N618GAT: signal is true;
	signal N620GAT: std_logic; attribute dont_touch of N620GAT: signal is true;
	signal N621GAT: std_logic; attribute dont_touch of N621GAT: signal is true;
	signal N622GAT: std_logic; attribute dont_touch of N622GAT: signal is true;
	signal N624GAT: std_logic; attribute dont_touch of N624GAT: signal is true;
	signal N625GAT: std_logic; attribute dont_touch of N625GAT: signal is true;
	signal N626GAT: std_logic; attribute dont_touch of N626GAT: signal is true;
	signal N628GAT: std_logic; attribute dont_touch of N628GAT: signal is true;
	signal N629GAT: std_logic; attribute dont_touch of N629GAT: signal is true;
	signal N630GAT: std_logic; attribute dont_touch of N630GAT: signal is true;
	signal N631GAT: std_logic; attribute dont_touch of N631GAT: signal is true;
	signal N632GAT: std_logic; attribute dont_touch of N632GAT: signal is true;
	signal N633GAT: std_logic; attribute dont_touch of N633GAT: signal is true;
	signal N634GAT: std_logic; attribute dont_touch of N634GAT: signal is true;
	signal N635GAT: std_logic; attribute dont_touch of N635GAT: signal is true;
	signal N636GAT: std_logic; attribute dont_touch of N636GAT: signal is true;
	signal N637GAT: std_logic; attribute dont_touch of N637GAT: signal is true;
	signal N638GAT: std_logic; attribute dont_touch of N638GAT: signal is true;
	signal N639GAT: std_logic; attribute dont_touch of N639GAT: signal is true;
	signal N640GAT: std_logic; attribute dont_touch of N640GAT: signal is true;
	signal N641GAT: std_logic; attribute dont_touch of N641GAT: signal is true;
	signal N642GAT: std_logic; attribute dont_touch of N642GAT: signal is true;
	signal N643GAT: std_logic; attribute dont_touch of N643GAT: signal is true;
	signal N644GAT: std_logic; attribute dont_touch of N644GAT: signal is true;
	signal N645GAT: std_logic; attribute dont_touch of N645GAT: signal is true;
	signal N646GAT: std_logic; attribute dont_touch of N646GAT: signal is true;
	signal N647GAT: std_logic; attribute dont_touch of N647GAT: signal is true;
	signal N648GAT: std_logic; attribute dont_touch of N648GAT: signal is true;
	signal N649GAT: std_logic; attribute dont_touch of N649GAT: signal is true;
	signal N650GAT: std_logic; attribute dont_touch of N650GAT: signal is true;
	signal N651GAT: std_logic; attribute dont_touch of N651GAT: signal is true;
	signal N652GAT: std_logic; attribute dont_touch of N652GAT: signal is true;
	signal N653GAT: std_logic; attribute dont_touch of N653GAT: signal is true;
	signal N654GAT: std_logic; attribute dont_touch of N654GAT: signal is true;
	signal N655GAT: std_logic; attribute dont_touch of N655GAT: signal is true;
	signal N656GAT: std_logic; attribute dont_touch of N656GAT: signal is true;
	signal N657GAT: std_logic; attribute dont_touch of N657GAT: signal is true;
	signal N658GAT: std_logic; attribute dont_touch of N658GAT: signal is true;
	signal N659GAT: std_logic; attribute dont_touch of N659GAT: signal is true;
	signal N661GAT: std_logic; attribute dont_touch of N661GAT: signal is true;
	signal N662GAT: std_logic; attribute dont_touch of N662GAT: signal is true;
	signal N663GAT: std_logic; attribute dont_touch of N663GAT: signal is true;
	signal N664GAT: std_logic; attribute dont_touch of N664GAT: signal is true;
	signal N665GAT: std_logic; attribute dont_touch of N665GAT: signal is true;
	signal N666GAT: std_logic; attribute dont_touch of N666GAT: signal is true;
	signal N667GAT: std_logic; attribute dont_touch of N667GAT: signal is true;
	signal N670GAT: std_logic; attribute dont_touch of N670GAT: signal is true;
	signal N671GAT: std_logic; attribute dont_touch of N671GAT: signal is true;
	signal N672GAT: std_logic; attribute dont_touch of N672GAT: signal is true;
	signal N673GAT: std_logic; attribute dont_touch of N673GAT: signal is true;
	signal N677GAT: std_logic; attribute dont_touch of N677GAT: signal is true;
	signal N678GAT: std_logic; attribute dont_touch of N678GAT: signal is true;
	signal N679GAT: std_logic; attribute dont_touch of N679GAT: signal is true;
	signal N680GAT: std_logic; attribute dont_touch of N680GAT: signal is true;
	signal N682GAT: std_logic; attribute dont_touch of N682GAT: signal is true;
	signal N683GAT: std_logic; attribute dont_touch of N683GAT: signal is true;
	signal N684GAT: std_logic; attribute dont_touch of N684GAT: signal is true;
	signal N686GAT: std_logic; attribute dont_touch of N686GAT: signal is true;
	signal N687GAT: std_logic; attribute dont_touch of N687GAT: signal is true;
	signal N688GAT: std_logic; attribute dont_touch of N688GAT: signal is true;
	signal N689GAT: std_logic; attribute dont_touch of N689GAT: signal is true;
	signal N690GAT: std_logic; attribute dont_touch of N690GAT: signal is true;
	signal N691GAT: std_logic; attribute dont_touch of N691GAT: signal is true;
	signal N692GAT: std_logic; attribute dont_touch of N692GAT: signal is true;
	signal N693GAT: std_logic; attribute dont_touch of N693GAT: signal is true;
	signal N694GAT: std_logic; attribute dont_touch of N694GAT: signal is true;
	signal N695GAT: std_logic; attribute dont_touch of N695GAT: signal is true;
	signal N696GAT: std_logic; attribute dont_touch of N696GAT: signal is true;
	signal N697GAT: std_logic; attribute dont_touch of N697GAT: signal is true;
	signal N698GAT: std_logic; attribute dont_touch of N698GAT: signal is true;
	signal N699GAT: std_logic; attribute dont_touch of N699GAT: signal is true;
	signal N701GAT: std_logic; attribute dont_touch of N701GAT: signal is true;
	signal N702GAT: std_logic; attribute dont_touch of N702GAT: signal is true;
	signal N703GAT: std_logic; attribute dont_touch of N703GAT: signal is true;
	signal N705GAT: std_logic; attribute dont_touch of N705GAT: signal is true;
	signal N706GAT: std_logic; attribute dont_touch of N706GAT: signal is true;
	signal N707GAT: std_logic; attribute dont_touch of N707GAT: signal is true;
	signal N709GAT: std_logic; attribute dont_touch of N709GAT: signal is true;
	signal N710GAT: std_logic; attribute dont_touch of N710GAT: signal is true;
	signal N711GAT: std_logic; attribute dont_touch of N711GAT: signal is true;
	signal N712GAT: std_logic; attribute dont_touch of N712GAT: signal is true;
	signal N713GAT: std_logic; attribute dont_touch of N713GAT: signal is true;
	signal N714GAT: std_logic; attribute dont_touch of N714GAT: signal is true;
	signal N715GAT: std_logic; attribute dont_touch of N715GAT: signal is true;
	signal N716GAT: std_logic; attribute dont_touch of N716GAT: signal is true;
	signal N717GAT: std_logic; attribute dont_touch of N717GAT: signal is true;
	signal N718GAT: std_logic; attribute dont_touch of N718GAT: signal is true;
	signal N719GAT: std_logic; attribute dont_touch of N719GAT: signal is true;
	signal N720GAT: std_logic; attribute dont_touch of N720GAT: signal is true;
	signal N721GAT: std_logic; attribute dont_touch of N721GAT: signal is true;
	signal N722GAT: std_logic; attribute dont_touch of N722GAT: signal is true;
	signal N724GAT: std_logic; attribute dont_touch of N724GAT: signal is true;
	signal N725GAT: std_logic; attribute dont_touch of N725GAT: signal is true;
	signal N726GAT: std_logic; attribute dont_touch of N726GAT: signal is true;
	signal N728GAT: std_logic; attribute dont_touch of N728GAT: signal is true;
	signal N729GAT: std_logic; attribute dont_touch of N729GAT: signal is true;
	signal N730GAT: std_logic; attribute dont_touch of N730GAT: signal is true;
	signal N731GAT: std_logic; attribute dont_touch of N731GAT: signal is true;
	signal N732GAT: std_logic; attribute dont_touch of N732GAT: signal is true;
	signal N733GAT: std_logic; attribute dont_touch of N733GAT: signal is true;
	signal N734GAT: std_logic; attribute dont_touch of N734GAT: signal is true;
	signal N735GAT: std_logic; attribute dont_touch of N735GAT: signal is true;
	signal N736GAT: std_logic; attribute dont_touch of N736GAT: signal is true;
	signal N737GAT: std_logic; attribute dont_touch of N737GAT: signal is true;
	signal N738GAT: std_logic; attribute dont_touch of N738GAT: signal is true;
	signal N739GAT: std_logic; attribute dont_touch of N739GAT: signal is true;
	signal N740GAT: std_logic; attribute dont_touch of N740GAT: signal is true;
	signal N741GAT: std_logic; attribute dont_touch of N741GAT: signal is true;
	signal N743GAT: std_logic; attribute dont_touch of N743GAT: signal is true;
	signal N745GAT: std_logic; attribute dont_touch of N745GAT: signal is true;
	signal N746GAT: std_logic; attribute dont_touch of N746GAT: signal is true;
	signal N747GAT: std_logic; attribute dont_touch of N747GAT: signal is true;
	signal N748GAT: std_logic; attribute dont_touch of N748GAT: signal is true;
	signal N749GAT: std_logic; attribute dont_touch of N749GAT: signal is true;
	signal N750GAT: std_logic; attribute dont_touch of N750GAT: signal is true;
	signal N751GAT: std_logic; attribute dont_touch of N751GAT: signal is true;
	signal N752GAT: std_logic; attribute dont_touch of N752GAT: signal is true;
	signal N753GAT: std_logic; attribute dont_touch of N753GAT: signal is true;
	signal N754GAT: std_logic; attribute dont_touch of N754GAT: signal is true;
	signal N755GAT: std_logic; attribute dont_touch of N755GAT: signal is true;
	signal N756GAT: std_logic; attribute dont_touch of N756GAT: signal is true;
	signal N757GAT: std_logic; attribute dont_touch of N757GAT: signal is true;
	signal N758GAT: std_logic; attribute dont_touch of N758GAT: signal is true;
	signal N759GAT: std_logic; attribute dont_touch of N759GAT: signal is true;
	signal N760GAT: std_logic; attribute dont_touch of N760GAT: signal is true;
	signal N761GAT: std_logic; attribute dont_touch of N761GAT: signal is true;
	signal N762GAT: std_logic; attribute dont_touch of N762GAT: signal is true;
	signal N763GAT: std_logic; attribute dont_touch of N763GAT: signal is true;
	signal N764GAT: std_logic; attribute dont_touch of N764GAT: signal is true;
	signal N765GAT: std_logic; attribute dont_touch of N765GAT: signal is true;
	signal N766GAT: std_logic; attribute dont_touch of N766GAT: signal is true;
	signal N767GAT: std_logic; attribute dont_touch of N767GAT: signal is true;
	signal N768GAT: std_logic; attribute dont_touch of N768GAT: signal is true;
	signal N769GAT: std_logic; attribute dont_touch of N769GAT: signal is true;
	signal N771GAT: std_logic; attribute dont_touch of N771GAT: signal is true;
	signal N772GAT: std_logic; attribute dont_touch of N772GAT: signal is true;
	signal N773GAT: std_logic; attribute dont_touch of N773GAT: signal is true;
	signal N774GAT: std_logic; attribute dont_touch of N774GAT: signal is true;
	signal N775GAT: std_logic; attribute dont_touch of N775GAT: signal is true;
	signal N776GAT: std_logic; attribute dont_touch of N776GAT: signal is true;
	signal N777GAT: std_logic; attribute dont_touch of N777GAT: signal is true;
	signal N779GAT: std_logic; attribute dont_touch of N779GAT: signal is true;
	signal N780GAT: std_logic; attribute dont_touch of N780GAT: signal is true;
	signal N781GAT: std_logic; attribute dont_touch of N781GAT: signal is true;
	signal N782GAT: std_logic; attribute dont_touch of N782GAT: signal is true;
	signal N783GAT: std_logic; attribute dont_touch of N783GAT: signal is true;
	signal N784GAT: std_logic; attribute dont_touch of N784GAT: signal is true;
	signal N785GAT: std_logic; attribute dont_touch of N785GAT: signal is true;
	signal N786GAT: std_logic; attribute dont_touch of N786GAT: signal is true;
	signal N787GAT: std_logic; attribute dont_touch of N787GAT: signal is true;
	signal N788GAT: std_logic; attribute dont_touch of N788GAT: signal is true;
	signal N789GAT: std_logic; attribute dont_touch of N789GAT: signal is true;
	signal N790GAT: std_logic; attribute dont_touch of N790GAT: signal is true;
	signal N791GAT: std_logic; attribute dont_touch of N791GAT: signal is true;
	signal N792GAT: std_logic; attribute dont_touch of N792GAT: signal is true;
	signal N793GAT: std_logic; attribute dont_touch of N793GAT: signal is true;
	signal N794GAT: std_logic; attribute dont_touch of N794GAT: signal is true;
	signal N795GAT: std_logic; attribute dont_touch of N795GAT: signal is true;
	signal N796GAT: std_logic; attribute dont_touch of N796GAT: signal is true;
	signal N797GAT: std_logic; attribute dont_touch of N797GAT: signal is true;
	signal N800GAT: std_logic; attribute dont_touch of N800GAT: signal is true;
	signal N801GAT: std_logic; attribute dont_touch of N801GAT: signal is true;
	signal N802GAT: std_logic; attribute dont_touch of N802GAT: signal is true;
	signal N803GAT: std_logic; attribute dont_touch of N803GAT: signal is true;
	signal N804GAT: std_logic; attribute dont_touch of N804GAT: signal is true;
	signal N805GAT: std_logic; attribute dont_touch of N805GAT: signal is true;
	signal N806GAT: std_logic; attribute dont_touch of N806GAT: signal is true;
	signal N807GAT: std_logic; attribute dont_touch of N807GAT: signal is true;
	signal N808GAT: std_logic; attribute dont_touch of N808GAT: signal is true;
	signal N809GAT: std_logic; attribute dont_touch of N809GAT: signal is true;
	signal N810GAT: std_logic; attribute dont_touch of N810GAT: signal is true;
	signal N811GAT: std_logic; attribute dont_touch of N811GAT: signal is true;
	signal N812GAT: std_logic; attribute dont_touch of N812GAT: signal is true;
	signal N813GAT: std_logic; attribute dont_touch of N813GAT: signal is true;
	signal N814GAT: std_logic; attribute dont_touch of N814GAT: signal is true;
	signal N815GAT: std_logic; attribute dont_touch of N815GAT: signal is true;
	signal N816GAT: std_logic; attribute dont_touch of N816GAT: signal is true;
	signal N818GAT: std_logic; attribute dont_touch of N818GAT: signal is true;
	signal N819GAT: std_logic; attribute dont_touch of N819GAT: signal is true;
	signal N820GAT: std_logic; attribute dont_touch of N820GAT: signal is true;
	signal N822GAT: std_logic; attribute dont_touch of N822GAT: signal is true;
	signal N823GAT: std_logic; attribute dont_touch of N823GAT: signal is true;
	signal N824GAT: std_logic; attribute dont_touch of N824GAT: signal is true;
	signal N827GAT: std_logic; attribute dont_touch of N827GAT: signal is true;
	signal N828GAT: std_logic; attribute dont_touch of N828GAT: signal is true;
	signal N829GAT: std_logic; attribute dont_touch of N829GAT: signal is true;
	signal N830GAT: std_logic; attribute dont_touch of N830GAT: signal is true;
	signal N832GAT: std_logic; attribute dont_touch of N832GAT: signal is true;
	signal N833GAT: std_logic; attribute dont_touch of N833GAT: signal is true;
	signal N834GAT: std_logic; attribute dont_touch of N834GAT: signal is true;
	signal N836GAT: std_logic; attribute dont_touch of N836GAT: signal is true;
	signal N837GAT: std_logic; attribute dont_touch of N837GAT: signal is true;
	signal N838GAT: std_logic; attribute dont_touch of N838GAT: signal is true;
	signal N840GAT: std_logic; attribute dont_touch of N840GAT: signal is true;
	signal N841GAT: std_logic; attribute dont_touch of N841GAT: signal is true;
	signal N842GAT: std_logic; attribute dont_touch of N842GAT: signal is true;
	signal N844GAT: std_logic; attribute dont_touch of N844GAT: signal is true;
	signal N845GAT: std_logic; attribute dont_touch of N845GAT: signal is true;
	signal N846GAT: std_logic; attribute dont_touch of N846GAT: signal is true;
	signal N848GAT: std_logic; attribute dont_touch of N848GAT: signal is true;
	signal N849GAT: std_logic; attribute dont_touch of N849GAT: signal is true;
	signal N850GAT: std_logic; attribute dont_touch of N850GAT: signal is true;
	signal N851GAT: std_logic; attribute dont_touch of N851GAT: signal is true;
	signal N852GAT: std_logic; attribute dont_touch of N852GAT: signal is true;
	signal N853GAT: std_logic; attribute dont_touch of N853GAT: signal is true;
	signal N854GAT: std_logic; attribute dont_touch of N854GAT: signal is true;
	signal N855GAT: std_logic; attribute dont_touch of N855GAT: signal is true;
	signal N856GAT: std_logic; attribute dont_touch of N856GAT: signal is true;
	signal N857GAT: std_logic; attribute dont_touch of N857GAT: signal is true;
	signal N858GAT: std_logic; attribute dont_touch of N858GAT: signal is true;
	signal N859GAT: std_logic; attribute dont_touch of N859GAT: signal is true;
	signal N860GAT: std_logic; attribute dont_touch of N860GAT: signal is true;
	signal N861GAT: std_logic; attribute dont_touch of N861GAT: signal is true;
	signal N863GAT: std_logic; attribute dont_touch of N863GAT: signal is true;
	signal N864GAT: std_logic; attribute dont_touch of N864GAT: signal is true;
	signal N865GAT: std_logic; attribute dont_touch of N865GAT: signal is true;
	signal N867GAT: std_logic; attribute dont_touch of N867GAT: signal is true;
	signal N868GAT: std_logic; attribute dont_touch of N868GAT: signal is true;
	signal N869GAT: std_logic; attribute dont_touch of N869GAT: signal is true;
	signal N870GAT: std_logic; attribute dont_touch of N870GAT: signal is true;
	signal N871GAT: std_logic; attribute dont_touch of N871GAT: signal is true;
	signal N872GAT: std_logic; attribute dont_touch of N872GAT: signal is true;
	signal N873GAT: std_logic; attribute dont_touch of N873GAT: signal is true;
	signal N874GAT: std_logic; attribute dont_touch of N874GAT: signal is true;
	signal N875GAT: std_logic; attribute dont_touch of N875GAT: signal is true;
	signal N876GAT: std_logic; attribute dont_touch of N876GAT: signal is true;
	signal N877GAT: std_logic; attribute dont_touch of N877GAT: signal is true;
	signal N878GAT: std_logic; attribute dont_touch of N878GAT: signal is true;
	signal N879GAT: std_logic; attribute dont_touch of N879GAT: signal is true;
	signal N880GAT: std_logic; attribute dont_touch of N880GAT: signal is true;
	signal N881GAT: std_logic; attribute dont_touch of N881GAT: signal is true;
	signal N882GAT: std_logic; attribute dont_touch of N882GAT: signal is true;
	signal N883GAT: std_logic; attribute dont_touch of N883GAT: signal is true;
	signal N885GAT: std_logic; attribute dont_touch of N885GAT: signal is true;
	signal N886GAT: std_logic; attribute dont_touch of N886GAT: signal is true;
	signal N887GAT: std_logic; attribute dont_touch of N887GAT: signal is true;
	signal N888GAT: std_logic; attribute dont_touch of N888GAT: signal is true;
	signal N889GAT: std_logic; attribute dont_touch of N889GAT: signal is true;
	signal N890GAT: std_logic; attribute dont_touch of N890GAT: signal is true;
	signal N891GAT: std_logic; attribute dont_touch of N891GAT: signal is true;
	signal N892GAT: std_logic; attribute dont_touch of N892GAT: signal is true;
	signal N893GAT: std_logic; attribute dont_touch of N893GAT: signal is true;
	signal N894GAT: std_logic; attribute dont_touch of N894GAT: signal is true;
	signal N895GAT: std_logic; attribute dont_touch of N895GAT: signal is true;
	signal N896GAT: std_logic; attribute dont_touch of N896GAT: signal is true;
	signal N897GAT: std_logic; attribute dont_touch of N897GAT: signal is true;
	signal N898GAT: std_logic; attribute dont_touch of N898GAT: signal is true;
	signal N899GAT: std_logic; attribute dont_touch of N899GAT: signal is true;
	signal N900GAT: std_logic; attribute dont_touch of N900GAT: signal is true;
	signal N901GAT: std_logic; attribute dont_touch of N901GAT: signal is true;
	signal N902GAT: std_logic; attribute dont_touch of N902GAT: signal is true;
	signal N903GAT: std_logic; attribute dont_touch of N903GAT: signal is true;
	signal N904GAT: std_logic; attribute dont_touch of N904GAT: signal is true;
	signal N905GAT: std_logic; attribute dont_touch of N905GAT: signal is true;
	signal N906GAT: std_logic; attribute dont_touch of N906GAT: signal is true;
	signal N907GAT: std_logic; attribute dont_touch of N907GAT: signal is true;
	signal N908GAT: std_logic; attribute dont_touch of N908GAT: signal is true;
	signal N909GAT: std_logic; attribute dont_touch of N909GAT: signal is true;
	signal N910GAT: std_logic; attribute dont_touch of N910GAT: signal is true;
	signal N911GAT: std_logic; attribute dont_touch of N911GAT: signal is true;
	signal N912GAT: std_logic; attribute dont_touch of N912GAT: signal is true;
	signal N913GAT: std_logic; attribute dont_touch of N913GAT: signal is true;
	signal N914GAT: std_logic; attribute dont_touch of N914GAT: signal is true;
	signal N915GAT: std_logic; attribute dont_touch of N915GAT: signal is true;
	signal N916GAT: std_logic; attribute dont_touch of N916GAT: signal is true;
	signal N917GAT: std_logic; attribute dont_touch of N917GAT: signal is true;
	signal N918GAT: std_logic; attribute dont_touch of N918GAT: signal is true;
	signal N919GAT: std_logic; attribute dont_touch of N919GAT: signal is true;
	signal N921GAT: std_logic; attribute dont_touch of N921GAT: signal is true;
	signal N922GAT: std_logic; attribute dont_touch of N922GAT: signal is true;
	signal N923GAT: std_logic; attribute dont_touch of N923GAT: signal is true;
	signal N924GAT: std_logic; attribute dont_touch of N924GAT: signal is true;
	signal N925GAT: std_logic; attribute dont_touch of N925GAT: signal is true;
	signal N926GAT: std_logic; attribute dont_touch of N926GAT: signal is true;
	signal N927GAT: std_logic; attribute dont_touch of N927GAT: signal is true;
	signal N928GAT: std_logic; attribute dont_touch of N928GAT: signal is true;
	signal N929GAT: std_logic; attribute dont_touch of N929GAT: signal is true;
	signal N930GAT: std_logic; attribute dont_touch of N930GAT: signal is true;
	signal N931GAT: std_logic; attribute dont_touch of N931GAT: signal is true;
	signal N933GAT: std_logic; attribute dont_touch of N933GAT: signal is true;
	signal N934GAT: std_logic; attribute dont_touch of N934GAT: signal is true;
	signal N935GAT: std_logic; attribute dont_touch of N935GAT: signal is true;
	signal N936GAT: std_logic; attribute dont_touch of N936GAT: signal is true;
	signal N937GAT: std_logic; attribute dont_touch of N937GAT: signal is true;
	signal N938GAT: std_logic; attribute dont_touch of N938GAT: signal is true;
	signal N939GAT: std_logic; attribute dont_touch of N939GAT: signal is true;
	signal N940GAT: std_logic; attribute dont_touch of N940GAT: signal is true;
	signal N941GAT: std_logic; attribute dont_touch of N941GAT: signal is true;
	signal N942GAT: std_logic; attribute dont_touch of N942GAT: signal is true;
	signal N943GAT: std_logic; attribute dont_touch of N943GAT: signal is true;
	signal N944GAT: std_logic; attribute dont_touch of N944GAT: signal is true;
	signal N945GAT: std_logic; attribute dont_touch of N945GAT: signal is true;
	signal N946GAT: std_logic; attribute dont_touch of N946GAT: signal is true;
	signal N947GAT: std_logic; attribute dont_touch of N947GAT: signal is true;
	signal N948GAT: std_logic; attribute dont_touch of N948GAT: signal is true;
	signal N949GAT: std_logic; attribute dont_touch of N949GAT: signal is true;
	signal N950GAT: std_logic; attribute dont_touch of N950GAT: signal is true;
	signal N951GAT: std_logic; attribute dont_touch of N951GAT: signal is true;
	signal N952GAT: std_logic; attribute dont_touch of N952GAT: signal is true;
	signal N953GAT: std_logic; attribute dont_touch of N953GAT: signal is true;
	signal N954GAT: std_logic; attribute dont_touch of N954GAT: signal is true;
	signal N955GAT: std_logic; attribute dont_touch of N955GAT: signal is true;
	signal N956GAT: std_logic; attribute dont_touch of N956GAT: signal is true;
	signal N957GAT: std_logic; attribute dont_touch of N957GAT: signal is true;
	signal N959GAT: std_logic; attribute dont_touch of N959GAT: signal is true;
	signal N960GAT: std_logic; attribute dont_touch of N960GAT: signal is true;
	signal N961GAT: std_logic; attribute dont_touch of N961GAT: signal is true;
	signal N962GAT: std_logic; attribute dont_touch of N962GAT: signal is true;
	signal N963GAT: std_logic; attribute dont_touch of N963GAT: signal is true;
	signal N964GAT: std_logic; attribute dont_touch of N964GAT: signal is true;
	signal N965GAT: std_logic; attribute dont_touch of N965GAT: signal is true;
	signal N966GAT: std_logic; attribute dont_touch of N966GAT: signal is true;
	signal N967GAT: std_logic; attribute dont_touch of N967GAT: signal is true;
	signal N968GAT: std_logic; attribute dont_touch of N968GAT: signal is true;
	signal N969GAT: std_logic; attribute dont_touch of N969GAT: signal is true;
	signal N970GAT: std_logic; attribute dont_touch of N970GAT: signal is true;
	signal N971GAT: std_logic; attribute dont_touch of N971GAT: signal is true;
	signal N972GAT: std_logic; attribute dont_touch of N972GAT: signal is true;
	signal N973GAT: std_logic; attribute dont_touch of N973GAT: signal is true;
	signal N974GAT: std_logic; attribute dont_touch of N974GAT: signal is true;
	signal N975GAT: std_logic; attribute dont_touch of N975GAT: signal is true;
	signal N976GAT: std_logic; attribute dont_touch of N976GAT: signal is true;
	signal N977GAT: std_logic; attribute dont_touch of N977GAT: signal is true;
	signal N978GAT: std_logic; attribute dont_touch of N978GAT: signal is true;
	signal N979GAT: std_logic; attribute dont_touch of N979GAT: signal is true;
	signal N980GAT: std_logic; attribute dont_touch of N980GAT: signal is true;
	signal N981GAT: std_logic; attribute dont_touch of N981GAT: signal is true;
	signal N982GAT: std_logic; attribute dont_touch of N982GAT: signal is true;
	signal N983GAT: std_logic; attribute dont_touch of N983GAT: signal is true;
	signal N984GAT: std_logic; attribute dont_touch of N984GAT: signal is true;
	signal N985GAT: std_logic; attribute dont_touch of N985GAT: signal is true;
	signal N986GAT: std_logic; attribute dont_touch of N986GAT: signal is true;
	signal N987GAT: std_logic; attribute dont_touch of N987GAT: signal is true;
	signal N988GAT: std_logic; attribute dont_touch of N988GAT: signal is true;
	signal N989GAT: std_logic; attribute dont_touch of N989GAT: signal is true;
	signal N990GAT: std_logic; attribute dont_touch of N990GAT: signal is true;
	signal N991GAT: std_logic; attribute dont_touch of N991GAT: signal is true;
	signal N992GAT: std_logic; attribute dont_touch of N992GAT: signal is true;
	signal N993GAT: std_logic; attribute dont_touch of N993GAT: signal is true;
	signal N994GAT: std_logic; attribute dont_touch of N994GAT: signal is true;
	signal N995GAT: std_logic; attribute dont_touch of N995GAT: signal is true;
	signal N996GAT: std_logic; attribute dont_touch of N996GAT: signal is true;
	signal N997GAT: std_logic; attribute dont_touch of N997GAT: signal is true;
	signal N998GAT: std_logic; attribute dont_touch of N998GAT: signal is true;
	signal N999GAT: std_logic; attribute dont_touch of N999GAT: signal is true;
	signal N1000GAT: std_logic; attribute dont_touch of N1000GAT: signal is true;
	signal N1001GAT: std_logic; attribute dont_touch of N1001GAT: signal is true;
	signal N1002GAT: std_logic; attribute dont_touch of N1002GAT: signal is true;
	signal N1003GAT: std_logic; attribute dont_touch of N1003GAT: signal is true;
	signal N1004GAT: std_logic; attribute dont_touch of N1004GAT: signal is true;
	signal N1005GAT: std_logic; attribute dont_touch of N1005GAT: signal is true;
	signal N1006GAT: std_logic; attribute dont_touch of N1006GAT: signal is true;
	signal N1007GAT: std_logic; attribute dont_touch of N1007GAT: signal is true;
	signal N1008GAT: std_logic; attribute dont_touch of N1008GAT: signal is true;
	signal N1009GAT: std_logic; attribute dont_touch of N1009GAT: signal is true;
	signal N1010GAT: std_logic; attribute dont_touch of N1010GAT: signal is true;
	signal N1011GAT: std_logic; attribute dont_touch of N1011GAT: signal is true;
	signal N1012GAT: std_logic; attribute dont_touch of N1012GAT: signal is true;
	signal N1013GAT: std_logic; attribute dont_touch of N1013GAT: signal is true;
	signal N1014GAT: std_logic; attribute dont_touch of N1014GAT: signal is true;
	signal N1015GAT: std_logic; attribute dont_touch of N1015GAT: signal is true;
	signal N1016GAT: std_logic; attribute dont_touch of N1016GAT: signal is true;
	signal N1017GAT: std_logic; attribute dont_touch of N1017GAT: signal is true;
	signal N1018GAT: std_logic; attribute dont_touch of N1018GAT: signal is true;
	signal N1019GAT: std_logic; attribute dont_touch of N1019GAT: signal is true;
	signal N1020GAT: std_logic; attribute dont_touch of N1020GAT: signal is true;
	signal N1021GAT: std_logic; attribute dont_touch of N1021GAT: signal is true;
	signal N1022GAT: std_logic; attribute dont_touch of N1022GAT: signal is true;
	signal N1023GAT: std_logic; attribute dont_touch of N1023GAT: signal is true;
	signal N1024GAT: std_logic; attribute dont_touch of N1024GAT: signal is true;
	signal N1025GAT: std_logic; attribute dont_touch of N1025GAT: signal is true;
	signal N1026GAT: std_logic; attribute dont_touch of N1026GAT: signal is true;
	signal N1028GAT: std_logic; attribute dont_touch of N1028GAT: signal is true;
	signal N1029GAT: std_logic; attribute dont_touch of N1029GAT: signal is true;
	signal N1030GAT: std_logic; attribute dont_touch of N1030GAT: signal is true;
	signal N1031GAT: std_logic; attribute dont_touch of N1031GAT: signal is true;
	signal N1032GAT: std_logic; attribute dont_touch of N1032GAT: signal is true;
	signal N1033GAT: std_logic; attribute dont_touch of N1033GAT: signal is true;
	signal N1034GAT: std_logic; attribute dont_touch of N1034GAT: signal is true;
	signal N1035GAT: std_logic; attribute dont_touch of N1035GAT: signal is true;
	signal N1043GAT: std_logic; attribute dont_touch of N1043GAT: signal is true;
	signal N1044GAT: std_logic; attribute dont_touch of N1044GAT: signal is true;
	signal N1045GAT: std_logic; attribute dont_touch of N1045GAT: signal is true;
	signal N1050GAT: std_logic; attribute dont_touch of N1050GAT: signal is true;
	signal N1051GAT: std_logic; attribute dont_touch of N1051GAT: signal is true;
	signal N1052GAT: std_logic; attribute dont_touch of N1052GAT: signal is true;
	signal N1053GAT: std_logic; attribute dont_touch of N1053GAT: signal is true;
	signal N1054GAT: std_logic; attribute dont_touch of N1054GAT: signal is true;
	signal N1055GAT: std_logic; attribute dont_touch of N1055GAT: signal is true;
	signal N1056GAT: std_logic; attribute dont_touch of N1056GAT: signal is true;
	signal N1057GAT: std_logic; attribute dont_touch of N1057GAT: signal is true;
	signal N1058GAT: std_logic; attribute dont_touch of N1058GAT: signal is true;
	signal N1059GAT: std_logic; attribute dont_touch of N1059GAT: signal is true;
	signal N1060GAT: std_logic; attribute dont_touch of N1060GAT: signal is true;
	signal N1066GAT: std_logic; attribute dont_touch of N1066GAT: signal is true;
	signal N1067GAT: std_logic; attribute dont_touch of N1067GAT: signal is true;
	signal N1068GAT: std_logic; attribute dont_touch of N1068GAT: signal is true;
	signal N1070GAT: std_logic; attribute dont_touch of N1070GAT: signal is true;
	signal N1071GAT: std_logic; attribute dont_touch of N1071GAT: signal is true;
	signal N1072GAT: std_logic; attribute dont_touch of N1072GAT: signal is true;
	signal N1074GAT: std_logic; attribute dont_touch of N1074GAT: signal is true;
	signal N1075GAT: std_logic; attribute dont_touch of N1075GAT: signal is true;
	signal N1076GAT: std_logic; attribute dont_touch of N1076GAT: signal is true;
	signal N1077GAT: std_logic; attribute dont_touch of N1077GAT: signal is true;
	signal N1078GAT: std_logic; attribute dont_touch of N1078GAT: signal is true;
	signal N1079GAT: std_logic; attribute dont_touch of N1079GAT: signal is true;
	signal N1080GAT: std_logic; attribute dont_touch of N1080GAT: signal is true;
	signal N1082GAT: std_logic; attribute dont_touch of N1082GAT: signal is true;
	signal N1083GAT: std_logic; attribute dont_touch of N1083GAT: signal is true;
	signal N1084GAT: std_logic; attribute dont_touch of N1084GAT: signal is true;
	signal N1085GAT: std_logic; attribute dont_touch of N1085GAT: signal is true;
	signal N1086GAT: std_logic; attribute dont_touch of N1086GAT: signal is true;
	signal N1087GAT: std_logic; attribute dont_touch of N1087GAT: signal is true;
	signal N1088GAT: std_logic; attribute dont_touch of N1088GAT: signal is true;
	signal N1089GAT: std_logic; attribute dont_touch of N1089GAT: signal is true;
	signal N1090GAT: std_logic; attribute dont_touch of N1090GAT: signal is true;
	signal N1091GAT: std_logic; attribute dont_touch of N1091GAT: signal is true;
	signal N1092GAT: std_logic; attribute dont_touch of N1092GAT: signal is true;
	signal N1093GAT: std_logic; attribute dont_touch of N1093GAT: signal is true;
	signal N1094GAT: std_logic; attribute dont_touch of N1094GAT: signal is true;
	signal N1095GAT: std_logic; attribute dont_touch of N1095GAT: signal is true;
	signal N1096GAT: std_logic; attribute dont_touch of N1096GAT: signal is true;
	signal N1097GAT: std_logic; attribute dont_touch of N1097GAT: signal is true;
	signal N1098GAT: std_logic; attribute dont_touch of N1098GAT: signal is true;
	signal N1099GAT: std_logic; attribute dont_touch of N1099GAT: signal is true;
	signal N1100GAT: std_logic; attribute dont_touch of N1100GAT: signal is true;
	signal N1101GAT: std_logic; attribute dont_touch of N1101GAT: signal is true;
	signal N1102GAT: std_logic; attribute dont_touch of N1102GAT: signal is true;
	signal N1103GAT: std_logic; attribute dont_touch of N1103GAT: signal is true;
	signal N1104GAT: std_logic; attribute dont_touch of N1104GAT: signal is true;
	signal N1105GAT: std_logic; attribute dont_touch of N1105GAT: signal is true;
	signal N1106GAT: std_logic; attribute dont_touch of N1106GAT: signal is true;
	signal N1111GAT: std_logic; attribute dont_touch of N1111GAT: signal is true;
	signal N1112GAT: std_logic; attribute dont_touch of N1112GAT: signal is true;
	signal N1113GAT: std_logic; attribute dont_touch of N1113GAT: signal is true;
	signal N1114GAT: std_logic; attribute dont_touch of N1114GAT: signal is true;
	signal N1115GAT: std_logic; attribute dont_touch of N1115GAT: signal is true;
	signal N1116GAT: std_logic; attribute dont_touch of N1116GAT: signal is true;
	signal N1117GAT: std_logic; attribute dont_touch of N1117GAT: signal is true;
	signal N1118GAT: std_logic; attribute dont_touch of N1118GAT: signal is true;
	signal N1119GAT: std_logic; attribute dont_touch of N1119GAT: signal is true;
	signal N1120GAT: std_logic; attribute dont_touch of N1120GAT: signal is true;
	signal N1121GAT: std_logic; attribute dont_touch of N1121GAT: signal is true;
	signal N1123GAT: std_logic; attribute dont_touch of N1123GAT: signal is true;
	signal N1133GAT: std_logic; attribute dont_touch of N1133GAT: signal is true;
	signal N1134GAT: std_logic; attribute dont_touch of N1134GAT: signal is true;
	signal N1135GAT: std_logic; attribute dont_touch of N1135GAT: signal is true;
	signal N1146GAT: std_logic; attribute dont_touch of N1146GAT: signal is true;
	signal N1147GAT: std_logic; attribute dont_touch of N1147GAT: signal is true;
	signal N1148GAT: std_logic; attribute dont_touch of N1148GAT: signal is true;
	signal N1150GAT: std_logic; attribute dont_touch of N1150GAT: signal is true;
	signal N1151GAT: std_logic; attribute dont_touch of N1151GAT: signal is true;
	signal N1152GAT: std_logic; attribute dont_touch of N1152GAT: signal is true;
	signal N1153GAT: std_logic; attribute dont_touch of N1153GAT: signal is true;
	signal N1154GAT: std_logic; attribute dont_touch of N1154GAT: signal is true;
	signal N1155GAT: std_logic; attribute dont_touch of N1155GAT: signal is true;
	signal N1156GAT: std_logic; attribute dont_touch of N1156GAT: signal is true;
	signal N1157GAT: std_logic; attribute dont_touch of N1157GAT: signal is true;
	signal N1158GAT: std_logic; attribute dont_touch of N1158GAT: signal is true;
	signal N1159GAT: std_logic; attribute dont_touch of N1159GAT: signal is true;
	signal N1160GAT: std_logic; attribute dont_touch of N1160GAT: signal is true;
	signal N1161GAT: std_logic; attribute dont_touch of N1161GAT: signal is true;
	signal N1162GAT: std_logic; attribute dont_touch of N1162GAT: signal is true;
	signal N1163GAT: std_logic; attribute dont_touch of N1163GAT: signal is true;
	signal N1164GAT: std_logic; attribute dont_touch of N1164GAT: signal is true;
	signal N1171GAT: std_logic; attribute dont_touch of N1171GAT: signal is true;
	signal N1172GAT: std_logic; attribute dont_touch of N1172GAT: signal is true;
	signal N1173GAT: std_logic; attribute dont_touch of N1173GAT: signal is true;
	signal N1174GAT: std_logic; attribute dont_touch of N1174GAT: signal is true;
	signal N1175GAT: std_logic; attribute dont_touch of N1175GAT: signal is true;
	signal N1176GAT: std_logic; attribute dont_touch of N1176GAT: signal is true;
	signal N1177GAT: std_logic; attribute dont_touch of N1177GAT: signal is true;
	signal N1178GAT: std_logic; attribute dont_touch of N1178GAT: signal is true;
	signal N1179GAT: std_logic; attribute dont_touch of N1179GAT: signal is true;
	signal N1180GAT: std_logic; attribute dont_touch of N1180GAT: signal is true;
	signal N1181GAT: std_logic; attribute dont_touch of N1181GAT: signal is true;
	signal N1182GAT: std_logic; attribute dont_touch of N1182GAT: signal is true;
	signal N1183GAT: std_logic; attribute dont_touch of N1183GAT: signal is true;
	signal N1184GAT: std_logic; attribute dont_touch of N1184GAT: signal is true;
	signal N1185GAT: std_logic; attribute dont_touch of N1185GAT: signal is true;
	signal N1186GAT: std_logic; attribute dont_touch of N1186GAT: signal is true;
	signal N1187GAT: std_logic; attribute dont_touch of N1187GAT: signal is true;
	signal N1188GAT: std_logic; attribute dont_touch of N1188GAT: signal is true;
	signal N1189GAT: std_logic; attribute dont_touch of N1189GAT: signal is true;
	signal N1190GAT: std_logic; attribute dont_touch of N1190GAT: signal is true;
	signal N1191GAT: std_logic; attribute dont_touch of N1191GAT: signal is true;
	signal N1192GAT: std_logic; attribute dont_touch of N1192GAT: signal is true;
	signal N1193GAT: std_logic; attribute dont_touch of N1193GAT: signal is true;
	signal N1194GAT: std_logic; attribute dont_touch of N1194GAT: signal is true;
	signal N1195GAT: std_logic; attribute dont_touch of N1195GAT: signal is true;
	signal N1196GAT: std_logic; attribute dont_touch of N1196GAT: signal is true;
	signal N1197GAT: std_logic; attribute dont_touch of N1197GAT: signal is true;
	signal N1199GAT: std_logic; attribute dont_touch of N1199GAT: signal is true;
	signal N1200GAT: std_logic; attribute dont_touch of N1200GAT: signal is true;
	signal N1201GAT: std_logic; attribute dont_touch of N1201GAT: signal is true;
	signal N1202GAT: std_logic; attribute dont_touch of N1202GAT: signal is true;
	signal N1203GAT: std_logic; attribute dont_touch of N1203GAT: signal is true;
	signal N1204GAT: std_logic; attribute dont_touch of N1204GAT: signal is true;
	signal N1205GAT: std_logic; attribute dont_touch of N1205GAT: signal is true;
	signal N1206GAT: std_logic; attribute dont_touch of N1206GAT: signal is true;
	signal N1207GAT: std_logic; attribute dont_touch of N1207GAT: signal is true;
	signal N1208GAT: std_logic; attribute dont_touch of N1208GAT: signal is true;
	signal N1209GAT: std_logic; attribute dont_touch of N1209GAT: signal is true;
	signal N1210GAT: std_logic; attribute dont_touch of N1210GAT: signal is true;
	signal N1211GAT: std_logic; attribute dont_touch of N1211GAT: signal is true;
	signal N1212GAT: std_logic; attribute dont_touch of N1212GAT: signal is true;
	signal N1213GAT: std_logic; attribute dont_touch of N1213GAT: signal is true;
	signal N1214GAT: std_logic; attribute dont_touch of N1214GAT: signal is true;
	signal N1215GAT: std_logic; attribute dont_touch of N1215GAT: signal is true;
	signal N1216GAT: std_logic; attribute dont_touch of N1216GAT: signal is true;
	signal N1217GAT: std_logic; attribute dont_touch of N1217GAT: signal is true;
	signal N1218GAT: std_logic; attribute dont_touch of N1218GAT: signal is true;
	signal N1219GAT: std_logic; attribute dont_touch of N1219GAT: signal is true;
	signal N1220GAT: std_logic; attribute dont_touch of N1220GAT: signal is true;
	signal N1221GAT: std_logic; attribute dont_touch of N1221GAT: signal is true;
	signal N1222GAT: std_logic; attribute dont_touch of N1222GAT: signal is true;
	signal N1223GAT: std_logic; attribute dont_touch of N1223GAT: signal is true;
	signal N1224GAT: std_logic; attribute dont_touch of N1224GAT: signal is true;
	signal N1225GAT: std_logic; attribute dont_touch of N1225GAT: signal is true;
	signal N1226GAT: std_logic; attribute dont_touch of N1226GAT: signal is true;
	signal N1228GAT: std_logic; attribute dont_touch of N1228GAT: signal is true;
	signal N1229GAT: std_logic; attribute dont_touch of N1229GAT: signal is true;
	signal N1230GAT: std_logic; attribute dont_touch of N1230GAT: signal is true;
	signal N1231GAT: std_logic; attribute dont_touch of N1231GAT: signal is true;
	signal N1232GAT: std_logic; attribute dont_touch of N1232GAT: signal is true;
	signal N1233GAT: std_logic; attribute dont_touch of N1233GAT: signal is true;
	signal N1234GAT: std_logic; attribute dont_touch of N1234GAT: signal is true;
	signal N1235GAT: std_logic; attribute dont_touch of N1235GAT: signal is true;
	signal N1236GAT: std_logic; attribute dont_touch of N1236GAT: signal is true;
	signal N1237GAT: std_logic; attribute dont_touch of N1237GAT: signal is true;
	signal N1238GAT: std_logic; attribute dont_touch of N1238GAT: signal is true;
	signal N1239GAT: std_logic; attribute dont_touch of N1239GAT: signal is true;
	signal N1240GAT: std_logic; attribute dont_touch of N1240GAT: signal is true;
	signal N1241GAT: std_logic; attribute dont_touch of N1241GAT: signal is true;
	signal N1243GAT: std_logic; attribute dont_touch of N1243GAT: signal is true;
	signal N1244GAT: std_logic; attribute dont_touch of N1244GAT: signal is true;
	signal N1245GAT: std_logic; attribute dont_touch of N1245GAT: signal is true;
	signal N1246GAT: std_logic; attribute dont_touch of N1246GAT: signal is true;
	signal N1247GAT: std_logic; attribute dont_touch of N1247GAT: signal is true;
	signal N1248GAT: std_logic; attribute dont_touch of N1248GAT: signal is true;
	signal N1249GAT: std_logic; attribute dont_touch of N1249GAT: signal is true;
	signal N1250GAT: std_logic; attribute dont_touch of N1250GAT: signal is true;
	signal N1251GAT: std_logic; attribute dont_touch of N1251GAT: signal is true;
	signal N1252GAT: std_logic; attribute dont_touch of N1252GAT: signal is true;
	signal N1253GAT: std_logic; attribute dont_touch of N1253GAT: signal is true;
	signal N1254GAT: std_logic; attribute dont_touch of N1254GAT: signal is true;
	signal N1255GAT: std_logic; attribute dont_touch of N1255GAT: signal is true;
	signal N1256GAT: std_logic; attribute dont_touch of N1256GAT: signal is true;
	signal N1257GAT: std_logic; attribute dont_touch of N1257GAT: signal is true;
	signal N1258GAT: std_logic; attribute dont_touch of N1258GAT: signal is true;
	signal N1259GAT: std_logic; attribute dont_touch of N1259GAT: signal is true;
	signal N1260GAT: std_logic; attribute dont_touch of N1260GAT: signal is true;
	signal N1261GAT: std_logic; attribute dont_touch of N1261GAT: signal is true;
	signal N1262GAT: std_logic; attribute dont_touch of N1262GAT: signal is true;
	signal N1263GAT: std_logic; attribute dont_touch of N1263GAT: signal is true;
	signal N1264GAT: std_logic; attribute dont_touch of N1264GAT: signal is true;
	signal N1265GAT: std_logic; attribute dont_touch of N1265GAT: signal is true;
	signal N1266GAT: std_logic; attribute dont_touch of N1266GAT: signal is true;
	signal N1267GAT: std_logic; attribute dont_touch of N1267GAT: signal is true;
	signal N1268GAT: std_logic; attribute dont_touch of N1268GAT: signal is true;
	signal N1269GAT: std_logic; attribute dont_touch of N1269GAT: signal is true;
	signal N1270GAT: std_logic; attribute dont_touch of N1270GAT: signal is true;
	signal N1271GAT: std_logic; attribute dont_touch of N1271GAT: signal is true;
	signal N1272GAT: std_logic; attribute dont_touch of N1272GAT: signal is true;
	signal N1273GAT: std_logic; attribute dont_touch of N1273GAT: signal is true;
	signal N1274GAT: std_logic; attribute dont_touch of N1274GAT: signal is true;
	signal N1275GAT: std_logic; attribute dont_touch of N1275GAT: signal is true;
	signal N1276GAT: std_logic; attribute dont_touch of N1276GAT: signal is true;
	signal N1277GAT: std_logic; attribute dont_touch of N1277GAT: signal is true;
	signal N1278GAT: std_logic; attribute dont_touch of N1278GAT: signal is true;
	signal N1279GAT: std_logic; attribute dont_touch of N1279GAT: signal is true;
	signal N1280GAT: std_logic; attribute dont_touch of N1280GAT: signal is true;
	signal N1281GAT: std_logic; attribute dont_touch of N1281GAT: signal is true;
	signal N1282GAT: std_logic; attribute dont_touch of N1282GAT: signal is true;
	signal N1284GAT: std_logic; attribute dont_touch of N1284GAT: signal is true;
	signal N1285GAT: std_logic; attribute dont_touch of N1285GAT: signal is true;
	signal N1286GAT: std_logic; attribute dont_touch of N1286GAT: signal is true;
	signal N1287GAT: std_logic; attribute dont_touch of N1287GAT: signal is true;
	signal N1291GAT: std_logic; attribute dont_touch of N1291GAT: signal is true;
	signal N1292GAT: std_logic; attribute dont_touch of N1292GAT: signal is true;
	signal N1293GAT: std_logic; attribute dont_touch of N1293GAT: signal is true;
	signal N1294GAT: std_logic; attribute dont_touch of N1294GAT: signal is true;
	signal N1296GAT: std_logic; attribute dont_touch of N1296GAT: signal is true;
	signal N1297GAT: std_logic; attribute dont_touch of N1297GAT: signal is true;
	signal N1298GAT: std_logic; attribute dont_touch of N1298GAT: signal is true;
	signal N1300GAT: std_logic; attribute dont_touch of N1300GAT: signal is true;
	signal N1301GAT: std_logic; attribute dont_touch of N1301GAT: signal is true;
	signal N1302GAT: std_logic; attribute dont_touch of N1302GAT: signal is true;
	signal N1303GAT: std_logic; attribute dont_touch of N1303GAT: signal is true;
	signal N1304GAT: std_logic; attribute dont_touch of N1304GAT: signal is true;
	signal N1305GAT: std_logic; attribute dont_touch of N1305GAT: signal is true;
	signal N1306GAT: std_logic; attribute dont_touch of N1306GAT: signal is true;
	signal N1307GAT: std_logic; attribute dont_touch of N1307GAT: signal is true;
	signal N1308GAT: std_logic; attribute dont_touch of N1308GAT: signal is true;
	signal N1309GAT: std_logic; attribute dont_touch of N1309GAT: signal is true;
	signal N1310GAT: std_logic; attribute dont_touch of N1310GAT: signal is true;
	signal N1311GAT: std_logic; attribute dont_touch of N1311GAT: signal is true;
	signal N1312GAT: std_logic; attribute dont_touch of N1312GAT: signal is true;
	signal N1314GAT: std_logic; attribute dont_touch of N1314GAT: signal is true;
	signal N1315GAT: std_logic; attribute dont_touch of N1315GAT: signal is true;
	signal N1316GAT: std_logic; attribute dont_touch of N1316GAT: signal is true;
	signal N1318GAT: std_logic; attribute dont_touch of N1318GAT: signal is true;
	signal N1319GAT: std_logic; attribute dont_touch of N1319GAT: signal is true;
	signal N1320GAT: std_logic; attribute dont_touch of N1320GAT: signal is true;
	signal N1321GAT: std_logic; attribute dont_touch of N1321GAT: signal is true;
	signal N1322GAT: std_logic; attribute dont_touch of N1322GAT: signal is true;
	signal N1323GAT: std_logic; attribute dont_touch of N1323GAT: signal is true;
	signal N1324GAT: std_logic; attribute dont_touch of N1324GAT: signal is true;
	signal N1325GAT: std_logic; attribute dont_touch of N1325GAT: signal is true;
	signal N1326GAT: std_logic; attribute dont_touch of N1326GAT: signal is true;
	signal N1327GAT: std_logic; attribute dont_touch of N1327GAT: signal is true;
	signal N1328GAT: std_logic; attribute dont_touch of N1328GAT: signal is true;
	signal N1329GAT: std_logic; attribute dont_touch of N1329GAT: signal is true;
	signal N1330GAT: std_logic; attribute dont_touch of N1330GAT: signal is true;
	signal N1332GAT: std_logic; attribute dont_touch of N1332GAT: signal is true;
	signal N1334GAT: std_logic; attribute dont_touch of N1334GAT: signal is true;
	signal N1336GAT: std_logic; attribute dont_touch of N1336GAT: signal is true;
	signal N1338GAT: std_logic; attribute dont_touch of N1338GAT: signal is true;
	signal N1339GAT: std_logic; attribute dont_touch of N1339GAT: signal is true;
	signal N1340GAT: std_logic; attribute dont_touch of N1340GAT: signal is true;
	signal N1347GAT: std_logic; attribute dont_touch of N1347GAT: signal is true;
	signal N1348GAT: std_logic; attribute dont_touch of N1348GAT: signal is true;
	signal N1349GAT: std_logic; attribute dont_touch of N1349GAT: signal is true;
	signal N1350GAT: std_logic; attribute dont_touch of N1350GAT: signal is true;
	signal N1351GAT: std_logic; attribute dont_touch of N1351GAT: signal is true;
	signal N1352GAT: std_logic; attribute dont_touch of N1352GAT: signal is true;
	signal N1353GAT: std_logic; attribute dont_touch of N1353GAT: signal is true;
	signal N1354GAT: std_logic; attribute dont_touch of N1354GAT: signal is true;
	signal N1355GAT: std_logic; attribute dont_touch of N1355GAT: signal is true;
	signal N1356GAT: std_logic; attribute dont_touch of N1356GAT: signal is true;
	signal N1357GAT: std_logic; attribute dont_touch of N1357GAT: signal is true;
	signal N1358GAT: std_logic; attribute dont_touch of N1358GAT: signal is true;
	signal N1359GAT: std_logic; attribute dont_touch of N1359GAT: signal is true;
	signal N1360GAT: std_logic; attribute dont_touch of N1360GAT: signal is true;
	signal N1361GAT: std_logic; attribute dont_touch of N1361GAT: signal is true;
	signal N1363GAT: std_logic; attribute dont_touch of N1363GAT: signal is true;
	signal N1365GAT: std_logic; attribute dont_touch of N1365GAT: signal is true;
	signal N1366GAT: std_logic; attribute dont_touch of N1366GAT: signal is true;
	signal N1367GAT: std_logic; attribute dont_touch of N1367GAT: signal is true;
	signal N1368GAT: std_logic; attribute dont_touch of N1368GAT: signal is true;
	signal N1369GAT: std_logic; attribute dont_touch of N1369GAT: signal is true;
	signal N1370GAT: std_logic; attribute dont_touch of N1370GAT: signal is true;
	signal N1371GAT: std_logic; attribute dont_touch of N1371GAT: signal is true;
	signal N1372GAT: std_logic; attribute dont_touch of N1372GAT: signal is true;
	signal N1373GAT: std_logic; attribute dont_touch of N1373GAT: signal is true;
	signal N1374GAT: std_logic; attribute dont_touch of N1374GAT: signal is true;
	signal N1375GAT: std_logic; attribute dont_touch of N1375GAT: signal is true;
	signal N1376GAT: std_logic; attribute dont_touch of N1376GAT: signal is true;
	signal N1377GAT: std_logic; attribute dont_touch of N1377GAT: signal is true;
	signal N1378GAT: std_logic; attribute dont_touch of N1378GAT: signal is true;
	signal N1379GAT: std_logic; attribute dont_touch of N1379GAT: signal is true;
	signal N1380GAT: std_logic; attribute dont_touch of N1380GAT: signal is true;
	signal N1381GAT: std_logic; attribute dont_touch of N1381GAT: signal is true;
	signal N1382GAT: std_logic; attribute dont_touch of N1382GAT: signal is true;
	signal N1383GAT: std_logic; attribute dont_touch of N1383GAT: signal is true;
	signal N1384GAT: std_logic; attribute dont_touch of N1384GAT: signal is true;
	signal N1387GAT: std_logic; attribute dont_touch of N1387GAT: signal is true;
	signal N1389GAT: std_logic; attribute dont_touch of N1389GAT: signal is true;
	signal N1391GAT: std_logic; attribute dont_touch of N1391GAT: signal is true;
	signal N1392GAT: std_logic; attribute dont_touch of N1392GAT: signal is true;
	signal N1393GAT: std_logic; attribute dont_touch of N1393GAT: signal is true;
	signal N1394GAT: std_logic; attribute dont_touch of N1394GAT: signal is true;
	signal N1396GAT: std_logic; attribute dont_touch of N1396GAT: signal is true;
	signal N1397GAT: std_logic; attribute dont_touch of N1397GAT: signal is true;
	signal N1398GAT: std_logic; attribute dont_touch of N1398GAT: signal is true;
	signal N1399GAT: std_logic; attribute dont_touch of N1399GAT: signal is true;
	signal N1400GAT: std_logic; attribute dont_touch of N1400GAT: signal is true;
	signal N1401GAT: std_logic; attribute dont_touch of N1401GAT: signal is true;
	signal N1402GAT: std_logic; attribute dont_touch of N1402GAT: signal is true;
	signal N1403GAT: std_logic; attribute dont_touch of N1403GAT: signal is true;
	signal N1406GAT: std_logic; attribute dont_touch of N1406GAT: signal is true;
	signal N1407GAT: std_logic; attribute dont_touch of N1407GAT: signal is true;
	signal N1408GAT: std_logic; attribute dont_touch of N1408GAT: signal is true;
	signal N1409GAT: std_logic; attribute dont_touch of N1409GAT: signal is true;
	signal N1410GAT: std_logic; attribute dont_touch of N1410GAT: signal is true;
	signal N1411GAT: std_logic; attribute dont_touch of N1411GAT: signal is true;
	signal N1412GAT: std_logic; attribute dont_touch of N1412GAT: signal is true;
	signal N1413GAT: std_logic; attribute dont_touch of N1413GAT: signal is true;
	signal N1414GAT: std_logic; attribute dont_touch of N1414GAT: signal is true;
	signal N1415GAT: std_logic; attribute dont_touch of N1415GAT: signal is true;
	signal N1416GAT: std_logic; attribute dont_touch of N1416GAT: signal is true;
	signal N1417GAT: std_logic; attribute dont_touch of N1417GAT: signal is true;
	signal N1418GAT: std_logic; attribute dont_touch of N1418GAT: signal is true;
	signal N1419GAT: std_logic; attribute dont_touch of N1419GAT: signal is true;
	signal N1420GAT: std_logic; attribute dont_touch of N1420GAT: signal is true;
	signal N1421GAT: std_logic; attribute dont_touch of N1421GAT: signal is true;
	signal N1422GAT: std_logic; attribute dont_touch of N1422GAT: signal is true;
	signal N1423GAT: std_logic; attribute dont_touch of N1423GAT: signal is true;
	signal N1424GAT: std_logic; attribute dont_touch of N1424GAT: signal is true;
	signal N1425GAT: std_logic; attribute dont_touch of N1425GAT: signal is true;
	signal N1426GAT: std_logic; attribute dont_touch of N1426GAT: signal is true;
	signal N1427GAT: std_logic; attribute dont_touch of N1427GAT: signal is true;
	signal N1428GAT: std_logic; attribute dont_touch of N1428GAT: signal is true;
	signal N1430GAT: std_logic; attribute dont_touch of N1430GAT: signal is true;
	signal N1431GAT: std_logic; attribute dont_touch of N1431GAT: signal is true;
	signal N1433GAT: std_logic; attribute dont_touch of N1433GAT: signal is true;
	signal N1435GAT: std_logic; attribute dont_touch of N1435GAT: signal is true;
	signal N1436GAT: std_logic; attribute dont_touch of N1436GAT: signal is true;
	signal N1437GAT: std_logic; attribute dont_touch of N1437GAT: signal is true;
	signal N1438GAT: std_logic; attribute dont_touch of N1438GAT: signal is true;
	signal N1439GAT: std_logic; attribute dont_touch of N1439GAT: signal is true;
	signal N1440GAT: std_logic; attribute dont_touch of N1440GAT: signal is true;
	signal N1441GAT: std_logic; attribute dont_touch of N1441GAT: signal is true;
	signal N1442GAT: std_logic; attribute dont_touch of N1442GAT: signal is true;
	signal N1443GAT: std_logic; attribute dont_touch of N1443GAT: signal is true;
	signal N1444GAT: std_logic; attribute dont_touch of N1444GAT: signal is true;
	signal N1446GAT: std_logic; attribute dont_touch of N1446GAT: signal is true;
	signal N1447GAT: std_logic; attribute dont_touch of N1447GAT: signal is true;
	signal N1448GAT: std_logic; attribute dont_touch of N1448GAT: signal is true;
	signal N1449GAT: std_logic; attribute dont_touch of N1449GAT: signal is true;
	signal N1450GAT: std_logic; attribute dont_touch of N1450GAT: signal is true;
	signal N1451GAT: std_logic; attribute dont_touch of N1451GAT: signal is true;
	signal N1452GAT: std_logic; attribute dont_touch of N1452GAT: signal is true;
	signal N1453GAT: std_logic; attribute dont_touch of N1453GAT: signal is true;
	signal N1454GAT: std_logic; attribute dont_touch of N1454GAT: signal is true;
	signal N1455GAT: std_logic; attribute dont_touch of N1455GAT: signal is true;
	signal N1456GAT: std_logic; attribute dont_touch of N1456GAT: signal is true;
	signal N1458GAT: std_logic; attribute dont_touch of N1458GAT: signal is true;
	signal N1459GAT: std_logic; attribute dont_touch of N1459GAT: signal is true;
	signal N1460GAT: std_logic; attribute dont_touch of N1460GAT: signal is true;
	signal N1461GAT: std_logic; attribute dont_touch of N1461GAT: signal is true;
	signal N1462GAT: std_logic; attribute dont_touch of N1462GAT: signal is true;
	signal N1466GAT: std_logic; attribute dont_touch of N1466GAT: signal is true;
	signal N1467GAT: std_logic; attribute dont_touch of N1467GAT: signal is true;
	signal N1468GAT: std_logic; attribute dont_touch of N1468GAT: signal is true;
	signal N1469GAT: std_logic; attribute dont_touch of N1469GAT: signal is true;
	signal N1470GAT: std_logic; attribute dont_touch of N1470GAT: signal is true;
	signal N1471GAT: std_logic; attribute dont_touch of N1471GAT: signal is true;
	signal N1472GAT: std_logic; attribute dont_touch of N1472GAT: signal is true;
	signal N1476GAT: std_logic; attribute dont_touch of N1476GAT: signal is true;
	signal N1477GAT: std_logic; attribute dont_touch of N1477GAT: signal is true;
	signal N1478GAT: std_logic; attribute dont_touch of N1478GAT: signal is true;
	signal N1479GAT: std_logic; attribute dont_touch of N1479GAT: signal is true;
	signal N1480GAT: std_logic; attribute dont_touch of N1480GAT: signal is true;
	signal N1481GAT: std_logic; attribute dont_touch of N1481GAT: signal is true;
	signal N1482GAT: std_logic; attribute dont_touch of N1482GAT: signal is true;
	signal N1483GAT: std_logic; attribute dont_touch of N1483GAT: signal is true;
	signal N1484GAT: std_logic; attribute dont_touch of N1484GAT: signal is true;
	signal N1485GAT: std_logic; attribute dont_touch of N1485GAT: signal is true;
	signal N1486GAT: std_logic; attribute dont_touch of N1486GAT: signal is true;
	signal N1487GAT: std_logic; attribute dont_touch of N1487GAT: signal is true;
	signal N1490GAT: std_logic; attribute dont_touch of N1490GAT: signal is true;
	signal N1494GAT: std_logic; attribute dont_touch of N1494GAT: signal is true;
	signal N1495GAT: std_logic; attribute dont_touch of N1495GAT: signal is true;
	signal N1496GAT: std_logic; attribute dont_touch of N1496GAT: signal is true;
	signal N1498GAT: std_logic; attribute dont_touch of N1498GAT: signal is true;
	signal N1499GAT: std_logic; attribute dont_touch of N1499GAT: signal is true;
	signal N1500GAT: std_logic; attribute dont_touch of N1500GAT: signal is true;
	signal N1501GAT: std_logic; attribute dont_touch of N1501GAT: signal is true;
	signal N1502GAT: std_logic; attribute dont_touch of N1502GAT: signal is true;
	signal N1503GAT: std_logic; attribute dont_touch of N1503GAT: signal is true;
	signal N1504GAT: std_logic; attribute dont_touch of N1504GAT: signal is true;
	signal N1505GAT: std_logic; attribute dont_touch of N1505GAT: signal is true;
	signal N1507GAT: std_logic; attribute dont_touch of N1507GAT: signal is true;
	signal N1508GAT: std_logic; attribute dont_touch of N1508GAT: signal is true;
	signal N1510GAT: std_logic; attribute dont_touch of N1510GAT: signal is true;
	signal N1513GAT: std_logic; attribute dont_touch of N1513GAT: signal is true;
	signal N1515GAT: std_logic; attribute dont_touch of N1515GAT: signal is true;
	signal N1516GAT: std_logic; attribute dont_touch of N1516GAT: signal is true;
	signal N1517GAT: std_logic; attribute dont_touch of N1517GAT: signal is true;
	signal N1518GAT: std_logic; attribute dont_touch of N1518GAT: signal is true;
	signal N1519GAT: std_logic; attribute dont_touch of N1519GAT: signal is true;
	signal N1520GAT: std_logic; attribute dont_touch of N1520GAT: signal is true;
	signal N1521GAT: std_logic; attribute dont_touch of N1521GAT: signal is true;
	signal N1523GAT: std_logic; attribute dont_touch of N1523GAT: signal is true;
	signal N1524GAT: std_logic; attribute dont_touch of N1524GAT: signal is true;
	signal N1525GAT: std_logic; attribute dont_touch of N1525GAT: signal is true;
	signal N1528GAT: std_logic; attribute dont_touch of N1528GAT: signal is true;
	signal N1529GAT: std_logic; attribute dont_touch of N1529GAT: signal is true;
	signal N1530GAT: std_logic; attribute dont_touch of N1530GAT: signal is true;
	signal N1531GAT: std_logic; attribute dont_touch of N1531GAT: signal is true;
	signal N1532GAT: std_logic; attribute dont_touch of N1532GAT: signal is true;
	signal N1533GAT: std_logic; attribute dont_touch of N1533GAT: signal is true;
	signal N1543GAT: std_logic; attribute dont_touch of N1543GAT: signal is true;
	signal N1544GAT: std_logic; attribute dont_touch of N1544GAT: signal is true;
	signal N1546GAT: std_logic; attribute dont_touch of N1546GAT: signal is true;
	signal N1548GAT: std_logic; attribute dont_touch of N1548GAT: signal is true;
	signal N1549GAT: std_logic; attribute dont_touch of N1549GAT: signal is true;
	signal N1550GAT: std_logic; attribute dont_touch of N1550GAT: signal is true;
	signal N1551GAT: std_logic; attribute dont_touch of N1551GAT: signal is true;
	signal N1552GAT: std_logic; attribute dont_touch of N1552GAT: signal is true;
	signal N1553GAT: std_logic; attribute dont_touch of N1553GAT: signal is true;
	signal N1554GAT: std_logic; attribute dont_touch of N1554GAT: signal is true;
	signal N1555GAT: std_logic; attribute dont_touch of N1555GAT: signal is true;
	signal N1556GAT: std_logic; attribute dont_touch of N1556GAT: signal is true;
	signal N1557GAT: std_logic; attribute dont_touch of N1557GAT: signal is true;
	signal N1558GAT: std_logic; attribute dont_touch of N1558GAT: signal is true;
	signal N1559GAT: std_logic; attribute dont_touch of N1559GAT: signal is true;
	signal N1560GAT: std_logic; attribute dont_touch of N1560GAT: signal is true;
	signal N1561GAT: std_logic; attribute dont_touch of N1561GAT: signal is true;
	signal N1562GAT: std_logic; attribute dont_touch of N1562GAT: signal is true;
	signal N1563GAT: std_logic; attribute dont_touch of N1563GAT: signal is true;
	signal N1564GAT: std_logic; attribute dont_touch of N1564GAT: signal is true;
	signal N1565GAT: std_logic; attribute dont_touch of N1565GAT: signal is true;
	signal N1566GAT: std_logic; attribute dont_touch of N1566GAT: signal is true;
	signal N1567GAT: std_logic; attribute dont_touch of N1567GAT: signal is true;
	signal N1568GAT: std_logic; attribute dont_touch of N1568GAT: signal is true;
	signal N1569GAT: std_logic; attribute dont_touch of N1569GAT: signal is true;
	signal N1570GAT: std_logic; attribute dont_touch of N1570GAT: signal is true;
	signal N1571GAT: std_logic; attribute dont_touch of N1571GAT: signal is true;
	signal N1572GAT: std_logic; attribute dont_touch of N1572GAT: signal is true;
	signal N1573GAT: std_logic; attribute dont_touch of N1573GAT: signal is true;
	signal N1574GAT: std_logic; attribute dont_touch of N1574GAT: signal is true;
	signal N1575GAT: std_logic; attribute dont_touch of N1575GAT: signal is true;
	signal N1576GAT: std_logic; attribute dont_touch of N1576GAT: signal is true;
	signal N1577GAT: std_logic; attribute dont_touch of N1577GAT: signal is true;
	signal N1578GAT: std_logic; attribute dont_touch of N1578GAT: signal is true;
	signal N1580GAT: std_logic; attribute dont_touch of N1580GAT: signal is true;
	signal N1581GAT: std_logic; attribute dont_touch of N1581GAT: signal is true;
	signal N1582GAT: std_logic; attribute dont_touch of N1582GAT: signal is true;
	signal N1584GAT: std_logic; attribute dont_touch of N1584GAT: signal is true;
	signal N1586GAT: std_logic; attribute dont_touch of N1586GAT: signal is true;
	signal N1587GAT: std_logic; attribute dont_touch of N1587GAT: signal is true;
	signal N1588GAT: std_logic; attribute dont_touch of N1588GAT: signal is true;
	signal N1590GAT: std_logic; attribute dont_touch of N1590GAT: signal is true;
	signal N1591GAT: std_logic; attribute dont_touch of N1591GAT: signal is true;
	signal N1592GAT: std_logic; attribute dont_touch of N1592GAT: signal is true;
	signal N1593GAT: std_logic; attribute dont_touch of N1593GAT: signal is true;
	signal N1594GAT: std_logic; attribute dont_touch of N1594GAT: signal is true;
	signal N1595GAT: std_logic; attribute dont_touch of N1595GAT: signal is true;
	signal N1596GAT: std_logic; attribute dont_touch of N1596GAT: signal is true;
	signal N1598GAT: std_logic; attribute dont_touch of N1598GAT: signal is true;
	signal N1599GAT: std_logic; attribute dont_touch of N1599GAT: signal is true;
	signal N1600GAT: std_logic; attribute dont_touch of N1600GAT: signal is true;
	signal N1601GAT: std_logic; attribute dont_touch of N1601GAT: signal is true;
	signal N1602GAT: std_logic; attribute dont_touch of N1602GAT: signal is true;
	signal N1603GAT: std_logic; attribute dont_touch of N1603GAT: signal is true;
	signal N1604GAT: std_logic; attribute dont_touch of N1604GAT: signal is true;
	signal N1605GAT: std_logic; attribute dont_touch of N1605GAT: signal is true;
	signal N1606GAT: std_logic; attribute dont_touch of N1606GAT: signal is true;
	signal N1607GAT: std_logic; attribute dont_touch of N1607GAT: signal is true;
	signal N1608GAT: std_logic; attribute dont_touch of N1608GAT: signal is true;
	signal N1609GAT: std_logic; attribute dont_touch of N1609GAT: signal is true;
	signal N1610GAT: std_logic; attribute dont_touch of N1610GAT: signal is true;
	signal N1613GAT: std_logic; attribute dont_touch of N1613GAT: signal is true;
	signal N1614GAT: std_logic; attribute dont_touch of N1614GAT: signal is true;
	signal N1615GAT: std_logic; attribute dont_touch of N1615GAT: signal is true;
	signal N1616GAT: std_logic; attribute dont_touch of N1616GAT: signal is true;
	signal N1617GAT: std_logic; attribute dont_touch of N1617GAT: signal is true;
	signal N1618GAT: std_logic; attribute dont_touch of N1618GAT: signal is true;
	signal N1619GAT: std_logic; attribute dont_touch of N1619GAT: signal is true;
	signal N1620GAT: std_logic; attribute dont_touch of N1620GAT: signal is true;
	signal N1621GAT: std_logic; attribute dont_touch of N1621GAT: signal is true;
	signal N1622GAT: std_logic; attribute dont_touch of N1622GAT: signal is true;
	signal N1623GAT: std_logic; attribute dont_touch of N1623GAT: signal is true;
	signal N1624GAT: std_logic; attribute dont_touch of N1624GAT: signal is true;
	signal N1625GAT: std_logic; attribute dont_touch of N1625GAT: signal is true;
	signal N1626GAT: std_logic; attribute dont_touch of N1626GAT: signal is true;
	signal N1627GAT: std_logic; attribute dont_touch of N1627GAT: signal is true;
	signal N1628GAT: std_logic; attribute dont_touch of N1628GAT: signal is true;
	signal N1629GAT: std_logic; attribute dont_touch of N1629GAT: signal is true;
	signal N1630GAT: std_logic; attribute dont_touch of N1630GAT: signal is true;
	signal N1631GAT: std_logic; attribute dont_touch of N1631GAT: signal is true;
	signal N1632GAT: std_logic; attribute dont_touch of N1632GAT: signal is true;
	signal N1633GAT: std_logic; attribute dont_touch of N1633GAT: signal is true;
	signal N1634GAT: std_logic; attribute dont_touch of N1634GAT: signal is true;
	signal N1635GAT: std_logic; attribute dont_touch of N1635GAT: signal is true;
	signal N1636GAT: std_logic; attribute dont_touch of N1636GAT: signal is true;
	signal N1639GAT: std_logic; attribute dont_touch of N1639GAT: signal is true;
	signal N1640GAT: std_logic; attribute dont_touch of N1640GAT: signal is true;
	signal N1641GAT: std_logic; attribute dont_touch of N1641GAT: signal is true;
	signal N1642GAT: std_logic; attribute dont_touch of N1642GAT: signal is true;
	signal N1643GAT: std_logic; attribute dont_touch of N1643GAT: signal is true;
	signal N1644GAT: std_logic; attribute dont_touch of N1644GAT: signal is true;
	signal N1645GAT: std_logic; attribute dont_touch of N1645GAT: signal is true;
	signal N1646GAT: std_logic; attribute dont_touch of N1646GAT: signal is true;
	signal N1647GAT: std_logic; attribute dont_touch of N1647GAT: signal is true;
	signal N1648GAT: std_logic; attribute dont_touch of N1648GAT: signal is true;
	signal N1649GAT: std_logic; attribute dont_touch of N1649GAT: signal is true;
	signal N1650GAT: std_logic; attribute dont_touch of N1650GAT: signal is true;
	signal N1651GAT: std_logic; attribute dont_touch of N1651GAT: signal is true;
	signal N1652GAT: std_logic; attribute dont_touch of N1652GAT: signal is true;
	signal N1653GAT: std_logic; attribute dont_touch of N1653GAT: signal is true;
	signal N1654GAT: std_logic; attribute dont_touch of N1654GAT: signal is true;
	signal N1655GAT: std_logic; attribute dont_touch of N1655GAT: signal is true;
	signal N1656GAT: std_logic; attribute dont_touch of N1656GAT: signal is true;
	signal N1657GAT: std_logic; attribute dont_touch of N1657GAT: signal is true;
	signal N1658GAT: std_logic; attribute dont_touch of N1658GAT: signal is true;
	signal N1659GAT: std_logic; attribute dont_touch of N1659GAT: signal is true;
	signal N1660GAT: std_logic; attribute dont_touch of N1660GAT: signal is true;
	signal N1661GAT: std_logic; attribute dont_touch of N1661GAT: signal is true;
	signal N1662GAT: std_logic; attribute dont_touch of N1662GAT: signal is true;
	signal N1663GAT: std_logic; attribute dont_touch of N1663GAT: signal is true;
	signal N1665GAT: std_logic; attribute dont_touch of N1665GAT: signal is true;
	signal N1666GAT: std_logic; attribute dont_touch of N1666GAT: signal is true;
	signal N1667GAT: std_logic; attribute dont_touch of N1667GAT: signal is true;
	signal N1668GAT: std_logic; attribute dont_touch of N1668GAT: signal is true;
	signal N1669GAT: std_logic; attribute dont_touch of N1669GAT: signal is true;
	signal N1670GAT: std_logic; attribute dont_touch of N1670GAT: signal is true;
	signal N1671GAT: std_logic; attribute dont_touch of N1671GAT: signal is true;
	signal N1673GAT: std_logic; attribute dont_touch of N1673GAT: signal is true;
	signal N1674GAT: std_logic; attribute dont_touch of N1674GAT: signal is true;
	signal N1675GAT: std_logic; attribute dont_touch of N1675GAT: signal is true;
	signal N1677GAT: std_logic; attribute dont_touch of N1677GAT: signal is true;
	signal N1678GAT: std_logic; attribute dont_touch of N1678GAT: signal is true;
	signal N1681GAT: std_logic; attribute dont_touch of N1681GAT: signal is true;
	signal N1683GAT: std_logic; attribute dont_touch of N1683GAT: signal is true;
	signal N1684GAT: std_logic; attribute dont_touch of N1684GAT: signal is true;
	signal N1685GAT: std_logic; attribute dont_touch of N1685GAT: signal is true;
	signal N1686GAT: std_logic; attribute dont_touch of N1686GAT: signal is true;
	signal N1690GAT: std_logic; attribute dont_touch of N1690GAT: signal is true;
	signal N1691GAT: std_logic; attribute dont_touch of N1691GAT: signal is true;
	signal N1692GAT: std_logic; attribute dont_touch of N1692GAT: signal is true;
	signal N1693GAT: std_logic; attribute dont_touch of N1693GAT: signal is true;
	signal N1694GAT: std_logic; attribute dont_touch of N1694GAT: signal is true;
	signal N1695GAT: std_logic; attribute dont_touch of N1695GAT: signal is true;
	signal N1696GAT: std_logic; attribute dont_touch of N1696GAT: signal is true;
	signal N1698GAT: std_logic; attribute dont_touch of N1698GAT: signal is true;
	signal N1699GAT: std_logic; attribute dont_touch of N1699GAT: signal is true;
	signal N1700GAT: std_logic; attribute dont_touch of N1700GAT: signal is true;
	signal N1701GAT: std_logic; attribute dont_touch of N1701GAT: signal is true;
	signal N1702GAT: std_logic; attribute dont_touch of N1702GAT: signal is true;
	signal N1703GAT: std_logic; attribute dont_touch of N1703GAT: signal is true;
	signal N1704GAT: std_logic; attribute dont_touch of N1704GAT: signal is true;
	signal N1705GAT: std_logic; attribute dont_touch of N1705GAT: signal is true;
	signal N1706GAT: std_logic; attribute dont_touch of N1706GAT: signal is true;
	signal N1707GAT: std_logic; attribute dont_touch of N1707GAT: signal is true;
	signal N1708GAT: std_logic; attribute dont_touch of N1708GAT: signal is true;
	signal N1709GAT: std_logic; attribute dont_touch of N1709GAT: signal is true;
	signal N1710GAT: std_logic; attribute dont_touch of N1710GAT: signal is true;
	signal N1711GAT: std_logic; attribute dont_touch of N1711GAT: signal is true;
	signal N1712GAT: std_logic; attribute dont_touch of N1712GAT: signal is true;
	signal N1713GAT: std_logic; attribute dont_touch of N1713GAT: signal is true;
	signal N1714GAT: std_logic; attribute dont_touch of N1714GAT: signal is true;
	signal N1716GAT: std_logic; attribute dont_touch of N1716GAT: signal is true;
	signal N1717GAT: std_logic; attribute dont_touch of N1717GAT: signal is true;
	signal N1718GAT: std_logic; attribute dont_touch of N1718GAT: signal is true;
	signal N1719GAT: std_logic; attribute dont_touch of N1719GAT: signal is true;
	signal N1721GAT: std_logic; attribute dont_touch of N1721GAT: signal is true;
	signal N1722GAT: std_logic; attribute dont_touch of N1722GAT: signal is true;
	signal N1723GAT: std_logic; attribute dont_touch of N1723GAT: signal is true;
	signal N1724GAT: std_logic; attribute dont_touch of N1724GAT: signal is true;
	signal N1725GAT: std_logic; attribute dont_touch of N1725GAT: signal is true;
	signal N1726GAT: std_logic; attribute dont_touch of N1726GAT: signal is true;
	signal N1727GAT: std_logic; attribute dont_touch of N1727GAT: signal is true;
	signal N1728GAT: std_logic; attribute dont_touch of N1728GAT: signal is true;
	signal N1729GAT: std_logic; attribute dont_touch of N1729GAT: signal is true;
	signal N1730GAT: std_logic; attribute dont_touch of N1730GAT: signal is true;
	signal N1731GAT: std_logic; attribute dont_touch of N1731GAT: signal is true;
	signal N1732GAT: std_logic; attribute dont_touch of N1732GAT: signal is true;
	signal N1733GAT: std_logic; attribute dont_touch of N1733GAT: signal is true;
	signal N1734GAT: std_logic; attribute dont_touch of N1734GAT: signal is true;
	signal N1735GAT: std_logic; attribute dont_touch of N1735GAT: signal is true;
	signal N1736GAT: std_logic; attribute dont_touch of N1736GAT: signal is true;
	signal N1737GAT: std_logic; attribute dont_touch of N1737GAT: signal is true;
	signal N1738GAT: std_logic; attribute dont_touch of N1738GAT: signal is true;
	signal N1739GAT: std_logic; attribute dont_touch of N1739GAT: signal is true;
	signal N1740GAT: std_logic; attribute dont_touch of N1740GAT: signal is true;
	signal N1742GAT: std_logic; attribute dont_touch of N1742GAT: signal is true;
	signal N1743GAT: std_logic; attribute dont_touch of N1743GAT: signal is true;
	signal N1745GAT: std_logic; attribute dont_touch of N1745GAT: signal is true;
	signal N1747GAT: std_logic; attribute dont_touch of N1747GAT: signal is true;
	signal N1748GAT: std_logic; attribute dont_touch of N1748GAT: signal is true;
	signal N1754GAT: std_logic; attribute dont_touch of N1754GAT: signal is true;
	signal N1755GAT: std_logic; attribute dont_touch of N1755GAT: signal is true;
	signal N1756GAT: std_logic; attribute dont_touch of N1756GAT: signal is true;
	signal N1757GAT: std_logic; attribute dont_touch of N1757GAT: signal is true;
	signal N1758GAT: std_logic; attribute dont_touch of N1758GAT: signal is true;
	signal N1759GAT: std_logic; attribute dont_touch of N1759GAT: signal is true;
	signal N1760GAT: std_logic; attribute dont_touch of N1760GAT: signal is true;
	signal N1761GAT: std_logic; attribute dont_touch of N1761GAT: signal is true;
	signal N1762GAT: std_logic; attribute dont_touch of N1762GAT: signal is true;
	signal N1763GAT: std_logic; attribute dont_touch of N1763GAT: signal is true;
	signal N1765GAT: std_logic; attribute dont_touch of N1765GAT: signal is true;
	signal N1767GAT: std_logic; attribute dont_touch of N1767GAT: signal is true;
	signal N1769GAT: std_logic; attribute dont_touch of N1769GAT: signal is true;
	signal N1771GAT: std_logic; attribute dont_touch of N1771GAT: signal is true;
	signal N1773GAT: std_logic; attribute dont_touch of N1773GAT: signal is true;
	signal N1774GAT: std_logic; attribute dont_touch of N1774GAT: signal is true;
	signal N1775GAT: std_logic; attribute dont_touch of N1775GAT: signal is true;
	signal N1777GAT: std_logic; attribute dont_touch of N1777GAT: signal is true;
	signal N1778GAT: std_logic; attribute dont_touch of N1778GAT: signal is true;
	signal N1779GAT: std_logic; attribute dont_touch of N1779GAT: signal is true;
	signal N1780GAT: std_logic; attribute dont_touch of N1780GAT: signal is true;
	signal N1781GAT: std_logic; attribute dont_touch of N1781GAT: signal is true;
	signal N1782GAT: std_logic; attribute dont_touch of N1782GAT: signal is true;
	signal N1783GAT: std_logic; attribute dont_touch of N1783GAT: signal is true;
	signal N1784GAT: std_logic; attribute dont_touch of N1784GAT: signal is true;
	signal N1785GAT: std_logic; attribute dont_touch of N1785GAT: signal is true;
	signal N1786GAT: std_logic; attribute dont_touch of N1786GAT: signal is true;
	signal N1787GAT: std_logic; attribute dont_touch of N1787GAT: signal is true;
	signal N1788GAT: std_logic; attribute dont_touch of N1788GAT: signal is true;
	signal N1790GAT: std_logic; attribute dont_touch of N1790GAT: signal is true;
	signal N1791GAT: std_logic; attribute dont_touch of N1791GAT: signal is true;
	signal N1792GAT: std_logic; attribute dont_touch of N1792GAT: signal is true;
	signal N1793GAT: std_logic; attribute dont_touch of N1793GAT: signal is true;
	signal N1794GAT: std_logic; attribute dont_touch of N1794GAT: signal is true;
	signal N1796GAT: std_logic; attribute dont_touch of N1796GAT: signal is true;
	signal N1797GAT: std_logic; attribute dont_touch of N1797GAT: signal is true;
	signal N1798GAT: std_logic; attribute dont_touch of N1798GAT: signal is true;
	signal N1800GAT: std_logic; attribute dont_touch of N1800GAT: signal is true;
	signal N1801GAT: std_logic; attribute dont_touch of N1801GAT: signal is true;
	signal N1806GAT: std_logic; attribute dont_touch of N1806GAT: signal is true;
	signal N1807GAT: std_logic; attribute dont_touch of N1807GAT: signal is true;
	signal N1816GAT: std_logic; attribute dont_touch of N1816GAT: signal is true;
	signal N1817GAT: std_logic; attribute dont_touch of N1817GAT: signal is true;
	signal N1818GAT: std_logic; attribute dont_touch of N1818GAT: signal is true;
	signal N1819GAT: std_logic; attribute dont_touch of N1819GAT: signal is true;
	signal N1821GAT: std_logic; attribute dont_touch of N1821GAT: signal is true;
	signal N1823GAT: std_logic; attribute dont_touch of N1823GAT: signal is true;
	signal N1825GAT: std_logic; attribute dont_touch of N1825GAT: signal is true;
	signal N1827GAT: std_logic; attribute dont_touch of N1827GAT: signal is true;
	signal N1828GAT: std_logic; attribute dont_touch of N1828GAT: signal is true;
	signal N1829GAT: std_logic; attribute dont_touch of N1829GAT: signal is true;
	signal N1831GAT: std_logic; attribute dont_touch of N1831GAT: signal is true;
	signal N1832GAT: std_logic; attribute dont_touch of N1832GAT: signal is true;
	signal N1834GAT: std_logic; attribute dont_touch of N1834GAT: signal is true;
	signal N1836GAT: std_logic; attribute dont_touch of N1836GAT: signal is true;
	signal N1838GAT: std_logic; attribute dont_touch of N1838GAT: signal is true;
	signal N1839GAT: std_logic; attribute dont_touch of N1839GAT: signal is true;
	signal N1840GAT: std_logic; attribute dont_touch of N1840GAT: signal is true;
	signal N1841GAT: std_logic; attribute dont_touch of N1841GAT: signal is true;
	signal N1842GAT: std_logic; attribute dont_touch of N1842GAT: signal is true;
	signal N1845GAT: std_logic; attribute dont_touch of N1845GAT: signal is true;
	signal N1846GAT: std_logic; attribute dont_touch of N1846GAT: signal is true;
	signal N1847GAT: std_logic; attribute dont_touch of N1847GAT: signal is true;
	signal N1848GAT: std_logic; attribute dont_touch of N1848GAT: signal is true;
	signal N1849GAT: std_logic; attribute dont_touch of N1849GAT: signal is true;
	signal N1850GAT: std_logic; attribute dont_touch of N1850GAT: signal is true;
	signal N1855GAT: std_logic; attribute dont_touch of N1855GAT: signal is true;
	signal N1858GAT: std_logic; attribute dont_touch of N1858GAT: signal is true;
	signal N1859GAT: std_logic; attribute dont_touch of N1859GAT: signal is true;
	signal N1860GAT: std_logic; attribute dont_touch of N1860GAT: signal is true;
	signal N1861GAT: std_logic; attribute dont_touch of N1861GAT: signal is true;
	signal N1862GAT: std_logic; attribute dont_touch of N1862GAT: signal is true;
	signal N1863GAT: std_logic; attribute dont_touch of N1863GAT: signal is true;
	signal N1864GAT: std_logic; attribute dont_touch of N1864GAT: signal is true;
	signal N1865GAT: std_logic; attribute dont_touch of N1865GAT: signal is true;
	signal N1866GAT: std_logic; attribute dont_touch of N1866GAT: signal is true;
	signal N1869GAT: std_logic; attribute dont_touch of N1869GAT: signal is true;
	signal N1870GAT: std_logic; attribute dont_touch of N1870GAT: signal is true;
	signal N1871GAT: std_logic; attribute dont_touch of N1871GAT: signal is true;
	signal N1878GAT: std_logic; attribute dont_touch of N1878GAT: signal is true;
	signal N1879GAT: std_logic; attribute dont_touch of N1879GAT: signal is true;
	signal N1880GAT: std_logic; attribute dont_touch of N1880GAT: signal is true;
	signal N1882GAT: std_logic; attribute dont_touch of N1882GAT: signal is true;
	signal N1884GAT: std_logic; attribute dont_touch of N1884GAT: signal is true;
	signal N1885GAT: std_logic; attribute dont_touch of N1885GAT: signal is true;
	signal N1886GAT: std_logic; attribute dont_touch of N1886GAT: signal is true;
	signal N1887GAT: std_logic; attribute dont_touch of N1887GAT: signal is true;
	signal N1888GAT: std_logic; attribute dont_touch of N1888GAT: signal is true;
	signal N1889GAT: std_logic; attribute dont_touch of N1889GAT: signal is true;
	signal N1890GAT: std_logic; attribute dont_touch of N1890GAT: signal is true;
	signal N1891GAT: std_logic; attribute dont_touch of N1891GAT: signal is true;
	signal N1892GAT: std_logic; attribute dont_touch of N1892GAT: signal is true;
	signal N1893GAT: std_logic; attribute dont_touch of N1893GAT: signal is true;
	signal N1894GAT: std_logic; attribute dont_touch of N1894GAT: signal is true;
	signal N1895GAT: std_logic; attribute dont_touch of N1895GAT: signal is true;
	signal N1896GAT: std_logic; attribute dont_touch of N1896GAT: signal is true;
	signal N1897GAT: std_logic; attribute dont_touch of N1897GAT: signal is true;
	signal N1898GAT: std_logic; attribute dont_touch of N1898GAT: signal is true;
	signal N1899GAT: std_logic; attribute dont_touch of N1899GAT: signal is true;
	signal N1915GAT: std_logic; attribute dont_touch of N1915GAT: signal is true;
	signal N1916GAT: std_logic; attribute dont_touch of N1916GAT: signal is true;
	signal N1917GAT: std_logic; attribute dont_touch of N1917GAT: signal is true;
	signal N1918GAT: std_logic; attribute dont_touch of N1918GAT: signal is true;
	signal N1919GAT: std_logic; attribute dont_touch of N1919GAT: signal is true;
	signal N1920GAT: std_logic; attribute dont_touch of N1920GAT: signal is true;
	signal N1921GAT: std_logic; attribute dont_touch of N1921GAT: signal is true;
	signal N1922GAT: std_logic; attribute dont_touch of N1922GAT: signal is true;
	signal N1923GAT: std_logic; attribute dont_touch of N1923GAT: signal is true;
	signal N1924GAT: std_logic; attribute dont_touch of N1924GAT: signal is true;
	signal N1925GAT: std_logic; attribute dont_touch of N1925GAT: signal is true;
	signal N1926GAT: std_logic; attribute dont_touch of N1926GAT: signal is true;
	signal N1927GAT: std_logic; attribute dont_touch of N1927GAT: signal is true;
	signal N1929GAT: std_logic; attribute dont_touch of N1929GAT: signal is true;
	signal N1934GAT: std_logic; attribute dont_touch of N1934GAT: signal is true;
	signal N1935GAT: std_logic; attribute dont_touch of N1935GAT: signal is true;
	signal N1945GAT: std_logic; attribute dont_touch of N1945GAT: signal is true;
	signal N1954GAT: std_logic; attribute dont_touch of N1954GAT: signal is true;
	signal N1955GAT: std_logic; attribute dont_touch of N1955GAT: signal is true;
	signal N1956GAT: std_logic; attribute dont_touch of N1956GAT: signal is true;
	signal N1957GAT: std_logic; attribute dont_touch of N1957GAT: signal is true;
	signal N1958GAT: std_logic; attribute dont_touch of N1958GAT: signal is true;
	signal N1959GAT: std_logic; attribute dont_touch of N1959GAT: signal is true;
	signal N1960GAT: std_logic; attribute dont_touch of N1960GAT: signal is true;
	signal N1961GAT: std_logic; attribute dont_touch of N1961GAT: signal is true;
	signal N1962GAT: std_logic; attribute dont_touch of N1962GAT: signal is true;
	signal N1963GAT: std_logic; attribute dont_touch of N1963GAT: signal is true;
	signal N1964GAT: std_logic; attribute dont_touch of N1964GAT: signal is true;
	signal N1967GAT: std_logic; attribute dont_touch of N1967GAT: signal is true;
	signal N1968GAT: std_logic; attribute dont_touch of N1968GAT: signal is true;
	signal N1969GAT: std_logic; attribute dont_touch of N1969GAT: signal is true;
	signal N1970GAT: std_logic; attribute dont_touch of N1970GAT: signal is true;
	signal N1971GAT: std_logic; attribute dont_touch of N1971GAT: signal is true;
	signal N1972GAT: std_logic; attribute dont_touch of N1972GAT: signal is true;
	signal N1973GAT: std_logic; attribute dont_touch of N1973GAT: signal is true;
	signal N1974GAT: std_logic; attribute dont_touch of N1974GAT: signal is true;
	signal N1975GAT: std_logic; attribute dont_touch of N1975GAT: signal is true;
	signal N1978GAT: std_logic; attribute dont_touch of N1978GAT: signal is true;
	signal N1986GAT: std_logic; attribute dont_touch of N1986GAT: signal is true;
	signal N1988GAT: std_logic; attribute dont_touch of N1988GAT: signal is true;
	signal N1989GAT: std_logic; attribute dont_touch of N1989GAT: signal is true;
	signal N1990GAT: std_logic; attribute dont_touch of N1990GAT: signal is true;
	signal N1991GAT: std_logic; attribute dont_touch of N1991GAT: signal is true;
	signal N1994GAT: std_logic; attribute dont_touch of N1994GAT: signal is true;
	signal N1999GAT: std_logic; attribute dont_touch of N1999GAT: signal is true;
	signal N2000GAT: std_logic; attribute dont_touch of N2000GAT: signal is true;
	signal N2001GAT: std_logic; attribute dont_touch of N2001GAT: signal is true;
	signal N2002GAT: std_logic; attribute dont_touch of N2002GAT: signal is true;
	signal N2004GAT: std_logic; attribute dont_touch of N2004GAT: signal is true;
	signal N2005GAT: std_logic; attribute dont_touch of N2005GAT: signal is true;
	signal N2008GAT: std_logic; attribute dont_touch of N2008GAT: signal is true;
	signal N2009GAT: std_logic; attribute dont_touch of N2009GAT: signal is true;
	signal N2011GAT: std_logic; attribute dont_touch of N2011GAT: signal is true;
	signal N2012GAT: std_logic; attribute dont_touch of N2012GAT: signal is true;
	signal N2013GAT: std_logic; attribute dont_touch of N2013GAT: signal is true;
	signal N2014GAT: std_logic; attribute dont_touch of N2014GAT: signal is true;
	signal N2015GAT: std_logic; attribute dont_touch of N2015GAT: signal is true;
	signal N2016GAT: std_logic; attribute dont_touch of N2016GAT: signal is true;
	signal N2017GAT: std_logic; attribute dont_touch of N2017GAT: signal is true;
	signal N2018GAT: std_logic; attribute dont_touch of N2018GAT: signal is true;
	signal N2019GAT: std_logic; attribute dont_touch of N2019GAT: signal is true;
	signal N2021GAT: std_logic; attribute dont_touch of N2021GAT: signal is true;
	signal N2023GAT: std_logic; attribute dont_touch of N2023GAT: signal is true;
	signal N2025GAT: std_logic; attribute dont_touch of N2025GAT: signal is true;
	signal N2027GAT: std_logic; attribute dont_touch of N2027GAT: signal is true;
	signal N2029GAT: std_logic; attribute dont_touch of N2029GAT: signal is true;
	signal N2031GAT: std_logic; attribute dont_touch of N2031GAT: signal is true;
	signal N2033GAT: std_logic; attribute dont_touch of N2033GAT: signal is true;
	signal N2035GAT: std_logic; attribute dont_touch of N2035GAT: signal is true;
	signal N2037GAT: std_logic; attribute dont_touch of N2037GAT: signal is true;
	signal N2039GAT: std_logic; attribute dont_touch of N2039GAT: signal is true;
	signal N2040GAT: std_logic; attribute dont_touch of N2040GAT: signal is true;
	signal N2042GAT: std_logic; attribute dont_touch of N2042GAT: signal is true;
	signal N2044GAT: std_logic; attribute dont_touch of N2044GAT: signal is true;
	signal N2046GAT: std_logic; attribute dont_touch of N2046GAT: signal is true;
	signal N2047GAT: std_logic; attribute dont_touch of N2047GAT: signal is true;
	signal N2048GAT: std_logic; attribute dont_touch of N2048GAT: signal is true;
	signal N2049GAT: std_logic; attribute dont_touch of N2049GAT: signal is true;
	signal N2050GAT: std_logic; attribute dont_touch of N2050GAT: signal is true;
	signal N2051GAT: std_logic; attribute dont_touch of N2051GAT: signal is true;
	signal N2052GAT: std_logic; attribute dont_touch of N2052GAT: signal is true;
	signal N2053GAT: std_logic; attribute dont_touch of N2053GAT: signal is true;
	signal N2054GAT: std_logic; attribute dont_touch of N2054GAT: signal is true;
	signal N2055GAT: std_logic; attribute dont_touch of N2055GAT: signal is true;
	signal N2056GAT: std_logic; attribute dont_touch of N2056GAT: signal is true;
	signal N2057GAT: std_logic; attribute dont_touch of N2057GAT: signal is true;
	signal N2058GAT: std_logic; attribute dont_touch of N2058GAT: signal is true;
	signal N2059GAT: std_logic; attribute dont_touch of N2059GAT: signal is true;
	signal N2060GAT: std_logic; attribute dont_touch of N2060GAT: signal is true;
	signal N2061GAT: std_logic; attribute dont_touch of N2061GAT: signal is true;
	signal N2073GAT: std_logic; attribute dont_touch of N2073GAT: signal is true;
	signal N2078GAT: std_logic; attribute dont_touch of N2078GAT: signal is true;
	signal N2079GAT: std_logic; attribute dont_touch of N2079GAT: signal is true;
	signal N2081GAT: std_logic; attribute dont_touch of N2081GAT: signal is true;
	signal N2082GAT: std_logic; attribute dont_touch of N2082GAT: signal is true;
	signal N2084GAT: std_logic; attribute dont_touch of N2084GAT: signal is true;
	signal N2090GAT: std_logic; attribute dont_touch of N2090GAT: signal is true;
	signal N2091GAT: std_logic; attribute dont_touch of N2091GAT: signal is true;
	signal N2093GAT: std_logic; attribute dont_touch of N2093GAT: signal is true;
	signal N2095GAT: std_logic; attribute dont_touch of N2095GAT: signal is true;
	signal N2097GAT: std_logic; attribute dont_touch of N2097GAT: signal is true;
	signal N2099GAT: std_logic; attribute dont_touch of N2099GAT: signal is true;
	signal N2101GAT: std_logic; attribute dont_touch of N2101GAT: signal is true;
	signal N2102GAT: std_logic; attribute dont_touch of N2102GAT: signal is true;
	signal N2108GAT: std_logic; attribute dont_touch of N2108GAT: signal is true;
	signal N2110GAT: std_logic; attribute dont_touch of N2110GAT: signal is true;
	signal N2115GAT: std_logic; attribute dont_touch of N2115GAT: signal is true;
	signal N2117GAT: std_logic; attribute dont_touch of N2117GAT: signal is true;
	signal N2119GAT: std_logic; attribute dont_touch of N2119GAT: signal is true;
	signal N2121GAT: std_logic; attribute dont_touch of N2121GAT: signal is true;
	signal N2123GAT: std_logic; attribute dont_touch of N2123GAT: signal is true;
	signal N2124GAT: std_logic; attribute dont_touch of N2124GAT: signal is true;
	signal N2125GAT: std_logic; attribute dont_touch of N2125GAT: signal is true;
	signal N2127GAT: std_logic; attribute dont_touch of N2127GAT: signal is true;
	signal N2128GAT: std_logic; attribute dont_touch of N2128GAT: signal is true;
	signal N2129GAT: std_logic; attribute dont_touch of N2129GAT: signal is true;
	signal N2130GAT: std_logic; attribute dont_touch of N2130GAT: signal is true;
	signal N2131GAT: std_logic; attribute dont_touch of N2131GAT: signal is true;
	signal N2132GAT: std_logic; attribute dont_touch of N2132GAT: signal is true;
	signal N2133GAT: std_logic; attribute dont_touch of N2133GAT: signal is true;
	signal N2134GAT: std_logic; attribute dont_touch of N2134GAT: signal is true;
	signal N2135GAT: std_logic; attribute dont_touch of N2135GAT: signal is true;
	signal N2137GAT: std_logic; attribute dont_touch of N2137GAT: signal is true;
	signal N2138GAT: std_logic; attribute dont_touch of N2138GAT: signal is true;
	signal N2139GAT: std_logic; attribute dont_touch of N2139GAT: signal is true;
	signal N2141GAT: std_logic; attribute dont_touch of N2141GAT: signal is true;
	signal N2142GAT: std_logic; attribute dont_touch of N2142GAT: signal is true;
	signal N2143GAT: std_logic; attribute dont_touch of N2143GAT: signal is true;
	signal N2146GAT: std_logic; attribute dont_touch of N2146GAT: signal is true;
	signal N2147GAT: std_logic; attribute dont_touch of N2147GAT: signal is true;
	signal N2148GAT: std_logic; attribute dont_touch of N2148GAT: signal is true;
	signal N2149GAT: std_logic; attribute dont_touch of N2149GAT: signal is true;
	signal N2150GAT: std_logic; attribute dont_touch of N2150GAT: signal is true;
	signal N2151GAT: std_logic; attribute dont_touch of N2151GAT: signal is true;
	signal N2152GAT: std_logic; attribute dont_touch of N2152GAT: signal is true;
	signal N2153GAT: std_logic; attribute dont_touch of N2153GAT: signal is true;
	signal N2154GAT: std_logic; attribute dont_touch of N2154GAT: signal is true;
	signal N2155GAT: std_logic; attribute dont_touch of N2155GAT: signal is true;
	signal N2158GAT: std_logic; attribute dont_touch of N2158GAT: signal is true;
	signal N2159GAT: std_logic; attribute dont_touch of N2159GAT: signal is true;
	signal N2162GAT: std_logic; attribute dont_touch of N2162GAT: signal is true;
	signal N2163GAT: std_logic; attribute dont_touch of N2163GAT: signal is true;
	signal N2167GAT: std_logic; attribute dont_touch of N2167GAT: signal is true;
	signal N2168GAT: std_logic; attribute dont_touch of N2168GAT: signal is true;
	signal N2169GAT: std_logic; attribute dont_touch of N2169GAT: signal is true;
	signal N2174GAT: std_logic; attribute dont_touch of N2174GAT: signal is true;
	signal N2176GAT: std_logic; attribute dont_touch of N2176GAT: signal is true;
	signal N2178GAT: std_logic; attribute dont_touch of N2178GAT: signal is true;
	signal N2179GAT: std_logic; attribute dont_touch of N2179GAT: signal is true;
	signal N2181GAT: std_logic; attribute dont_touch of N2181GAT: signal is true;
	signal N2182GAT: std_logic; attribute dont_touch of N2182GAT: signal is true;
	signal N2184GAT: std_logic; attribute dont_touch of N2184GAT: signal is true;
	signal N2185GAT: std_logic; attribute dont_touch of N2185GAT: signal is true;
	signal N2186GAT: std_logic; attribute dont_touch of N2186GAT: signal is true;
	signal N2187GAT: std_logic; attribute dont_touch of N2187GAT: signal is true;
	signal N2188GAT: std_logic; attribute dont_touch of N2188GAT: signal is true;
	signal N2189GAT: std_logic; attribute dont_touch of N2189GAT: signal is true;
	signal N2190GAT: std_logic; attribute dont_touch of N2190GAT: signal is true;
	signal N2192GAT: std_logic; attribute dont_touch of N2192GAT: signal is true;
	signal N2193GAT: std_logic; attribute dont_touch of N2193GAT: signal is true;
	signal N2194GAT: std_logic; attribute dont_touch of N2194GAT: signal is true;
	signal N2195GAT: std_logic; attribute dont_touch of N2195GAT: signal is true;
	signal N2196GAT: std_logic; attribute dont_touch of N2196GAT: signal is true;
	signal N2197GAT: std_logic; attribute dont_touch of N2197GAT: signal is true;
	signal N2198GAT: std_logic; attribute dont_touch of N2198GAT: signal is true;
	signal N2199GAT: std_logic; attribute dont_touch of N2199GAT: signal is true;
	signal N2200GAT: std_logic; attribute dont_touch of N2200GAT: signal is true;
	signal N2201GAT: std_logic; attribute dont_touch of N2201GAT: signal is true;
	signal N2202GAT: std_logic; attribute dont_touch of N2202GAT: signal is true;
	signal N2203GAT: std_logic; attribute dont_touch of N2203GAT: signal is true;
	signal N2205GAT: std_logic; attribute dont_touch of N2205GAT: signal is true;
	signal N2206GAT: std_logic; attribute dont_touch of N2206GAT: signal is true;
	signal N2207GAT: std_logic; attribute dont_touch of N2207GAT: signal is true;
	signal N2209GAT: std_logic; attribute dont_touch of N2209GAT: signal is true;
	signal N2210GAT: std_logic; attribute dont_touch of N2210GAT: signal is true;
	signal N2211GAT: std_logic; attribute dont_touch of N2211GAT: signal is true;
	signal N2212GAT: std_logic; attribute dont_touch of N2212GAT: signal is true;
	signal N2213GAT: std_logic; attribute dont_touch of N2213GAT: signal is true;
	signal N2214GAT: std_logic; attribute dont_touch of N2214GAT: signal is true;
	signal N2215GAT: std_logic; attribute dont_touch of N2215GAT: signal is true;
	signal N2216GAT: std_logic; attribute dont_touch of N2216GAT: signal is true;
	signal N2217GAT: std_logic; attribute dont_touch of N2217GAT: signal is true;
	signal N2218GAT: std_logic; attribute dont_touch of N2218GAT: signal is true;
	signal N2219GAT: std_logic; attribute dont_touch of N2219GAT: signal is true;
	signal N2220GAT: std_logic; attribute dont_touch of N2220GAT: signal is true;
	signal N2223GAT: std_logic; attribute dont_touch of N2223GAT: signal is true;
	signal N2237GAT: std_logic; attribute dont_touch of N2237GAT: signal is true;
	signal N2238GAT: std_logic; attribute dont_touch of N2238GAT: signal is true;
	signal N2239GAT: std_logic; attribute dont_touch of N2239GAT: signal is true;
	signal N2243GAT: std_logic; attribute dont_touch of N2243GAT: signal is true;
	signal N2244GAT: std_logic; attribute dont_touch of N2244GAT: signal is true;
	signal N2245GAT: std_logic; attribute dont_touch of N2245GAT: signal is true;
	signal N2246GAT: std_logic; attribute dont_touch of N2246GAT: signal is true;
	signal N2248GAT: std_logic; attribute dont_touch of N2248GAT: signal is true;
	signal N2249GAT: std_logic; attribute dont_touch of N2249GAT: signal is true;
	signal N2250GAT: std_logic; attribute dont_touch of N2250GAT: signal is true;
	signal N2251GAT: std_logic; attribute dont_touch of N2251GAT: signal is true;
	signal N2252GAT: std_logic; attribute dont_touch of N2252GAT: signal is true;
	signal N2253GAT: std_logic; attribute dont_touch of N2253GAT: signal is true;
	signal N2255GAT: std_logic; attribute dont_touch of N2255GAT: signal is true;
	signal N2256GAT: std_logic; attribute dont_touch of N2256GAT: signal is true;
	signal N2257GAT: std_logic; attribute dont_touch of N2257GAT: signal is true;
	signal N2258GAT: std_logic; attribute dont_touch of N2258GAT: signal is true;
	signal N2259GAT: std_logic; attribute dont_touch of N2259GAT: signal is true;
	signal N2260GAT: std_logic; attribute dont_touch of N2260GAT: signal is true;
	signal N2261GAT: std_logic; attribute dont_touch of N2261GAT: signal is true;
	signal N2262GAT: std_logic; attribute dont_touch of N2262GAT: signal is true;
	signal N2264GAT: std_logic; attribute dont_touch of N2264GAT: signal is true;
	signal N2265GAT: std_logic; attribute dont_touch of N2265GAT: signal is true;
	signal N2266GAT: std_logic; attribute dont_touch of N2266GAT: signal is true;
	signal N2268GAT: std_logic; attribute dont_touch of N2268GAT: signal is true;
	signal N2269GAT: std_logic; attribute dont_touch of N2269GAT: signal is true;
	signal N2270GAT: std_logic; attribute dont_touch of N2270GAT: signal is true;
	signal N2281GAT: std_logic; attribute dont_touch of N2281GAT: signal is true;
	signal N2282GAT: std_logic; attribute dont_touch of N2282GAT: signal is true;
	signal N2283GAT: std_logic; attribute dont_touch of N2283GAT: signal is true;
	signal N2284GAT: std_logic; attribute dont_touch of N2284GAT: signal is true;
	signal N2285GAT: std_logic; attribute dont_touch of N2285GAT: signal is true;
	signal N2286GAT: std_logic; attribute dont_touch of N2286GAT: signal is true;
	signal N2288GAT: std_logic; attribute dont_touch of N2288GAT: signal is true;
	signal N2289GAT: std_logic; attribute dont_touch of N2289GAT: signal is true;
	signal N2290GAT: std_logic; attribute dont_touch of N2290GAT: signal is true;
	signal N2291GAT: std_logic; attribute dont_touch of N2291GAT: signal is true;
	signal N2292GAT: std_logic; attribute dont_touch of N2292GAT: signal is true;
	signal N2293GAT: std_logic; attribute dont_touch of N2293GAT: signal is true;
	signal N2306GAT: std_logic; attribute dont_touch of N2306GAT: signal is true;
	signal N2307GAT: std_logic; attribute dont_touch of N2307GAT: signal is true;
	signal N2309GAT: std_logic; attribute dont_touch of N2309GAT: signal is true;
	signal N2317GAT: std_logic; attribute dont_touch of N2317GAT: signal is true;
	signal N2319GAT: std_logic; attribute dont_touch of N2319GAT: signal is true;
	signal N2325GAT: std_logic; attribute dont_touch of N2325GAT: signal is true;
	signal N2328GAT: std_logic; attribute dont_touch of N2328GAT: signal is true;
	signal N2329GAT: std_logic; attribute dont_touch of N2329GAT: signal is true;
	signal N2330GAT: std_logic; attribute dont_touch of N2330GAT: signal is true;
	signal N2331GAT: std_logic; attribute dont_touch of N2331GAT: signal is true;
	signal N2332GAT: std_logic; attribute dont_touch of N2332GAT: signal is true;
	signal N2333GAT: std_logic; attribute dont_touch of N2333GAT: signal is true;
	signal N2337GAT: std_logic; attribute dont_touch of N2337GAT: signal is true;
	signal N2338GAT: std_logic; attribute dont_touch of N2338GAT: signal is true;
	signal N2339GAT: std_logic; attribute dont_touch of N2339GAT: signal is true;
	signal N2341GAT: std_logic; attribute dont_touch of N2341GAT: signal is true;
	signal N2342GAT: std_logic; attribute dont_touch of N2342GAT: signal is true;
	signal N2343GAT: std_logic; attribute dont_touch of N2343GAT: signal is true;
	signal N2345GAT: std_logic; attribute dont_touch of N2345GAT: signal is true;
	signal N2346GAT: std_logic; attribute dont_touch of N2346GAT: signal is true;
	signal N2347GAT: std_logic; attribute dont_touch of N2347GAT: signal is true;
	signal N2349GAT: std_logic; attribute dont_touch of N2349GAT: signal is true;
	signal N2350GAT: std_logic; attribute dont_touch of N2350GAT: signal is true;
	signal N2351GAT: std_logic; attribute dont_touch of N2351GAT: signal is true;
	signal N2352GAT: std_logic; attribute dont_touch of N2352GAT: signal is true;
	signal N2353GAT: std_logic; attribute dont_touch of N2353GAT: signal is true;
	signal N2354GAT: std_logic; attribute dont_touch of N2354GAT: signal is true;
	signal N2355GAT: std_logic; attribute dont_touch of N2355GAT: signal is true;
	signal N2356GAT: std_logic; attribute dont_touch of N2356GAT: signal is true;
	signal N2357GAT: std_logic; attribute dont_touch of N2357GAT: signal is true;
	signal N2358GAT: std_logic; attribute dont_touch of N2358GAT: signal is true;
	signal N2359GAT: std_logic; attribute dont_touch of N2359GAT: signal is true;
	signal N2363GAT: std_logic; attribute dont_touch of N2363GAT: signal is true;
	signal N2364GAT: std_logic; attribute dont_touch of N2364GAT: signal is true;
	signal N2384GAT: std_logic; attribute dont_touch of N2384GAT: signal is true;
	signal N2385GAT: std_logic; attribute dont_touch of N2385GAT: signal is true;
	signal N2387GAT: std_logic; attribute dont_touch of N2387GAT: signal is true;
	signal N2388GAT: std_logic; attribute dont_touch of N2388GAT: signal is true;
	signal N2389GAT: std_logic; attribute dont_touch of N2389GAT: signal is true;
	signal N2390GAT: std_logic; attribute dont_touch of N2390GAT: signal is true;
	signal N2392GAT: std_logic; attribute dont_touch of N2392GAT: signal is true;
	signal N2393GAT: std_logic; attribute dont_touch of N2393GAT: signal is true;
	signal N2394GAT: std_logic; attribute dont_touch of N2394GAT: signal is true;
	signal N2396GAT: std_logic; attribute dont_touch of N2396GAT: signal is true;
	signal N2397GAT: std_logic; attribute dont_touch of N2397GAT: signal is true;
	signal N2398GAT: std_logic; attribute dont_touch of N2398GAT: signal is true;
	signal N2399GAT: std_logic; attribute dont_touch of N2399GAT: signal is true;
	signal N2401GAT: std_logic; attribute dont_touch of N2401GAT: signal is true;
	signal N2402GAT: std_logic; attribute dont_touch of N2402GAT: signal is true;
	signal N2403GAT: std_logic; attribute dont_touch of N2403GAT: signal is true;
	signal N2405GAT: std_logic; attribute dont_touch of N2405GAT: signal is true;
	signal N2406GAT: std_logic; attribute dont_touch of N2406GAT: signal is true;
	signal N2407GAT: std_logic; attribute dont_touch of N2407GAT: signal is true;
	signal N2409GAT: std_logic; attribute dont_touch of N2409GAT: signal is true;
	signal N2410GAT: std_logic; attribute dont_touch of N2410GAT: signal is true;
	signal N2411GAT: std_logic; attribute dont_touch of N2411GAT: signal is true;
	signal N2412GAT: std_logic; attribute dont_touch of N2412GAT: signal is true;
	signal N2413GAT: std_logic; attribute dont_touch of N2413GAT: signal is true;
	signal N2414GAT: std_logic; attribute dont_touch of N2414GAT: signal is true;
	signal N2415GAT: std_logic; attribute dont_touch of N2415GAT: signal is true;
	signal N2416GAT: std_logic; attribute dont_touch of N2416GAT: signal is true;
	signal N2417GAT: std_logic; attribute dont_touch of N2417GAT: signal is true;
	signal N2418GAT: std_logic; attribute dont_touch of N2418GAT: signal is true;
	signal N2419GAT: std_logic; attribute dont_touch of N2419GAT: signal is true;
	signal N2421GAT: std_logic; attribute dont_touch of N2421GAT: signal is true;
	signal N2422GAT: std_logic; attribute dont_touch of N2422GAT: signal is true;
	signal N2423GAT: std_logic; attribute dont_touch of N2423GAT: signal is true;
	signal N2426GAT: std_logic; attribute dont_touch of N2426GAT: signal is true;
	signal N2427GAT: std_logic; attribute dont_touch of N2427GAT: signal is true;
	signal N2428GAT: std_logic; attribute dont_touch of N2428GAT: signal is true;
	signal N2429GAT: std_logic; attribute dont_touch of N2429GAT: signal is true;
	signal N2430GAT: std_logic; attribute dont_touch of N2430GAT: signal is true;
	signal N2432GAT: std_logic; attribute dont_touch of N2432GAT: signal is true;
	signal N2433GAT: std_logic; attribute dont_touch of N2433GAT: signal is true;
	signal N2436GAT: std_logic; attribute dont_touch of N2436GAT: signal is true;
	signal N2437GAT: std_logic; attribute dont_touch of N2437GAT: signal is true;
	signal N2438GAT: std_logic; attribute dont_touch of N2438GAT: signal is true;
	signal N2439GAT: std_logic; attribute dont_touch of N2439GAT: signal is true;
	signal N2440GAT: std_logic; attribute dont_touch of N2440GAT: signal is true;
	signal N2442GAT: std_logic; attribute dont_touch of N2442GAT: signal is true;
	signal N2443GAT: std_logic; attribute dont_touch of N2443GAT: signal is true;
	signal N2444GAT: std_logic; attribute dont_touch of N2444GAT: signal is true;
	signal N2446GAT: std_logic; attribute dont_touch of N2446GAT: signal is true;
	signal N2448GAT: std_logic; attribute dont_touch of N2448GAT: signal is true;
	signal N2449GAT: std_logic; attribute dont_touch of N2449GAT: signal is true;
	signal N2450GAT: std_logic; attribute dont_touch of N2450GAT: signal is true;
	signal N2452GAT: std_logic; attribute dont_touch of N2452GAT: signal is true;
	signal N2454GAT: std_logic; attribute dont_touch of N2454GAT: signal is true;
	signal N2456GAT: std_logic; attribute dont_touch of N2456GAT: signal is true;
	signal N2458GAT: std_logic; attribute dont_touch of N2458GAT: signal is true;
	signal N2460GAT: std_logic; attribute dont_touch of N2460GAT: signal is true;
	signal N2461GAT: std_logic; attribute dont_touch of N2461GAT: signal is true;
	signal N2462GAT: std_logic; attribute dont_touch of N2462GAT: signal is true;
	signal N2464GAT: std_logic; attribute dont_touch of N2464GAT: signal is true;
	signal N2466GAT: std_logic; attribute dont_touch of N2466GAT: signal is true;
	signal N2468GAT: std_logic; attribute dont_touch of N2468GAT: signal is true;
	signal N2470GAT: std_logic; attribute dont_touch of N2470GAT: signal is true;
	signal N2472GAT: std_logic; attribute dont_touch of N2472GAT: signal is true;
	signal N2474GAT: std_logic; attribute dont_touch of N2474GAT: signal is true;
	signal N2476GAT: std_logic; attribute dont_touch of N2476GAT: signal is true;
	signal N2478GAT: std_logic; attribute dont_touch of N2478GAT: signal is true;
	signal N2480GAT: std_logic; attribute dont_touch of N2480GAT: signal is true;
	signal N2482GAT: std_logic; attribute dont_touch of N2482GAT: signal is true;
	signal N2483GAT: std_logic; attribute dont_touch of N2483GAT: signal is true;
	signal N2486GAT: std_logic; attribute dont_touch of N2486GAT: signal is true;
	signal N2487GAT: std_logic; attribute dont_touch of N2487GAT: signal is true;
	signal N2488GAT: std_logic; attribute dont_touch of N2488GAT: signal is true;
	signal N2489GAT: std_logic; attribute dont_touch of N2489GAT: signal is true;
	signal N2490GAT: std_logic; attribute dont_touch of N2490GAT: signal is true;
	signal N2492GAT: std_logic; attribute dont_touch of N2492GAT: signal is true;
	signal N2493GAT: std_logic; attribute dont_touch of N2493GAT: signal is true;
	signal N2494GAT: std_logic; attribute dont_touch of N2494GAT: signal is true;
	signal N2495GAT: std_logic; attribute dont_touch of N2495GAT: signal is true;
	signal N2498GAT: std_logic; attribute dont_touch of N2498GAT: signal is true;
	signal N2499GAT: std_logic; attribute dont_touch of N2499GAT: signal is true;
	signal N2500GAT: std_logic; attribute dont_touch of N2500GAT: signal is true;
	signal N2502GAT: std_logic; attribute dont_touch of N2502GAT: signal is true;
	signal N2504GAT: std_logic; attribute dont_touch of N2504GAT: signal is true;
	signal N2506GAT: std_logic; attribute dont_touch of N2506GAT: signal is true;
	signal N2508GAT: std_logic; attribute dont_touch of N2508GAT: signal is true;
	signal N2510GAT: std_logic; attribute dont_touch of N2510GAT: signal is true;
	signal N2512GAT: std_logic; attribute dont_touch of N2512GAT: signal is true;
	signal N2514GAT: std_logic; attribute dont_touch of N2514GAT: signal is true;
	signal N2516GAT: std_logic; attribute dont_touch of N2516GAT: signal is true;
	signal N2518GAT: std_logic; attribute dont_touch of N2518GAT: signal is true;
	signal N2520GAT: std_logic; attribute dont_touch of N2520GAT: signal is true;
	signal N2522GAT: std_logic; attribute dont_touch of N2522GAT: signal is true;
	signal N2524GAT: std_logic; attribute dont_touch of N2524GAT: signal is true;
	signal N2526GAT: std_logic; attribute dont_touch of N2526GAT: signal is true;
	signal N2530GAT: std_logic; attribute dont_touch of N2530GAT: signal is true;
	signal N2531GAT: std_logic; attribute dont_touch of N2531GAT: signal is true;
	signal N2532GAT: std_logic; attribute dont_touch of N2532GAT: signal is true;
	signal N2533GAT: std_logic; attribute dont_touch of N2533GAT: signal is true;
	signal N2534GAT: std_logic; attribute dont_touch of N2534GAT: signal is true;
	signal N2536GAT: std_logic; attribute dont_touch of N2536GAT: signal is true;
	signal N2537GAT: std_logic; attribute dont_touch of N2537GAT: signal is true;
	signal N2538GAT: std_logic; attribute dont_touch of N2538GAT: signal is true;
	signal N2539GAT: std_logic; attribute dont_touch of N2539GAT: signal is true;
	signal N2540GAT: std_logic; attribute dont_touch of N2540GAT: signal is true;
	signal N2541GAT: std_logic; attribute dont_touch of N2541GAT: signal is true;
	signal N2542GAT: std_logic; attribute dont_touch of N2542GAT: signal is true;
	signal N2543GAT: std_logic; attribute dont_touch of N2543GAT: signal is true;
	signal N2545GAT: std_logic; attribute dont_touch of N2545GAT: signal is true;
	signal N2546GAT: std_logic; attribute dont_touch of N2546GAT: signal is true;
	signal N2547GAT: std_logic; attribute dont_touch of N2547GAT: signal is true;
	signal N2548GAT: std_logic; attribute dont_touch of N2548GAT: signal is true;
	signal N2549GAT: std_logic; attribute dont_touch of N2549GAT: signal is true;
	signal N2550GAT: std_logic; attribute dont_touch of N2550GAT: signal is true;
	signal N2551GAT: std_logic; attribute dont_touch of N2551GAT: signal is true;
	signal N2552GAT: std_logic; attribute dont_touch of N2552GAT: signal is true;
	signal N2553GAT: std_logic; attribute dont_touch of N2553GAT: signal is true;
	signal N2554GAT: std_logic; attribute dont_touch of N2554GAT: signal is true;
	signal N2555GAT: std_logic; attribute dont_touch of N2555GAT: signal is true;
	signal N2556GAT: std_logic; attribute dont_touch of N2556GAT: signal is true;
	signal N2557GAT: std_logic; attribute dont_touch of N2557GAT: signal is true;
	signal N2558GAT: std_logic; attribute dont_touch of N2558GAT: signal is true;
	signal N2559GAT: std_logic; attribute dont_touch of N2559GAT: signal is true;
	signal N2560GAT: std_logic; attribute dont_touch of N2560GAT: signal is true;
	signal N2561GAT: std_logic; attribute dont_touch of N2561GAT: signal is true;
	signal N2562GAT: std_logic; attribute dont_touch of N2562GAT: signal is true;
	signal N2564GAT: std_logic; attribute dont_touch of N2564GAT: signal is true;
	signal N2565GAT: std_logic; attribute dont_touch of N2565GAT: signal is true;
	signal N2566GAT: std_logic; attribute dont_touch of N2566GAT: signal is true;
	signal N2567GAT: std_logic; attribute dont_touch of N2567GAT: signal is true;
	signal N2568GAT: std_logic; attribute dont_touch of N2568GAT: signal is true;
	signal N2569GAT: std_logic; attribute dont_touch of N2569GAT: signal is true;
	signal N2570GAT: std_logic; attribute dont_touch of N2570GAT: signal is true;
	signal N2571GAT: std_logic; attribute dont_touch of N2571GAT: signal is true;
	signal N2572GAT: std_logic; attribute dont_touch of N2572GAT: signal is true;
	signal N2573GAT: std_logic; attribute dont_touch of N2573GAT: signal is true;
	signal N2574GAT: std_logic; attribute dont_touch of N2574GAT: signal is true;
	signal N2575GAT: std_logic; attribute dont_touch of N2575GAT: signal is true;
	signal N2576GAT: std_logic; attribute dont_touch of N2576GAT: signal is true;
	signal N2577GAT: std_logic; attribute dont_touch of N2577GAT: signal is true;
	signal N2578GAT: std_logic; attribute dont_touch of N2578GAT: signal is true;
	signal N2579GAT: std_logic; attribute dont_touch of N2579GAT: signal is true;
	signal N2580GAT: std_logic; attribute dont_touch of N2580GAT: signal is true;
	signal N2581GAT: std_logic; attribute dont_touch of N2581GAT: signal is true;
	signal N2582GAT: std_logic; attribute dont_touch of N2582GAT: signal is true;
	signal N2583GAT: std_logic; attribute dont_touch of N2583GAT: signal is true;
	signal N2585GAT: std_logic; attribute dont_touch of N2585GAT: signal is true;
	signal N2586GAT: std_logic; attribute dont_touch of N2586GAT: signal is true;
	signal N2588GAT: std_logic; attribute dont_touch of N2588GAT: signal is true;
	signal N2590GAT: std_logic; attribute dont_touch of N2590GAT: signal is true;
	signal N2591GAT: std_logic; attribute dont_touch of N2591GAT: signal is true;
	signal N2592GAT: std_logic; attribute dont_touch of N2592GAT: signal is true;
	signal N2594GAT: std_logic; attribute dont_touch of N2594GAT: signal is true;
	signal N2595GAT: std_logic; attribute dont_touch of N2595GAT: signal is true;
	signal N2596GAT: std_logic; attribute dont_touch of N2596GAT: signal is true;
	signal N2597GAT: std_logic; attribute dont_touch of N2597GAT: signal is true;
	signal N2599GAT: std_logic; attribute dont_touch of N2599GAT: signal is true;
	signal N2601GAT: std_logic; attribute dont_touch of N2601GAT: signal is true;
	signal N2602GAT: std_logic; attribute dont_touch of N2602GAT: signal is true;
	signal N2603GAT: std_logic; attribute dont_touch of N2603GAT: signal is true;
	signal N2604GAT: std_logic; attribute dont_touch of N2604GAT: signal is true;
	signal N2605GAT: std_logic; attribute dont_touch of N2605GAT: signal is true;
	signal N2606GAT: std_logic; attribute dont_touch of N2606GAT: signal is true;
	signal N2607GAT: std_logic; attribute dont_touch of N2607GAT: signal is true;
	signal N2608GAT: std_logic; attribute dont_touch of N2608GAT: signal is true;
	signal N2609GAT: std_logic; attribute dont_touch of N2609GAT: signal is true;
	signal N2610GAT: std_logic; attribute dont_touch of N2610GAT: signal is true;
	signal N2611GAT: std_logic; attribute dont_touch of N2611GAT: signal is true;
	signal N2612GAT: std_logic; attribute dont_touch of N2612GAT: signal is true;
	signal N2613GAT: std_logic; attribute dont_touch of N2613GAT: signal is true;
	signal N2614GAT: std_logic; attribute dont_touch of N2614GAT: signal is true;
	signal N2615GAT: std_logic; attribute dont_touch of N2615GAT: signal is true;
	signal N2616GAT: std_logic; attribute dont_touch of N2616GAT: signal is true;
	signal N2617GAT: std_logic; attribute dont_touch of N2617GAT: signal is true;
	signal N2619GAT: std_logic; attribute dont_touch of N2619GAT: signal is true;
	signal N2620GAT: std_logic; attribute dont_touch of N2620GAT: signal is true;
	signal N2621GAT: std_logic; attribute dont_touch of N2621GAT: signal is true;
	signal N2622GAT: std_logic; attribute dont_touch of N2622GAT: signal is true;
	signal N2624GAT: std_logic; attribute dont_touch of N2624GAT: signal is true;
	signal N2625GAT: std_logic; attribute dont_touch of N2625GAT: signal is true;
	signal N2626GAT: std_logic; attribute dont_touch of N2626GAT: signal is true;
	signal N2628GAT: std_logic; attribute dont_touch of N2628GAT: signal is true;
	signal N2629GAT: std_logic; attribute dont_touch of N2629GAT: signal is true;
	signal N2630GAT: std_logic; attribute dont_touch of N2630GAT: signal is true;
	signal N2632GAT: std_logic; attribute dont_touch of N2632GAT: signal is true;
	signal N2633GAT: std_logic; attribute dont_touch of N2633GAT: signal is true;
	signal N2634GAT: std_logic; attribute dont_touch of N2634GAT: signal is true;
	signal N2636GAT: std_logic; attribute dont_touch of N2636GAT: signal is true;
	signal N2637GAT: std_logic; attribute dont_touch of N2637GAT: signal is true;
	signal N2638GAT: std_logic; attribute dont_touch of N2638GAT: signal is true;
	signal N2639GAT: std_logic; attribute dont_touch of N2639GAT: signal is true;
	signal N2640GAT: std_logic; attribute dont_touch of N2640GAT: signal is true;
	signal N2642GAT: std_logic; attribute dont_touch of N2642GAT: signal is true;
	signal N2643GAT: std_logic; attribute dont_touch of N2643GAT: signal is true;
	signal N2644GAT: std_logic; attribute dont_touch of N2644GAT: signal is true;
	signal N2646GAT: std_logic; attribute dont_touch of N2646GAT: signal is true;
	signal N2647GAT: std_logic; attribute dont_touch of N2647GAT: signal is true;
	signal N2648GAT: std_logic; attribute dont_touch of N2648GAT: signal is true;
	signal N2649GAT: std_logic; attribute dont_touch of N2649GAT: signal is true;
	signal N2650GAT: std_logic; attribute dont_touch of N2650GAT: signal is true;
	signal N2652GAT: std_logic; attribute dont_touch of N2652GAT: signal is true;
	signal N2655GAT: std_logic; attribute dont_touch of N2655GAT: signal is true;
	signal N2656GAT: std_logic; attribute dont_touch of N2656GAT: signal is true;
	signal N2658GAT: std_logic; attribute dont_touch of N2658GAT: signal is true;
	signal N2660GAT: std_logic; attribute dont_touch of N2660GAT: signal is true;
	signal N2661GAT: std_logic; attribute dont_touch of N2661GAT: signal is true;
	signal N2662GAT: std_logic; attribute dont_touch of N2662GAT: signal is true;
	signal N2663GAT: std_logic; attribute dont_touch of N2663GAT: signal is true;
	signal N2664GAT: std_logic; attribute dont_touch of N2664GAT: signal is true;
	signal N2665GAT: std_logic; attribute dont_touch of N2665GAT: signal is true;
	signal N2666GAT: std_logic; attribute dont_touch of N2666GAT: signal is true;
	signal N2667GAT: std_logic; attribute dont_touch of N2667GAT: signal is true;
	signal N2668GAT: std_logic; attribute dont_touch of N2668GAT: signal is true;
	signal N2669GAT: std_logic; attribute dont_touch of N2669GAT: signal is true;
	signal N2670GAT: std_logic; attribute dont_touch of N2670GAT: signal is true;
	signal N2671GAT: std_logic; attribute dont_touch of N2671GAT: signal is true;
	signal N2672GAT: std_logic; attribute dont_touch of N2672GAT: signal is true;
	signal N2673GAT: std_logic; attribute dont_touch of N2673GAT: signal is true;
	signal N2674GAT: std_logic; attribute dont_touch of N2674GAT: signal is true;
	signal N2677GAT: std_logic; attribute dont_touch of N2677GAT: signal is true;
	signal N2678GAT: std_logic; attribute dont_touch of N2678GAT: signal is true;
	signal N2679GAT: std_logic; attribute dont_touch of N2679GAT: signal is true;
	signal N2680GAT: std_logic; attribute dont_touch of N2680GAT: signal is true;
	signal N2681GAT: std_logic; attribute dont_touch of N2681GAT: signal is true;
	signal N2682GAT: std_logic; attribute dont_touch of N2682GAT: signal is true;
	signal N2683GAT: std_logic; attribute dont_touch of N2683GAT: signal is true;
	signal N2684GAT: std_logic; attribute dont_touch of N2684GAT: signal is true;
	signal N2685GAT: std_logic; attribute dont_touch of N2685GAT: signal is true;
	signal N2686GAT: std_logic; attribute dont_touch of N2686GAT: signal is true;
	signal N2687GAT: std_logic; attribute dont_touch of N2687GAT: signal is true;
	signal N2688GAT: std_logic; attribute dont_touch of N2688GAT: signal is true;
	signal N2689GAT: std_logic; attribute dont_touch of N2689GAT: signal is true;
	signal N2690GAT: std_logic; attribute dont_touch of N2690GAT: signal is true;
	signal N2691GAT: std_logic; attribute dont_touch of N2691GAT: signal is true;
	signal N2692GAT: std_logic; attribute dont_touch of N2692GAT: signal is true;
	signal N2693GAT: std_logic; attribute dont_touch of N2693GAT: signal is true;
	signal N2694GAT: std_logic; attribute dont_touch of N2694GAT: signal is true;
	signal N2695GAT: std_logic; attribute dont_touch of N2695GAT: signal is true;
	signal N2696GAT: std_logic; attribute dont_touch of N2696GAT: signal is true;
	signal N2697GAT: std_logic; attribute dont_touch of N2697GAT: signal is true;
	signal N2698GAT: std_logic; attribute dont_touch of N2698GAT: signal is true;
	signal N2699GAT: std_logic; attribute dont_touch of N2699GAT: signal is true;
	signal N2700GAT: std_logic; attribute dont_touch of N2700GAT: signal is true;
	signal N2701GAT: std_logic; attribute dont_touch of N2701GAT: signal is true;
	signal N2702GAT: std_logic; attribute dont_touch of N2702GAT: signal is true;
	signal N2703GAT: std_logic; attribute dont_touch of N2703GAT: signal is true;
	signal N2704GAT: std_logic; attribute dont_touch of N2704GAT: signal is true;
	signal N2705GAT: std_logic; attribute dont_touch of N2705GAT: signal is true;
	signal N2706GAT: std_logic; attribute dont_touch of N2706GAT: signal is true;
	signal N2707GAT: std_logic; attribute dont_touch of N2707GAT: signal is true;
	signal N2708GAT: std_logic; attribute dont_touch of N2708GAT: signal is true;
	signal N2709GAT: std_logic; attribute dont_touch of N2709GAT: signal is true;
	signal N2710GAT: std_logic; attribute dont_touch of N2710GAT: signal is true;
	signal N2711GAT: std_logic; attribute dont_touch of N2711GAT: signal is true;
	signal N2712GAT: std_logic; attribute dont_touch of N2712GAT: signal is true;
	signal N2715GAT: std_logic; attribute dont_touch of N2715GAT: signal is true;
	signal N2716GAT: std_logic; attribute dont_touch of N2716GAT: signal is true;
	signal N2717GAT: std_logic; attribute dont_touch of N2717GAT: signal is true;
	signal N2718GAT: std_logic; attribute dont_touch of N2718GAT: signal is true;
	signal N2719GAT: std_logic; attribute dont_touch of N2719GAT: signal is true;
	signal N2720GAT: std_logic; attribute dont_touch of N2720GAT: signal is true;
	signal N2721GAT: std_logic; attribute dont_touch of N2721GAT: signal is true;
	signal N2722GAT: std_logic; attribute dont_touch of N2722GAT: signal is true;
	signal N2723GAT: std_logic; attribute dont_touch of N2723GAT: signal is true;
	signal N2724GAT: std_logic; attribute dont_touch of N2724GAT: signal is true;
	signal N2725GAT: std_logic; attribute dont_touch of N2725GAT: signal is true;
	signal N2726GAT: std_logic; attribute dont_touch of N2726GAT: signal is true;
	signal N2727GAT: std_logic; attribute dont_touch of N2727GAT: signal is true;
	signal N2728GAT: std_logic; attribute dont_touch of N2728GAT: signal is true;
	signal N2729GAT: std_logic; attribute dont_touch of N2729GAT: signal is true;
	signal N2730GAT: std_logic; attribute dont_touch of N2730GAT: signal is true;
	signal N2731GAT: std_logic; attribute dont_touch of N2731GAT: signal is true;
	signal N2732GAT: std_logic; attribute dont_touch of N2732GAT: signal is true;
	signal N2733GAT: std_logic; attribute dont_touch of N2733GAT: signal is true;
	signal N2734GAT: std_logic; attribute dont_touch of N2734GAT: signal is true;
	signal N2735GAT: std_logic; attribute dont_touch of N2735GAT: signal is true;
	signal N2736GAT: std_logic; attribute dont_touch of N2736GAT: signal is true;
	signal N2737GAT: std_logic; attribute dont_touch of N2737GAT: signal is true;
	signal N2738GAT: std_logic; attribute dont_touch of N2738GAT: signal is true;
	signal N2739GAT: std_logic; attribute dont_touch of N2739GAT: signal is true;
	signal N2740GAT: std_logic; attribute dont_touch of N2740GAT: signal is true;
	signal N2741GAT: std_logic; attribute dont_touch of N2741GAT: signal is true;
	signal N2742GAT: std_logic; attribute dont_touch of N2742GAT: signal is true;
	signal N2743GAT: std_logic; attribute dont_touch of N2743GAT: signal is true;
	signal N2744GAT: std_logic; attribute dont_touch of N2744GAT: signal is true;
	signal N2745GAT: std_logic; attribute dont_touch of N2745GAT: signal is true;
	signal N2746GAT: std_logic; attribute dont_touch of N2746GAT: signal is true;
	signal N2747GAT: std_logic; attribute dont_touch of N2747GAT: signal is true;
	signal N2748GAT: std_logic; attribute dont_touch of N2748GAT: signal is true;
	signal N2749GAT: std_logic; attribute dont_touch of N2749GAT: signal is true;
	signal N2750GAT: std_logic; attribute dont_touch of N2750GAT: signal is true;
	signal N2751GAT: std_logic; attribute dont_touch of N2751GAT: signal is true;
	signal N2752GAT: std_logic; attribute dont_touch of N2752GAT: signal is true;
	signal N2753GAT: std_logic; attribute dont_touch of N2753GAT: signal is true;
	signal N2754GAT: std_logic; attribute dont_touch of N2754GAT: signal is true;
	signal N2755GAT: std_logic; attribute dont_touch of N2755GAT: signal is true;
	signal N2756GAT: std_logic; attribute dont_touch of N2756GAT: signal is true;
	signal N2757GAT: std_logic; attribute dont_touch of N2757GAT: signal is true;
	signal N2758GAT: std_logic; attribute dont_touch of N2758GAT: signal is true;
	signal N2759GAT: std_logic; attribute dont_touch of N2759GAT: signal is true;
	signal N2760GAT: std_logic; attribute dont_touch of N2760GAT: signal is true;
	signal N2761GAT: std_logic; attribute dont_touch of N2761GAT: signal is true;
	signal N2762GAT: std_logic; attribute dont_touch of N2762GAT: signal is true;
	signal N2763GAT: std_logic; attribute dont_touch of N2763GAT: signal is true;
	signal N2764GAT: std_logic; attribute dont_touch of N2764GAT: signal is true;
	signal N2765GAT: std_logic; attribute dont_touch of N2765GAT: signal is true;
	signal N2766GAT: std_logic; attribute dont_touch of N2766GAT: signal is true;
	signal N2767GAT: std_logic; attribute dont_touch of N2767GAT: signal is true;
	signal N2768GAT: std_logic; attribute dont_touch of N2768GAT: signal is true;
	signal N2775GAT: std_logic; attribute dont_touch of N2775GAT: signal is true;
	signal N2776GAT: std_logic; attribute dont_touch of N2776GAT: signal is true;
	signal N2777GAT: std_logic; attribute dont_touch of N2777GAT: signal is true;
	signal N2778GAT: std_logic; attribute dont_touch of N2778GAT: signal is true;
	signal N2779GAT: std_logic; attribute dont_touch of N2779GAT: signal is true;
	signal N2780GAT: std_logic; attribute dont_touch of N2780GAT: signal is true;
	signal N2781GAT: std_logic; attribute dont_touch of N2781GAT: signal is true;
	signal N2782GAT: std_logic; attribute dont_touch of N2782GAT: signal is true;
	signal N2783GAT: std_logic; attribute dont_touch of N2783GAT: signal is true;
	signal N2784GAT: std_logic; attribute dont_touch of N2784GAT: signal is true;
	signal N2785GAT: std_logic; attribute dont_touch of N2785GAT: signal is true;
	signal N2786GAT: std_logic; attribute dont_touch of N2786GAT: signal is true;
	signal N2789GAT: std_logic; attribute dont_touch of N2789GAT: signal is true;
	signal N2790GAT: std_logic; attribute dont_touch of N2790GAT: signal is true;
	signal N2791GAT: std_logic; attribute dont_touch of N2791GAT: signal is true;
	signal N2792GAT: std_logic; attribute dont_touch of N2792GAT: signal is true;
	signal N2793GAT: std_logic; attribute dont_touch of N2793GAT: signal is true;
	signal N2794GAT: std_logic; attribute dont_touch of N2794GAT: signal is true;
	signal N2795GAT: std_logic; attribute dont_touch of N2795GAT: signal is true;
	signal N2796GAT: std_logic; attribute dont_touch of N2796GAT: signal is true;
	signal N2797GAT: std_logic; attribute dont_touch of N2797GAT: signal is true;
	signal N2798GAT: std_logic; attribute dont_touch of N2798GAT: signal is true;
	signal N2799GAT: std_logic; attribute dont_touch of N2799GAT: signal is true;
	signal N2800GAT: std_logic; attribute dont_touch of N2800GAT: signal is true;
	signal N2801GAT: std_logic; attribute dont_touch of N2801GAT: signal is true;
	signal N2802GAT: std_logic; attribute dont_touch of N2802GAT: signal is true;
	signal N2803GAT: std_logic; attribute dont_touch of N2803GAT: signal is true;
	signal N2804GAT: std_logic; attribute dont_touch of N2804GAT: signal is true;
	signal N2805GAT: std_logic; attribute dont_touch of N2805GAT: signal is true;
	signal N2806GAT: std_logic; attribute dont_touch of N2806GAT: signal is true;
	signal N2807GAT: std_logic; attribute dont_touch of N2807GAT: signal is true;
	signal N2808GAT: std_logic; attribute dont_touch of N2808GAT: signal is true;
	signal N2809GAT: std_logic; attribute dont_touch of N2809GAT: signal is true;
	signal N2810GAT: std_logic; attribute dont_touch of N2810GAT: signal is true;
	signal N2811GAT: std_logic; attribute dont_touch of N2811GAT: signal is true;
	signal N2812GAT: std_logic; attribute dont_touch of N2812GAT: signal is true;
	signal N2813GAT: std_logic; attribute dont_touch of N2813GAT: signal is true;
	signal N2814GAT: std_logic; attribute dont_touch of N2814GAT: signal is true;
	signal N2815GAT: std_logic; attribute dont_touch of N2815GAT: signal is true;
	signal N2816GAT: std_logic; attribute dont_touch of N2816GAT: signal is true;
	signal N2817GAT: std_logic; attribute dont_touch of N2817GAT: signal is true;
	signal N2818GAT: std_logic; attribute dont_touch of N2818GAT: signal is true;
	signal N2819GAT: std_logic; attribute dont_touch of N2819GAT: signal is true;
	signal N2820GAT: std_logic; attribute dont_touch of N2820GAT: signal is true;
	signal N2821GAT: std_logic; attribute dont_touch of N2821GAT: signal is true;
	signal N2822GAT: std_logic; attribute dont_touch of N2822GAT: signal is true;
	signal N2823GAT: std_logic; attribute dont_touch of N2823GAT: signal is true;
	signal N2824GAT: std_logic; attribute dont_touch of N2824GAT: signal is true;
	signal N2825GAT: std_logic; attribute dont_touch of N2825GAT: signal is true;
	signal N2826GAT: std_logic; attribute dont_touch of N2826GAT: signal is true;
	signal N2827GAT: std_logic; attribute dont_touch of N2827GAT: signal is true;
	signal N2828GAT: std_logic; attribute dont_touch of N2828GAT: signal is true;
	signal N2829GAT: std_logic; attribute dont_touch of N2829GAT: signal is true;
	signal N2830GAT: std_logic; attribute dont_touch of N2830GAT: signal is true;
	signal N2831GAT: std_logic; attribute dont_touch of N2831GAT: signal is true;
	signal N2832GAT: std_logic; attribute dont_touch of N2832GAT: signal is true;
	signal N2836GAT: std_logic; attribute dont_touch of N2836GAT: signal is true;
	signal N2837GAT: std_logic; attribute dont_touch of N2837GAT: signal is true;
	signal N2838GAT: std_logic; attribute dont_touch of N2838GAT: signal is true;
	signal N2839GAT: std_logic; attribute dont_touch of N2839GAT: signal is true;
	signal N2840GAT: std_logic; attribute dont_touch of N2840GAT: signal is true;
	signal N2841GAT: std_logic; attribute dont_touch of N2841GAT: signal is true;
	signal N2842GAT: std_logic; attribute dont_touch of N2842GAT: signal is true;
	signal N2843GAT: std_logic; attribute dont_touch of N2843GAT: signal is true;
	signal N2844GAT: std_logic; attribute dont_touch of N2844GAT: signal is true;
	signal N2845GAT: std_logic; attribute dont_touch of N2845GAT: signal is true;
	signal N2846GAT: std_logic; attribute dont_touch of N2846GAT: signal is true;
	signal N2847GAT: std_logic; attribute dont_touch of N2847GAT: signal is true;
	signal N2850GAT: std_logic; attribute dont_touch of N2850GAT: signal is true;
	signal N2851GAT: std_logic; attribute dont_touch of N2851GAT: signal is true;
	signal N2852GAT: std_logic; attribute dont_touch of N2852GAT: signal is true;
	signal N2853GAT: std_logic; attribute dont_touch of N2853GAT: signal is true;
	signal N2854GAT: std_logic; attribute dont_touch of N2854GAT: signal is true;
	signal N2855GAT: std_logic; attribute dont_touch of N2855GAT: signal is true;
	signal N2856GAT: std_logic; attribute dont_touch of N2856GAT: signal is true;
	signal N2857GAT: std_logic; attribute dont_touch of N2857GAT: signal is true;
	signal N2858GAT: std_logic; attribute dont_touch of N2858GAT: signal is true;
	signal N2859GAT: std_logic; attribute dont_touch of N2859GAT: signal is true;
	signal N2860GAT: std_logic; attribute dont_touch of N2860GAT: signal is true;
	signal N2861GAT: std_logic; attribute dont_touch of N2861GAT: signal is true;
	signal N2862GAT: std_logic; attribute dont_touch of N2862GAT: signal is true;
	signal N2863GAT: std_logic; attribute dont_touch of N2863GAT: signal is true;
	signal N2864GAT: std_logic; attribute dont_touch of N2864GAT: signal is true;
	signal N2867GAT: std_logic; attribute dont_touch of N2867GAT: signal is true;
	signal N2868GAT: std_logic; attribute dont_touch of N2868GAT: signal is true;
	signal N2869GAT: std_logic; attribute dont_touch of N2869GAT: signal is true;
	signal N2874GAT: std_logic; attribute dont_touch of N2874GAT: signal is true;
	signal N2875GAT: std_logic; attribute dont_touch of N2875GAT: signal is true;
	signal N2876GAT: std_logic; attribute dont_touch of N2876GAT: signal is true;
	signal N2877GAT: std_logic; attribute dont_touch of N2877GAT: signal is true;
	signal N2878GAT: std_logic; attribute dont_touch of N2878GAT: signal is true;
	signal N2879GAT: std_logic; attribute dont_touch of N2879GAT: signal is true;
	signal N2880GAT: std_logic; attribute dont_touch of N2880GAT: signal is true;
	signal N2881GAT: std_logic; attribute dont_touch of N2881GAT: signal is true;
	signal N2882GAT: std_logic; attribute dont_touch of N2882GAT: signal is true;
	signal N2883GAT: std_logic; attribute dont_touch of N2883GAT: signal is true;
	signal N2884GAT: std_logic; attribute dont_touch of N2884GAT: signal is true;
	signal N2885GAT: std_logic; attribute dont_touch of N2885GAT: signal is true;
	signal N2886GAT: std_logic; attribute dont_touch of N2886GAT: signal is true;
	signal N2887GAT: std_logic; attribute dont_touch of N2887GAT: signal is true;
	signal N2888GAT: std_logic; attribute dont_touch of N2888GAT: signal is true;
	signal N2889GAT: std_logic; attribute dont_touch of N2889GAT: signal is true;
	signal N2890GAT: std_logic; attribute dont_touch of N2890GAT: signal is true;
	signal N2891GAT: std_logic; attribute dont_touch of N2891GAT: signal is true;
	signal N2892GAT: std_logic; attribute dont_touch of N2892GAT: signal is true;
	signal N2893GAT: std_logic; attribute dont_touch of N2893GAT: signal is true;
	signal N2894GAT: std_logic; attribute dont_touch of N2894GAT: signal is true;
	signal N2895GAT: std_logic; attribute dont_touch of N2895GAT: signal is true;
	signal N2896GAT: std_logic; attribute dont_touch of N2896GAT: signal is true;
	signal N2897GAT: std_logic; attribute dont_touch of N2897GAT: signal is true;
	signal N2898GAT: std_logic; attribute dont_touch of N2898GAT: signal is true;
	signal N2899GAT: std_logic; attribute dont_touch of N2899GAT: signal is true;
	signal N2900GAT: std_logic; attribute dont_touch of N2900GAT: signal is true;
	signal N2901GAT: std_logic; attribute dont_touch of N2901GAT: signal is true;
	signal N2902GAT: std_logic; attribute dont_touch of N2902GAT: signal is true;
	signal N2903GAT: std_logic; attribute dont_touch of N2903GAT: signal is true;
	signal N2904GAT: std_logic; attribute dont_touch of N2904GAT: signal is true;
	signal N2905GAT: std_logic; attribute dont_touch of N2905GAT: signal is true;
	signal N2906GAT: std_logic; attribute dont_touch of N2906GAT: signal is true;
	signal N2907GAT: std_logic; attribute dont_touch of N2907GAT: signal is true;
	signal N2908GAT: std_logic; attribute dont_touch of N2908GAT: signal is true;
	signal N2909GAT: std_logic; attribute dont_touch of N2909GAT: signal is true;
	signal N2910GAT: std_logic; attribute dont_touch of N2910GAT: signal is true;
	signal N2911GAT: std_logic; attribute dont_touch of N2911GAT: signal is true;
	signal N2912GAT: std_logic; attribute dont_touch of N2912GAT: signal is true;
	signal N2913GAT: std_logic; attribute dont_touch of N2913GAT: signal is true;
	signal N2914GAT: std_logic; attribute dont_touch of N2914GAT: signal is true;
	signal N2915GAT: std_logic; attribute dont_touch of N2915GAT: signal is true;
	signal N2916GAT: std_logic; attribute dont_touch of N2916GAT: signal is true;
	signal N2917GAT: std_logic; attribute dont_touch of N2917GAT: signal is true;
	signal N2918GAT: std_logic; attribute dont_touch of N2918GAT: signal is true;
	signal N2919GAT: std_logic; attribute dont_touch of N2919GAT: signal is true;
	signal N2920GAT: std_logic; attribute dont_touch of N2920GAT: signal is true;
	signal N2921GAT: std_logic; attribute dont_touch of N2921GAT: signal is true;
	signal N2922GAT: std_logic; attribute dont_touch of N2922GAT: signal is true;
	signal N2923GAT: std_logic; attribute dont_touch of N2923GAT: signal is true;
	signal N2924GAT: std_logic; attribute dont_touch of N2924GAT: signal is true;
	signal N2925GAT: std_logic; attribute dont_touch of N2925GAT: signal is true;
	signal N2926GAT: std_logic; attribute dont_touch of N2926GAT: signal is true;
	signal N2927GAT: std_logic; attribute dont_touch of N2927GAT: signal is true;
	signal N2928GAT: std_logic; attribute dont_touch of N2928GAT: signal is true;
	signal N2929GAT: std_logic; attribute dont_touch of N2929GAT: signal is true;
	signal N2930GAT: std_logic; attribute dont_touch of N2930GAT: signal is true;
	signal N2931GAT: std_logic; attribute dont_touch of N2931GAT: signal is true;
	signal N2932GAT: std_logic; attribute dont_touch of N2932GAT: signal is true;
	signal N2933GAT: std_logic; attribute dont_touch of N2933GAT: signal is true;
	signal N2934GAT: std_logic; attribute dont_touch of N2934GAT: signal is true;
	signal N2935GAT: std_logic; attribute dont_touch of N2935GAT: signal is true;
	signal N2936GAT: std_logic; attribute dont_touch of N2936GAT: signal is true;
	signal N2937GAT: std_logic; attribute dont_touch of N2937GAT: signal is true;
	signal N2938GAT: std_logic; attribute dont_touch of N2938GAT: signal is true;
	signal N2939GAT: std_logic; attribute dont_touch of N2939GAT: signal is true;
	signal N2940GAT: std_logic; attribute dont_touch of N2940GAT: signal is true;
	signal N2941GAT: std_logic; attribute dont_touch of N2941GAT: signal is true;
	signal N2942GAT: std_logic; attribute dont_touch of N2942GAT: signal is true;
	signal N2943GAT: std_logic; attribute dont_touch of N2943GAT: signal is true;
	signal N2944GAT: std_logic; attribute dont_touch of N2944GAT: signal is true;
	signal N2945GAT: std_logic; attribute dont_touch of N2945GAT: signal is true;
	signal N2946GAT: std_logic; attribute dont_touch of N2946GAT: signal is true;
	signal N2947GAT: std_logic; attribute dont_touch of N2947GAT: signal is true;
	signal N2948GAT: std_logic; attribute dont_touch of N2948GAT: signal is true;
	signal N2949GAT: std_logic; attribute dont_touch of N2949GAT: signal is true;
	signal N2950GAT: std_logic; attribute dont_touch of N2950GAT: signal is true;
	signal N2951GAT: std_logic; attribute dont_touch of N2951GAT: signal is true;
	signal N2952GAT: std_logic; attribute dont_touch of N2952GAT: signal is true;
	signal N2953GAT: std_logic; attribute dont_touch of N2953GAT: signal is true;
	signal N2954GAT: std_logic; attribute dont_touch of N2954GAT: signal is true;
	signal N2955GAT: std_logic; attribute dont_touch of N2955GAT: signal is true;
	signal N2956GAT: std_logic; attribute dont_touch of N2956GAT: signal is true;
	signal N2957GAT: std_logic; attribute dont_touch of N2957GAT: signal is true;
	signal N2958GAT: std_logic; attribute dont_touch of N2958GAT: signal is true;
	signal N2959GAT: std_logic; attribute dont_touch of N2959GAT: signal is true;
	signal N2960GAT: std_logic; attribute dont_touch of N2960GAT: signal is true;
	signal N2961GAT: std_logic; attribute dont_touch of N2961GAT: signal is true;
	signal N2962GAT: std_logic; attribute dont_touch of N2962GAT: signal is true;
	signal N2963GAT: std_logic; attribute dont_touch of N2963GAT: signal is true;
	signal N2964GAT: std_logic; attribute dont_touch of N2964GAT: signal is true;
	signal N2965GAT: std_logic; attribute dont_touch of N2965GAT: signal is true;
	signal N2966GAT: std_logic; attribute dont_touch of N2966GAT: signal is true;
	signal N2967GAT: std_logic; attribute dont_touch of N2967GAT: signal is true;
	signal N2968GAT: std_logic; attribute dont_touch of N2968GAT: signal is true;
	signal N2969GAT: std_logic; attribute dont_touch of N2969GAT: signal is true;
	signal N2970GAT: std_logic; attribute dont_touch of N2970GAT: signal is true;
	signal N2971GAT: std_logic; attribute dont_touch of N2971GAT: signal is true;
	signal N2973GAT: std_logic; attribute dont_touch of N2973GAT: signal is true;
	signal N2974GAT: std_logic; attribute dont_touch of N2974GAT: signal is true;
	signal N2975GAT: std_logic; attribute dont_touch of N2975GAT: signal is true;
	signal N2977GAT: std_logic; attribute dont_touch of N2977GAT: signal is true;
	signal N2978GAT: std_logic; attribute dont_touch of N2978GAT: signal is true;
	signal N2979GAT: std_logic; attribute dont_touch of N2979GAT: signal is true;
	signal N2980GAT: std_logic; attribute dont_touch of N2980GAT: signal is true;
	signal N2981GAT: std_logic; attribute dont_touch of N2981GAT: signal is true;
	signal N2982GAT: std_logic; attribute dont_touch of N2982GAT: signal is true;
	signal N2983GAT: std_logic; attribute dont_touch of N2983GAT: signal is true;
	signal N2984GAT: std_logic; attribute dont_touch of N2984GAT: signal is true;
	signal N2985GAT: std_logic; attribute dont_touch of N2985GAT: signal is true;
	signal N2986GAT: std_logic; attribute dont_touch of N2986GAT: signal is true;
	signal N2987GAT: std_logic; attribute dont_touch of N2987GAT: signal is true;
	signal N2988GAT: std_logic; attribute dont_touch of N2988GAT: signal is true;
	signal N2989GAT: std_logic; attribute dont_touch of N2989GAT: signal is true;
	signal N2990GAT: std_logic; attribute dont_touch of N2990GAT: signal is true;
	signal N2991GAT: std_logic; attribute dont_touch of N2991GAT: signal is true;
	signal N2992GAT: std_logic; attribute dont_touch of N2992GAT: signal is true;
	signal N2993GAT: std_logic; attribute dont_touch of N2993GAT: signal is true;
	signal N2994GAT: std_logic; attribute dont_touch of N2994GAT: signal is true;
	signal N2995GAT: std_logic; attribute dont_touch of N2995GAT: signal is true;
	signal N2996GAT: std_logic; attribute dont_touch of N2996GAT: signal is true;
	signal N2997GAT: std_logic; attribute dont_touch of N2997GAT: signal is true;
	signal N2998GAT: std_logic; attribute dont_touch of N2998GAT: signal is true;
	signal N2999GAT: std_logic; attribute dont_touch of N2999GAT: signal is true;
	signal N3000GAT: std_logic; attribute dont_touch of N3000GAT: signal is true;
	signal N3001GAT: std_logic; attribute dont_touch of N3001GAT: signal is true;
	signal N3002GAT: std_logic; attribute dont_touch of N3002GAT: signal is true;
	signal N3003GAT: std_logic; attribute dont_touch of N3003GAT: signal is true;
	signal N3004GAT: std_logic; attribute dont_touch of N3004GAT: signal is true;
	signal N3005GAT: std_logic; attribute dont_touch of N3005GAT: signal is true;
	signal N3006GAT: std_logic; attribute dont_touch of N3006GAT: signal is true;
	signal N3007GAT: std_logic; attribute dont_touch of N3007GAT: signal is true;
	signal N3008GAT: std_logic; attribute dont_touch of N3008GAT: signal is true;
	signal N3009GAT: std_logic; attribute dont_touch of N3009GAT: signal is true;
	signal N3010GAT: std_logic; attribute dont_touch of N3010GAT: signal is true;
	signal N3011GAT: std_logic; attribute dont_touch of N3011GAT: signal is true;
	signal N3013GAT: std_logic; attribute dont_touch of N3013GAT: signal is true;
	signal N3014GAT: std_logic; attribute dont_touch of N3014GAT: signal is true;
	signal N3015GAT: std_logic; attribute dont_touch of N3015GAT: signal is true;
	signal N3016GAT: std_logic; attribute dont_touch of N3016GAT: signal is true;
	signal N3017GAT: std_logic; attribute dont_touch of N3017GAT: signal is true;
	signal N3018GAT: std_logic; attribute dont_touch of N3018GAT: signal is true;
	signal N3019GAT: std_logic; attribute dont_touch of N3019GAT: signal is true;
	signal N3020GAT: std_logic; attribute dont_touch of N3020GAT: signal is true;
	signal N3021GAT: std_logic; attribute dont_touch of N3021GAT: signal is true;
	signal N3022GAT: std_logic; attribute dont_touch of N3022GAT: signal is true;
	signal N3023GAT: std_logic; attribute dont_touch of N3023GAT: signal is true;
	signal N3024GAT: std_logic; attribute dont_touch of N3024GAT: signal is true;
	signal N3025GAT: std_logic; attribute dont_touch of N3025GAT: signal is true;
	signal N3026GAT: std_logic; attribute dont_touch of N3026GAT: signal is true;
	signal N3027GAT: std_logic; attribute dont_touch of N3027GAT: signal is true;
	signal N3028GAT: std_logic; attribute dont_touch of N3028GAT: signal is true;
	signal N3029GAT: std_logic; attribute dont_touch of N3029GAT: signal is true;
	signal N3030GAT: std_logic; attribute dont_touch of N3030GAT: signal is true;
	signal N3031GAT: std_logic; attribute dont_touch of N3031GAT: signal is true;
	signal N3032GAT: std_logic; attribute dont_touch of N3032GAT: signal is true;
	signal N3033GAT: std_logic; attribute dont_touch of N3033GAT: signal is true;
	signal N3034GAT: std_logic; attribute dont_touch of N3034GAT: signal is true;
	signal N3035GAT: std_logic; attribute dont_touch of N3035GAT: signal is true;
	signal N3036GAT: std_logic; attribute dont_touch of N3036GAT: signal is true;
	signal N3037GAT: std_logic; attribute dont_touch of N3037GAT: signal is true;
	signal N3038GAT: std_logic; attribute dont_touch of N3038GAT: signal is true;
	signal N3039GAT: std_logic; attribute dont_touch of N3039GAT: signal is true;
	signal N3040GAT: std_logic; attribute dont_touch of N3040GAT: signal is true;
	signal N3041GAT: std_logic; attribute dont_touch of N3041GAT: signal is true;
	signal N3042GAT: std_logic; attribute dont_touch of N3042GAT: signal is true;
	signal N3043GAT: std_logic; attribute dont_touch of N3043GAT: signal is true;
	signal N3044GAT: std_logic; attribute dont_touch of N3044GAT: signal is true;
	signal N3045GAT: std_logic; attribute dont_touch of N3045GAT: signal is true;
	signal N3046GAT: std_logic; attribute dont_touch of N3046GAT: signal is true;
	signal N3047GAT: std_logic; attribute dont_touch of N3047GAT: signal is true;
	signal N3048GAT: std_logic; attribute dont_touch of N3048GAT: signal is true;
	signal N3049GAT: std_logic; attribute dont_touch of N3049GAT: signal is true;
	signal N3050GAT: std_logic; attribute dont_touch of N3050GAT: signal is true;
	signal N3051GAT: std_logic; attribute dont_touch of N3051GAT: signal is true;
	signal N3052GAT: std_logic; attribute dont_touch of N3052GAT: signal is true;
	signal N3053GAT: std_logic; attribute dont_touch of N3053GAT: signal is true;
	signal N3054GAT: std_logic; attribute dont_touch of N3054GAT: signal is true;
	signal N3055GAT: std_logic; attribute dont_touch of N3055GAT: signal is true;
	signal N3056GAT: std_logic; attribute dont_touch of N3056GAT: signal is true;
	signal N3057GAT: std_logic; attribute dont_touch of N3057GAT: signal is true;
	signal N3058GAT: std_logic; attribute dont_touch of N3058GAT: signal is true;
	signal N3059GAT: std_logic; attribute dont_touch of N3059GAT: signal is true;
	signal N3060GAT: std_logic; attribute dont_touch of N3060GAT: signal is true;
	signal N3061GAT: std_logic; attribute dont_touch of N3061GAT: signal is true;
	signal N3062GAT: std_logic; attribute dont_touch of N3062GAT: signal is true;
	signal N3063GAT: std_logic; attribute dont_touch of N3063GAT: signal is true;
	signal N3064GAT: std_logic; attribute dont_touch of N3064GAT: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			N148GAT<=N832GAT;
			N152GAT<=N705GAT;
			N156GAT<=N612GAT;
			N160GAT<=N2776GAT;
			N165GAT<=N2776GAT;
			N256GAT<=N836GAT;
			N271GAT<=N2732GAT;
			N275GAT<=N2779GAT;
			N279GAT<=N2735GAT;
			N283GAT<=N2732GAT;
			N314GAT<=N2886GAT;
			N318GAT<=N2887GAT;
			N322GAT<=N2888GAT;
			N327GAT<=N682GAT;
			N331GAT<=N822GAT;
			N337GAT<=N2735GAT;
			N341GAT<=N2779GAT;
			N366GAT<=N2890GAT;
			N384GAT<=N697GAT;
			N388GAT<=N881GAT;
			N394GAT<=N2782GAT;
			N398GAT<=N2782GAT;
			N402GAT<=N2790GAT;
			N463GAT<=N818GAT;
			N470GAT<=N828GAT;
			N491GAT<=N2782GAT;
			N553GAT<=N2903GAT;
			N561GAT<=N2901GAT;
			N580GAT<=N2905GAT;
			N584GAT<=N2898GAT;
			N614GAT<=N3056GAT;
			N618GAT<=N2790GAT;
			N622GAT<=N2793GAT;
			N626GAT<=N2670GAT;
			N659GAT<=N2891GAT;
			N667GAT<=N2904GAT;
			N673GAT<=N2897GAT;
			N680GAT<=N2913GAT;
			N684GAT<=N3060GAT;
			N699GAT<=N3061GAT;
			N703GAT<=N2790GAT;
			N707GAT<=N3055GAT;
			N722GAT<=N2670GAT;
			N726GAT<=N2793GAT;
			N777GAT<=N2915GAT;
			N816GAT<=N2920GAT;
			N820GAT<=N3059GAT;
			N824GAT<=N3057GAT;
			N830GAT<=N3062GAT;
			N834GAT<=N3064GAT;
			N838GAT<=N3063GAT;
			N842GAT<=N2673GAT;
			N846GAT<=N2793GAT;
			N861GAT<=N2927GAT;
			N865GAT<=N2894GAT;
			N883GAT<=N3058GAT;
			N919GAT<=N2670GAT;
			N931GAT<=N2911GAT;
			N957GAT<=N2928GAT;
			N1026GAT<=N2673GAT;
			N1035GAT<=N2918GAT;
			N1045GAT<=N2909GAT;
			N1068GAT<=N2914GAT;
			N1072GAT<=N2919GAT;
			N1080GAT<=N2921GAT;
			N1121GAT<=N2952GAT;
			N1135GAT<=N2912GAT;
			N1148GAT<=N2895GAT;
			N1197GAT<=N2908GAT;
			N1226GAT<=N2907GAT;
			N1241GAT<=N2922GAT;
			N1282GAT<=N2910GAT;
			N1294GAT<=N2896GAT;
			N1298GAT<=N2897GAT;
			N1312GAT<=N1361GAT;
			N1316GAT<=N1431GAT;
			N1332GAT<=N1565GAT;
			N1336GAT<=N1391GAT;
			N1340GAT<=N1567GAT;
			N1363GAT<=N1314GAT;
			N1389GAT<=N1793GAT;
			N1394GAT<=N1516GAT;
			N1433GAT<=N2983GAT;
			N1456GAT<=N1564GAT;
			N1462GAT<=N1915GAT;
			N1496GAT<=N1392GAT;
			N1508GAT<=N1636GAT;
			N1525GAT<=N1632GAT;
			N1588GAT<=N1593GAT;
			N1596GAT<=N1800GAT;
			N1675GAT<=N1713GAT;
			N1678GAT<=N1712GAT;
			N1740GAT<=N1330GAT;
			N1748GAT<=N1927GAT;
			N1763GAT<=N1610GAT;
			N1767GAT<=N1626GAT;
			N1771GAT<=N1613GAT;
			N1775GAT<=N1696GAT;
			N1807GAT<=N1717GAT;
			N1821GAT<=N1827GAT;
			N1825GAT<=N1827GAT;
			N1829GAT<=N2027GAT;
			N1834GAT<=N1625GAT;
			N1850GAT<=N2628GAT;
			N1871GAT<=N2009GAT;
			N1880GAT<=N3052GAT;
			N1899GAT<=N2532GAT;
			N1975GAT<=N2632GAT;
			N2021GAT<=N1781GAT;
			N2025GAT<=N2017GAT;
			N2029GAT<=N1816GAT;
			N2033GAT<=N2035GAT;
			N2037GAT<=N2042GAT;
			N2040GAT<=N1777GAT;
			N2044GAT<=N2015GAT;
			N2061GAT<=N2557GAT;
			N2084GAT<=N1603GAT;
			N2091GAT<=N1685GAT;
			N2095GAT<=N827GAT;
			N2099GAT<=N2023GAT;
			N2102GAT<=N1606GAT;
			N2110GAT<=N2031GAT;
			N2117GAT<=N2119GAT;
			N2121GAT<=N2123GAT;
			N2125GAT<=N2108GAT;
			N2135GAT<=N2337GAT;
			N2139GAT<=N2487GAT;
			N2143GAT<=N2541GAT;
			N2155GAT<=N1858GAT;
			N2169GAT<=N2174GAT;
			N2176GAT<=N2093GAT;
			N2179GAT<=N1945GAT;
			N2182GAT<=N1836GAT;
			N2190GAT<=N2268GAT;
			N2203GAT<=N3051GAT;
			N2207GAT<=N3050GAT;
			N2262GAT<=N2388GAT;
			N2266GAT<=N2493GAT;
			N2270GAT<=N3031GAT;
			N2309GAT<=N3000GAT;
			N2319GAT<=N2470GAT;
			N2339GAT<=N3035GAT;
			N2343GAT<=N3049GAT;
			N2347GAT<=N2201GAT;
			N2390GAT<=N3034GAT;
			N2394GAT<=N2341GAT;
			N2399GAT<=N3048GAT;
			N2403GAT<=N2397GAT;
			N2407GAT<=N2205GAT;
			N2440GAT<=N2560GAT;
			N2446GAT<=N2661GAT;
			N2450GAT<=N2307GAT;
			N2454GAT<=N2163GAT;
			N2458GAT<=N2590GAT;
			N2464GAT<=N567GAT;
			N2468GAT<=N933GAT;
			N2472GAT<=N1620GAT;
			N2476GAT<=N55GAT;
			N2490GAT<=N3044GAT;
			N2495GAT<=N3036GAT;
			N2502GAT<=N2646GAT;
			N2506GAT<=N2613GAT;
			N2510GAT<=N748GAT;
			N2514GAT<=N2456GAT;
			N2518GAT<=N2971GAT;
			N2522GAT<=N43GAT;
			N2526GAT<=N504GAT;
			N2543GAT<=N3041GAT;
			N2562GAT<=N3047GAT;
			N2588GAT<=N3016GAT;
			N2592GAT<=N1773GAT;
			N2599GAT<=N3010GAT;
			N2622GAT<=N3042GAT;
			N2626GAT<=N3040GAT;
			N2630GAT<=N3037GAT;
			N2634GAT<=N3053GAT;
			N2640GAT<=N3054GAT;
			N2644GAT<=N2638GAT;
			N2658GAT<=N2579GAT;
		end if;
	end process;
	I1<= not N3088GAT;
	I5<= not N3087GAT;
	I11<= not N3093GAT;
	I14<= not N2768GAT;
	I18<= not N3072GAT;
	I23<= not N3081GAT;
	I27<= not N3095GAT;
	I30<= not N2668GAT;
	I44<= not N673GAT;
	I47<= not N3069GAT;
	I50<= not N2783GAT;
	I62<= not N3070GAT;
	I65<= not N2791GAT;
	I76<= not N402GAT;
	I81<= not N2671GAT;
	I92<= not N919GAT;
	I97<= not N3071GAT;
	I100<= not N2794GAT;
	I111<= not N846GAT;
	I149<= not N703GAT;
	I171<= not N726GAT;
	I178<= not N722GAT;
	I192<= not N3083GAT;
	I196<= not N2854GAT;
	I199<= not N3085GAT;
	I203<= not N2859GAT;
	I206<= not N3084GAT;
	I210<= not N2862GAT;
	I214<= not N2861GAT;
	I217<= not N2860GAT;
	I220<= not N2864GAT;
	I223<= not N2863GAT;
	I227<= not N2856GAT;
	I230<= not N2855GAT;
	I237<= not N640GAT;
	I240<= not N2717GAT;
	I243<= not N3089GAT;
	I248<= not N2869GAT;
	I253<= not N2906GAT;
	I256<= not N2725GAT;
	I259<= not N3086GAT;
	I264<= not N2728GAT;
	I270<= not N422GAT;
	I275<= not N747GAT;
	I278<= not N2889GAT;
	I282<= not N1213GAT;
	I297<= not N3065GAT;
	I300<= not N2733GAT;
	I311<= not N271GAT;
	I314<= not N270GAT;
	I317<= not N3067GAT;
	I320<= not N2777GAT;
	I331<= not N160GAT;
	I334<= not N159GAT;
	I337<= not N3066GAT;
	I340<= not N2736GAT;
	I351<= not N337GAT;
	I354<= not N336GAT;
	I359<= not N158GAT;
	I363<= not N335GAT;
	I368<= not N269GAT;
	I375<= not N41GAT;
	I378<= not N725GAT;
	I381<= not N3073GAT;
	I384<= not N2674GAT;
	I395<= not N842GAT;
	I398<= not N841GAT;
	I401<= not N721GAT;
	I406<= not N840GAT;
	I409<= not N720GAT;
	I414<= not N724GAT;
	I420<= not N1013GAT;
	I423<= not N3068GAT;
	I426<= not N2780GAT;
	I437<= not N341GAT;
	I440<= not N340GAT;
	I443<= not N702GAT;
	I446<= not N394GAT;
	I449<= not N393GAT;
	I453<= not N701GAT;
	I456<= not N392GAT;
	I461<= not N339GAT;
	I468<= not N42GAT;
	I473<= not N162GAT;
	I476<= not N475GAT;
	I480<= not N258GAT;
	I509<= not N3099GAT;
	I512<= not N2730GAT;
	I572<= not N1829GAT;
	I576<= not N3100GAT;
	I579<= not N2851GAT;
	I583<= not N2786GAT;
	I591<= not N3094GAT;
	I594<= not N2722GAT;
	I606<= not N283GAT;
	I609<= not N282GAT;
	I620<= not N165GAT;
	I623<= not N164GAT;
	I634<= not N279GAT;
	I637<= not N278GAT;
	I642<= not N163GAT;
	I646<= not N277GAT;
	I651<= not N281GAT;
	I658<= not N54GAT;
	I661<= not N845GAT;
	I672<= not N1026GAT;
	I675<= not N1025GAT;
	I678<= not N918GAT;
	I683<= not N1024GAT;
	I687<= not N917GAT;
	I692<= not N844GAT;
	I698<= not N906GAT;
	I709<= not N275GAT;
	I712<= not N274GAT;
	I715<= not N401GAT;
	I718<= not N398GAT;
	I721<= not N397GAT;
	I726<= not N400GAT;
	I729<= not N396GAT;
	I734<= not N273GAT;
	I741<= not N178GAT;
	I746<= not N66GAT;
	I749<= not N343GAT;
	I753<= not N167GAT;
	I768<= not N3090GAT;
	I771<= not N2832GAT;
	I776<= not N3074GAT;
	I790<= not N1068GAT;
	I793<= not N1067GAT;
	I796<= not N3076GAT;
	I812<= not N957GAT;
	I815<= not N956GAT;
	I818<= not N3075GAT;
	I834<= not N861GAT;
	I837<= not N860GAT;
	I842<= not N955GAT;
	I846<= not N859GAT;
	I851<= not N1066GAT;
	I858<= not N857GAT;
	I863<= not N3080GAT;
	I877<= not N1294GAT;
	I880<= not N1293GAT;
	I885<= not N3082GAT;
	I899<= not N1241GAT;
	I902<= not N1240GAT;
	I913<= not N1298GAT;
	I916<= not N1297GAT;
	I921<= not N1239GAT;
	I925<= not N1296GAT;
	I930<= not N1292GAT;
	I936<= not N1228GAT;
	I941<= not N3077GAT;
	I955<= not N865GAT;
	I958<= not N864GAT;
	I963<= not N3079GAT;
	I977<= not N1080GAT;
	I980<= not N1079GAT;
	I985<= not N3078GAT;
	I999<= not N1148GAT;
	I1002<= not N1147GAT;
	I1007<= not N1078GAT;
	I1011<= not N1146GAT;
	I1016<= not N863GAT;
	I1023<= not N928GAT;
	I1028<= not N858GAT;
	I1031<= not N1050GAT;
	I1035<= not N944GAT;
	I1067<= not N616GAT;
	I1079<= not N489GAT;
	I1082<= not N618GAT;
	I1085<= not N617GAT;
	I1088<= not N491GAT;
	I1091<= not N490GAT;
	I1103<= not N620GAT;
	I1115<= not N624GAT;
	I1118<= not N622GAT;
	I1121<= not N621GAT;
	I1124<= not N626GAT;
	I1127<= not N625GAT;
	I1138<= not N834GAT;
	I1141<= not N833GAT;
	I1152<= not N707GAT;
	I1155<= not N706GAT;
	I1166<= not N838GAT;
	I1169<= not N837GAT;
	I1174<= not N705GAT;
	I1178<= not N836GAT;
	I1183<= not N832GAT;
	I1190<= not N515GAT;
	I1201<= not N830GAT;
	I1204<= not N829GAT;
	I1209<= not N828GAT;
	I1216<= not N728GAT;
	I1227<= not N614GAT;
	I1230<= not N613GAT;
	I1236<= not N612GAT;
	I1243<= not N404GAT;
	I1248<= not N405GAT;
	I1251<= not N493GAT;
	I1255<= not N709GAT;
	I1302<= not N680GAT;
	I1305<= not N679GAT;
	I1319<= not N816GAT;
	I1322<= not N815GAT;
	I1336<= not N580GAT;
	I1339<= not N579GAT;
	I1344<= not N814GAT;
	I1348<= not N578GAT;
	I1353<= not N678GAT;
	I1360<= not N677GAT;
	I1371<= not N824GAT;
	I1374<= not N823GAT;
	I1385<= not N820GAT;
	I1388<= not N819GAT;
	I1399<= not N883GAT;
	I1402<= not N882GAT;
	I1407<= not N818GAT;
	I1411<= not N881GAT;
	I1416<= not N822GAT;
	I1422<= not N586GAT;
	I1436<= not N584GAT;
	I1439<= not N583GAT;
	I1450<= not N684GAT;
	I1453<= not N683GAT;
	I1464<= not N699GAT;
	I1467<= not N698GAT;
	I1472<= not N682GAT;
	I1476<= not N697GAT;
	I1481<= not N582GAT;
	I1488<= not N456GAT;
	I1493<= not N565GAT;
	I1496<= not N686GAT;
	I1500<= not N803GAT;
	I1538<= not N2399GAT;
	I1550<= not N2343GAT;
	I1606<= not N2490GAT;
	I1617<= not N2622GAT;
	I1630<= not N2630GAT;
	I1655<= not N2102GAT;
	I1667<= not N1880GAT;
	I1683<= not N1763GAT;
	I1698<= not N2155GAT;
	I1703<= not N2626GAT;
	I1708<= not N2543GAT;
	I1719<= not N2562GAT;
	I1749<= not N1035GAT;
	I1752<= not N1034GAT;
	I1766<= not N1121GAT;
	I1769<= not N1120GAT;
	I1783<= not N1072GAT;
	I1786<= not N1071GAT;
	I1791<= not N1119GAT;
	I1795<= not N1070GAT;
	I1800<= not N1033GAT;
	I1807<= not N1183GAT;
	I1833<= not N1226GAT;
	I1837<= not N1282GAT;
	I1843<= not N2970GAT;
	I1857<= not N931GAT;
	I1860<= not N930GAT;
	I1874<= not N1135GAT;
	I1877<= not N1134GAT;
	I1891<= not N1045GAT;
	I1894<= not N1044GAT;
	I1899<= not N1133GAT;
	I1903<= not N1043GAT;
	I1908<= not N929GAT;
	I1915<= not N1268GAT;
	I1920<= not N1329GAT;
	I1923<= not N1201GAT;
	I1927<= not N1184GAT;
	I1947<= not N1197GAT;
	I1961<= not N2516GAT;
	I1981<= not N667GAT;
	I1996<= not N659GAT;
	I1999<= not N658GAT;
	I2014<= not N553GAT;
	I2017<= not N552GAT;
	I2032<= not N777GAT;
	I2035<= not N776GAT;
	I2040<= not N551GAT;
	I2044<= not N775GAT;
	I2049<= not N657GAT;
	I2056<= not N35GAT;
	I2084<= not N366GAT;
	I2088<= not N561GAT;
	I2094<= not N2876GAT;
	I2109<= not N322GAT;
	I2112<= not N321GAT;
	I2127<= not N318GAT;
	I2130<= not N317GAT;
	I2145<= not N314GAT;
	I2148<= not N313GAT;
	I2153<= not N316GAT;
	I2157<= not N312GAT;
	I2162<= not N320GAT;
	I2169<= not N34GAT;
	I2174<= not N133GAT;
	I2177<= not N221GAT;
	I2181<= not N779GAT;
	I2213<= not N2342GAT;
	I2225<= not N2638GAT;
	I2228<= not N2561GAT;
	I2232<= not N2640GAT;
	I2235<= not N2639GAT;
	I2238<= not N2560GAT;
	I2242<= not N2341GAT;
	I2248<= not N2568GAT;
	I2251<= not N2207GAT;
	I2254<= not N2206GAT;
	I2257<= not N2398GAT;
	I2260<= not N2203GAT;
	I2263<= not N2202GAT;
	I2268<= not N2397GAT;
	I2271<= not N2201GAT;
	I2275<= not N2205GAT;
	I2281<= not N2409GAT;
	I2316<= not N2390GAT;
	I2319<= not N2495GAT;
	I2324<= not N3014GAT;
	I2344<= not N2339GAT;
	I2349<= not N2270GAT;
	I2354<= not N2880GAT;
	I2372<= not N2612GAT;
	I2376<= not N2532GAT;
	I2380<= not N2540GAT;
	I2385<= not N2536GAT;
	I2389<= not N2487GAT;
	I2394<= not N2557GAT;
	I2400<= not N2601GAT;
	I2403<= not N2629GAT;
	I2414<= not N2634GAT;
	I2417<= not N2633GAT;
	I2420<= not N2542GAT;
	I2425<= not N2632GAT;
	I2428<= not N2541GAT;
	I2433<= not N2628GAT;
	I2439<= not N2545GAT;
	I2672<= not N2143GAT;
	I2684<= not N2061GAT;
	I2696<= not N2139GAT;
	I2731<= not N1850GAT;
	I2771<= not N2440GAT;
	I2785<= not N2407GAT;
	I2837<= not N2347GAT;
	I2843<= not N2403GAT;
	I2847<= not N2394GAT;
	I2873<= not N1496GAT;
	I2885<= not N2091GAT;
	I2915<= not N1740GAT;
	I2953<= not N2179GAT;
	I2978<= not N2190GAT;
	I2989<= not N2135GAT;
	I3000<= not N2262GAT;
	I3016<= not N2182GAT;
	I3056<= not N1312GAT;
	I3143<= not N2592GAT;
	I3163<= not N1508GAT;
	I3168<= not N1394GAT;
	I3174<= not N1899GAT;
	I3191<= not N1678GAT;
	I3211<= not N2663GAT;
	I3235<= not N2238GAT;
	I3273<= not N2169GAT;
	I3287<= not N1691GAT;
	I3290<= not N1691GAT;
	I3293<= not N1691GAT;
	I3297<= not N1699GAT;
	I3300<= not N1699GAT;
	I3303<= not N1691GAT;
	I3306<= not N1699GAT;
	I3309<= not N1699GAT;
	I3312<= not N1699GAT;
	I3315<= not N1869GAT;
	I3318<= not N1869GAT;
	I3336<= not N2040GAT;
	I3339<= not N1775GAT;
	I3342<= not N1316GAT;
	I3387<= not N2194GAT;
	I3390<= not N2261GAT;
	I3394<= not N2260GAT;
	I3401<= not N2192GAT;
	I3412<= not N2057GAT;
	I3429<= not N2266GAT;
	I3436<= not N2492GAT;
	I3457<= not N2556GAT;
	I3461<= not N1956GAT;
	I3465<= not N1886GAT;
	I3472<= not N2539GAT;
	I3483<= not N2436GAT;
	I3491<= not N2387GAT;
	I3494<= not N1963GAT;
	I3504<= not N2330GAT;
	I3509<= not N2438GAT;
	I3513<= not N2439GAT;
	I3520<= not N2498GAT;
	I3530<= not N2396GAT;
	I3539<= not N2198GAT;
	I3549<= not N2197GAT;
	I3558<= not N2196GAT;
	I3587<= not N2125GAT;
	I3610<= not N1882GAT;
	I3621<= not N1975GAT;
	I3635<= not N2558GAT;
	I3646<= not N2644GAT;
	I3660<= not N2636GAT;
	I3677<= not N156GAT;
	I3691<= not N152GAT;
	I3703<= not N2917GAT;
	I3713<= not N2892GAT;
	I3736<= not N388GAT;
	I3742<= not N331GAT;
	I3754<= not N2900GAT;
	I3765<= not N2929GAT;
	I3777<= not N463GAT;
	I3801<= not N2925GAT;
	I3808<= not N327GAT;
	I3817<= not N2916GAT;
	I3831<= not N384GAT;
	I3841<= not N2899GAT;
	I3867<= not N470GAT;
	I3876<= not N2926GAT;
	I3882<= not N256GAT;
	I3891<= not N2924GAT;
	I3904<= not N148GAT;
	I3914<= not N2923GAT;
	I3923<= not N2710GAT;
	I3935<= not N2704GAT;
	I3941<= not N2684GAT;
	I3945<= not N1350GAT;
	I3948<= not N2696GAT;
	I3951<= not N2448GAT;
	I3954<= not N2683GAT;
	I3957<= not N2450GAT;
	I3962<= not N2830GAT;
	I4014<= not N2744GAT;
	I4020<= not N2800GAT;
	I4055<= not N1748GAT;
	I4067<= not N1675GAT;
	I4081<= not N1807GAT;
	I4105<= not N1456GAT;
	I4108<= not N1340GAT;
	I4117<= not N1505GAT;
	I4122<= not N1546GAT;
	I4129<= not N3097GAT;
	I4135<= not N3098GAT;
	I4138<= not N2766GAT;
	I4157<= not N1525GAT;
	I4185<= not N1596GAT;
	I4194<= not N1462GAT;
	I4212<= not N1588GAT;
	I4222<= not N1761GAT;
	I4227<= not N1760GAT;
	I4233<= not N1721GAT;
	I4236<= not N2808GAT;
	I4309<= not N2941GAT;
	I4312<= not N2814GAT;
	I4329<= not N2950GAT;
	I4332<= not N2813GAT;
	I4349<= not N2935GAT;
	I4352<= not N2818GAT;
	I4369<= not N2937GAT;
	I4372<= not N2817GAT;
	I4389<= not N2956GAT;
	I4392<= not N2824GAT;
	I4409<= not N2938GAT;
	I4412<= not N2823GAT;
	I4429<= not N2936GAT;
	I4432<= not N2829GAT;
	I4449<= not N2955GAT;
	I4452<= not N2828GAT;
	I4475<= not N2951GAT;
	I4478<= not N2807GAT;
	I4482<= not N2127GAT;
	I4485<= not N2682GAT;
	I4489<= not N2046GAT;
	I4492<= not N2681GAT;
	I4496<= not N1708GAT;
	I4499<= not N2688GAT;
	I4506<= not N2764GAT;
	I4512<= not N2762GAT;
	I4518<= not N2761GAT;
	I4524<= not N2757GAT;
	I4530<= not N2756GAT;
	I4536<= not N2750GAT;
	I4542<= not N2749GAT;
	I4548<= not N2742GAT;
	I4554<= not N2741GAT;
	I4558<= not N1286GAT;
	I4566<= not N2694GAT;
	I4573<= not N2693GAT;
	I4580<= not N2702GAT;
	I4587<= not N2701GAT;
	I4594<= not N2709GAT;
	I4601<= not N2708GAT;
	I4608<= not N2799GAT;
	I4615<= not N2798GAT;
	I4620<= not N1745GAT;
	I4623<= not N2806GAT;
	I4626<= not N1871GAT;
	I4630<= not N1086GAT;
	I4633<= not N2805GAT;
	I4642<= not N2812GAT;
	I4651<= not N2822GAT;
	I4654<= not N2819GAT;
	I4657<= not N2809GAT;
	I4660<= not N2801GAT;
	I4663<= not N2802GAT;
	I4666<= not N2795GAT;
	I4669<= not N2796GAT;
	I4672<= not N2705GAT;
	I4675<= not N2706GAT;
	I4678<= not N2697GAT;
	I4681<= not N2698GAT;
	I4684<= not N2689GAT;
	I4687<= not N2690GAT;
	I4690<= not N2685GAT;
	I4693<= not N2737GAT;
	I4696<= not N2738GAT;
	I4699<= not N2745GAT;
	I4702<= not N2746GAT;
	I4705<= not N2753GAT;
	I4708<= not N2754GAT;
	I4711<= not N2759GAT;
	I4714<= not N2760GAT;
	I4717<= not N2763GAT;
	I4720<= not N2686GAT;
	I4723<= not N2677GAT;
	I4726<= not N2678GAT;
	I4729<= not N2803GAT;
	I4732<= not N2825GAT;
	I4735<= not N2826GAT;
	I4738<= not N2820GAT;
	I4741<= not N2821GAT;
	I4744<= not N2815GAT;
	I4747<= not N2816GAT;
	I4750<= not N2810GAT;
	I4753<= not N2811GAT;
	I4756<= not N2804GAT;
	I4759<= not N2739GAT;
	I4762<= not N2747GAT;
	I4765<= not N2748GAT;
	I4768<= not N2755GAT;
	I4771<= not N2797GAT;
	I4774<= not N2740GAT;
	I4777<= not N2699GAT;
	I4780<= not N2691GAT;
	I4783<= not N2827GAT;
	I4786<= not N2679GAT;
	I4789<= not N2692GAT;
	I4792<= not N2680GAT;
	I4795<= not N2700GAT;
	I4798<= not N2707GAT;
	N11GAT<= not N12GAT;
	N14GAT<= not N186GAT;
	N16GAT<= not N564GAT;
	N17GAT<= not N564GAT;
	N21GAT<= not N15GAT;
	N34GAT<= not N221GAT;
	N35GAT<= not N779GAT;
	N41GAT<= not N258GAT;
	N42GAT<= not N475GAT;
	N48GAT<= not I375;
	N49GAT<= not I420;
	N50GAT<= not I468;
	N51GAT<= not I473;
	N52GAT<= not I476;
	N53GAT<= not I480;
	N54GAT<= not N167GAT;
	N60GAT<= not I658;
	N61GAT<= not I698;
	N62GAT<= not I741;
	N63GAT<= not I746;
	N64GAT<= not I749;
	N65GAT<= not I753;
	N66GAT<= not N906GAT;
	N67GAT<= not N85GAT;
	N69GAT<= not N68GAT;
	N71GAT<= not N180GAT;
	N72GAT<= not N181GAT;
	N76GAT<= not N82GAT;
	N79GAT<= not N86GAT;
	N88GAT<= not N84GAT;
	N92GAT<= not N2785GAT;
	N111GAT<= not N182GAT;
	N125GAT<= not I2056;
	N126GAT<= not I2094;
	N127GAT<= not I2169;
	N128GAT<= not I2174;
	N129GAT<= not I2177;
	N130GAT<= not I2181;
	N133GAT<= not N2876GAT;
	N134GAT<= not N2875GAT;
	N144GAT<= not N247GAT;
	N146GAT<= not N148GAT;
	N147GAT<= not I3904;
	N150GAT<= not N152GAT;
	N151GAT<= not I3691;
	N154GAT<= not N156GAT;
	N155GAT<= not I3677;
	N158GAT<= not N160GAT;
	N159GAT<= not I331;
	N162GAT<= not N1013GAT;
	N163GAT<= not N165GAT;
	N164GAT<= not I620;
	N172GAT<= not I609;
	N173GAT<= not I623;
	N174GAT<= not I637;
	N175GAT<= not I642;
	N176GAT<= not I646;
	N177GAT<= not I651;
	N178GAT<= not N343GAT;
	N179GAT<= not N287GAT;
	N188GAT<= not N288GAT;
	N189GAT<= not N286GAT;
	N194GAT<= not N187GAT;
	N195GAT<= not N184GAT;
	N199GAT<= not N87GAT;
	N219GAT<= not N78GAT;
	N226GAT<= not I2112;
	N227GAT<= not I2130;
	N228GAT<= not I2148;
	N229GAT<= not I2153;
	N230GAT<= not I2157;
	N231GAT<= not I2162;
	N233GAT<= not N243GAT;
	N235GAT<= not N2878GAT;
	N241GAT<= not N140GAT;
	N243GAT<= not N1702GAT;
	N252GAT<= not N2877GAT;
	N253GAT<= not N1702GAT;
	N254GAT<= not N256GAT;
	N255GAT<= not I3882;
	N263GAT<= not I314;
	N264GAT<= not I334;
	N265GAT<= not I354;
	N266GAT<= not I359;
	N267GAT<= not I363;
	N268GAT<= not I368;
	N269GAT<= not N271GAT;
	N270GAT<= not I311;
	N273GAT<= not N275GAT;
	N274GAT<= not I709;
	N277GAT<= not N279GAT;
	N278GAT<= not I634;
	N281GAT<= not N283GAT;
	N282GAT<= not I606;
	N289GAT<= not N563GAT;
	N290GAT<= not N525GAT;
	N293GAT<= not N361GAT;
	N294GAT<= not N360GAT;
	N295GAT<= not N357GAT;
	N296GAT<= not N421GAT;
	N297GAT<= not N2721GAT;
	N312GAT<= not N314GAT;
	N313GAT<= not I2145;
	N316GAT<= not N318GAT;
	N317GAT<= not I2127;
	N320GAT<= not N322GAT;
	N321GAT<= not I2109;
	N325GAT<= not N327GAT;
	N326GAT<= not I3808;
	N329GAT<= not N331GAT;
	N330GAT<= not I3742;
	N333GAT<= not N2883GAT;
	N334GAT<= not N1700GAT;
	N335GAT<= not N337GAT;
	N336GAT<= not I351;
	N339GAT<= not N341GAT;
	N340GAT<= not I437;
	N348GAT<= not I712;
	N349GAT<= not I715;
	N350GAT<= not I721;
	N351GAT<= not I726;
	N352GAT<= not I729;
	N353GAT<= not I734;
	N358GAT<= not N532GAT;
	N364GAT<= not N366GAT;
	N365GAT<= not I2084;
	N368GAT<= not N1725GAT;
	N369GAT<= not N1725GAT;
	N370GAT<= not N1725GAT;
	N371GAT<= not N1725GAT;
	N372GAT<= not N212GAT;
	N373GAT<= not N2767GAT;
	N374GAT<= not N2767GAT;
	N375GAT<= not N110GAT;
	N380GAT<= not N2881GAT;
	N381GAT<= not N2893GAT;
	N382GAT<= not N384GAT;
	N383GAT<= not I3831;
	N386GAT<= not N388GAT;
	N387GAT<= not I3736;
	N392GAT<= not N394GAT;
	N393GAT<= not I446;
	N396GAT<= not N398GAT;
	N397GAT<= not I718;
	N400GAT<= not N402GAT;
	N401GAT<= not I76;
	N404GAT<= not N493GAT;
	N405GAT<= not N728GAT;
	N406GAT<= not N516GAT;
	N407GAT<= not N355GAT;
	N412GAT<= not N522GAT;
	N413GAT<= not N411GAT;
	N416GAT<= not N415GAT;
	N417GAT<= not N418GAT;
	N422GAT<= not N2889GAT;
	N452GAT<= not N2885GAT;
	N455GAT<= not N291GAT;
	N456GAT<= not N686GAT;
	N457GAT<= not N2884GAT;
	N458GAT<= not N2902GAT;
	N461GAT<= not N463GAT;
	N462GAT<= not I3777;
	N468GAT<= not N470GAT;
	N469GAT<= not I3867;
	N480GAT<= not I440;
	N481GAT<= not I443;
	N482GAT<= not I449;
	N483GAT<= not I453;
	N484GAT<= not I456;
	N485GAT<= not I461;
	N489GAT<= not N491GAT;
	N490GAT<= not I1088;
	N498GAT<= not I1230;
	N499GAT<= not I1085;
	N500GAT<= not I1091;
	N501GAT<= not I1067;
	N502GAT<= not I1079;
	N503GAT<= not I1236;
	N509GAT<= not I1190;
	N510GAT<= not I1216;
	N511GAT<= not I1243;
	N512GAT<= not I1248;
	N513GAT<= not I1251;
	N514GAT<= not I1255;
	N515GAT<= not N709GAT;
	N517GAT<= not N518GAT;
	N524GAT<= not N414GAT;
	N527GAT<= not N356GAT;
	N528GAT<= not N521GAT;
	N551GAT<= not N553GAT;
	N552GAT<= not I2014;
	N558GAT<= not N1725GAT;
	N559GAT<= not N561GAT;
	N560GAT<= not I2088;
	N563GAT<= not I1278;
	N565GAT<= not N586GAT;
	N566GAT<= not N364GAT;
	N572GAT<= not I1360;
	N573GAT<= not I1422;
	N574GAT<= not I1488;
	N575GAT<= not I1493;
	N576GAT<= not I1496;
	N577GAT<= not I1500;
	N578GAT<= not N580GAT;
	N579GAT<= not I1336;
	N582GAT<= not N584GAT;
	N583GAT<= not I1436;
	N591GAT<= not I1374;
	N592GAT<= not I1388;
	N593GAT<= not I1402;
	N594GAT<= not I1407;
	N595GAT<= not I1411;
	N596GAT<= not I1416;
	N612GAT<= not N614GAT;
	N613GAT<= not I1227;
	N616GAT<= not N618GAT;
	N617GAT<= not I1082;
	N620GAT<= not N622GAT;
	N621GAT<= not I1118;
	N624GAT<= not N626GAT;
	N625GAT<= not I1124;
	N628GAT<= not N631GAT;
	N633GAT<= not N634GAT;
	N637GAT<= not N529GAT;
	N639GAT<= not N523GAT;
	N640GAT<= not N1213GAT;
	N641GAT<= not N855GAT;
	N642GAT<= not N855GAT;
	N643GAT<= not N855GAT;
	N644GAT<= not N855GAT;
	N657GAT<= not N659GAT;
	N658GAT<= not I1996;
	N661GAT<= not N1725GAT;
	N662GAT<= not N1725GAT;
	N663GAT<= not N1725GAT;
	N664GAT<= not N1725GAT;
	N665GAT<= not N667GAT;
	N666GAT<= not I1981;
	N670GAT<= not N636GAT;
	N671GAT<= not N673GAT;
	N672GAT<= not I44;
	N677GAT<= not N803GAT;
	N678GAT<= not N680GAT;
	N679GAT<= not I1302;
	N682GAT<= not N684GAT;
	N683GAT<= not I1450;
	N691GAT<= not I1439;
	N692GAT<= not I1453;
	N693GAT<= not I1467;
	N694GAT<= not I1472;
	N695GAT<= not I1476;
	N696GAT<= not I1481;
	N697GAT<= not N699GAT;
	N698GAT<= not I1464;
	N701GAT<= not N703GAT;
	N702GAT<= not I149;
	N705GAT<= not N707GAT;
	N706GAT<= not I1152;
	N714GAT<= not I1141;
	N715GAT<= not I1155;
	N716GAT<= not I1169;
	N717GAT<= not I1174;
	N718GAT<= not I1178;
	N719GAT<= not I1183;
	N720GAT<= not N722GAT;
	N721GAT<= not I178;
	N724GAT<= not N726GAT;
	N725GAT<= not I171;
	N733GAT<= not I1121;
	N734GAT<= not I1204;
	N735GAT<= not I1127;
	N736GAT<= not I1209;
	N737GAT<= not I1115;
	N738GAT<= not I1103;
	N739GAT<= not N850GAT;
	N740GAT<= not N2667GAT;
	N741GAT<= not N629GAT;
	N743GAT<= not N746GAT;
	N747GAT<= not N2906GAT;
	N753GAT<= not I237;
	N754GAT<= not I253;
	N755GAT<= not I270;
	N756GAT<= not I275;
	N757GAT<= not I278;
	N758GAT<= not I282;
	N759GAT<= not N855GAT;
	N760GAT<= not N855GAT;
	N761GAT<= not N855GAT;
	N762GAT<= not N855GAT;
	N775GAT<= not N777GAT;
	N776GAT<= not I2032;
	N784GAT<= not I1999;
	N785GAT<= not I2017;
	N786GAT<= not I2035;
	N787GAT<= not I2040;
	N788GAT<= not I2044;
	N789GAT<= not I2049;
	N800GAT<= not N2874GAT;
	N802GAT<= not N2882GAT;
	N808GAT<= not I1305;
	N809GAT<= not I1322;
	N810GAT<= not I1339;
	N811GAT<= not I1344;
	N812GAT<= not I1348;
	N813GAT<= not I1353;
	N814GAT<= not N816GAT;
	N815GAT<= not I1319;
	N818GAT<= not N820GAT;
	N819GAT<= not I1385;
	N822GAT<= not N824GAT;
	N823GAT<= not I1371;
	N827GAT<= not N204GAT;
	N828GAT<= not N830GAT;
	N829GAT<= not I1201;
	N832GAT<= not N834GAT;
	N833GAT<= not I1138;
	N836GAT<= not N838GAT;
	N837GAT<= not I1166;
	N840GAT<= not N842GAT;
	N841GAT<= not I395;
	N844GAT<= not N846GAT;
	N845GAT<= not I111;
	N848GAT<= not N922GAT;
	N849GAT<= not N924GAT;
	N850GAT<= not N929GAT;
	N851GAT<= not N853GAT;
	N852GAT<= not N854GAT;
	N855GAT<= not N2148GAT;
	N856GAT<= not N2667GAT;
	N857GAT<= not N944GAT;
	N858GAT<= not N1228GAT;
	N859GAT<= not N861GAT;
	N860GAT<= not I834;
	N863GAT<= not N865GAT;
	N864GAT<= not I955;
	N873GAT<= not N316GAT;
	N875GAT<= not N559GAT;
	N876GAT<= not N1347GAT;
	N878GAT<= not N2879GAT;
	N881GAT<= not N883GAT;
	N882GAT<= not I1399;
	N888GAT<= not N2933GAT;
	N894GAT<= not N2932GAT;
	N897GAT<= not N2939GAT;
	N898GAT<= not N2940GAT;
	N911GAT<= not I661;
	N912GAT<= not I675;
	N913GAT<= not I678;
	N914GAT<= not I683;
	N915GAT<= not I687;
	N916GAT<= not I692;
	N917GAT<= not N919GAT;
	N918GAT<= not I92;
	N921GAT<= not N923GAT;
	N922GAT<= not N1119GAT;
	N923GAT<= not N1043GAT;
	N924GAT<= not N1070GAT;
	N925GAT<= not N927GAT;
	N926GAT<= not N632GAT;
	N927GAT<= not N1133GAT;
	N928GAT<= not N1050GAT;
	N929GAT<= not N931GAT;
	N930GAT<= not I1857;
	N938GAT<= not I858;
	N939GAT<= not I936;
	N940GAT<= not I1023;
	N941GAT<= not I1028;
	N942GAT<= not I1031;
	N943GAT<= not I1035;
	N949GAT<= not I793;
	N950GAT<= not I815;
	N951GAT<= not I837;
	N952GAT<= not I842;
	N953GAT<= not I846;
	N954GAT<= not I851;
	N955GAT<= not N957GAT;
	N956GAT<= not I812;
	N976GAT<= not N628GAT;
	N983GAT<= not N320GAT;
	N985GAT<= not N775GAT;
	N1002GAT<= not N2946GAT;
	N1006GAT<= not N630GAT;
	N1007GAT<= not N635GAT;
	N1018GAT<= not I378;
	N1019GAT<= not I398;
	N1020GAT<= not I401;
	N1021GAT<= not I406;
	N1022GAT<= not I409;
	N1023GAT<= not I414;
	N1024GAT<= not N1026GAT;
	N1025GAT<= not I672;
	N1032GAT<= not N1118GAT;
	N1033GAT<= not N1035GAT;
	N1034GAT<= not I1749;
	N1043GAT<= not N1045GAT;
	N1044GAT<= not I1891;
	N1055GAT<= not I958;
	N1056GAT<= not I980;
	N1057GAT<= not I1002;
	N1058GAT<= not I1007;
	N1059GAT<= not I1011;
	N1060GAT<= not I1016;
	N1066GAT<= not N1068GAT;
	N1067GAT<= not I790;
	N1070GAT<= not N1072GAT;
	N1071GAT<= not I1783;
	N1075GAT<= not N855GAT;
	N1078GAT<= not N1080GAT;
	N1079GAT<= not I977;
	N1084GAT<= not N657GAT;
	N1085GAT<= not N551GAT;
	N1086GAT<= not N1870GAT;
	N1105GAT<= not N2934GAT;
	N1106GAT<= not N2949GAT;
	N1111GAT<= not N635GAT;
	N1112GAT<= not N630GAT;
	N1118GAT<= not N1033GAT;
	N1119GAT<= not N1121GAT;
	N1120GAT<= not I1766;
	N1123GAT<= not N632GAT;
	N1133GAT<= not N1135GAT;
	N1134GAT<= not I1874;
	N1146GAT<= not N1148GAT;
	N1147GAT<= not I999;
	N1150GAT<= not N312GAT;
	N1157GAT<= not N1483GAT;
	N1160GAT<= not N1484GAT;
	N1164GAT<= not N2953GAT;
	N1179GAT<= not N2947GAT;
	N1180GAT<= not N2948GAT;
	N1183GAT<= not N1184GAT;
	N1189GAT<= not I1752;
	N1190GAT<= not I1769;
	N1191GAT<= not I1786;
	N1192GAT<= not I1791;
	N1193GAT<= not I1795;
	N1194GAT<= not I1800;
	N1195GAT<= not N1197GAT;
	N1196GAT<= not I1947;
	N1206GAT<= not I1860;
	N1207GAT<= not I1877;
	N1208GAT<= not I1894;
	N1209GAT<= not I1899;
	N1210GAT<= not I1903;
	N1211GAT<= not I1908;
	N1218GAT<= not I196;
	N1219GAT<= not I203;
	N1220GAT<= not I210;
	N1221GAT<= not I217;
	N1222GAT<= not I223;
	N1223GAT<= not I230;
	N1224GAT<= not N1226GAT;
	N1225GAT<= not I1833;
	N1233GAT<= not I880;
	N1234GAT<= not I902;
	N1235GAT<= not I916;
	N1236GAT<= not I921;
	N1237GAT<= not I925;
	N1238GAT<= not I930;
	N1239GAT<= not N1241GAT;
	N1240GAT<= not I899;
	N1247GAT<= not N2958GAT;
	N1248GAT<= not N2954GAT;
	N1268GAT<= not N1201GAT;
	N1274GAT<= not I1807;
	N1275GAT<= not I1843;
	N1276GAT<= not I1915;
	N1277GAT<= not I1920;
	N1278GAT<= not I1923;
	N1279GAT<= not I1927;
	N1280GAT<= not N1282GAT;
	N1281GAT<= not I1837;
	N1284GAT<= not N1269GAT;
	N1286GAT<= not N1269GAT;
	N1292GAT<= not N1294GAT;
	N1293GAT<= not I877;
	N1296GAT<= not N1298GAT;
	N1297GAT<= not I913;
	N1300GAT<= not N2963GAT;
	N1301GAT<= not N1416GAT;
	N1306GAT<= not N2964GAT;
	N1307GAT<= not N1308GAT;
	N1309GAT<= not N2959GAT;
	N1310GAT<= not N1312GAT;
	N1311GAT<= not I3056;
	N1314GAT<= not N1316GAT;
	N1315GAT<= not I3342;
	N1319GAT<= not N1256GAT;
	N1322GAT<= not N2974GAT;
	N1328GAT<= not N1224GAT;
	N1329GAT<= not N2970GAT;
	N1330GAT<= not N1332GAT;
	N1334GAT<= not N1336GAT;
	N1338GAT<= not N1340GAT;
	N1339GAT<= not I4108;
	N1348GAT<= not N1349GAT;
	N1350GAT<= not N1831GAT;
	N1353GAT<= not N1419GAT;
	N1355GAT<= not N1422GAT;
	N1356GAT<= not N1354GAT;
	N1361GAT<= not N1363GAT;
	N1366GAT<= not N1365GAT;
	N1369GAT<= not N2966GAT;
	N1370GAT<= not N1426GAT;
	N1374GAT<= not N2979GAT;
	N1378GAT<= not N2975GAT;
	N1379GAT<= not N1377GAT;
	N1380GAT<= not N1114GAT;
	N1381GAT<= not N1328GAT;
	N1382GAT<= not N1280GAT;
	N1384GAT<= not N2184GAT;
	N1387GAT<= not N1389GAT;
	N1392GAT<= not N1394GAT;
	N1393GAT<= not I3168;
	N1396GAT<= not N1401GAT;
	N1403GAT<= not N1402GAT;
	N1409GAT<= not N1476GAT;
	N1410GAT<= not N2357GAT;
	N1414GAT<= not N1415GAT;
	N1418GAT<= not N1417GAT;
	N1424GAT<= not N1420GAT;
	N1425GAT<= not N1421GAT;
	N1427GAT<= not N1608GAT;
	N1430GAT<= not N1700GAT;
	N1431GAT<= not N1433GAT;
	N1436GAT<= not N1435GAT;
	N1437GAT<= not N1438GAT;
	N1439GAT<= not N1486GAT;
	N1442GAT<= not N1831GAT;
	N1444GAT<= not N1442GAT;
	N1446GAT<= not N1318GAT;
	N1447GAT<= not N1117GAT;
	N1448GAT<= not N1376GAT;
	N1449GAT<= not N1494GAT;
	N1450GAT<= not N1423GAT;
	N1451GAT<= not N1382GAT;
	N1452GAT<= not N2049GAT;
	N1453GAT<= not N2187GAT;
	N1454GAT<= not N1469GAT;
	N1455GAT<= not I4105;
	N1460GAT<= not N1462GAT;
	N1461GAT<= not I4194;
	N1468GAT<= not N1519GAT;
	N1477GAT<= not N2984GAT;
	N1478GAT<= not N1481GAT;
	N1479GAT<= not N2291GAT;
	N1480GAT<= not N2292GAT;
	N1482GAT<= not N2363GAT;
	N1487GAT<= not N1485GAT;
	N1490GAT<= not N1430GAT;
	N1495GAT<= not I2873;
	N1500GAT<= not N1113GAT;
	N1503GAT<= not N1501GAT;
	N1505GAT<= not N2980GAT;
	N1507GAT<= not I3163;
	N1513GAT<= not N2288GAT;
	N1515GAT<= not N1521GAT;
	N1517GAT<= not N1578GAT;
	N1518GAT<= not N1694GAT;
	N1520GAT<= not N1582GAT;
	N1523GAT<= not N2219GAT;
	N1524GAT<= not I4157;
	N1528GAT<= not N2293GAT;
	N1530GAT<= not N2364GAT;
	N1543GAT<= not N1606GAT;
	N1544GAT<= not N1625GAT;
	N1546GAT<= not N2980GAT;
	N1548GAT<= not I2721;
	N1549GAT<= not I2832;
	N1550GAT<= not I2890;
	N1551GAT<= not N1549GAT;
	N1552GAT<= not N1550GAT;
	N1553GAT<= not N1616GAT;
	N1554GAT<= not N1555GAT;
	N1559GAT<= not N1614GAT;
	N1560GAT<= not N1557GAT;
	N1561GAT<= not N1571GAT;
	N1562GAT<= not N1556GAT;
	N1566GAT<= not N1605GAT;
	N1568GAT<= not N1575GAT;
	N1569GAT<= not N1570GAT;
	N1572GAT<= not N1576GAT;
	N1580GAT<= not N1577GAT;
	N1584GAT<= not N2989GAT;
	N1587GAT<= not I4212;
	N1590GAT<= not N1603GAT;
	N1591GAT<= not N2223GAT;
	N1592GAT<= not N1529GAT;
	N1594GAT<= not N1596GAT;
	N1595GAT<= not I4185;
	N1601GAT<= not N120GAT;
	N1603GAT<= not N1831GAT;
	N1615GAT<= not N1624GAT;
	N1627GAT<= not N1618GAT;
	N1628GAT<= not N1621GAT;
	N1629GAT<= not N1895GAT;
	N1631GAT<= not N1848GAT;
	N1632GAT<= not I4145;
	N1633GAT<= not N2137GAT;
	N1634GAT<= not N1712GAT;
	N1635GAT<= not N1716GAT;
	N1640GAT<= not N1639GAT;
	N1643GAT<= not N1641GAT;
	N1645GAT<= not N1499GAT;
	N1648GAT<= not N1729GAT;
	N1651GAT<= not N1642GAT;
	N1652GAT<= not N1657GAT;
	N1656GAT<= not N1655GAT;
	N1658GAT<= not N2216GAT;
	N1659GAT<= not N2987GAT;
	N1661GAT<= not N1660GAT;
	N1662GAT<= not N1663GAT;
	N1665GAT<= not N1666GAT;
	N1668GAT<= not N1734GAT;
	N1670GAT<= not N1667GAT;
	N1671GAT<= not N1669GAT;
	N1673GAT<= not N2989GAT;
	N1674GAT<= not I4067;
	N1677GAT<= not I3191;
	N1681GAT<= not I4217;
	N1683GAT<= not N1756GAT;
	N1684GAT<= not N1759GAT;
	N1685GAT<= not N1604GAT;
	N1691GAT<= not N2452GAT;
	N1693GAT<= not N2101GAT;
	N1694GAT<= not I2813;
	N1698GAT<= not N1934GAT;
	N1699GAT<= not N2452GAT;
	N1701GAT<= not N1617GAT;
	N1705GAT<= not N1619GAT;
	N1706GAT<= not N1622GAT;
	N1707GAT<= not N1626GAT;
	N1708GAT<= not N2338GAT;
	N1709GAT<= not N1849GAT;
	N1711GAT<= not N2990GAT;
	N1712GAT<= not I3179;
	N1713GAT<= not I2935;
	N1714GAT<= not I3149;
	N1716GAT<= not I2736;
	N1717GAT<= not I2926;
	N1718GAT<= not N1714GAT;
	N1719GAT<= not N1548GAT;
	N1722GAT<= not N1558GAT;
	N1724GAT<= not N1732GAT;
	N1725GAT<= not N2148GAT;
	N1727GAT<= not N1728GAT;
	N1730GAT<= not N1731GAT;
	N1735GAT<= not N1861GAT;
	N1736GAT<= not N1737GAT;
	N1738GAT<= not N1740GAT;
	N1739GAT<= not I2915;
	N1742GAT<= not N2216GAT;
	N1743GAT<= not N1713GAT;
	N1747GAT<= not I4055;
	N1754GAT<= not N2449GAT;
	N1762GAT<= not I1683;
	N1765GAT<= not N1767GAT;
	N1769GAT<= not N1771GAT;
	N1773GAT<= not N1775GAT;
	N1774GAT<= not I3339;
	N1777GAT<= not N1694GAT;
	N1779GAT<= not N1623GAT;
	N1781GAT<= not N1780GAT;
	N1782GAT<= not N2971GAT;
	N1783GAT<= not N1848GAT;
	N1784GAT<= not N1849GAT;
	N1785GAT<= not N2059GAT;
	N1786GAT<= not N2060GAT;
	N1787GAT<= not N2141GAT;
	N1788GAT<= not N2142GAT;
	N1790GAT<= not N1726GAT;
	N1791GAT<= not N2013GAT;
	N1797GAT<= not N1801GAT;
	N1806GAT<= not I4081;
	N1816GAT<= not N1817GAT;
	N1819GAT<= not N1821GAT;
	N1823GAT<= not N1825GAT;
	N1828GAT<= not I572;
	N1832GAT<= not N1834GAT;
	N1836GAT<= not N1695GAT;
	N1838GAT<= not N1898GAT;
	N1839GAT<= not N2138GAT;
	N1840GAT<= not N1892GAT;
	N1841GAT<= not N2058GAT;
	N1842GAT<= not N1711GAT;
	N1845GAT<= not N2141GAT;
	N1848GAT<= not N1850GAT;
	N1849GAT<= not I2731;
	N1855GAT<= not N2014GAT;
	N1858GAT<= not N1673GAT;
	N1859GAT<= not N1717GAT;
	N1862GAT<= not N1863GAT;
	N1866GAT<= not N1865GAT;
	N1869GAT<= not N1871GAT;
	N1870GAT<= not I4626;
	N1878GAT<= not N1880GAT;
	N1879GAT<= not I1667;
	N1884GAT<= not N1897GAT;
	N1885GAT<= not N2048GAT;
	N1886GAT<= not N1897GAT;
	N1887GAT<= not N2138GAT;
	N1888GAT<= not N3039GAT;
	N1889GAT<= not N1961GAT;
	N1890GAT<= not N2328GAT;
	N1891GAT<= not N2059GAT;
	N1892GAT<= not N2993GAT;
	N1893GAT<= not N2060GAT;
	N1897GAT<= not N1899GAT;
	N1898GAT<= not I3174;
	N1917GAT<= not N1921GAT;
	N1918GAT<= not N2392GAT;
	N1919GAT<= not N1860GAT;
	N1922GAT<= not N1798GAT;
	N1923GAT<= not N1864GAT;
	N1925GAT<= not N1920GAT;
	N1945GAT<= not N1690GAT;
	N1954GAT<= not N3038GAT;
	N1955GAT<= not N1956GAT;
	N1956GAT<= not N1898GAT;
	N1960GAT<= not N3043GAT;
	N1961GAT<= not N2996GAT;
	N1963GAT<= not N2137GAT;
	N1968GAT<= not N1958GAT;
	N1969GAT<= not N2142GAT;
	N1970GAT<= not N1896GAT;
	N1973GAT<= not N1975GAT;
	N1974GAT<= not I3621;
	N1978GAT<= not N2286GAT;
	N1986GAT<= not N2439GAT;
	N1988GAT<= not N2345GAT;
	N1989GAT<= not N2401GAT;
	N1990GAT<= not N2988GAT;
	N1991GAT<= not N2393GAT;
	N1999GAT<= not N2001GAT;
	N2000GAT<= not N1412GAT;
	N2001GAT<= not N1412GAT;
	N2002GAT<= not N2008GAT;
	N2004GAT<= not N1929GAT;
	N2011GAT<= not N2306GAT;
	N2012GAT<= not N2016GAT;
	N2013GAT<= not I4000;
	N2019GAT<= not N2021GAT;
	N2023GAT<= not N2025GAT;
	N2027GAT<= not N2029GAT;
	N2031GAT<= not N2033GAT;
	N2035GAT<= not N2037GAT;
	N2039GAT<= not I3336;
	N2042GAT<= not N2044GAT;
	N2046GAT<= not N2269GAT;
	N2047GAT<= not N2209GAT;
	N2048GAT<= not N2994GAT;
	N2049GAT<= not N3001GAT;
	N2050GAT<= not N2146GAT;
	N2051GAT<= not N2056GAT;
	N2052GAT<= not N2393GAT;
	N2054GAT<= not N2281GAT;
	N2056GAT<= not N2998GAT;
	N2058GAT<= not N2997GAT;
	N2059GAT<= not N2061GAT;
	N2060GAT<= not I2684;
	N2081GAT<= not N2218GAT;
	N2082GAT<= not N2084GAT;
	N2090GAT<= not I2885;
	N2093GAT<= not N2095GAT;
	N2097GAT<= not N2099GAT;
	N2101GAT<= not I1655;
	N2108GAT<= not N2110GAT;
	N2115GAT<= not N2117GAT;
	N2119GAT<= not N2121GAT;
	N2123GAT<= not N2125GAT;
	N2124GAT<= not I3587;
	N2127GAT<= not N2389GAT;
	N2128GAT<= not N2129GAT;
	N2131GAT<= not N2185GAT;
	N2133GAT<= not N2135GAT;
	N2134GAT<= not I2989;
	N2137GAT<= not N2139GAT;
	N2138GAT<= not I2696;
	N2141GAT<= not N2143GAT;
	N2142GAT<= not I2672;
	N2146GAT<= not N3002GAT;
	N2148GAT<= not I1734;
	N2151GAT<= not N2193GAT;
	N2152GAT<= not N2346GAT;
	N2153GAT<= not N2155GAT;
	N2154GAT<= not I1698;
	N2158GAT<= not N1412GAT;
	N2159GAT<= not N1412GAT;
	N2162GAT<= not N2220GAT;
	N2167GAT<= not N2169GAT;
	N2168GAT<= not I3273;
	N2174GAT<= not N2176GAT;
	N2178GAT<= not I2953;
	N2181GAT<= not I3016;
	N2184GAT<= not N3003GAT;
	N2186GAT<= not N2613GAT;
	N2187GAT<= not N3004GAT;
	N2188GAT<= not N2190GAT;
	N2189GAT<= not I2978;
	N2199GAT<= not N2147GAT;
	N2200GAT<= not N2078GAT;
	N2201GAT<= not N2203GAT;
	N2202GAT<= not I2260;
	N2205GAT<= not N2207GAT;
	N2206GAT<= not I2251;
	N2209GAT<= not N3005GAT;
	N2212GAT<= not N2402GAT;
	N2214GAT<= not N2205GAT;
	N2216GAT<= not N2406GAT;
	N2217GAT<= not N2206GAT;
	N2237GAT<= not N2646GAT;
	N2243GAT<= not N55GAT;
	N2244GAT<= not N567GAT;
	N2245GAT<= not N504GAT;
	N2246GAT<= not N933GAT;
	N2248GAT<= not N3006GAT;
	N2251GAT<= not N3033GAT;
	N2252GAT<= not N2260GAT;
	N2253GAT<= not N2189GAT;
	N2256GAT<= not N3032GAT;
	N2257GAT<= not N2189GAT;
	N2259GAT<= not N3046GAT;
	N2260GAT<= not N2262GAT;
	N2261GAT<= not I3000;
	N2264GAT<= not N2266GAT;
	N2265GAT<= not I3429;
	N2268GAT<= not N2270GAT;
	N2269GAT<= not I2349;
	N2281GAT<= not N3009GAT;
	N2283GAT<= not N2438GAT;
	N2284GAT<= not N2342GAT;
	N2285GAT<= not N2397GAT;
	N2286GAT<= not I1585;
	N2288GAT<= not I4024;
	N2289GAT<= not I1724;
	N2290GAT<= not N2202GAT;
	N2307GAT<= not N2309GAT;
	N2317GAT<= not N2319GAT;
	N2325GAT<= not N3010GAT;
	N2328GAT<= not N3008GAT;
	N2332GAT<= not N3045GAT;
	N2333GAT<= not N2438GAT;
	N2337GAT<= not N2339GAT;
	N2338GAT<= not I2344;
	N2341GAT<= not N2343GAT;
	N2342GAT<= not I1550;
	N2345GAT<= not N2347GAT;
	N2346GAT<= not I2837;
	N2349GAT<= not N2215GAT;
	N2351GAT<= not N2405GAT;
	N2353GAT<= not N2398GAT;
	N2354GAT<= not N2201GAT;
	N2355GAT<= not N2341GAT;
	N2356GAT<= not N2560GAT;
	N2359GAT<= not N2358GAT;
	N2384GAT<= not N43GAT;
	N2385GAT<= not N748GAT;
	N2388GAT<= not N2390GAT;
	N2389GAT<= not I2316;
	N2392GAT<= not N2394GAT;
	N2393GAT<= not I2847;
	N2397GAT<= not N2399GAT;
	N2398GAT<= not I1538;
	N2401GAT<= not N2403GAT;
	N2402GAT<= not I2843;
	N2405GAT<= not N2407GAT;
	N2406GAT<= not I2785;
	N2414GAT<= not I2254;
	N2415GAT<= not I2257;
	N2416GAT<= not I2263;
	N2417GAT<= not I2268;
	N2418GAT<= not I2271;
	N2419GAT<= not I2275;
	N2422GAT<= not N3013GAT;
	N2426GAT<= not N2480GAT;
	N2429GAT<= not N2541GAT;
	N2432GAT<= not N2430GAT;
	N2437GAT<= not N2195GAT;
	N2438GAT<= not N2440GAT;
	N2439GAT<= not I2771;
	N2442GAT<= not N2483GAT;
	N2443GAT<= not N2561GAT;
	N2444GAT<= not N2446GAT;
	N2448GAT<= not N2450GAT;
	N2449GAT<= not I3957;
	N2452GAT<= not N2454GAT;
	N2456GAT<= not N2458GAT;
	N2462GAT<= not N2464GAT;
	N2466GAT<= not N2468GAT;
	N2470GAT<= not N2472GAT;
	N2474GAT<= not N2476GAT;
	N2478GAT<= not N2579GAT;
	N2482GAT<= not N2542GAT;
	N2486GAT<= not N2629GAT;
	N2487GAT<= not N2489GAT;
	N2488GAT<= not N2490GAT;
	N2489GAT<= not I1606;
	N2492GAT<= not N2329GAT;
	N2493GAT<= not N2495GAT;
	N2494GAT<= not I2319;
	N2500GAT<= not N2502GAT;
	N2504GAT<= not N2506GAT;
	N2508GAT<= not N2510GAT;
	N2512GAT<= not N2514GAT;
	N2516GAT<= not N2518GAT;
	N2520GAT<= not N2522GAT;
	N2524GAT<= not N2526GAT;
	N2530GAT<= not N2531GAT;
	N2532GAT<= not N2625GAT;
	N2533GAT<= not N2534GAT;
	N2536GAT<= not N2624GAT;
	N2537GAT<= not N2538GAT;
	N2540GAT<= not N2488GAT;
	N2541GAT<= not N2543GAT;
	N2542GAT<= not I1708;
	N2550GAT<= not I2403;
	N2551GAT<= not I2417;
	N2552GAT<= not I2420;
	N2553GAT<= not I2425;
	N2554GAT<= not I2428;
	N2555GAT<= not I2433;
	N2557GAT<= not N2621GAT;
	N2558GAT<= not N2559GAT;
	N2560GAT<= not N2562GAT;
	N2561GAT<= not I1719;
	N2564GAT<= not N2352GAT;
	N2573GAT<= not I2213;
	N2574GAT<= not I2225;
	N2575GAT<= not I2228;
	N2576GAT<= not I2235;
	N2577GAT<= not I2238;
	N2578GAT<= not I2242;
	N2582GAT<= not I2248;
	N2585GAT<= not I2281;
	N2586GAT<= not N2588GAT;
	N2590GAT<= not N2592GAT;
	N2591GAT<= not I3143;
	N2595GAT<= not N2594GAT;
	N2596GAT<= not N2665GAT;
	N2597GAT<= not N2599GAT;
	N2606GAT<= not I2372;
	N2607GAT<= not I2376;
	N2608GAT<= not I2380;
	N2609GAT<= not I2385;
	N2610GAT<= not I2389;
	N2611GAT<= not I2394;
	N2612GAT<= not N2620GAT;
	N2616GAT<= not I2400;
	N2619GAT<= not I2439;
	N2620GAT<= not N2622GAT;
	N2621GAT<= not I1617;
	N2624GAT<= not N2626GAT;
	N2625GAT<= not I1703;
	N2628GAT<= not N2630GAT;
	N2629GAT<= not I1630;
	N2632GAT<= not N2634GAT;
	N2633GAT<= not I2414;
	N2636GAT<= not N2637GAT;
	N2638GAT<= not N2640GAT;
	N2639GAT<= not I2232;
	N2642GAT<= not N2644GAT;
	N2643GAT<= not I3646;
	N2649GAT<= not I2324;
	N2652GAT<= not I2354;
	N2656GAT<= not N2658GAT;
	N2660GAT<= not N2655GAT;
	N2661GAT<= not N2662GAT;
	N2665GAT<= not I1516;
	N2666GAT<= not N1704GAT;
	N2667GAT<= not I30;
	N2668GAT<= not I27;
	N2669GAT<= not N2671GAT;
	N2670GAT<= not I81;
	N2671GAT<= not I18;
	N2672GAT<= not N2674GAT;
	N2673GAT<= not I384;
	N2674GAT<= not I381;
	N2677GAT<= not I4492;
	N2678GAT<= not I4485;
	N2679GAT<= not I3954;
	N2680GAT<= not I3941;
	N2681GAT<= not I4489;
	N2682GAT<= not I4482;
	N2683GAT<= not I3951;
	N2685GAT<= not N2687GAT;
	N2686GAT<= not I4499;
	N2687GAT<= not I4558;
	N2688GAT<= not I4496;
	N2689GAT<= not I4573;
	N2690GAT<= not I4566;
	N2691GAT<= not N2695GAT;
	N2692GAT<= not I3948;
	N2696GAT<= not I3945;
	N2697GAT<= not I4587;
	N2698GAT<= not I4580;
	N2699GAT<= not N2703GAT;
	N2700GAT<= not I3935;
	N2705GAT<= not I4601;
	N2706GAT<= not I4594;
	N2707GAT<= not I3923;
	N2711GAT<= not N2712GAT;
	N2712GAT<= not I818;
	N2715GAT<= not N2717GAT;
	N2716GAT<= not I240;
	N2717GAT<= not I1;
	N2718GAT<= not N2719GAT;
	N2719GAT<= not I776;
	N2720GAT<= not N2722GAT;
	N2721GAT<= not I594;
	N2722GAT<= not I591;
	N2723GAT<= not N2725GAT;
	N2724GAT<= not I256;
	N2725GAT<= not I5;
	N2726GAT<= not N2728GAT;
	N2727GAT<= not I264;
	N2728GAT<= not I259;
	N2729GAT<= not I512;
	N2730GAT<= not I509;
	N2731GAT<= not N2733GAT;
	N2732GAT<= not I300;
	N2733GAT<= not I297;
	N2734GAT<= not N2736GAT;
	N2735GAT<= not I340;
	N2736GAT<= not I337;
	N2737GAT<= not I4554;
	N2738GAT<= not I4548;
	N2739GAT<= not N2743GAT;
	N2740GAT<= not I4014;
	N2743GAT<= not I4227;
	N2745GAT<= not I4542;
	N2746GAT<= not I4536;
	N2747GAT<= not N2751GAT;
	N2748GAT<= not N2752GAT;
	N2751GAT<= not I4222;
	N2752GAT<= not I4122;
	N2753GAT<= not I4530;
	N2754GAT<= not I4524;
	N2755GAT<= not N2758GAT;
	N2758GAT<= not I4117;
	N2759GAT<= not I4518;
	N2760GAT<= not I4512;
	N2763GAT<= not I4506;
	N2765GAT<= not I4138;
	N2766GAT<= not I4135;
	N2767GAT<= not I14;
	N2768GAT<= not I11;
	N2775GAT<= not N2777GAT;
	N2776GAT<= not I320;
	N2777GAT<= not I317;
	N2778GAT<= not N2780GAT;
	N2779GAT<= not I426;
	N2780GAT<= not I423;
	N2781GAT<= not N2783GAT;
	N2782GAT<= not I50;
	N2783GAT<= not I47;
	N2784GAT<= not N2786GAT;
	N2785GAT<= not I583;
	N2789GAT<= not N2791GAT;
	N2790GAT<= not I65;
	N2791GAT<= not I62;
	N2792GAT<= not N2794GAT;
	N2793GAT<= not I100;
	N2794GAT<= not I97;
	N2795GAT<= not I4615;
	N2796GAT<= not I4608;
	N2797GAT<= not I4020;
	N2801GAT<= not I4633;
	N2802GAT<= not I4623;
	N2803GAT<= not I4478;
	N2804GAT<= not I4236;
	N2805GAT<= not I4630;
	N2806GAT<= not I4620;
	N2807GAT<= not I4475;
	N2808GAT<= not I4233;
	N2809GAT<= not I4642;
	N2810GAT<= not I4332;
	N2811GAT<= not I4312;
	N2813GAT<= not I4329;
	N2814GAT<= not I4309;
	N2815GAT<= not I4372;
	N2816GAT<= not I4352;
	N2817GAT<= not I4369;
	N2818GAT<= not I4349;
	N2819GAT<= not I4651;
	N2820GAT<= not I4412;
	N2821GAT<= not I4392;
	N2823GAT<= not I4409;
	N2824GAT<= not I4389;
	N2825GAT<= not I4452;
	N2826GAT<= not I4432;
	N2827GAT<= not I3962;
	N2828GAT<= not I4449;
	N2829GAT<= not I4429;
	N2831GAT<= not I771;
	N2832GAT<= not I768;
	N2836GAT<= not N2837GAT;
	N2837GAT<= not I941;
	N2838GAT<= not N2839GAT;
	N2839GAT<= not I796;
	N2840GAT<= not N2841GAT;
	N2841GAT<= not I963;
	N2842GAT<= not N2843GAT;
	N2843GAT<= not I985;
	N2844GAT<= not N2845GAT;
	N2845GAT<= not I23;
	N2846GAT<= not N2847GAT;
	N2847GAT<= not I863;
	N2850GAT<= not I579;
	N2851GAT<= not I576;
	N2852GAT<= not N2853GAT;
	N2853GAT<= not I885;
	N2854GAT<= not N2856GAT;
	N2855GAT<= not I227;
	N2856GAT<= not I192;
	N2857GAT<= not N2858GAT;
	N2858GAT<= not I4129;
	N2859GAT<= not N2861GAT;
	N2860GAT<= not I214;
	N2861GAT<= not I199;
	N2862GAT<= not N2864GAT;
	N2863GAT<= not I220;
	N2864GAT<= not I206;
	N2867GAT<= not N2869GAT;
	N2868GAT<= not I248;
	N2869GAT<= not I243;
	N3017GAT<= not I1961;
	N3018GAT<= not I3211;
	N3019GAT<= not I3235;
	N3020GAT<= not I3287;
	N3021GAT<= not I3290;
	N3022GAT<= not I3293;
	N3023GAT<= not I3297;
	N3024GAT<= not I3300;
	N3025GAT<= not I3303;
	N3026GAT<= not I3306;
	N3027GAT<= not I3309;
	N3028GAT<= not I3312;
	N3029GAT<= not I3315;
	N3030GAT<= not I3318;
	N3031GAT<= not I3387;
	N3032GAT<= not I3390;
	N3033GAT<= not I3394;
	N3034GAT<= not I3401;
	N3035GAT<= not I3412;
	N3036GAT<= not I3436;
	N3037GAT<= not I3457;
	N3038GAT<= not I3461;
	N3039GAT<= not I3465;
	N3040GAT<= not I3472;
	N3041GAT<= not I3483;
	N3042GAT<= not I3491;
	N3043GAT<= not I3494;
	N3044GAT<= not I3504;
	N3045GAT<= not I3509;
	N3046GAT<= not I3513;
	N3047GAT<= not I3520;
	N3048GAT<= not I3530;
	N3049GAT<= not I3539;
	N3050GAT<= not I3549;
	N3051GAT<= not I3558;
	N3052GAT<= not I3610;
	N3053GAT<= not I3635;
	N3054GAT<= not I3660;
	N3055GAT<= not I3703;
	N3056GAT<= not I3713;
	N3057GAT<= not I3754;
	N3058GAT<= not I3765;
	N3059GAT<= not I3801;
	N3060GAT<= not I3817;
	N3061GAT<= not I3841;
	N3062GAT<= not I3876;
	N3063GAT<= not I3891;
	N3064GAT<= not I3914;
	N3104GAT<= not I4654;
	N3105GAT<= not I4657;
	N3106GAT<= not I4660;
	N3107GAT<= not I4663;
	N3108GAT<= not I4666;
	N3109GAT<= not I4669;
	N3110GAT<= not I4672;
	N3111GAT<= not I4675;
	N3112GAT<= not I4678;
	N3113GAT<= not I4681;
	N3114GAT<= not I4684;
	N3115GAT<= not I4687;
	N3116GAT<= not I4690;
	N3117GAT<= not I4693;
	N3118GAT<= not I4696;
	N3119GAT<= not I4699;
	N3120GAT<= not I4702;
	N3121GAT<= not I4705;
	N3122GAT<= not I4708;
	N3123GAT<= not I4711;
	N3124GAT<= not I4714;
	N3125GAT<= not I4717;
	N3126GAT<= not I4720;
	N3127GAT<= not I4723;
	N3128GAT<= not I4726;
	N3129GAT<= not I4729;
	N3130GAT<= not I4732;
	N3131GAT<= not I4735;
	N3132GAT<= not I4738;
	N3133GAT<= not I4741;
	N3134GAT<= not I4744;
	N3135GAT<= not I4747;
	N3136GAT<= not I4750;
	N3137GAT<= not I4753;
	N3138GAT<= not I4756;
	N3139GAT<= not I4759;
	N3140GAT<= not I4762;
	N3141GAT<= not I4765;
	N3142GAT<= not I4768;
	N3143GAT<= not I4771;
	N3144GAT<= not I4774;
	N3145GAT<= not I4777;
	N3146GAT<= not I4780;
	N3147GAT<= not I4783;
	N3148GAT<= not I4786;
	N3149GAT<= not I4789;
	N3150GAT<= not I4792;
	N3151GAT<= not I4795;
	N3152GAT<= not I4798;
	I1277<=N2860GAT or N2855GAT or N2863GAT;
	I1278<=N740GAT or N3030GAT or I1277;
	I1515<=N2474GAT or N2524GAT or N2831GAT;
	I1516<=N2466GAT or N2462GAT or I1515;
	I1584<=N2353GAT or N2284GAT or N2354GAT;
	I1585<=N2356GAT or N2214GAT or I1584;
	I1723<=N2354GAT or N2353GAT or N2214GAT;
	I1724<=N2355GAT or N2443GAT or I1723;
	I1733<=N2286GAT or N2428GAT or N2289GAT;
	I1734<=N1604GAT or N2214GAT or I1733;
	I2720<=N1788GAT or N1786GAT or N1839GAT;
	I2721<=N1884GAT or N1783GAT or I2720;
	I2735<=N1788GAT or N1884GAT or N1633GAT;
	I2736<=N1785GAT or N1784GAT or I2735;
	I2812<=N1703GAT or N1704GAT or N1778GAT;
	I2813<=N1609GAT or N1702GAT or N1700GAT or I2812;
	I2831<=N1839GAT or N1786GAT or N1788GAT;
	I2832<=N1884GAT or N1784GAT or I2831;
	I2889<=N1784GAT or N1633GAT or N1884GAT;
	I2890<=N1788GAT or N1786GAT or I2889;
	I2925<=N1784GAT or N1785GAT or N1633GAT;
	I2926<=N1884GAT or N1787GAT or I2925;
	I2934<=N1784GAT or N1839GAT or N1788GAT;
	I2935<=N1785GAT or N1884GAT or I2934;
	I3148<=N1839GAT or N1884GAT or N1784GAT;
	I3149<=N1786GAT or N1787GAT or I3148;
	I3178<=N1838GAT or N1785GAT or N1788GAT;
	I3179<=N1839GAT or N1784GAT or I3178;
	I3999<=N2167GAT or N2031GAT or N2174GAT;
	I4000<=N2108GAT or N2093GAT or N2035GAT or I3999;
	I4023<=N2443GAT or N2290GAT or N2214GAT;
	I4024<=N2353GAT or N2284GAT or I4023;
	I4144<=N1633GAT or N1838GAT or N1786GAT;
	I4145<=N1788GAT or N1784GAT or I4144;
	I4216<=N1427GAT or N1595GAT or N1677GAT;
	I4217<=N1392GAT or N2989GAT or I4216;
	N43GAT<=N44GAT or N45GAT or N46GAT or N47GAT;
	N55GAT<=N56GAT or N57GAT or N58GAT or N59GAT;
	N120GAT<=N121GAT or N122GAT or N123GAT or N124GAT;
	N167GAT<=N168GAT or N169GAT or N170GAT or N171GAT;
	N221GAT<=N222GAT or N223GAT or N224GAT or N225GAT;
	N258GAT<=N259GAT or N260GAT or N261GAT or N262GAT;
	N343GAT<=N344GAT or N345GAT or N346GAT or N347GAT;
	N475GAT<=N476GAT or N477GAT or N478GAT or N479GAT;
	N493GAT<=N494GAT or N495GAT or N496GAT or N497GAT;
	N504GAT<=N505GAT or N506GAT or N507GAT or N508GAT;
	N567GAT<=N568GAT or N569GAT or N570GAT or N571GAT;
	N586GAT<=N587GAT or N588GAT or N589GAT or N590GAT;
	N686GAT<=N687GAT or N688GAT or N689GAT or N690GAT;
	N709GAT<=N710GAT or N711GAT or N712GAT or N713GAT;
	N728GAT<=N729GAT or N730GAT or N731GAT or N732GAT;
	N748GAT<=N749GAT or N750GAT or N751GAT or N752GAT;
	N779GAT<=N780GAT or N781GAT or N782GAT or N783GAT;
	N803GAT<=N804GAT or N805GAT or N806GAT or N807GAT;
	N906GAT<=N907GAT or N908GAT or N909GAT or N910GAT;
	N933GAT<=N934GAT or N935GAT or N936GAT or N937GAT;
	N944GAT<=N945GAT or N946GAT or N947GAT or N948GAT;
	N1013GAT<=N1014GAT or N1015GAT or N1016GAT or N1017GAT;
	N1050GAT<=N1051GAT or N1052GAT or N1053GAT or N1054GAT;
	N1184GAT<=N1185GAT or N1186GAT or N1187GAT or N1188GAT;
	N1201GAT<=N1202GAT or N1203GAT or N1204GAT or N1205GAT;
	N1213GAT<=N1214GAT or N1215GAT or N1216GAT or N1217GAT;
	N1228GAT<=N1229GAT or N1230GAT or N1231GAT or N1232GAT;
	N1269GAT<=N1270GAT or N1271GAT or N1272GAT or N1273GAT;
	N2409GAT<=N2410GAT or N2411GAT or N2412GAT or N2413GAT;
	N2545GAT<=N2546GAT or N2547GAT or N2548GAT or N2549GAT;
	N2568GAT<=N2569GAT or N2570GAT or N2571GAT or N2572GAT;
	N2579GAT<=N2580GAT or N2581GAT;
	N2601GAT<=N2602GAT or N2603GAT or N2604GAT or N2605GAT;
	N2613GAT<=N2614GAT or N2615GAT;
	N2646GAT<=N2647GAT or N2648GAT;
	N2684GAT<=N1599GAT or N2051GAT;
	N2693GAT<=N1451GAT or N1453GAT;
	N2694GAT<=N1381GAT or N1384GAT;
	N2695GAT<=N1586GAT or N1791GAT;
	N2701GAT<=N921GAT or N1890GAT;
	N2702GAT<=N925GAT or N1452GAT;
	N2703GAT<=N1755GAT or N1518GAT;
	N2704GAT<=N11GAT or N1889GAT;
	N2708GAT<=N848GAT or N2047GAT;
	N2709GAT<=N739GAT or N1841GAT;
	N2710GAT<=N69GAT or N1885GAT;
	N2741GAT<=N1182GAT or N2385GAT;
	N2742GAT<=N1005GAT or N2384GAT;
	N2744GAT<=N2159GAT or N2478GAT;
	N2749GAT<=N1010GAT or N2246GAT;
	N2750GAT<=N1181GAT or N2243GAT;
	N2756GAT<=N1011GAT or N2244GAT;
	N2757GAT<=N1030GAT or N2245GAT;
	N2761GAT<=N1031GAT or N2325GAT;
	N2762GAT<=N1028GAT or N1782GAT;
	N2764GAT<=N1029GAT or N2237GAT;
	N2786GAT<=N3091GAT or N3092GAT;
	N2798GAT<=N1032GAT or N2054GAT;
	N2799GAT<=N849GAT or N2050GAT;
	N2800GAT<=N2158GAT or N2186GAT;
	N2812GAT<=N73GAT or N70GAT or N1840GAT;
	N2822GAT<=N77GAT or N13GAT or N1842GAT;
	N2830GAT<=N2444GAT or N1754GAT;
	N2874GAT<=N141GAT or N38GAT or N37GAT;
	N2875GAT<=N142GAT or N40GAT or N39GAT;
	N2876GAT<=N874GAT or N132GAT;
	N2877GAT<=N139GAT or N136GAT;
	N2878GAT<=N234GAT or N137GAT;
	N2879GAT<=N145GAT or N143GAT;
	N2880GAT<=N299GAT or N207GAT;
	N2881GAT<=N324GAT or N238GAT or N237GAT;
	N2882GAT<=N242GAT or N240GAT;
	N2883GAT<=N251GAT or N244GAT;
	N2884GAT<=N246GAT or N245GAT;
	N2885GAT<=N250GAT or N249GAT or N248GAT;
	N2886GAT<=N774GAT or N764GAT or N369GAT;
	N2887GAT<=N791GAT or N650GAT or N370GAT;
	N2888GAT<=N663GAT or N649GAT or N449GAT;
	N2889GAT<=N423GAT or N362GAT;
	N2890GAT<=N654GAT or N557GAT or N371GAT;
	N2891GAT<=N795GAT or N656GAT or N368GAT;
	N2892GAT<=N378GAT or N377GAT;
	N2893GAT<=N391GAT or N390GAT;
	N2894GAT<=N443GAT or N439GAT;
	N2895GAT<=N444GAT or N440GAT;
	N2896GAT<=N647GAT or N441GAT;
	N2897GAT<=N648GAT or N442GAT;
	N2898GAT<=N447GAT or N445GAT;
	N2899GAT<=N772GAT or N451GAT or N446GAT;
	N2900GAT<=N869GAT or N453GAT or N448GAT;
	N2901GAT<=N558GAT or N555GAT or N450GAT;
	N2902GAT<=N460GAT or N459GAT;
	N2903GAT<=N794GAT or N773GAT or N662GAT;
	N2904GAT<=N793GAT or N664GAT or N556GAT;
	N2905GAT<=N964GAT or N961GAT;
	N2906GAT<=N745GAT or N638GAT;
	N2907GAT<=N646GAT or N641GAT;
	N2908GAT<=N763GAT or N642GAT;
	N2909GAT<=N765GAT or N643GAT;
	N2910GAT<=N645GAT or N644GAT;
	N2911GAT<=N761GAT or N651GAT;
	N2912GAT<=N762GAT or N652GAT;
	N2913GAT<=N767GAT or N653GAT;
	N2914GAT<=N768GAT or N655GAT;
	N2915GAT<=N965GAT or N960GAT or N661GAT;
	N2916GAT<=N971GAT or N970GAT or N968GAT;
	N2917GAT<=N1074GAT or N872GAT;
	N2918GAT<=N769GAT or N759GAT;
	N2919GAT<=N766GAT or N760GAT;
	N2920GAT<=N867GAT or N771GAT;
	N2921GAT<=N966GAT or N790GAT;
	N2922GAT<=N967GAT or N792GAT;
	N2923GAT<=N1082GAT or N796GAT;
	N2924GAT<=N871GAT or N797GAT;
	N2925GAT<=N975GAT or N972GAT or N969GAT;
	N2926GAT<=N1083GAT or N1077GAT;
	N2927GAT<=N962GAT or N959GAT;
	N2928GAT<=N963GAT or N868GAT;
	N2929GAT<=N974GAT or N973GAT or N870GAT;
	N2930GAT<=N1153GAT or N1151GAT or N982GAT or N877GAT;
	N2931GAT<=N1100GAT or N994GAT or N989GAT or N880GAT;
	N2932GAT<=N1098GAT or N1090GAT or N986GAT or N885GAT;
	N2933GAT<=N981GAT or N890GAT or N889GAT or N886GAT;
	N2934GAT<=N1104GAT or N887GAT;
	N2935GAT<=N892GAT or N891GAT;
	N2936GAT<=N901GAT or N893GAT;
	N2937GAT<=N900GAT or N895GAT;
	N2938GAT<=N899GAT or N896GAT;
	N2939GAT<=N1091GAT or N1088GAT or N992GAT or N987GAT;
	N2940GAT<=N1152GAT or N1092GAT or N997GAT or N993GAT;
	N2941GAT<=N1003GAT or N902GAT;
	N2942GAT<=N904GAT or N903GAT;
	N2943GAT<=N1012GAT or N905GAT;
	N2944GAT<=N977GAT or N976GAT;
	N2945GAT<=N1096GAT or N1095GAT or N990GAT or N979GAT;
	N2946GAT<=N1099GAT or N998GAT or N995GAT or N980GAT;
	N2947GAT<=N1094GAT or N1093GAT or N988GAT or N984GAT;
	N2948GAT<=N1097GAT or N1089GAT or N1087GAT or N991GAT;
	N2949GAT<=N1101GAT or N996GAT;
	N2950GAT<=N1001GAT or N999GAT;
	N2951GAT<=N1004GAT or N1000GAT;
	N2952GAT<=N1076GAT or N1075GAT;
	N2953GAT<=N1163GAT or N1102GAT;
	N2954GAT<=N1250GAT or N1103GAT;
	N2955GAT<=N1177GAT or N1115GAT;
	N2956GAT<=N1178GAT or N1116GAT;
	N2957GAT<=N1159GAT or N1158GAT or N1156GAT or N1155GAT;
	N2958GAT<=N1246GAT or N1161GAT;
	N2959GAT<=N1305GAT or N1162GAT;
	N2960GAT<=N1175GAT or N1174GAT;
	N2961GAT<=N1375GAT or N1324GAT;
	N2962GAT<=N1176GAT or N1173GAT;
	N2963GAT<=N1291GAT or N1245GAT;
	N2964GAT<=N1304GAT or N1249GAT;
	N2965GAT<=N1267GAT or N1257GAT;
	N2966GAT<=N1368GAT or N1258GAT;
	N2967GAT<=N1262GAT or N1260GAT;
	N2968GAT<=N1326GAT or N1261GAT;
	N2969GAT<=N1323GAT or N1264GAT;
	N2970GAT<=N1383GAT or N1327GAT;
	N2971GAT<=N1287GAT or N1285GAT;
	N2973GAT<=N1352GAT or N1351GAT or N1303GAT or N1302GAT;
	N2974GAT<=N1321GAT or N1320GAT;
	N2975GAT<=N1443GAT or N1325GAT;
	N2977GAT<=N1360GAT or N1359GAT or N1358GAT or N1357GAT;
	N2978GAT<=N1441GAT or N1440GAT or N1371GAT or N1367GAT;
	N2979GAT<=N1373GAT or N1372GAT;
	N2980GAT<=N1470GAT or N1400GAT or N1399GAT or N1398GAT;
	N2981GAT<=N1413GAT or N1408GAT or N1407GAT;
	N2982GAT<=N1504GAT or N1502GAT;
	N2983GAT<=N2079GAT or N2073GAT;
	N2984GAT<=N1467GAT or N1466GAT;
	N2985GAT<=N1686GAT or N1533GAT or N1532GAT or N1531GAT;
	N2986GAT<=N1650GAT or N1649GAT or N1563GAT;
	N2987GAT<=N1574GAT or N1573GAT;
	N2988GAT<=N1733GAT or N1581GAT;
	N2989GAT<=N1693GAT or N1692GAT;
	N2990GAT<=N1710GAT or N1630GAT;
	N2991GAT<=N1654GAT or N1653GAT or N1644GAT;
	N2992GAT<=N1723GAT or N1647GAT or N1646GAT;
	N2993GAT<=N1894GAT or N1847GAT or N1846GAT;
	N2994GAT<=N1954GAT or N1888GAT;
	N2995GAT<=N1962GAT or N1955GAT;
	N2996GAT<=N1960GAT or N1959GAT or N1957GAT;
	N2997GAT<=N2053GAT or N2052GAT or N1964GAT;
	N2998GAT<=N2055GAT or N1967GAT;
	N2999GAT<=N1972GAT or N1971GAT;
	N3000GAT<=N2000GAT or N1999GAT;
	N3001GAT<=N2132GAT or N2130GAT;
	N3002GAT<=N2213GAT or N2150GAT or N2149GAT;
	N3003GAT<=N2256GAT or N2251GAT;
	N3004GAT<=N2258GAT or N2257GAT or N2255GAT;
	N3005GAT<=N2211GAT or N2210GAT;
	N3006GAT<=N2253GAT or N2252GAT;
	N3007GAT<=N2250GAT or N2249GAT;
	N3008GAT<=N2332GAT or N2259GAT;
	N3009GAT<=N2350GAT or N2282GAT;
	N3010GAT<=N2460GAT or N2423GAT;
	N3011GAT<=N2333GAT or N2331GAT;
	N3013GAT<=N2461GAT or N2421GAT;
	N3014GAT<=N2567GAT or N2499GAT;
	N3015GAT<=N2566GAT or N2565GAT;
	N3016GAT<=N2596GAT or N2595GAT;
	N12GAT<= not (N186GAT or N82GAT);
	N13GAT<= not (N2720GAT or N14GAT);
	N15GAT<= not (N637GAT or N17GAT or N293GAT);
	N22GAT<= not (N92GAT or N21GAT);
	N37GAT<= not (N151GAT or N154GAT);
	N38GAT<= not (N151GAT or N233GAT);
	N39GAT<= not (N383GAT or N247GAT);
	N40GAT<= not (N325GAT or N383GAT);
	N44GAT<= not (N48GAT or N49GAT or N50GAT);
	N45GAT<= not (N48GAT or N51GAT or N52GAT);
	N46GAT<= not (N53GAT or N49GAT or N52GAT);
	N47GAT<= not (N53GAT or N51GAT or N50GAT);
	N56GAT<= not (N60GAT or N61GAT or N62GAT);
	N57GAT<= not (N60GAT or N63GAT or N64GAT);
	N58GAT<= not (N65GAT or N61GAT or N64GAT);
	N59GAT<= not (N65GAT or N63GAT or N62GAT);
	N68GAT<= not (N85GAT or N180GAT);
	N70GAT<= not (N71GAT or N2720GAT);
	N73GAT<= not (N67GAT or N2784GAT);
	N77GAT<= not (N76GAT or N2784GAT);
	N78GAT<= not (N2784GAT or N79GAT);
	N82GAT<= not (N16GAT or N295GAT or N637GAT);
	N84GAT<= not (N296GAT or N17GAT or N294GAT);
	N85GAT<= not (N17GAT or N294GAT or N637GAT);
	N86GAT<= not (N743GAT or N294GAT or N17GAT);
	N87GAT<= not (N743GAT or N17GAT or N293GAT);
	N89GAT<= not (N88GAT or N2784GAT);
	N93GAT<= not (N197GAT or N22GAT);
	N110GAT<= not (N182GAT or N89GAT);
	N121GAT<= not (N125GAT or N126GAT or N127GAT);
	N122GAT<= not (N125GAT or N128GAT or N129GAT);
	N123GAT<= not (N130GAT or N126GAT or N129GAT);
	N124GAT<= not (N130GAT or N128GAT or N127GAT);
	N132GAT<= not (N560GAT or N364GAT);
	N136GAT<= not (N253GAT or N154GAT);
	N137GAT<= not (N154GAT or N253GAT);
	N139GAT<= not (N253GAT or N151GAT or N254GAT);
	N140GAT<= not (N151GAT or N253GAT or N155GAT);
	N141GAT<= not (N155GAT or N253GAT or N150GAT);
	N142GAT<= not (N382GAT or N326GAT or N144GAT);
	N143GAT<= not (N326GAT or N247GAT);
	N145GAT<= not (N144GAT or N325GAT);
	N168GAT<= not (N172GAT or N173GAT or N174GAT);
	N169GAT<= not (N172GAT or N175GAT or N176GAT);
	N170GAT<= not (N177GAT or N173GAT or N176GAT);
	N171GAT<= not (N177GAT or N175GAT or N174GAT);
	N180GAT<= not (N286GAT or N188GAT or N287GAT);
	N181GAT<= not (N286GAT or N179GAT or N188GAT);
	N182GAT<= not (N72GAT or N2720GAT);
	N184GAT<= not (N189GAT or N188GAT or N179GAT);
	N186GAT<= not (N189GAT or N287GAT or N288GAT);
	N187GAT<= not (N189GAT or N287GAT or N188GAT);
	N196GAT<= not (N297GAT or N195GAT);
	N197GAT<= not (N194GAT or N297GAT);
	N200GAT<= not (N199GAT or N92GAT);
	N204GAT<= not (N200GAT or N196GAT);
	N207GAT<= not (N2337GAT or N2269GAT);
	N212GAT<= not (N182GAT or N78GAT);
	N222GAT<= not (N226GAT or N227GAT or N228GAT);
	N223GAT<= not (N226GAT or N229GAT or N230GAT);
	N224GAT<= not (N231GAT or N227GAT or N230GAT);
	N225GAT<= not (N231GAT or N229GAT or N228GAT);
	N234GAT<= not (N155GAT or N233GAT);
	N237GAT<= not (N140GAT or N147GAT);
	N238GAT<= not (N147GAT or N254GAT);
	N240GAT<= not (N255GAT or N140GAT);
	N242GAT<= not (N254GAT or N241GAT);
	N244GAT<= not (N334GAT or N386GAT);
	N245GAT<= not (N386GAT or N334GAT);
	N246GAT<= not (N330GAT or N325GAT or N334GAT);
	N247GAT<= not (N334GAT or N387GAT or N330GAT);
	N248GAT<= not (N330GAT or N1490GAT);
	N249GAT<= not (N386GAT or N330GAT);
	N250GAT<= not (N329GAT or N387GAT or N334GAT);
	N251GAT<= not (N1490GAT or N387GAT);
	N259GAT<= not (N263GAT or N264GAT or N265GAT);
	N260GAT<= not (N263GAT or N266GAT or N267GAT);
	N261GAT<= not (N268GAT or N264GAT or N267GAT);
	N262GAT<= not (N268GAT or N266GAT or N265GAT);
	N286GAT<= not (N289GAT or N2723GAT);
	N287GAT<= not (N289GAT or N2715GAT);
	N288GAT<= not (N289GAT or N2726GAT);
	N291GAT<= not (N290GAT or N292GAT);
	N292GAT<= not (N415GAT or N356GAT);
	N299GAT<= not (N2268GAT or N2338GAT);
	N324GAT<= not (N255GAT or N146GAT or N241GAT);
	N344GAT<= not (N348GAT or N349GAT or N350GAT);
	N345GAT<= not (N348GAT or N351GAT or N352GAT);
	N346GAT<= not (N353GAT or N349GAT or N352GAT);
	N347GAT<= not (N353GAT or N351GAT or N350GAT);
	N354GAT<= not (N411GAT or N522GAT);
	N355GAT<= not (N517GAT or N410GAT or N354GAT);
	N356GAT<= not (N2726GAT or N740GAT);
	N357GAT<= not (N2726GAT or N2860GAT);
	N359GAT<= not (N290GAT or N358GAT);
	N360GAT<= not (N2859GAT or N2727GAT);
	N361GAT<= not (N2859GAT or N2726GAT);
	N362GAT<= not (N2723GAT or N2727GAT);
	N377GAT<= not (N110GAT or N2778GAT);
	N378GAT<= not (N375GAT or N235GAT);
	N390GAT<= not (N469GAT or N2877GAT);
	N391GAT<= not (N252GAT or N468GAT);
	N408GAT<= not (N516GAT or N407GAT);
	N409GAT<= not (N406GAT or N407GAT);
	N410GAT<= not (N417GAT or N413GAT or N412GAT or N406GAT);
	N411GAT<= not (N374GAT or N2726GAT);
	N414GAT<= not (N411GAT or N415GAT);
	N415GAT<= not (N2723GAT or N740GAT);
	N418GAT<= not (N374GAT or N2723GAT);
	N419GAT<= not (N409GAT or N291GAT);
	N420GAT<= not (N408GAT or N359GAT);
	N421GAT<= not (N2715GAT or N2723GAT);
	N423GAT<= not (N2724GAT or N2726GAT);
	N439GAT<= not (N856GAT or N2836GAT);
	N440GAT<= not (N856GAT or N2842GAT);
	N441GAT<= not (N856GAT or N2846GAT);
	N442GAT<= not (N2844GAT or N856GAT);
	N443GAT<= not (N2778GAT or N373GAT);
	N444GAT<= not (N373GAT or N2781GAT);
	N445GAT<= not (N2778GAT or N219GAT);
	N446GAT<= not (N219GAT or N2781GAT);
	N447GAT<= not (N2836GAT or N111GAT);
	N448GAT<= not (N111GAT or N2846GAT);
	N449GAT<= not (N2836GAT or N851GAT);
	N450GAT<= not (N851GAT or N2846GAT);
	N451GAT<= not (N134GAT or N372GAT);
	N453GAT<= not (N372GAT or N452GAT);
	N459GAT<= not (N457GAT or N461GAT);
	N460GAT<= not (N462GAT or N2884GAT);
	N476GAT<= not (N480GAT or N481GAT or N482GAT);
	N477GAT<= not (N480GAT or N483GAT or N484GAT);
	N478GAT<= not (N485GAT or N481GAT or N484GAT);
	N479GAT<= not (N485GAT or N483GAT or N482GAT);
	N494GAT<= not (N498GAT or N499GAT or N500GAT);
	N495GAT<= not (N498GAT or N501GAT or N502GAT);
	N496GAT<= not (N503GAT or N499GAT or N502GAT);
	N497GAT<= not (N503GAT or N501GAT or N500GAT);
	N505GAT<= not (N509GAT or N510GAT or N511GAT);
	N506GAT<= not (N509GAT or N512GAT or N513GAT);
	N507GAT<= not (N514GAT or N510GAT or N513GAT);
	N508GAT<= not (N514GAT or N512GAT or N511GAT);
	N516GAT<= not (N374GAT or N2715GAT);
	N518GAT<= not (N520GAT or N519GAT);
	N519GAT<= not (N2854GAT or N374GAT);
	N520GAT<= not (N374GAT or N2862GAT);
	N521GAT<= not (N740GAT or N2715GAT);
	N522GAT<= not (N374GAT or N2859GAT);
	N523GAT<= not (N522GAT or N356GAT);
	N525GAT<= not (N526GAT or N531GAT or N530GAT);
	N526GAT<= not (N2859GAT or N740GAT);
	N529GAT<= not (N2724GAT or N2715GAT);
	N530GAT<= not (N2862GAT or N740GAT);
	N531GAT<= not (N740GAT or N2854GAT);
	N532GAT<= not (N527GAT or N416GAT or N528GAT);
	N555GAT<= not (N852GAT or N2792GAT);
	N556GAT<= not (N2672GAT or N852GAT);
	N557GAT<= not (N2669GAT or N852GAT);
	N564GAT<= not (N3029GAT or N2863GAT or N2855GAT or N374GAT);
	N568GAT<= not (N572GAT or N573GAT or N574GAT);
	N569GAT<= not (N572GAT or N575GAT or N576GAT);
	N570GAT<= not (N577GAT or N573GAT or N576GAT);
	N571GAT<= not (N577GAT or N575GAT or N574GAT);
	N587GAT<= not (N591GAT or N592GAT or N593GAT);
	N588GAT<= not (N591GAT or N594GAT or N595GAT);
	N589GAT<= not (N596GAT or N592GAT or N595GAT);
	N590GAT<= not (N596GAT or N594GAT or N593GAT);
	N629GAT<= not (N414GAT or N634GAT or N523GAT);
	N630GAT<= not (N634GAT or N523GAT or N524GAT);
	N631GAT<= not (N523GAT or N633GAT or N524GAT);
	N632GAT<= not (N414GAT or N523GAT or N633GAT);
	N634GAT<= not (N418GAT or N521GAT);
	N635GAT<= not (N639GAT or N634GAT or N414GAT);
	N636GAT<= not (N414GAT or N633GAT or N639GAT);
	N638GAT<= not (N2715GAT or N2868GAT);
	N645GAT<= not (N2792GAT or N93GAT);
	N646GAT<= not (N93GAT or N2669GAT);
	N647GAT<= not (N2792GAT or N373GAT);
	N648GAT<= not (N373GAT or N2669GAT);
	N649GAT<= not (N2778GAT or N852GAT);
	N650GAT<= not (N852GAT or N2789GAT);
	N651GAT<= not (N93GAT or N2778GAT);
	N652GAT<= not (N2789GAT or N93GAT);
	N653GAT<= not (N2718GAT or N111GAT);
	N654GAT<= not (N851GAT or N2844GAT);
	N655GAT<= not (N856GAT or N2718GAT);
	N656GAT<= not (N851GAT or N2718GAT);
	N687GAT<= not (N691GAT or N692GAT or N693GAT);
	N688GAT<= not (N691GAT or N694GAT or N695GAT);
	N689GAT<= not (N696GAT or N692GAT or N695GAT);
	N690GAT<= not (N696GAT or N694GAT or N693GAT);
	N710GAT<= not (N714GAT or N715GAT or N716GAT);
	N711GAT<= not (N714GAT or N717GAT or N718GAT);
	N712GAT<= not (N719GAT or N715GAT or N718GAT);
	N713GAT<= not (N719GAT or N717GAT or N716GAT);
	N729GAT<= not (N733GAT or N734GAT or N735GAT);
	N730GAT<= not (N733GAT or N736GAT or N737GAT);
	N731GAT<= not (N738GAT or N734GAT or N737GAT);
	N732GAT<= not (N738GAT or N736GAT or N735GAT);
	N745GAT<= not (N2716GAT or N2867GAT);
	N746GAT<= not (N2716GAT or N2723GAT);
	N749GAT<= not (N753GAT or N754GAT or N755GAT);
	N750GAT<= not (N753GAT or N756GAT or N757GAT);
	N751GAT<= not (N758GAT or N754GAT or N757GAT);
	N752GAT<= not (N758GAT or N756GAT or N755GAT);
	N763GAT<= not (N2672GAT or N93GAT);
	N764GAT<= not (N852GAT or N2781GAT);
	N765GAT<= not (N2781GAT or N93GAT);
	N766GAT<= not (N93GAT or N2734GAT);
	N767GAT<= not (N219GAT or N2731GAT);
	N768GAT<= not (N373GAT or N2731GAT);
	N769GAT<= not (N93GAT or N2731GAT);
	N771GAT<= not (N2838GAT or N111GAT);
	N772GAT<= not (N111GAT or N2842GAT);
	N773GAT<= not (N851GAT or N2838GAT);
	N774GAT<= not (N2842GAT or N851GAT);
	N780GAT<= not (N784GAT or N785GAT or N786GAT);
	N781GAT<= not (N784GAT or N787GAT or N788GAT);
	N782GAT<= not (N789GAT or N785GAT or N788GAT);
	N783GAT<= not (N789GAT or N787GAT or N786GAT);
	N790GAT<= not (N856GAT or N2840GAT);
	N791GAT<= not (N851GAT or N2840GAT);
	N792GAT<= not (N2852GAT or N856GAT);
	N793GAT<= not (N2852GAT or N851GAT);
	N794GAT<= not (N852GAT or N2775GAT);
	N795GAT<= not (N2731GAT or N852GAT);
	N796GAT<= not (N2731GAT or N110GAT);
	N797GAT<= not (N110GAT or N2734GAT);
	N801GAT<= not (N672GAT or N670GAT);
	N804GAT<= not (N808GAT or N809GAT or N810GAT);
	N805GAT<= not (N808GAT or N811GAT or N812GAT);
	N806GAT<= not (N813GAT or N809GAT or N812GAT);
	N807GAT<= not (N813GAT or N811GAT or N810GAT);
	N853GAT<= not (N740GAT or N2148GAT);
	N854GAT<= not (N2148GAT or N374GAT);
	N867GAT<= not (N219GAT or N2775GAT);
	N868GAT<= not (N2775GAT or N373GAT);
	N869GAT<= not (N219GAT or N2792GAT);
	N870GAT<= not (N2669GAT or N219GAT);
	N871GAT<= not (N802GAT or N375GAT);
	N872GAT<= not (N375GAT or N800GAT);
	N874GAT<= not (N559GAT or N365GAT);
	N877GAT<= not (N875GAT or N876GAT);
	N879GAT<= not (N2931GAT or N801GAT);
	N880GAT<= not (N926GAT or N566GAT);
	N885GAT<= not (N579GAT or N1112GAT);
	N886GAT<= not (N683GAT or N1112GAT);
	N887GAT<= not (N1603GAT or N683GAT);
	N889GAT<= not (N1111GAT or N1079GAT);
	N890GAT<= not (N741GAT or N702GAT);
	N891GAT<= not (N420GAT or N888GAT);
	N892GAT<= not (N419GAT or N1265GAT);
	N893GAT<= not (N894GAT or N420GAT);
	N895GAT<= not (N420GAT or N898GAT);
	N896GAT<= not (N897GAT or N420GAT);
	N899GAT<= not (N419GAT or N1172GAT);
	N900GAT<= not (N419GAT or N1008GAT);
	N901GAT<= not (N419GAT or N1259GAT);
	N902GAT<= not (N1009GAT or N419GAT);
	N903GAT<= not (N1007GAT or N397GAT);
	N904GAT<= not (N1006GAT or N490GAT);
	N905GAT<= not (N625GAT or N1006GAT);
	N907GAT<= not (N911GAT or N912GAT or N913GAT);
	N908GAT<= not (N911GAT or N914GAT or N915GAT);
	N909GAT<= not (N916GAT or N912GAT or N915GAT);
	N910GAT<= not (N916GAT or N914GAT or N913GAT);
	N934GAT<= not (N938GAT or N939GAT or N940GAT);
	N935GAT<= not (N938GAT or N941GAT or N942GAT);
	N936GAT<= not (N943GAT or N939GAT or N942GAT);
	N937GAT<= not (N943GAT or N941GAT or N940GAT);
	N945GAT<= not (N949GAT or N950GAT or N951GAT);
	N946GAT<= not (N949GAT or N952GAT or N953GAT);
	N947GAT<= not (N954GAT or N950GAT or N953GAT);
	N948GAT<= not (N954GAT or N952GAT or N951GAT);
	N959GAT<= not (N373GAT or N2734GAT);
	N960GAT<= not (N2734GAT or N852GAT);
	N961GAT<= not (N219GAT or N2734GAT);
	N962GAT<= not (N856GAT or N2711GAT);
	N963GAT<= not (N856GAT or N2838GAT);
	N964GAT<= not (N111GAT or N2711GAT);
	N965GAT<= not (N2711GAT or N851GAT);
	N966GAT<= not (N2789GAT or N373GAT);
	N967GAT<= not (N373GAT or N2672GAT);
	N968GAT<= not (N2789GAT or N219GAT);
	N969GAT<= not (N219GAT or N2672GAT);
	N970GAT<= not (N372GAT or N878GAT);
	N971GAT<= not (N111GAT or N2840GAT);
	N972GAT<= not (N372GAT or N458GAT);
	N973GAT<= not (N372GAT or N333GAT);
	N974GAT<= not (N2844GAT or N111GAT);
	N975GAT<= not (N111GAT or N2852GAT);
	N977GAT<= not (N670GAT or N671GAT);
	N978GAT<= not (N2944GAT or N2945GAT);
	N979GAT<= not (N1601GAT or N926GAT);
	N980GAT<= not (N875GAT or N926GAT);
	N981GAT<= not (N926GAT or N873GAT);
	N982GAT<= not (N873GAT or N1478GAT);
	N984GAT<= not (N926GAT or N983GAT);
	N986GAT<= not (N985GAT or N926GAT);
	N987GAT<= not (N741GAT or N159GAT);
	N988GAT<= not (N340GAT or N741GAT);
	N989GAT<= not (N721GAT or N741GAT);
	N990GAT<= not (N841GAT or N741GAT);
	N991GAT<= not (N1112GAT or N679GAT);
	N992GAT<= not (N815GAT or N1112GAT);
	N993GAT<= not (N1112GAT or N698GAT);
	N994GAT<= not (N1112GAT or N882GAT);
	N995GAT<= not (N823GAT or N1112GAT);
	N996GAT<= not (N1603GAT or N823GAT);
	N997GAT<= not (N741GAT or N393GAT);
	N998GAT<= not (N725GAT or N741GAT);
	N999GAT<= not (N419GAT or N1171GAT);
	N1000GAT<= not (N419GAT or N1252GAT);
	N1001GAT<= not (N420GAT or N1002GAT);
	N1003GAT<= not (N420GAT or N879GAT);
	N1004GAT<= not (N978GAT or N420GAT);
	N1005GAT<= not (N894GAT or N455GAT);
	N1008GAT<= not (N2942GAT or N1254GAT);
	N1009GAT<= not (N1255GAT or N2943GAT);
	N1010GAT<= not (N897GAT or N455GAT);
	N1011GAT<= not (N455GAT or N898GAT);
	N1012GAT<= not (N1007GAT or N918GAT);
	N1014GAT<= not (N1018GAT or N1019GAT or N1020GAT);
	N1015GAT<= not (N1018GAT or N1021GAT or N1022GAT);
	N1016GAT<= not (N1023GAT or N1019GAT or N1022GAT);
	N1017GAT<= not (N1023GAT or N1021GAT or N1020GAT);
	N1028GAT<= not (N455GAT or N879GAT);
	N1029GAT<= not (N978GAT or N455GAT);
	N1030GAT<= not (N455GAT or N888GAT);
	N1031GAT<= not (N1002GAT or N455GAT);
	N1051GAT<= not (N1055GAT or N1056GAT or N1057GAT);
	N1052GAT<= not (N1055GAT or N1058GAT or N1059GAT);
	N1053GAT<= not (N1060GAT or N1056GAT or N1059GAT);
	N1054GAT<= not (N1060GAT or N1058GAT or N1057GAT);
	N1074GAT<= not (N2775GAT or N110GAT);
	N1076GAT<= not (N93GAT or N2775GAT);
	N1077GAT<= not (N110GAT or N2672GAT);
	N1082GAT<= not (N375GAT or N380GAT);
	N1083GAT<= not (N381GAT or N375GAT);
	N1087GAT<= not (N926GAT or N1084GAT);
	N1088GAT<= not (N1085GAT or N926GAT);
	N1089GAT<= not (N1067GAT or N1111GAT);
	N1090GAT<= not (N1111GAT or N860GAT);
	N1091GAT<= not (N1111GAT or N956GAT);
	N1092GAT<= not (N1147GAT or N1111GAT);
	N1093GAT<= not (N1111GAT or N864GAT);
	N1094GAT<= not (N1112GAT or N583GAT);
	N1095GAT<= not (N1240GAT or N1111GAT);
	N1096GAT<= not (N819GAT or N1112GAT);
	N1097GAT<= not (N270GAT or N741GAT);
	N1098GAT<= not (N336GAT or N741GAT);
	N1099GAT<= not (N1111GAT or N1293GAT);
	N1100GAT<= not (N1297GAT or N1111GAT);
	N1101GAT<= not (N1590GAT or N1293GAT);
	N1102GAT<= not (N1297GAT or N1590GAT);
	N1103GAT<= not (N956GAT or N1590GAT);
	N1104GAT<= not (N1079GAT or N1590GAT);
	N1113GAT<= not (N393GAT or N701GAT);
	N1114GAT<= not (N725GAT or N721GAT);
	N1115GAT<= not (N1263GAT or N419GAT);
	N1116GAT<= not (N419GAT or N1266GAT);
	N1117GAT<= not (N720GAT or N725GAT);
	N1151GAT<= not (N1301GAT or N1150GAT);
	N1152GAT<= not (N926GAT or N1150GAT);
	N1153GAT<= not (N1414GAT or N566GAT);
	N1154GAT<= not (N1598GAT or N2930GAT or N2957GAT);
	N1155GAT<= not (N1085GAT or N1348GAT);
	N1156GAT<= not (N985GAT or N1307GAT);
	N1158GAT<= not (N983GAT or N1157GAT);
	N1159GAT<= not (N1160GAT or N1084GAT);
	N1161GAT<= not (N583GAT or N1603GAT);
	N1162GAT<= not (N698GAT or N1603GAT);
	N1163GAT<= not (N882GAT or N1603GAT);
	N1171GAT<= not (N2960GAT or N1243GAT);
	N1172GAT<= not (N2961GAT or N1200GAT);
	N1173GAT<= not (N1007GAT or N1025GAT);
	N1174GAT<= not (N845GAT or N1007GAT);
	N1175GAT<= not (N621GAT or N1006GAT);
	N1176GAT<= not (N829GAT or N1006GAT);
	N1177GAT<= not (N1180GAT or N420GAT);
	N1178GAT<= not (N420GAT or N1179GAT);
	N1181GAT<= not (N455GAT or N1179GAT);
	N1182GAT<= not (N1180GAT or N455GAT);
	N1185GAT<= not (N1189GAT or N1190GAT or N1191GAT);
	N1186GAT<= not (N1189GAT or N1192GAT or N1193GAT);
	N1187GAT<= not (N1194GAT or N1190GAT or N1193GAT);
	N1188GAT<= not (N1194GAT or N1192GAT or N1191GAT);
	N1199GAT<= not (N1123GAT or N1284GAT);
	N1200GAT<= not (N1120GAT or N1123GAT);
	N1202GAT<= not (N1206GAT or N1207GAT or N1208GAT);
	N1203GAT<= not (N1206GAT or N1209GAT or N1210GAT);
	N1204GAT<= not (N1211GAT or N1207GAT or N1210GAT);
	N1205GAT<= not (N1211GAT or N1209GAT or N1208GAT);
	N1212GAT<= not (N1123GAT or N1034GAT);
	N1214GAT<= not (N1218GAT or N1219GAT or N1220GAT);
	N1215GAT<= not (N1218GAT or N1221GAT or N1222GAT);
	N1216GAT<= not (N1223GAT or N1219GAT or N1222GAT);
	N1217GAT<= not (N1223GAT or N1221GAT or N1220GAT);
	N1229GAT<= not (N1233GAT or N1234GAT or N1235GAT);
	N1230GAT<= not (N1233GAT or N1236GAT or N1237GAT);
	N1231GAT<= not (N1238GAT or N1234GAT or N1237GAT);
	N1232GAT<= not (N1238GAT or N1236GAT or N1235GAT);
	N1243GAT<= not (N1281GAT or N1123GAT);
	N1244GAT<= not (N1123GAT or N1134GAT);
	N1245GAT<= not (N1590GAT or N860GAT);
	N1246GAT<= not (N864GAT or N1590GAT);
	N1249GAT<= not (N679GAT or N1603GAT);
	N1250GAT<= not (N1603GAT or N815GAT);
	N1251GAT<= not (N1123GAT or N1071GAT);
	N1252GAT<= not (N1199GAT or N2962GAT);
	N1253GAT<= not (N930GAT or N1123GAT);
	N1254GAT<= not (N1123GAT or N1044GAT);
	N1255GAT<= not (N1123GAT or N1225GAT);
	N1256GAT<= not (N392GAT or N702GAT);
	N1257GAT<= not (N1007GAT or N274GAT);
	N1258GAT<= not (N274GAT or N1444GAT);
	N1259GAT<= not (N2967GAT or N1251GAT);
	N1260GAT<= not (N1007GAT or N278GAT);
	N1261GAT<= not (N833GAT or N1006GAT);
	N1262GAT<= not (N837GAT or N1006GAT);
	N1263GAT<= not (N1212GAT or N2968GAT);
	N1264GAT<= not (N1006GAT or N617GAT);
	N1265GAT<= not (N1244GAT or N2969GAT);
	N1266GAT<= not (N2965GAT or N1253GAT);
	N1267GAT<= not (N613GAT or N1006GAT);
	N1270GAT<= not (N1274GAT or N1275GAT or N1276GAT);
	N1271GAT<= not (N1274GAT or N1277GAT or N1278GAT);
	N1272GAT<= not (N1279GAT or N1275GAT or N1278GAT);
	N1273GAT<= not (N1279GAT or N1277GAT or N1276GAT);
	N1285GAT<= not (N1196GAT or N1269GAT);
	N1287GAT<= not (N1284GAT or N1195GAT);
	N1291GAT<= not (N1603GAT or N579GAT);
	N1302GAT<= not (N1300GAT or N1487GAT);
	N1303GAT<= not (N1247GAT or N1355GAT);
	N1304GAT<= not (N1590GAT or N1067GAT);
	N1305GAT<= not (N1147GAT or N1590GAT);
	N1308GAT<= not (N2081GAT or N1530GAT);
	N1318GAT<= not (N392GAT or N701GAT);
	N1320GAT<= not (N1444GAT or N278GAT);
	N1321GAT<= not (N1442GAT or N837GAT);
	N1323GAT<= not (N1007GAT or N401GAT);
	N1324GAT<= not (N164GAT or N1007GAT);
	N1325GAT<= not (N1444GAT or N164GAT);
	N1326GAT<= not (N1007GAT or N282GAT);
	N1327GAT<= not (N1281GAT or N1224GAT);
	N1347GAT<= not (N2081GAT or N1410GAT);
	N1349GAT<= not (N1479GAT or N2081GAT);
	N1351GAT<= not (N1306GAT or N1353GAT);
	N1352GAT<= not (N1248GAT or N1418GAT);
	N1354GAT<= not (N1591GAT or N1530GAT);
	N1357GAT<= not (N1424GAT or N1309GAT);
	N1358GAT<= not (N1425GAT or N1105GAT);
	N1359GAT<= not (N1436GAT or N1106GAT);
	N1360GAT<= not (N1164GAT or N1356GAT);
	N1365GAT<= not (N1479GAT or N1591GAT);
	N1367GAT<= not (N1366GAT or N1374GAT);
	N1368GAT<= not (N1442GAT or N613GAT);
	N1371GAT<= not (N1370GAT or N1369GAT);
	N1372GAT<= not (N282GAT or N1444GAT);
	N1373GAT<= not (N833GAT or N1442GAT);
	N1375GAT<= not (N1006GAT or N706GAT);
	N1376GAT<= not (N724GAT or N720GAT);
	N1377GAT<= not (N724GAT or N721GAT);
	N1383GAT<= not (N1280GAT or N1225GAT);
	N1391GAT<= not (N1513GAT or N2442GAT);
	N1397GAT<= not (N1519GAT or N1401GAT);
	N1398GAT<= not (N1455GAT or N1397GAT);
	N1399GAT<= not (N1806GAT or N1338GAT or N1584GAT);
	N1400GAT<= not (N1674GAT or N1403GAT);
	N1401GAT<= not (N1584GAT or N1590GAT);
	N1402GAT<= not (N1858GAT or N1393GAT or N1604GAT);
	N1406GAT<= not (N1428GAT or N1387GAT);
	N1407GAT<= not (N1393GAT or N1409GAT or N1677GAT);
	N1408GAT<= not (N1507GAT or N1396GAT or N1393GAT);
	N1411GAT<= not (N1154GAT or N1608GAT);
	N1412GAT<= not (N1411GAT or N1406GAT or N2981GAT);
	N1413GAT<= not (N1869GAT or N672GAT or N2591GAT);
	N1415GAT<= not (N2081GAT or N2359GAT);
	N1416GAT<= not (N2081GAT or N1480GAT);
	N1417GAT<= not (N2162GAT or N1480GAT);
	N1419GAT<= not (N2162GAT or N1479GAT);
	N1420GAT<= not (N1410GAT or N2162GAT);
	N1421GAT<= not (N2162GAT or N2359GAT);
	N1422GAT<= not (N2011GAT or N2162GAT);
	N1423GAT<= not (N2162GAT or N1530GAT);
	N1426GAT<= not (N2011GAT or N1591GAT);
	N1428GAT<= not (N2978GAT or N2982GAT or N2973GAT or N2977GAT);
	N1435GAT<= not (N1591GAT or N1528GAT);
	N1438GAT<= not (N1591GAT or N1480GAT);
	N1440GAT<= not (N1322GAT or N1439GAT);
	N1441GAT<= not (N1437GAT or N1378GAT);
	N1443GAT<= not (N1442GAT or N706GAT);
	N1458GAT<= not (N1510GAT or N1459GAT);
	N1459GAT<= not (N1595GAT or N1454GAT);
	N1466GAT<= not (N1392GAT or N1461GAT or N1396GAT);
	N1467GAT<= not (N2289GAT or N1468GAT);
	N1469GAT<= not (N1858GAT or N1608GAT);
	N1470GAT<= not (N1472GAT or N1747GAT);
	N1471GAT<= not (N1334GAT or N1858GAT or N1604GAT);
	N1472GAT<= not (N1476GAT or N1471GAT or N1469GAT);
	N1476GAT<= not (N1858GAT or N1590GAT);
	N1481GAT<= not (N2081GAT or N2011GAT);
	N1483GAT<= not (N2081GAT or N1482GAT);
	N1484GAT<= not (N2081GAT or N1528GAT);
	N1485GAT<= not (N1482GAT or N2162GAT);
	N1486GAT<= not (N1482GAT or N1591GAT);
	N1494GAT<= not (N1528GAT or N2162GAT);
	N1498GAT<= not (N1609GAT or N1427GAT);
	N1499GAT<= not (N396GAT or N401GAT);
	N1501GAT<= not (N1448GAT or N1500GAT);
	N1502GAT<= not (N1607GAT or N1449GAT);
	N1504GAT<= not (N1450GAT or N1498GAT);
	N1510GAT<= not (N1584GAT or N1460GAT);
	N1516GAT<= not (N1551GAT or N1517GAT);
	N1519GAT<= not (N1584GAT or N1339GAT or N1600GAT);
	N1521GAT<= not (N2283GAT or N1991GAT);
	N1529GAT<= not (N1528GAT or N1523GAT);
	N1531GAT<= not (N1507GAT or N1477GAT);
	N1532GAT<= not (N1677GAT or N1458GAT);
	N1533GAT<= not (N1524GAT or N1403GAT);
	N1555GAT<= not (N1616GAT or N1559GAT or N1499GAT);
	N1556GAT<= not (N1614GAT or N1645GAT or N1616GAT);
	N1557GAT<= not (N1553GAT or N1645GAT or N1614GAT);
	N1558GAT<= not (N1614GAT or N1553GAT or N1499GAT);
	N1563GAT<= not (N1561GAT or N1562GAT or N1659GAT);
	N1564GAT<= not (N1584GAT or N1719GAT or N1790GAT or N1576GAT);
	N1565GAT<= not (N1735GAT or N1552GAT);
	N1567GAT<= not (N1634GAT or N1735GAT);
	N1570GAT<= not (N1736GAT or N1658GAT or N1670GAT);
	N1571GAT<= not (N1670GAT or N1658GAT or N1797GAT);
	N1573GAT<= not (N1444GAT or N1858GAT or N1635GAT);
	N1574GAT<= not (N1719GAT or N1673GAT or N1444GAT);
	N1575GAT<= not (N1918GAT or N2283GAT);
	N1576GAT<= not (N2351GAT or N1988GAT or N1661GAT);
	N1577GAT<= not (N1520GAT or N2351GAT or N1988GAT);
	N1578GAT<= not (N2152GAT or N2351GAT or N1665GAT);
	N1581GAT<= not (N1858GAT or N1580GAT);
	N1582GAT<= not (N2283GAT or N1991GAT or N2212GAT);
	N1586GAT<= not (N1869GAT or N1683GAT);
	N1593GAT<= not (N1551GAT or N1310GAT);
	N1598GAT<= not (N1592GAT or N2422GAT);
	N1599GAT<= not (N1691GAT or N336GAT);
	N1600GAT<= not (N1685GAT or N1427GAT);
	N1602GAT<= not (N1594GAT or N1587GAT or N2989GAT);
	N1604GAT<= not (N1778GAT or N1609GAT or N1702GAT or N1700GAT);
	N1605GAT<= not (N1614GAT or N1616GAT or N1499GAT or N396GAT);
	N1606GAT<= not (N3020GAT or N270GAT);
	N1607GAT<= not (N2082GAT or N1609GAT);
	N1608GAT<= not (N1704GAT or N1703GAT);
	N1609GAT<= not (N1503GAT or N3025GAT);
	N1610GAT<= not (N1698GAT or N1543GAT);
	N1613GAT<= not (N1544GAT or N1698GAT);
	N1614GAT<= not (N396GAT or N845GAT);
	N1616GAT<= not (N918GAT or N396GAT);
	N1617GAT<= not (N1319GAT or N1448GAT);
	N1618GAT<= not (N1319GAT or N1447GAT);
	N1619GAT<= not (N1447GAT or N1446GAT);
	N1620GAT<= not (N1448GAT or N1446GAT);
	N1621GAT<= not (N1319GAT or N1380GAT);
	N1622GAT<= not (N1380GAT or N1446GAT);
	N1623GAT<= not (N1379GAT or N1446GAT);
	N1624GAT<= not (N1319GAT or N1379GAT);
	N1625GAT<= not (N3021GAT or N1628GAT);
	N1626GAT<= not (N1627GAT or N3022GAT);
	N1630GAT<= not (N1895GAT or N1631GAT);
	N1636GAT<= not (N1584GAT or N1718GAT);
	N1639GAT<= not (N1499GAT or N1559GAT or N1553GAT);
	N1641GAT<= not (N1645GAT or N1553GAT or N1559GAT);
	N1642GAT<= not (N1559GAT or N1616GAT or N1645GAT);
	N1644GAT<= not (N1643GAT or N1648GAT or N1659GAT);
	N1646GAT<= not (N1569GAT or N1659GAT or N1566GAT);
	N1647GAT<= not (N1656GAT or N1659GAT or N1554GAT);
	N1649GAT<= not (N1560GAT or N1659GAT or N1730GAT);
	N1650GAT<= not (N1727GAT or N1659GAT or N1640GAT);
	N1653GAT<= not (N1651GAT or N1652GAT or N1659GAT);
	N1654GAT<= not (N1671GAT or N1659GAT);
	N1655GAT<= not (N1736GAT or N1662GAT or N1658GAT);
	N1657GAT<= not (N1662GAT or N1797GAT or N1658GAT);
	N1660GAT<= not (N1918GAT or N1986GAT or N2212GAT);
	N1663GAT<= not (N1986GAT or N1918GAT);
	N1666GAT<= not (N1986GAT or N2212GAT or N1991GAT);
	N1667GAT<= not (N1991GAT or N1986GAT);
	N1669GAT<= not (N1668GAT or N1742GAT or N1670GAT);
	N1686GAT<= not (N1774GAT or N1869GAT or N1684GAT);
	N1690GAT<= not (N1700GAT or N1702GAT);
	N1692GAT<= not (N1879GAT or N1762GAT);
	N1695GAT<= not (N1609GAT or N1778GAT or N1704GAT or N1703GAT);
	N1696GAT<= not (N1707GAT or N1698GAT);
	N1700GAT<= not (N1701GAT or N3023GAT);
	N1702GAT<= not (N3024GAT or N1615GAT);
	N1703GAT<= not (N1705GAT or N3028GAT);
	N1704GAT<= not (N3027GAT or N1706GAT);
	N1710GAT<= not (N1709GAT or N1629GAT);
	N1721GAT<= not (N2442GAT or N1690GAT or N1978GAT);
	N1723GAT<= not (N1659GAT or N1722GAT or N1724GAT);
	N1726GAT<= not (N2992GAT or N2986GAT or N2991GAT);
	N1728GAT<= not (N1568GAT or N1736GAT or N1658GAT);
	N1729GAT<= not (N1658GAT or N1797GAT or N1568GAT);
	N1731GAT<= not (N1658GAT or N1515GAT or N1797GAT);
	N1732GAT<= not (N1515GAT or N1736GAT or N1658GAT);
	N1733GAT<= not (N1673GAT or N1572GAT);
	N1734GAT<= not (N1988GAT or N2212GAT);
	N1737GAT<= not (N2212GAT or N2152GAT);
	N1745GAT<= not (N1869GAT or N1757GAT);
	N1755GAT<= not (N1769GAT or N1773GAT or N2512GAT);
	N1756GAT<= not (N2512GAT or N1769GAT or N1773GAT);
	N1757GAT<= not (N1773GAT or N1769GAT);
	N1758GAT<= not (N1311GAT or N1773GAT);
	N1759GAT<= not (N1818GAT or N1935GAT or N2765GAT);
	N1760GAT<= not (N1681GAT or N1602GAT or N2985GAT);
	N1761GAT<= not (N2985GAT or N1602GAT or N1681GAT);
	N1778GAT<= not (N3026GAT or N1779GAT);
	N1780GAT<= not (N1777GAT or N1625GAT or N1626GAT);
	N1792GAT<= not (N1794GAT or N1796GAT);
	N1793GAT<= not (N1792GAT or N1735GAT);
	N1794GAT<= not (N1673GAT or N1719GAT);
	N1796GAT<= not (N1858GAT or N1635GAT);
	N1798GAT<= not (N1739GAT or N1673GAT);
	N1800GAT<= not (N1635GAT or N1919GAT);
	N1801GAT<= not (N2152GAT or N1989GAT);
	N1817GAT<= not (N1819GAT or N1823GAT);
	N1818GAT<= not (N1823GAT or N2005GAT);
	N1827GAT<= not (N2729GAT or N2317GAT);
	N1831GAT<= not (N1832GAT or N1765GAT or N1878GAT);
	N1846GAT<= not (N1845GAT or N1893GAT);
	N1847GAT<= not (N1958GAT or N1845GAT);
	N1860GAT<= not (N1988GAT or N2216GAT or N1862GAT);
	N1861GAT<= not (N1866GAT or N2216GAT or N1988GAT);
	N1863GAT<= not (N1991GAT or N2283GAT or N1989GAT);
	N1864GAT<= not (N1858GAT or N1495GAT or N2090GAT);
	N1865GAT<= not (N1989GAT or N1918GAT or N1986GAT);
	N1882GAT<= not (N2124GAT or N2115GAT or N2239GAT);
	N1894GAT<= not (N1968GAT or N1891GAT or N1969GAT);
	N1895GAT<= not (N1845GAT or N1891GAT or N1968GAT);
	N1896GAT<= not (N2995GAT or N1895GAT);
	N1915GAT<= not (N1859GAT or N1919GAT);
	N1916GAT<= not (N1917GAT or N1859GAT);
	N1920GAT<= not (N1864GAT or N1921GAT or N1798GAT);
	N1921GAT<= not (N1738GAT or N1673GAT);
	N1924GAT<= not (N1743GAT or N1923GAT);
	N1926GAT<= not (N1925GAT or N1635GAT);
	N1927GAT<= not (N1790GAT or N1635GAT);
	N1929GAT<= not (N1758GAT or N1790GAT);
	N1934GAT<= not (N2470GAT or N1935GAT or N2239GAT);
	N1935GAT<= not (N1816GAT or N1828GAT);
	N1957GAT<= not (N1886GAT or N1887GAT);
	N1958GAT<= not (N1963GAT or N1886GAT);
	N1959GAT<= not (N1956GAT or N1963GAT);
	N1962GAT<= not (N1963GAT or N1893GAT);
	N1964GAT<= not (N2392GAT or N2439GAT);
	N1967GAT<= not (N1893GAT or N1968GAT);
	N1971GAT<= not (N1896GAT or N1973GAT);
	N1972GAT<= not (N1974GAT or N1970GAT);
	N1994GAT<= not (N1719GAT or N1922GAT);
	N2005GAT<= not (N2002GAT or N2857GAT);
	N2008GAT<= not (N2012GAT or N1774GAT);
	N2009GAT<= not (N2016GAT or N2664GAT or N2004GAT);
	N2014GAT<= not (N2035GAT or N2093GAT or N2018GAT or N2664GAT);
	N2015GAT<= not (N2039GAT or N1774GAT or N1315GAT);
	N2016GAT<= not (N2019GAT or N1878GAT);
	N2017GAT<= not (N1790GAT or N2016GAT);
	N2018GAT<= not (N2016GAT or N2097GAT);
	N2053GAT<= not (N2393GAT or N2438GAT);
	N2055GAT<= not (N1891GAT or N1958GAT);
	N2057GAT<= not (N2049GAT or N1855GAT);
	N2073GAT<= not (N2078GAT or N1990GAT or N2181GAT);
	N2078GAT<= not (N1926GAT or N1916GAT or N1994GAT or N1924GAT);
	N2079GAT<= not (N2078GAT or N2178GAT or N1990GAT or N2128GAT);
	N2129GAT<= not (N2189GAT or N2134GAT or N2261GAT);
	N2130GAT<= not (N2134GAT or N2185GAT);
	N2132GAT<= not (N2133GAT or N2131GAT);
	N2147GAT<= not (N2988GAT or N1855GAT);
	N2149GAT<= not (N2193GAT or N2346GAT);
	N2150GAT<= not (N2401GAT or N2346GAT);
	N2163GAT<= not (N1790GAT or N1310GAT or N2664GAT or N2168GAT);
	N2185GAT<= not (N2261GAT or N2189GAT);
	N2192GAT<= not (N2184GAT or N1855GAT);
	N2193GAT<= not (N2393GAT or N2439GAT);
	N2194GAT<= not (N2187GAT or N1855GAT);
	N2195GAT<= not (N2200GAT or N1855GAT);
	N2196GAT<= not (N2199GAT or N2146GAT);
	N2197GAT<= not (N2199GAT or N2281GAT);
	N2198GAT<= not (N2199GAT or N2058GAT);
	N2210GAT<= not (N2401GAT or N2151GAT);
	N2211GAT<= not (N2193GAT or N2402GAT);
	N2213GAT<= not (N2402GAT or N2151GAT or N2345GAT);
	N2215GAT<= not (N2346GAT or N2151GAT or N2402GAT);
	N2218GAT<= not (N2214GAT or N2290GAT);
	N2219GAT<= not (N2354GAT or N2214GAT);
	N2220GAT<= not (N2290GAT or N2217GAT);
	N2223GAT<= not (N2354GAT or N2217GAT);
	N2238GAT<= not (N2448GAT or N2444GAT);
	N2239GAT<= not (N2850GAT or N3019GAT);
	N2249GAT<= not (N2265GAT or N3006GAT);
	N2250GAT<= not (N2248GAT or N2264GAT);
	N2255GAT<= not (N2261GAT or N2188GAT);
	N2258GAT<= not (N2260GAT or N2189GAT);
	N2282GAT<= not (N2406GAT or N2215GAT);
	N2291GAT<= not (N2353GAT or N2355GAT or N2443GAT);
	N2292GAT<= not (N2443GAT or N2284GAT or N2285GAT);
	N2293GAT<= not (N2353GAT or N2284GAT or N2443GAT);
	N2306GAT<= not (N2356GAT or N2284GAT or N2285GAT);
	N2329GAT<= not (N1855GAT or N3007GAT);
	N2330GAT<= not (N2437GAT or N1961GAT);
	N2331GAT<= not (N2393GAT or N2401GAT);
	N2350GAT<= not (N2405GAT or N2349GAT);
	N2352GAT<= not (N3011GAT or N2215GAT);
	N2357GAT<= not (N2285GAT or N2355GAT or N2443GAT);
	N2358GAT<= not (N2285GAT or N2356GAT or N2355GAT);
	N2363GAT<= not (N2353GAT or N2356GAT or N2355GAT);
	N2364GAT<= not (N2353GAT or N2284GAT or N2356GAT);
	N2387GAT<= not (N2056GAT or N2437GAT);
	N2396GAT<= not (N2199GAT or N2209GAT);
	N2410GAT<= not (N2414GAT or N2415GAT or N2416GAT);
	N2411GAT<= not (N2414GAT or N2417GAT or N2418GAT);
	N2412GAT<= not (N2419GAT or N2415GAT or N2418GAT);
	N2413GAT<= not (N2419GAT or N2417GAT or N2416GAT);
	N2421GAT<= not (N1601GAT or N1704GAT);
	N2423GAT<= not (N665GAT or N1601GAT);
	N2427GAT<= not (N2426GAT or N2153GAT);
	N2428GAT<= not (N2433GAT or N2427GAT);
	N2430GAT<= not (N2533GAT or N2486GAT or N2429GAT);
	N2433GAT<= not (N2432GAT or N2154GAT);
	N2436GAT<= not (N2437GAT or N1892GAT);
	N2460GAT<= not (N666GAT or N120GAT);
	N2461GAT<= not (N120GAT or N2666GAT);
	N2480GAT<= not (N2530GAT or N2482GAT or N2486GAT);
	N2483GAT<= not (N2537GAT or N2482GAT or N2486GAT);
	N2498GAT<= not (N2199GAT or N2328GAT);
	N2499GAT<= not (N2389GAT or N2494GAT);
	N2531GAT<= not (N2488GAT or N2625GAT or N2621GAT);
	N2534GAT<= not (N2624GAT or N2489GAT or N2621GAT);
	N2538GAT<= not (N2620GAT or N2625GAT or N2488GAT);
	N2539GAT<= not (N2048GAT or N2437GAT);
	N2546GAT<= not (N2550GAT or N2551GAT or N2552GAT);
	N2547GAT<= not (N2550GAT or N2553GAT or N2554GAT);
	N2548GAT<= not (N2555GAT or N2551GAT or N2554GAT);
	N2549GAT<= not (N2555GAT or N2553GAT or N2552GAT);
	N2556GAT<= not (N1711GAT or N2437GAT);
	N2559GAT<= not (N2999GAT or N2437GAT);
	N2565GAT<= not (N2352GAT or N2642GAT);
	N2566GAT<= not (N2643GAT or N2564GAT);
	N2567GAT<= not (N2493GAT or N2388GAT);
	N2569GAT<= not (N2573GAT or N2574GAT or N2575GAT);
	N2570GAT<= not (N2573GAT or N2576GAT or N2577GAT);
	N2571GAT<= not (N2578GAT or N2574GAT or N2577GAT);
	N2572GAT<= not (N2578GAT or N2576GAT or N2575GAT);
	N2580GAT<= not (N2582GAT or N2583GAT);
	N2581GAT<= not (N2583GAT or N2585GAT);
	N2583GAT<= not (N2582GAT or N2585GAT);
	N2594GAT<= not (N3017GAT or N2520GAT or N2597GAT);
	N2602GAT<= not (N2606GAT or N2607GAT or N2608GAT);
	N2603GAT<= not (N2606GAT or N2609GAT or N2610GAT);
	N2604GAT<= not (N2611GAT or N2607GAT or N2610GAT);
	N2605GAT<= not (N2611GAT or N2609GAT or N2608GAT);
	N2614GAT<= not (N2616GAT or N2617GAT);
	N2615GAT<= not (N2617GAT or N2619GAT);
	N2617GAT<= not (N2616GAT or N2619GAT);
	N2637GAT<= not (N3015GAT or N2199GAT);
	N2647GAT<= not (N2649GAT or N2650GAT);
	N2648GAT<= not (N2650GAT or N2652GAT);
	N2650GAT<= not (N2649GAT or N2652GAT);
	N2655GAT<= not (N2508GAT or N2656GAT or N2500GAT or N2504GAT);
	N2662GAT<= not (N2660GAT or N2586GAT);
	N2663GAT<= not (N2586GAT or N2660GAT or N2307GAT);
	N2664GAT<= not (N2850GAT or N3018GAT);
end RTL;
