-- File created by Bench2VHDL
-- Name: s838
-- File: bench/s838.bench
-- Timestamp: 2019-05-21T22:08:28.059388
--
-- Original File
-- =============
--	# s838
--	# 35 inputs
--	# 2 outputs
--	# 32 D-type flipflops
--	# 149 inverters
--	# 241 gates (58 ANDs + 89 NANDs + 16 ORs + 78 NORs)
--	
--	INPUT(X)
--	INPUT(Clear)
--	INPUT(C_32)
--	INPUT(C_31)
--	INPUT(C_30)
--	INPUT(C_29)
--	INPUT(C_28)
--	INPUT(C_27)
--	INPUT(C_26)
--	INPUT(C_25)
--	INPUT(C_24)
--	INPUT(C_23)
--	INPUT(C_22)
--	INPUT(C_21)
--	INPUT(C_20)
--	INPUT(C_19)
--	INPUT(C_18)
--	INPUT(C_17)
--	INPUT(C_16)
--	INPUT(C_15)
--	INPUT(C_14)
--	INPUT(C_13)
--	INPUT(C_12)
--	INPUT(C_11)
--	INPUT(C_10)
--	INPUT(C_9)
--	INPUT(C_8)
--	INPUT(C_7)
--	INPUT(C_6)
--	INPUT(C_5)
--	INPUT(C_4)
--	INPUT(C_3)
--	INPUT(C_2)
--	INPUT(C_1)
--	INPUT(C_0)
--	
--	OUTPUT(W)
--	OUTPUT(Z)
--	
--	Y_4 = DFF(II3)
--	Y_3 = DFF(II4)
--	Y_2 = DFF(II5)
--	Y_1 = DFF(II6)
--	Y_8 = DFF(II155)
--	Y_7 = DFF(II156)
--	Y_6 = DFF(II157)
--	Y_5 = DFF(II158)
--	Y_12 = DFF(II307)
--	Y_11 = DFF(II308)
--	Y_10 = DFF(II309)
--	Y_9 = DFF(II310)
--	Y_16 = DFF(II459)
--	Y_15 = DFF(II460)
--	Y_14 = DFF(II461)
--	Y_13 = DFF(II462)
--	Y_20 = DFF(II611)
--	Y_19 = DFF(II612)
--	Y_18 = DFF(II613)
--	Y_17 = DFF(II614)
--	Y_24 = DFF(II763)
--	Y_23 = DFF(II764)
--	Y_22 = DFF(II765)
--	Y_21 = DFF(II766)
--	Y_28 = DFF(II915)
--	Y_27 = DFF(II916)
--	Y_26 = DFF(II917)
--	Y_25 = DFF(II918)
--	Y_32 = DFF(II1067)
--	Y_31 = DFF(II1068)
--	Y_30 = DFF(II1069)
--	Y_29 = DFF(II1070)
--	
--	II6 = NOT(II104)
--	II50 = NOT(II92)
--	II40 = NOT(X)
--	II41 = NOT(Y_4)
--	II42 = NOT(Y_3)
--	II43 = NOT(Y_2)
--	II44 = NOT(Y_1)
--	II3 = NOT(II46)
--	II4 = NOT(II47)
--	II158 = NOT(II256)
--	II202 = NOT(II244)
--	II192 = NOT(II1_1)
--	II193 = NOT(Y_8)
--	II194 = NOT(Y_7)
--	II195 = NOT(Y_6)
--	II196 = NOT(Y_5)
--	II155 = NOT(II198)
--	II156 = NOT(II199)
--	II310 = NOT(II408)
--	II354 = NOT(II396)
--	II344 = NOT(II1_2)
--	II345 = NOT(Y_12)
--	II346 = NOT(Y_11)
--	II347 = NOT(Y_10)
--	II348 = NOT(Y_9)
--	II307 = NOT(II350)
--	II308 = NOT(II351)
--	II462 = NOT(II560)
--	II506 = NOT(II548)
--	II496 = NOT(II1_3)
--	II497 = NOT(Y_16)
--	II498 = NOT(Y_15)
--	II499 = NOT(Y_14)
--	II500 = NOT(Y_13)
--	II459 = NOT(II502)
--	II460 = NOT(II503)
--	II614 = NOT(II712)
--	II658 = NOT(II700)
--	II648 = NOT(II1_4)
--	II649 = NOT(Y_20)
--	II650 = NOT(Y_19)
--	II651 = NOT(Y_18)
--	II652 = NOT(Y_17)
--	II611 = NOT(II654)
--	II612 = NOT(II655)
--	II766 = NOT(II864)
--	II810 = NOT(II852)
--	II800 = NOT(II1_5)
--	II801 = NOT(Y_24)
--	II802 = NOT(Y_23)
--	II803 = NOT(Y_22)
--	II804 = NOT(Y_21)
--	II763 = NOT(II806)
--	II764 = NOT(II807)
--	II918 = NOT(II1016)
--	II962 = NOT(II1004)
--	II952 = NOT(II1_6)
--	II953 = NOT(Y_28)
--	II954 = NOT(Y_27)
--	II955 = NOT(Y_26)
--	II956 = NOT(Y_25)
--	II915 = NOT(II958)
--	II916 = NOT(II959)
--	II1070 = NOT(II1168)
--	II1114 = NOT(II1156)
--	II1104 = NOT(II1_7)
--	II1105 = NOT(Y_32)
--	II1106 = NOT(Y_31)
--	II1107 = NOT(Y_30)
--	II1108 = NOT(Y_29)
--	II1067 = NOT(II1110)
--	II1068 = NOT(II1111)
--	II1219_1 = NOT(II1253)
--	II1230 = NOT(II1253)
--	II1221 = NOT(Y_1)
--	II1222 = NOT(Y_2)
--	II1223 = NOT(Y_3)
--	P_1 = NOT(II1226)
--	P_3 = NOT(II1228)
--	P_4 = NOT(II1229)
--	II1219_2 = NOT(II1316)
--	II1290 = NOT(II1316)
--	II1280 = NOT(Y_4)
--	II1281 = NOT(Y_5)
--	II1282 = NOT(Y_6)
--	II1283 = NOT(Y_7)
--	P_7 = NOT(II1288)
--	P_8 = NOT(II1289)
--	II1329 = NOT(II1328)
--	II1219_3 = NOT(II1384)
--	II1358 = NOT(II1384)
--	II1348 = NOT(Y_8)
--	II1349 = NOT(Y_9)
--	II1350 = NOT(Y_10)
--	II1351 = NOT(Y_11)
--	P_11 = NOT(II1356)
--	P_12 = NOT(II1357)
--	II1397 = NOT(II1396)
--	II1219_4 = NOT(II1452)
--	II1426 = NOT(II1452)
--	II1416 = NOT(Y_12)
--	II1417 = NOT(Y_13)
--	II1418 = NOT(Y_14)
--	II1419 = NOT(Y_15)
--	P_15 = NOT(II1424)
--	P_16 = NOT(II1425)
--	II1465 = NOT(II1464)
--	II1219_5 = NOT(II1520)
--	II1494 = NOT(II1520)
--	II1484 = NOT(Y_16)
--	II1485 = NOT(Y_17)
--	II1486 = NOT(Y_18)
--	II1487 = NOT(Y_19)
--	P_19 = NOT(II1492)
--	P_20 = NOT(II1493)
--	II1533 = NOT(II1532)
--	II1219_6 = NOT(II1588)
--	II1562 = NOT(II1588)
--	II1552 = NOT(Y_20)
--	II1553 = NOT(Y_21)
--	II1554 = NOT(Y_22)
--	II1555 = NOT(Y_23)
--	P_23 = NOT(II1560)
--	P_24 = NOT(II1561)
--	II1601 = NOT(II1600)
--	II1219_7 = NOT(II1656)
--	II1630 = NOT(II1656)
--	II1620 = NOT(Y_24)
--	II1621 = NOT(Y_25)
--	II1622 = NOT(Y_26)
--	II1623 = NOT(Y_27)
--	P_27 = NOT(II1628)
--	P_28 = NOT(II1629)
--	II1669 = NOT(II1668)
--	II1688 = NOT(Y_28)
--	II1689 = NOT(Y_29)
--	II1690 = NOT(Y_30)
--	II1691 = NOT(Y_31)
--	II1692 = NOT(Y_32)
--	P_30 = NOT(II1694)
--	II1947 = NOT(II1948)
--	II1951 = NOT(II1952)
--	II1955 = NOT(II1956)
--	II1963 = NOT(II1964)
--	II1965 = NOT(II1966)
--	II1971 = NOT(II1972)
--	II1973 = NOT(II1974)
--	II1996 = NOT(II1995)
--	II2002 = NOT(II2001)
--	
--	II127_1 = AND(II41, Y_3, II109)
--	II127_2 = AND(II96, II113, Y_4)
--	II131_1 = AND(II113, II92, Y_3)
--	II131_2 = AND(II42, II109)
--	II279_1 = AND(II193, Y_7, II261)
--	II279_2 = AND(II248, II265, Y_8)
--	II283_1 = AND(II265, II244, Y_7)
--	II283_2 = AND(II194, II261)
--	II431_1 = AND(II345, Y_11, II413)
--	II431_2 = AND(II400, II417, Y_12)
--	II435_1 = AND(II417, II396, Y_11)
--	II435_2 = AND(II346, II413)
--	II583_1 = AND(II497, Y_15, II565)
--	II583_2 = AND(II552, II569, Y_16)
--	II587_1 = AND(II569, II548, Y_15)
--	II587_2 = AND(II498, II565)
--	II735_1 = AND(II649, Y_19, II717)
--	II735_2 = AND(II704, II721, Y_20)
--	II739_1 = AND(II721, II700, Y_19)
--	II739_2 = AND(II650, II717)
--	II887_1 = AND(II801, Y_23, II869)
--	II887_2 = AND(II856, II873, Y_24)
--	II891_1 = AND(II873, II852, Y_23)
--	II891_2 = AND(II802, II869)
--	II1039_1 = AND(II953, Y_27, II1021)
--	II1039_2 = AND(II1008, II1025, Y_28)
--	II1043_1 = AND(II1025, II1004, Y_27)
--	II1043_2 = AND(II954, II1021)
--	II1191_1 = AND(II1105, Y_31, II1173)
--	II1191_2 = AND(II1160, II1177, Y_32)
--	II1195_1 = AND(II1177, II1156, Y_31)
--	II1195_2 = AND(II1106, II1173)
--	II2017_1 = AND(P_29, C_29)
--	II2017_2 = AND(P_19, C_19)
--	II2021_1 = AND(P_30, C_30)
--	II2021_2 = AND(P_31, C_31)
--	II2025_1 = AND(P_32, C_32)
--	II2025_2 = AND(P_24, C_24)
--	II2029_1 = AND(P_23, C_23)
--	II2032_1 = AND(P_28, C_28)
--	II2032_2 = AND(P_11, C_11)
--	II2032_3 = AND(P_15, C_15)
--	II2037_1 = AND(P_14, C_14)
--	II2040_1 = AND(P_7, C_7)
--	II2043_1 = AND(P_18, C_18)
--	II2043_2 = AND(P_20, C_20)
--	II2047_1 = AND(P_10, C_10)
--	II2047_2 = AND(P_3, C_3)
--	II2051_1 = AND(P_8, C_8)
--	II2051_2 = AND(P_27, C_27)
--	II2055_1 = AND(P_26, C_26)
--	II2055_2 = AND(P_2, C_2)
--	II2059_1 = AND(X, C_0)
--	II2059_2 = AND(P_25, C_25)
--	II2063_1 = AND(P_16, C_16)
--	II2063_2 = AND(P_5, C_5)
--	II2070_1 = AND(P_13, C_13)
--	II2070_2 = AND(P_9, C_9)
--	
--	II135_1 = OR(II43, II104)
--	II135_2 = OR(Y_2, II100)
--	II287_1 = OR(II195, II256)
--	II287_2 = OR(Y_6, II252)
--	II439_1 = OR(II347, II408)
--	II439_2 = OR(Y_10, II404)
--	II591_1 = OR(II499, II560)
--	II591_2 = OR(Y_14, II556)
--	II743_1 = OR(II651, II712)
--	II743_2 = OR(Y_18, II708)
--	II895_1 = OR(II803, II864)
--	II895_2 = OR(Y_22, II860)
--	II1047_1 = OR(II955, II1016)
--	II1047_2 = OR(Y_26, II1012)
--	II1199_1 = OR(II1107, II1168)
--	II1199_2 = OR(Y_30, II1164)
--	
--	II5 = NAND(II135_1, II135_2)
--	II92 = NAND(Y_2, Y_1)
--	II96 = NAND(Y_3, II50)
--	II100 = NAND(Y_1, II113)
--	II104 = NAND(II44, II113)
--	II157 = NAND(II287_1, II287_2)
--	II244 = NAND(Y_6, Y_5)
--	II248 = NAND(Y_7, II202)
--	II252 = NAND(Y_5, II265)
--	II256 = NAND(II196, II265)
--	II309 = NAND(II439_1, II439_2)
--	II396 = NAND(Y_10, Y_9)
--	II400 = NAND(Y_11, II354)
--	II404 = NAND(Y_9, II417)
--	II408 = NAND(II348, II417)
--	II461 = NAND(II591_1, II591_2)
--	II548 = NAND(Y_14, Y_13)
--	II552 = NAND(Y_15, II506)
--	II556 = NAND(Y_13, II569)
--	II560 = NAND(II500, II569)
--	II613 = NAND(II743_1, II743_2)
--	II700 = NAND(Y_18, Y_17)
--	II704 = NAND(Y_19, II658)
--	II708 = NAND(Y_17, II721)
--	II712 = NAND(II652, II721)
--	II765 = NAND(II895_1, II895_2)
--	II852 = NAND(Y_22, Y_21)
--	II856 = NAND(Y_23, II810)
--	II860 = NAND(Y_21, II873)
--	II864 = NAND(II804, II873)
--	II917 = NAND(II1047_1, II1047_2)
--	II1004 = NAND(Y_26, Y_25)
--	II1008 = NAND(Y_27, II962)
--	II1012 = NAND(Y_25, II1025)
--	II1016 = NAND(II956, II1025)
--	II1069 = NAND(II1199_1, II1199_2)
--	II1156 = NAND(Y_30, Y_29)
--	II1160 = NAND(Y_31, II1114)
--	II1164 = NAND(Y_29, II1177)
--	II1168 = NAND(II1108, II1177)
--	II1226 = NAND(X, Y_1)
--	II1228 = NAND(Y_3, II1259)
--	II1229 = NAND(Y_4, II1230)
--	II1253 = NAND(II1223, II1259)
--	II1262 = NAND(X, II1221)
--	II1288 = NAND(Y_7, II1321)
--	II1289 = NAND(Y_8, II1290)
--	II1316 = NAND(II1283, II1321)
--	II1324 = NAND(II1281, II1329)
--	II1328 = NAND(II1219_1, II1280)
--	II1356 = NAND(Y_11, II1389)
--	II1357 = NAND(Y_12, II1358)
--	II1384 = NAND(II1351, II1389)
--	II1392 = NAND(II1349, II1397)
--	II1396 = NAND(II1219_2, II1348)
--	II1424 = NAND(Y_15, II1457)
--	II1425 = NAND(Y_16, II1426)
--	II1452 = NAND(II1419, II1457)
--	II1460 = NAND(II1417, II1465)
--	II1464 = NAND(II1219_3, II1416)
--	II1492 = NAND(Y_19, II1525)
--	II1493 = NAND(Y_20, II1494)
--	II1520 = NAND(II1487, II1525)
--	II1528 = NAND(II1485, II1533)
--	II1532 = NAND(II1219_4, II1484)
--	II1560 = NAND(Y_23, II1593)
--	II1561 = NAND(Y_24, II1562)
--	II1588 = NAND(II1555, II1593)
--	II1596 = NAND(II1553, II1601)
--	II1600 = NAND(II1219_5, II1552)
--	II1628 = NAND(Y_27, II1661)
--	II1629 = NAND(Y_28, II1630)
--	II1656 = NAND(II1623, II1661)
--	II1664 = NAND(II1621, II1669)
--	II1668 = NAND(II1219_6, II1620)
--	II1694 = NAND(Y_30, II1726)
--	II1698 = NAND(II1726, II1690)
--	II1729 = NAND(II1688, II1219_7)
--	Z = NAND(II2002, II2008, II1996, II1976)
--	II1821 = NAND(P_1, C_1)
--	II1833 = NAND(P_4, C_4)
--	II1841 = NAND(P_6, C_6)
--	II1865 = NAND(P_12, C_12)
--	II1885 = NAND(P_17, C_17)
--	II1901 = NAND(P_21, C_21)
--	II1905 = NAND(P_22, C_22)
--	II1995 = NAND(II1986, II1990, II1982, II1885)
--	II1997 = NAND(II1950, II1833, II1821, II1905)
--	II2001 = NAND(II1865, II1841, II1978, II1901)
--	
--	II1_1 = NOR(II41, II96)
--	II46 = NOR(II127_1, II127_2)
--	II47 = NOR(II131_1, II131_2)
--	II109 = NOR(II43, II100)
--	II113 = NOR(Clear, II40)
--	II1_2 = NOR(II193, II248)
--	II198 = NOR(II279_1, II279_2)
--	II199 = NOR(II283_1, II283_2)
--	II261 = NOR(II195, II252)
--	II265 = NOR(Clear, II192)
--	II1_3 = NOR(II345, II400)
--	II350 = NOR(II431_1, II431_2)
--	II351 = NOR(II435_1, II435_2)
--	II413 = NOR(II347, II404)
--	II417 = NOR(Clear, II344)
--	II1_4 = NOR(II497, II552)
--	II502 = NOR(II583_1, II583_2)
--	II503 = NOR(II587_1, II587_2)
--	II565 = NOR(II499, II556)
--	II569 = NOR(Clear, II496)
--	II1_5 = NOR(II649, II704)
--	II654 = NOR(II735_1, II735_2)
--	II655 = NOR(II739_1, II739_2)
--	II717 = NOR(II651, II708)
--	II721 = NOR(Clear, II648)
--	II1_6 = NOR(II801, II856)
--	II806 = NOR(II887_1, II887_2)
--	II807 = NOR(II891_1, II891_2)
--	II869 = NOR(II803, II860)
--	II873 = NOR(Clear, II800)
--	II1_7 = NOR(II953, II1008)
--	II958 = NOR(II1039_1, II1039_2)
--	II959 = NOR(II1043_1, II1043_2)
--	II1021 = NOR(II955, II1012)
--	II1025 = NOR(Clear, II952)
--	W = NOR(II1105, II1160)
--	II1110 = NOR(II1191_1, II1191_2)
--	II1111 = NOR(II1195_1, II1195_2)
--	II1173 = NOR(II1107, II1164)
--	II1177 = NOR(Clear, II1104)
--	P_2 = NOR(II1222, II1262)
--	II1259 = NOR(Y_2, II1262)
--	P_5 = NOR(II1281, II1328)
--	P_6 = NOR(II1282, II1324)
--	II1321 = NOR(Y_6, II1324)
--	P_9 = NOR(II1349, II1396)
--	P_10 = NOR(II1350, II1392)
--	II1389 = NOR(Y_10, II1392)
--	P_13 = NOR(II1417, II1464)
--	P_14 = NOR(II1418, II1460)
--	II1457 = NOR(Y_14, II1460)
--	P_17 = NOR(II1485, II1532)
--	P_18 = NOR(II1486, II1528)
--	II1525 = NOR(Y_18, II1528)
--	P_21 = NOR(II1553, II1600)
--	P_22 = NOR(II1554, II1596)
--	II1593 = NOR(Y_22, II1596)
--	P_25 = NOR(II1621, II1668)
--	P_26 = NOR(II1622, II1664)
--	II1661 = NOR(Y_26, II1664)
--	P_29 = NOR(II1689, II1729)
--	P_31 = NOR(II1691, II1698)
--	P_32 = NOR(Y_31, II1698, II1692)
--	II1726 = NOR(II1729, Y_29)
--	II1948 = NOR(II2017_1, II2017_2)
--	II1950 = NOR(II2021_1, II2021_2)
--	II1952 = NOR(II2025_1, II2025_2)
--	II1956 = NOR(II1951, II2029_1)
--	II1964 = NOR(II2032_1, II2032_2, II2032_3)
--	II1966 = NOR(II1955, II2037_1)
--	II1972 = NOR(II1947, II2040_1)
--	II1974 = NOR(II2043_1, II2043_2)
--	II1976 = NOR(II2047_1, II2047_2, II1963)
--	II1978 = NOR(II2051_1, II2051_2, II1971)
--	II1982 = NOR(II2055_1, II2055_2, II1965)
--	II1986 = NOR(II2059_1, II2059_2)
--	II1990 = NOR(II2063_1, II2063_2, II1973)
--	II2008 = NOR(II2070_1, II2070_2, II1997)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s838 is
	port (
		CLEAR: in std_logic;
		CLK: in std_logic;
		C_0: in std_logic;
		C_1: in std_logic;
		C_2: in std_logic;
		C_3: in std_logic;
		C_4: in std_logic;
		C_5: in std_logic;
		C_6: in std_logic;
		C_7: in std_logic;
		C_8: in std_logic;
		C_9: in std_logic;
		C_10: in std_logic;
		C_11: in std_logic;
		C_12: in std_logic;
		C_13: in std_logic;
		C_14: in std_logic;
		C_15: in std_logic;
		C_16: in std_logic;
		C_17: in std_logic;
		C_18: in std_logic;
		C_19: in std_logic;
		C_20: in std_logic;
		C_21: in std_logic;
		C_22: in std_logic;
		C_23: in std_logic;
		C_24: in std_logic;
		C_25: in std_logic;
		C_26: in std_logic;
		C_27: in std_logic;
		C_28: in std_logic;
		C_29: in std_logic;
		C_30: in std_logic;
		C_31: in std_logic;
		C_32: in std_logic;
		X: in std_logic;
		W: out std_logic;
		Z: out std_logic
	);
end entity;

architecture RTL of s838 is
	attribute dont_touch: boolean;

	signal II1_1: std_logic; attribute dont_touch of II1_1: signal is true;
	signal II1_2: std_logic; attribute dont_touch of II1_2: signal is true;
	signal II1_3: std_logic; attribute dont_touch of II1_3: signal is true;
	signal II1_4: std_logic; attribute dont_touch of II1_4: signal is true;
	signal II1_5: std_logic; attribute dont_touch of II1_5: signal is true;
	signal II1_6: std_logic; attribute dont_touch of II1_6: signal is true;
	signal II1_7: std_logic; attribute dont_touch of II1_7: signal is true;
	signal II3: std_logic; attribute dont_touch of II3: signal is true;
	signal II4: std_logic; attribute dont_touch of II4: signal is true;
	signal II5: std_logic; attribute dont_touch of II5: signal is true;
	signal II6: std_logic; attribute dont_touch of II6: signal is true;
	signal II40: std_logic; attribute dont_touch of II40: signal is true;
	signal II41: std_logic; attribute dont_touch of II41: signal is true;
	signal II42: std_logic; attribute dont_touch of II42: signal is true;
	signal II43: std_logic; attribute dont_touch of II43: signal is true;
	signal II44: std_logic; attribute dont_touch of II44: signal is true;
	signal II46: std_logic; attribute dont_touch of II46: signal is true;
	signal II47: std_logic; attribute dont_touch of II47: signal is true;
	signal II50: std_logic; attribute dont_touch of II50: signal is true;
	signal II92: std_logic; attribute dont_touch of II92: signal is true;
	signal II96: std_logic; attribute dont_touch of II96: signal is true;
	signal II100: std_logic; attribute dont_touch of II100: signal is true;
	signal II104: std_logic; attribute dont_touch of II104: signal is true;
	signal II109: std_logic; attribute dont_touch of II109: signal is true;
	signal II113: std_logic; attribute dont_touch of II113: signal is true;
	signal II127_1: std_logic; attribute dont_touch of II127_1: signal is true;
	signal II127_2: std_logic; attribute dont_touch of II127_2: signal is true;
	signal II131_1: std_logic; attribute dont_touch of II131_1: signal is true;
	signal II131_2: std_logic; attribute dont_touch of II131_2: signal is true;
	signal II135_1: std_logic; attribute dont_touch of II135_1: signal is true;
	signal II135_2: std_logic; attribute dont_touch of II135_2: signal is true;
	signal II155: std_logic; attribute dont_touch of II155: signal is true;
	signal II156: std_logic; attribute dont_touch of II156: signal is true;
	signal II157: std_logic; attribute dont_touch of II157: signal is true;
	signal II158: std_logic; attribute dont_touch of II158: signal is true;
	signal II192: std_logic; attribute dont_touch of II192: signal is true;
	signal II193: std_logic; attribute dont_touch of II193: signal is true;
	signal II194: std_logic; attribute dont_touch of II194: signal is true;
	signal II195: std_logic; attribute dont_touch of II195: signal is true;
	signal II196: std_logic; attribute dont_touch of II196: signal is true;
	signal II198: std_logic; attribute dont_touch of II198: signal is true;
	signal II199: std_logic; attribute dont_touch of II199: signal is true;
	signal II202: std_logic; attribute dont_touch of II202: signal is true;
	signal II244: std_logic; attribute dont_touch of II244: signal is true;
	signal II248: std_logic; attribute dont_touch of II248: signal is true;
	signal II252: std_logic; attribute dont_touch of II252: signal is true;
	signal II256: std_logic; attribute dont_touch of II256: signal is true;
	signal II261: std_logic; attribute dont_touch of II261: signal is true;
	signal II265: std_logic; attribute dont_touch of II265: signal is true;
	signal II279_1: std_logic; attribute dont_touch of II279_1: signal is true;
	signal II279_2: std_logic; attribute dont_touch of II279_2: signal is true;
	signal II283_1: std_logic; attribute dont_touch of II283_1: signal is true;
	signal II283_2: std_logic; attribute dont_touch of II283_2: signal is true;
	signal II287_1: std_logic; attribute dont_touch of II287_1: signal is true;
	signal II287_2: std_logic; attribute dont_touch of II287_2: signal is true;
	signal II307: std_logic; attribute dont_touch of II307: signal is true;
	signal II308: std_logic; attribute dont_touch of II308: signal is true;
	signal II309: std_logic; attribute dont_touch of II309: signal is true;
	signal II310: std_logic; attribute dont_touch of II310: signal is true;
	signal II344: std_logic; attribute dont_touch of II344: signal is true;
	signal II345: std_logic; attribute dont_touch of II345: signal is true;
	signal II346: std_logic; attribute dont_touch of II346: signal is true;
	signal II347: std_logic; attribute dont_touch of II347: signal is true;
	signal II348: std_logic; attribute dont_touch of II348: signal is true;
	signal II350: std_logic; attribute dont_touch of II350: signal is true;
	signal II351: std_logic; attribute dont_touch of II351: signal is true;
	signal II354: std_logic; attribute dont_touch of II354: signal is true;
	signal II396: std_logic; attribute dont_touch of II396: signal is true;
	signal II400: std_logic; attribute dont_touch of II400: signal is true;
	signal II404: std_logic; attribute dont_touch of II404: signal is true;
	signal II408: std_logic; attribute dont_touch of II408: signal is true;
	signal II413: std_logic; attribute dont_touch of II413: signal is true;
	signal II417: std_logic; attribute dont_touch of II417: signal is true;
	signal II431_1: std_logic; attribute dont_touch of II431_1: signal is true;
	signal II431_2: std_logic; attribute dont_touch of II431_2: signal is true;
	signal II435_1: std_logic; attribute dont_touch of II435_1: signal is true;
	signal II435_2: std_logic; attribute dont_touch of II435_2: signal is true;
	signal II439_1: std_logic; attribute dont_touch of II439_1: signal is true;
	signal II439_2: std_logic; attribute dont_touch of II439_2: signal is true;
	signal II459: std_logic; attribute dont_touch of II459: signal is true;
	signal II460: std_logic; attribute dont_touch of II460: signal is true;
	signal II461: std_logic; attribute dont_touch of II461: signal is true;
	signal II462: std_logic; attribute dont_touch of II462: signal is true;
	signal II496: std_logic; attribute dont_touch of II496: signal is true;
	signal II497: std_logic; attribute dont_touch of II497: signal is true;
	signal II498: std_logic; attribute dont_touch of II498: signal is true;
	signal II499: std_logic; attribute dont_touch of II499: signal is true;
	signal II500: std_logic; attribute dont_touch of II500: signal is true;
	signal II502: std_logic; attribute dont_touch of II502: signal is true;
	signal II503: std_logic; attribute dont_touch of II503: signal is true;
	signal II506: std_logic; attribute dont_touch of II506: signal is true;
	signal II548: std_logic; attribute dont_touch of II548: signal is true;
	signal II552: std_logic; attribute dont_touch of II552: signal is true;
	signal II556: std_logic; attribute dont_touch of II556: signal is true;
	signal II560: std_logic; attribute dont_touch of II560: signal is true;
	signal II565: std_logic; attribute dont_touch of II565: signal is true;
	signal II569: std_logic; attribute dont_touch of II569: signal is true;
	signal II583_1: std_logic; attribute dont_touch of II583_1: signal is true;
	signal II583_2: std_logic; attribute dont_touch of II583_2: signal is true;
	signal II587_1: std_logic; attribute dont_touch of II587_1: signal is true;
	signal II587_2: std_logic; attribute dont_touch of II587_2: signal is true;
	signal II591_1: std_logic; attribute dont_touch of II591_1: signal is true;
	signal II591_2: std_logic; attribute dont_touch of II591_2: signal is true;
	signal II611: std_logic; attribute dont_touch of II611: signal is true;
	signal II612: std_logic; attribute dont_touch of II612: signal is true;
	signal II613: std_logic; attribute dont_touch of II613: signal is true;
	signal II614: std_logic; attribute dont_touch of II614: signal is true;
	signal II648: std_logic; attribute dont_touch of II648: signal is true;
	signal II649: std_logic; attribute dont_touch of II649: signal is true;
	signal II650: std_logic; attribute dont_touch of II650: signal is true;
	signal II651: std_logic; attribute dont_touch of II651: signal is true;
	signal II652: std_logic; attribute dont_touch of II652: signal is true;
	signal II654: std_logic; attribute dont_touch of II654: signal is true;
	signal II655: std_logic; attribute dont_touch of II655: signal is true;
	signal II658: std_logic; attribute dont_touch of II658: signal is true;
	signal II700: std_logic; attribute dont_touch of II700: signal is true;
	signal II704: std_logic; attribute dont_touch of II704: signal is true;
	signal II708: std_logic; attribute dont_touch of II708: signal is true;
	signal II712: std_logic; attribute dont_touch of II712: signal is true;
	signal II717: std_logic; attribute dont_touch of II717: signal is true;
	signal II721: std_logic; attribute dont_touch of II721: signal is true;
	signal II735_1: std_logic; attribute dont_touch of II735_1: signal is true;
	signal II735_2: std_logic; attribute dont_touch of II735_2: signal is true;
	signal II739_1: std_logic; attribute dont_touch of II739_1: signal is true;
	signal II739_2: std_logic; attribute dont_touch of II739_2: signal is true;
	signal II743_1: std_logic; attribute dont_touch of II743_1: signal is true;
	signal II743_2: std_logic; attribute dont_touch of II743_2: signal is true;
	signal II763: std_logic; attribute dont_touch of II763: signal is true;
	signal II764: std_logic; attribute dont_touch of II764: signal is true;
	signal II765: std_logic; attribute dont_touch of II765: signal is true;
	signal II766: std_logic; attribute dont_touch of II766: signal is true;
	signal II800: std_logic; attribute dont_touch of II800: signal is true;
	signal II801: std_logic; attribute dont_touch of II801: signal is true;
	signal II802: std_logic; attribute dont_touch of II802: signal is true;
	signal II803: std_logic; attribute dont_touch of II803: signal is true;
	signal II804: std_logic; attribute dont_touch of II804: signal is true;
	signal II806: std_logic; attribute dont_touch of II806: signal is true;
	signal II807: std_logic; attribute dont_touch of II807: signal is true;
	signal II810: std_logic; attribute dont_touch of II810: signal is true;
	signal II852: std_logic; attribute dont_touch of II852: signal is true;
	signal II856: std_logic; attribute dont_touch of II856: signal is true;
	signal II860: std_logic; attribute dont_touch of II860: signal is true;
	signal II864: std_logic; attribute dont_touch of II864: signal is true;
	signal II869: std_logic; attribute dont_touch of II869: signal is true;
	signal II873: std_logic; attribute dont_touch of II873: signal is true;
	signal II887_1: std_logic; attribute dont_touch of II887_1: signal is true;
	signal II887_2: std_logic; attribute dont_touch of II887_2: signal is true;
	signal II891_1: std_logic; attribute dont_touch of II891_1: signal is true;
	signal II891_2: std_logic; attribute dont_touch of II891_2: signal is true;
	signal II895_1: std_logic; attribute dont_touch of II895_1: signal is true;
	signal II895_2: std_logic; attribute dont_touch of II895_2: signal is true;
	signal II915: std_logic; attribute dont_touch of II915: signal is true;
	signal II916: std_logic; attribute dont_touch of II916: signal is true;
	signal II917: std_logic; attribute dont_touch of II917: signal is true;
	signal II918: std_logic; attribute dont_touch of II918: signal is true;
	signal II952: std_logic; attribute dont_touch of II952: signal is true;
	signal II953: std_logic; attribute dont_touch of II953: signal is true;
	signal II954: std_logic; attribute dont_touch of II954: signal is true;
	signal II955: std_logic; attribute dont_touch of II955: signal is true;
	signal II956: std_logic; attribute dont_touch of II956: signal is true;
	signal II958: std_logic; attribute dont_touch of II958: signal is true;
	signal II959: std_logic; attribute dont_touch of II959: signal is true;
	signal II962: std_logic; attribute dont_touch of II962: signal is true;
	signal II1004: std_logic; attribute dont_touch of II1004: signal is true;
	signal II1008: std_logic; attribute dont_touch of II1008: signal is true;
	signal II1012: std_logic; attribute dont_touch of II1012: signal is true;
	signal II1016: std_logic; attribute dont_touch of II1016: signal is true;
	signal II1021: std_logic; attribute dont_touch of II1021: signal is true;
	signal II1025: std_logic; attribute dont_touch of II1025: signal is true;
	signal II1039_1: std_logic; attribute dont_touch of II1039_1: signal is true;
	signal II1039_2: std_logic; attribute dont_touch of II1039_2: signal is true;
	signal II1043_1: std_logic; attribute dont_touch of II1043_1: signal is true;
	signal II1043_2: std_logic; attribute dont_touch of II1043_2: signal is true;
	signal II1047_1: std_logic; attribute dont_touch of II1047_1: signal is true;
	signal II1047_2: std_logic; attribute dont_touch of II1047_2: signal is true;
	signal II1067: std_logic; attribute dont_touch of II1067: signal is true;
	signal II1068: std_logic; attribute dont_touch of II1068: signal is true;
	signal II1069: std_logic; attribute dont_touch of II1069: signal is true;
	signal II1070: std_logic; attribute dont_touch of II1070: signal is true;
	signal II1104: std_logic; attribute dont_touch of II1104: signal is true;
	signal II1105: std_logic; attribute dont_touch of II1105: signal is true;
	signal II1106: std_logic; attribute dont_touch of II1106: signal is true;
	signal II1107: std_logic; attribute dont_touch of II1107: signal is true;
	signal II1108: std_logic; attribute dont_touch of II1108: signal is true;
	signal II1110: std_logic; attribute dont_touch of II1110: signal is true;
	signal II1111: std_logic; attribute dont_touch of II1111: signal is true;
	signal II1114: std_logic; attribute dont_touch of II1114: signal is true;
	signal II1156: std_logic; attribute dont_touch of II1156: signal is true;
	signal II1160: std_logic; attribute dont_touch of II1160: signal is true;
	signal II1164: std_logic; attribute dont_touch of II1164: signal is true;
	signal II1168: std_logic; attribute dont_touch of II1168: signal is true;
	signal II1173: std_logic; attribute dont_touch of II1173: signal is true;
	signal II1177: std_logic; attribute dont_touch of II1177: signal is true;
	signal II1191_1: std_logic; attribute dont_touch of II1191_1: signal is true;
	signal II1191_2: std_logic; attribute dont_touch of II1191_2: signal is true;
	signal II1195_1: std_logic; attribute dont_touch of II1195_1: signal is true;
	signal II1195_2: std_logic; attribute dont_touch of II1195_2: signal is true;
	signal II1199_1: std_logic; attribute dont_touch of II1199_1: signal is true;
	signal II1199_2: std_logic; attribute dont_touch of II1199_2: signal is true;
	signal II1219_1: std_logic; attribute dont_touch of II1219_1: signal is true;
	signal II1219_2: std_logic; attribute dont_touch of II1219_2: signal is true;
	signal II1219_3: std_logic; attribute dont_touch of II1219_3: signal is true;
	signal II1219_4: std_logic; attribute dont_touch of II1219_4: signal is true;
	signal II1219_5: std_logic; attribute dont_touch of II1219_5: signal is true;
	signal II1219_6: std_logic; attribute dont_touch of II1219_6: signal is true;
	signal II1219_7: std_logic; attribute dont_touch of II1219_7: signal is true;
	signal II1221: std_logic; attribute dont_touch of II1221: signal is true;
	signal II1222: std_logic; attribute dont_touch of II1222: signal is true;
	signal II1223: std_logic; attribute dont_touch of II1223: signal is true;
	signal II1226: std_logic; attribute dont_touch of II1226: signal is true;
	signal II1228: std_logic; attribute dont_touch of II1228: signal is true;
	signal II1229: std_logic; attribute dont_touch of II1229: signal is true;
	signal II1230: std_logic; attribute dont_touch of II1230: signal is true;
	signal II1253: std_logic; attribute dont_touch of II1253: signal is true;
	signal II1259: std_logic; attribute dont_touch of II1259: signal is true;
	signal II1262: std_logic; attribute dont_touch of II1262: signal is true;
	signal II1280: std_logic; attribute dont_touch of II1280: signal is true;
	signal II1281: std_logic; attribute dont_touch of II1281: signal is true;
	signal II1282: std_logic; attribute dont_touch of II1282: signal is true;
	signal II1283: std_logic; attribute dont_touch of II1283: signal is true;
	signal II1288: std_logic; attribute dont_touch of II1288: signal is true;
	signal II1289: std_logic; attribute dont_touch of II1289: signal is true;
	signal II1290: std_logic; attribute dont_touch of II1290: signal is true;
	signal II1316: std_logic; attribute dont_touch of II1316: signal is true;
	signal II1321: std_logic; attribute dont_touch of II1321: signal is true;
	signal II1324: std_logic; attribute dont_touch of II1324: signal is true;
	signal II1328: std_logic; attribute dont_touch of II1328: signal is true;
	signal II1329: std_logic; attribute dont_touch of II1329: signal is true;
	signal II1348: std_logic; attribute dont_touch of II1348: signal is true;
	signal II1349: std_logic; attribute dont_touch of II1349: signal is true;
	signal II1350: std_logic; attribute dont_touch of II1350: signal is true;
	signal II1351: std_logic; attribute dont_touch of II1351: signal is true;
	signal II1356: std_logic; attribute dont_touch of II1356: signal is true;
	signal II1357: std_logic; attribute dont_touch of II1357: signal is true;
	signal II1358: std_logic; attribute dont_touch of II1358: signal is true;
	signal II1384: std_logic; attribute dont_touch of II1384: signal is true;
	signal II1389: std_logic; attribute dont_touch of II1389: signal is true;
	signal II1392: std_logic; attribute dont_touch of II1392: signal is true;
	signal II1396: std_logic; attribute dont_touch of II1396: signal is true;
	signal II1397: std_logic; attribute dont_touch of II1397: signal is true;
	signal II1416: std_logic; attribute dont_touch of II1416: signal is true;
	signal II1417: std_logic; attribute dont_touch of II1417: signal is true;
	signal II1418: std_logic; attribute dont_touch of II1418: signal is true;
	signal II1419: std_logic; attribute dont_touch of II1419: signal is true;
	signal II1424: std_logic; attribute dont_touch of II1424: signal is true;
	signal II1425: std_logic; attribute dont_touch of II1425: signal is true;
	signal II1426: std_logic; attribute dont_touch of II1426: signal is true;
	signal II1452: std_logic; attribute dont_touch of II1452: signal is true;
	signal II1457: std_logic; attribute dont_touch of II1457: signal is true;
	signal II1460: std_logic; attribute dont_touch of II1460: signal is true;
	signal II1464: std_logic; attribute dont_touch of II1464: signal is true;
	signal II1465: std_logic; attribute dont_touch of II1465: signal is true;
	signal II1484: std_logic; attribute dont_touch of II1484: signal is true;
	signal II1485: std_logic; attribute dont_touch of II1485: signal is true;
	signal II1486: std_logic; attribute dont_touch of II1486: signal is true;
	signal II1487: std_logic; attribute dont_touch of II1487: signal is true;
	signal II1492: std_logic; attribute dont_touch of II1492: signal is true;
	signal II1493: std_logic; attribute dont_touch of II1493: signal is true;
	signal II1494: std_logic; attribute dont_touch of II1494: signal is true;
	signal II1520: std_logic; attribute dont_touch of II1520: signal is true;
	signal II1525: std_logic; attribute dont_touch of II1525: signal is true;
	signal II1528: std_logic; attribute dont_touch of II1528: signal is true;
	signal II1532: std_logic; attribute dont_touch of II1532: signal is true;
	signal II1533: std_logic; attribute dont_touch of II1533: signal is true;
	signal II1552: std_logic; attribute dont_touch of II1552: signal is true;
	signal II1553: std_logic; attribute dont_touch of II1553: signal is true;
	signal II1554: std_logic; attribute dont_touch of II1554: signal is true;
	signal II1555: std_logic; attribute dont_touch of II1555: signal is true;
	signal II1560: std_logic; attribute dont_touch of II1560: signal is true;
	signal II1561: std_logic; attribute dont_touch of II1561: signal is true;
	signal II1562: std_logic; attribute dont_touch of II1562: signal is true;
	signal II1588: std_logic; attribute dont_touch of II1588: signal is true;
	signal II1593: std_logic; attribute dont_touch of II1593: signal is true;
	signal II1596: std_logic; attribute dont_touch of II1596: signal is true;
	signal II1600: std_logic; attribute dont_touch of II1600: signal is true;
	signal II1601: std_logic; attribute dont_touch of II1601: signal is true;
	signal II1620: std_logic; attribute dont_touch of II1620: signal is true;
	signal II1621: std_logic; attribute dont_touch of II1621: signal is true;
	signal II1622: std_logic; attribute dont_touch of II1622: signal is true;
	signal II1623: std_logic; attribute dont_touch of II1623: signal is true;
	signal II1628: std_logic; attribute dont_touch of II1628: signal is true;
	signal II1629: std_logic; attribute dont_touch of II1629: signal is true;
	signal II1630: std_logic; attribute dont_touch of II1630: signal is true;
	signal II1656: std_logic; attribute dont_touch of II1656: signal is true;
	signal II1661: std_logic; attribute dont_touch of II1661: signal is true;
	signal II1664: std_logic; attribute dont_touch of II1664: signal is true;
	signal II1668: std_logic; attribute dont_touch of II1668: signal is true;
	signal II1669: std_logic; attribute dont_touch of II1669: signal is true;
	signal II1688: std_logic; attribute dont_touch of II1688: signal is true;
	signal II1689: std_logic; attribute dont_touch of II1689: signal is true;
	signal II1690: std_logic; attribute dont_touch of II1690: signal is true;
	signal II1691: std_logic; attribute dont_touch of II1691: signal is true;
	signal II1692: std_logic; attribute dont_touch of II1692: signal is true;
	signal II1694: std_logic; attribute dont_touch of II1694: signal is true;
	signal II1698: std_logic; attribute dont_touch of II1698: signal is true;
	signal II1726: std_logic; attribute dont_touch of II1726: signal is true;
	signal II1729: std_logic; attribute dont_touch of II1729: signal is true;
	signal II1821: std_logic; attribute dont_touch of II1821: signal is true;
	signal II1833: std_logic; attribute dont_touch of II1833: signal is true;
	signal II1841: std_logic; attribute dont_touch of II1841: signal is true;
	signal II1865: std_logic; attribute dont_touch of II1865: signal is true;
	signal II1885: std_logic; attribute dont_touch of II1885: signal is true;
	signal II1901: std_logic; attribute dont_touch of II1901: signal is true;
	signal II1905: std_logic; attribute dont_touch of II1905: signal is true;
	signal II1947: std_logic; attribute dont_touch of II1947: signal is true;
	signal II1948: std_logic; attribute dont_touch of II1948: signal is true;
	signal II1950: std_logic; attribute dont_touch of II1950: signal is true;
	signal II1951: std_logic; attribute dont_touch of II1951: signal is true;
	signal II1952: std_logic; attribute dont_touch of II1952: signal is true;
	signal II1955: std_logic; attribute dont_touch of II1955: signal is true;
	signal II1956: std_logic; attribute dont_touch of II1956: signal is true;
	signal II1963: std_logic; attribute dont_touch of II1963: signal is true;
	signal II1964: std_logic; attribute dont_touch of II1964: signal is true;
	signal II1965: std_logic; attribute dont_touch of II1965: signal is true;
	signal II1966: std_logic; attribute dont_touch of II1966: signal is true;
	signal II1971: std_logic; attribute dont_touch of II1971: signal is true;
	signal II1972: std_logic; attribute dont_touch of II1972: signal is true;
	signal II1973: std_logic; attribute dont_touch of II1973: signal is true;
	signal II1974: std_logic; attribute dont_touch of II1974: signal is true;
	signal II1976: std_logic; attribute dont_touch of II1976: signal is true;
	signal II1978: std_logic; attribute dont_touch of II1978: signal is true;
	signal II1982: std_logic; attribute dont_touch of II1982: signal is true;
	signal II1986: std_logic; attribute dont_touch of II1986: signal is true;
	signal II1990: std_logic; attribute dont_touch of II1990: signal is true;
	signal II1995: std_logic; attribute dont_touch of II1995: signal is true;
	signal II1996: std_logic; attribute dont_touch of II1996: signal is true;
	signal II1997: std_logic; attribute dont_touch of II1997: signal is true;
	signal II2001: std_logic; attribute dont_touch of II2001: signal is true;
	signal II2002: std_logic; attribute dont_touch of II2002: signal is true;
	signal II2008: std_logic; attribute dont_touch of II2008: signal is true;
	signal II2017_1: std_logic; attribute dont_touch of II2017_1: signal is true;
	signal II2017_2: std_logic; attribute dont_touch of II2017_2: signal is true;
	signal II2021_1: std_logic; attribute dont_touch of II2021_1: signal is true;
	signal II2021_2: std_logic; attribute dont_touch of II2021_2: signal is true;
	signal II2025_1: std_logic; attribute dont_touch of II2025_1: signal is true;
	signal II2025_2: std_logic; attribute dont_touch of II2025_2: signal is true;
	signal II2029_1: std_logic; attribute dont_touch of II2029_1: signal is true;
	signal II2032_1: std_logic; attribute dont_touch of II2032_1: signal is true;
	signal II2032_2: std_logic; attribute dont_touch of II2032_2: signal is true;
	signal II2032_3: std_logic; attribute dont_touch of II2032_3: signal is true;
	signal II2037_1: std_logic; attribute dont_touch of II2037_1: signal is true;
	signal II2040_1: std_logic; attribute dont_touch of II2040_1: signal is true;
	signal II2043_1: std_logic; attribute dont_touch of II2043_1: signal is true;
	signal II2043_2: std_logic; attribute dont_touch of II2043_2: signal is true;
	signal II2047_1: std_logic; attribute dont_touch of II2047_1: signal is true;
	signal II2047_2: std_logic; attribute dont_touch of II2047_2: signal is true;
	signal II2051_1: std_logic; attribute dont_touch of II2051_1: signal is true;
	signal II2051_2: std_logic; attribute dont_touch of II2051_2: signal is true;
	signal II2055_1: std_logic; attribute dont_touch of II2055_1: signal is true;
	signal II2055_2: std_logic; attribute dont_touch of II2055_2: signal is true;
	signal II2059_1: std_logic; attribute dont_touch of II2059_1: signal is true;
	signal II2059_2: std_logic; attribute dont_touch of II2059_2: signal is true;
	signal II2063_1: std_logic; attribute dont_touch of II2063_1: signal is true;
	signal II2063_2: std_logic; attribute dont_touch of II2063_2: signal is true;
	signal II2070_1: std_logic; attribute dont_touch of II2070_1: signal is true;
	signal II2070_2: std_logic; attribute dont_touch of II2070_2: signal is true;
	signal P_1: std_logic; attribute dont_touch of P_1: signal is true;
	signal P_2: std_logic; attribute dont_touch of P_2: signal is true;
	signal P_3: std_logic; attribute dont_touch of P_3: signal is true;
	signal P_4: std_logic; attribute dont_touch of P_4: signal is true;
	signal P_5: std_logic; attribute dont_touch of P_5: signal is true;
	signal P_6: std_logic; attribute dont_touch of P_6: signal is true;
	signal P_7: std_logic; attribute dont_touch of P_7: signal is true;
	signal P_8: std_logic; attribute dont_touch of P_8: signal is true;
	signal P_9: std_logic; attribute dont_touch of P_9: signal is true;
	signal P_10: std_logic; attribute dont_touch of P_10: signal is true;
	signal P_11: std_logic; attribute dont_touch of P_11: signal is true;
	signal P_12: std_logic; attribute dont_touch of P_12: signal is true;
	signal P_13: std_logic; attribute dont_touch of P_13: signal is true;
	signal P_14: std_logic; attribute dont_touch of P_14: signal is true;
	signal P_15: std_logic; attribute dont_touch of P_15: signal is true;
	signal P_16: std_logic; attribute dont_touch of P_16: signal is true;
	signal P_17: std_logic; attribute dont_touch of P_17: signal is true;
	signal P_18: std_logic; attribute dont_touch of P_18: signal is true;
	signal P_19: std_logic; attribute dont_touch of P_19: signal is true;
	signal P_20: std_logic; attribute dont_touch of P_20: signal is true;
	signal P_21: std_logic; attribute dont_touch of P_21: signal is true;
	signal P_22: std_logic; attribute dont_touch of P_22: signal is true;
	signal P_23: std_logic; attribute dont_touch of P_23: signal is true;
	signal P_24: std_logic; attribute dont_touch of P_24: signal is true;
	signal P_25: std_logic; attribute dont_touch of P_25: signal is true;
	signal P_26: std_logic; attribute dont_touch of P_26: signal is true;
	signal P_27: std_logic; attribute dont_touch of P_27: signal is true;
	signal P_28: std_logic; attribute dont_touch of P_28: signal is true;
	signal P_29: std_logic; attribute dont_touch of P_29: signal is true;
	signal P_30: std_logic; attribute dont_touch of P_30: signal is true;
	signal P_31: std_logic; attribute dont_touch of P_31: signal is true;
	signal P_32: std_logic; attribute dont_touch of P_32: signal is true;
	signal Y_1: std_logic; attribute dont_touch of Y_1: signal is true;
	signal Y_2: std_logic; attribute dont_touch of Y_2: signal is true;
	signal Y_3: std_logic; attribute dont_touch of Y_3: signal is true;
	signal Y_4: std_logic; attribute dont_touch of Y_4: signal is true;
	signal Y_5: std_logic; attribute dont_touch of Y_5: signal is true;
	signal Y_6: std_logic; attribute dont_touch of Y_6: signal is true;
	signal Y_7: std_logic; attribute dont_touch of Y_7: signal is true;
	signal Y_8: std_logic; attribute dont_touch of Y_8: signal is true;
	signal Y_9: std_logic; attribute dont_touch of Y_9: signal is true;
	signal Y_10: std_logic; attribute dont_touch of Y_10: signal is true;
	signal Y_11: std_logic; attribute dont_touch of Y_11: signal is true;
	signal Y_12: std_logic; attribute dont_touch of Y_12: signal is true;
	signal Y_13: std_logic; attribute dont_touch of Y_13: signal is true;
	signal Y_14: std_logic; attribute dont_touch of Y_14: signal is true;
	signal Y_15: std_logic; attribute dont_touch of Y_15: signal is true;
	signal Y_16: std_logic; attribute dont_touch of Y_16: signal is true;
	signal Y_17: std_logic; attribute dont_touch of Y_17: signal is true;
	signal Y_18: std_logic; attribute dont_touch of Y_18: signal is true;
	signal Y_19: std_logic; attribute dont_touch of Y_19: signal is true;
	signal Y_20: std_logic; attribute dont_touch of Y_20: signal is true;
	signal Y_21: std_logic; attribute dont_touch of Y_21: signal is true;
	signal Y_22: std_logic; attribute dont_touch of Y_22: signal is true;
	signal Y_23: std_logic; attribute dont_touch of Y_23: signal is true;
	signal Y_24: std_logic; attribute dont_touch of Y_24: signal is true;
	signal Y_25: std_logic; attribute dont_touch of Y_25: signal is true;
	signal Y_26: std_logic; attribute dont_touch of Y_26: signal is true;
	signal Y_27: std_logic; attribute dont_touch of Y_27: signal is true;
	signal Y_28: std_logic; attribute dont_touch of Y_28: signal is true;
	signal Y_29: std_logic; attribute dont_touch of Y_29: signal is true;
	signal Y_30: std_logic; attribute dont_touch of Y_30: signal is true;
	signal Y_31: std_logic; attribute dont_touch of Y_31: signal is true;
	signal Y_32: std_logic; attribute dont_touch of Y_32: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			Y_1<=II6;
			Y_2<=II5;
			Y_3<=II4;
			Y_4<=II3;
			Y_5<=II158;
			Y_6<=II157;
			Y_7<=II156;
			Y_8<=II155;
			Y_9<=II310;
			Y_10<=II309;
			Y_11<=II308;
			Y_12<=II307;
			Y_13<=II462;
			Y_14<=II461;
			Y_15<=II460;
			Y_16<=II459;
			Y_17<=II614;
			Y_18<=II613;
			Y_19<=II612;
			Y_20<=II611;
			Y_21<=II766;
			Y_22<=II765;
			Y_23<=II764;
			Y_24<=II763;
			Y_25<=II918;
			Y_26<=II917;
			Y_27<=II916;
			Y_28<=II915;
			Y_29<=II1070;
			Y_30<=II1069;
			Y_31<=II1068;
			Y_32<=II1067;
		end if;
	end process;
	II3<= not II46;
	II4<= not II47;
	II6<= not II104;
	II40<= not X;
	II41<= not Y_4;
	II42<= not Y_3;
	II43<= not Y_2;
	II44<= not Y_1;
	II50<= not II92;
	II155<= not II198;
	II156<= not II199;
	II158<= not II256;
	II192<= not II1_1;
	II193<= not Y_8;
	II194<= not Y_7;
	II195<= not Y_6;
	II196<= not Y_5;
	II202<= not II244;
	II307<= not II350;
	II308<= not II351;
	II310<= not II408;
	II344<= not II1_2;
	II345<= not Y_12;
	II346<= not Y_11;
	II347<= not Y_10;
	II348<= not Y_9;
	II354<= not II396;
	II459<= not II502;
	II460<= not II503;
	II462<= not II560;
	II496<= not II1_3;
	II497<= not Y_16;
	II498<= not Y_15;
	II499<= not Y_14;
	II500<= not Y_13;
	II506<= not II548;
	II611<= not II654;
	II612<= not II655;
	II614<= not II712;
	II648<= not II1_4;
	II649<= not Y_20;
	II650<= not Y_19;
	II651<= not Y_18;
	II652<= not Y_17;
	II658<= not II700;
	II763<= not II806;
	II764<= not II807;
	II766<= not II864;
	II800<= not II1_5;
	II801<= not Y_24;
	II802<= not Y_23;
	II803<= not Y_22;
	II804<= not Y_21;
	II810<= not II852;
	II915<= not II958;
	II916<= not II959;
	II918<= not II1016;
	II952<= not II1_6;
	II953<= not Y_28;
	II954<= not Y_27;
	II955<= not Y_26;
	II956<= not Y_25;
	II962<= not II1004;
	II1067<= not II1110;
	II1068<= not II1111;
	II1070<= not II1168;
	II1104<= not II1_7;
	II1105<= not Y_32;
	II1106<= not Y_31;
	II1107<= not Y_30;
	II1108<= not Y_29;
	II1114<= not II1156;
	II1219_1<= not II1253;
	II1219_2<= not II1316;
	II1219_3<= not II1384;
	II1219_4<= not II1452;
	II1219_5<= not II1520;
	II1219_6<= not II1588;
	II1219_7<= not II1656;
	II1221<= not Y_1;
	II1222<= not Y_2;
	II1223<= not Y_3;
	II1230<= not II1253;
	II1280<= not Y_4;
	II1281<= not Y_5;
	II1282<= not Y_6;
	II1283<= not Y_7;
	II1290<= not II1316;
	II1329<= not II1328;
	II1348<= not Y_8;
	II1349<= not Y_9;
	II1350<= not Y_10;
	II1351<= not Y_11;
	II1358<= not II1384;
	II1397<= not II1396;
	II1416<= not Y_12;
	II1417<= not Y_13;
	II1418<= not Y_14;
	II1419<= not Y_15;
	II1426<= not II1452;
	II1465<= not II1464;
	II1484<= not Y_16;
	II1485<= not Y_17;
	II1486<= not Y_18;
	II1487<= not Y_19;
	II1494<= not II1520;
	II1533<= not II1532;
	II1552<= not Y_20;
	II1553<= not Y_21;
	II1554<= not Y_22;
	II1555<= not Y_23;
	II1562<= not II1588;
	II1601<= not II1600;
	II1620<= not Y_24;
	II1621<= not Y_25;
	II1622<= not Y_26;
	II1623<= not Y_27;
	II1630<= not II1656;
	II1669<= not II1668;
	II1688<= not Y_28;
	II1689<= not Y_29;
	II1690<= not Y_30;
	II1691<= not Y_31;
	II1692<= not Y_32;
	II1947<= not II1948;
	II1951<= not II1952;
	II1955<= not II1956;
	II1963<= not II1964;
	II1965<= not II1966;
	II1971<= not II1972;
	II1973<= not II1974;
	II1996<= not II1995;
	II2002<= not II2001;
	P_1<= not II1226;
	P_3<= not II1228;
	P_4<= not II1229;
	P_7<= not II1288;
	P_8<= not II1289;
	P_11<= not II1356;
	P_12<= not II1357;
	P_15<= not II1424;
	P_16<= not II1425;
	P_19<= not II1492;
	P_20<= not II1493;
	P_23<= not II1560;
	P_24<= not II1561;
	P_27<= not II1628;
	P_28<= not II1629;
	P_30<= not II1694;
	II127_1<=II41 and Y_3 and II109;
	II127_2<=II96 and II113 and Y_4;
	II131_1<=II113 and II92 and Y_3;
	II131_2<=II42 and II109;
	II279_1<=II193 and Y_7 and II261;
	II279_2<=II248 and II265 and Y_8;
	II283_1<=II265 and II244 and Y_7;
	II283_2<=II194 and II261;
	II431_1<=II345 and Y_11 and II413;
	II431_2<=II400 and II417 and Y_12;
	II435_1<=II417 and II396 and Y_11;
	II435_2<=II346 and II413;
	II583_1<=II497 and Y_15 and II565;
	II583_2<=II552 and II569 and Y_16;
	II587_1<=II569 and II548 and Y_15;
	II587_2<=II498 and II565;
	II735_1<=II649 and Y_19 and II717;
	II735_2<=II704 and II721 and Y_20;
	II739_1<=II721 and II700 and Y_19;
	II739_2<=II650 and II717;
	II887_1<=II801 and Y_23 and II869;
	II887_2<=II856 and II873 and Y_24;
	II891_1<=II873 and II852 and Y_23;
	II891_2<=II802 and II869;
	II1039_1<=II953 and Y_27 and II1021;
	II1039_2<=II1008 and II1025 and Y_28;
	II1043_1<=II1025 and II1004 and Y_27;
	II1043_2<=II954 and II1021;
	II1191_1<=II1105 and Y_31 and II1173;
	II1191_2<=II1160 and II1177 and Y_32;
	II1195_1<=II1177 and II1156 and Y_31;
	II1195_2<=II1106 and II1173;
	II2017_1<=P_29 and C_29;
	II2017_2<=P_19 and C_19;
	II2021_1<=P_30 and C_30;
	II2021_2<=P_31 and C_31;
	II2025_1<=P_32 and C_32;
	II2025_2<=P_24 and C_24;
	II2029_1<=P_23 and C_23;
	II2032_1<=P_28 and C_28;
	II2032_2<=P_11 and C_11;
	II2032_3<=P_15 and C_15;
	II2037_1<=P_14 and C_14;
	II2040_1<=P_7 and C_7;
	II2043_1<=P_18 and C_18;
	II2043_2<=P_20 and C_20;
	II2047_1<=P_10 and C_10;
	II2047_2<=P_3 and C_3;
	II2051_1<=P_8 and C_8;
	II2051_2<=P_27 and C_27;
	II2055_1<=P_26 and C_26;
	II2055_2<=P_2 and C_2;
	II2059_1<=X and C_0;
	II2059_2<=P_25 and C_25;
	II2063_1<=P_16 and C_16;
	II2063_2<=P_5 and C_5;
	II2070_1<=P_13 and C_13;
	II2070_2<=P_9 and C_9;
	II5<= not (II135_1 and II135_2);
	II92<= not (Y_2 and Y_1);
	II96<= not (Y_3 and II50);
	II100<= not (Y_1 and II113);
	II104<= not (II44 and II113);
	II157<= not (II287_1 and II287_2);
	II244<= not (Y_6 and Y_5);
	II248<= not (Y_7 and II202);
	II252<= not (Y_5 and II265);
	II256<= not (II196 and II265);
	II309<= not (II439_1 and II439_2);
	II396<= not (Y_10 and Y_9);
	II400<= not (Y_11 and II354);
	II404<= not (Y_9 and II417);
	II408<= not (II348 and II417);
	II461<= not (II591_1 and II591_2);
	II548<= not (Y_14 and Y_13);
	II552<= not (Y_15 and II506);
	II556<= not (Y_13 and II569);
	II560<= not (II500 and II569);
	II613<= not (II743_1 and II743_2);
	II700<= not (Y_18 and Y_17);
	II704<= not (Y_19 and II658);
	II708<= not (Y_17 and II721);
	II712<= not (II652 and II721);
	II765<= not (II895_1 and II895_2);
	II852<= not (Y_22 and Y_21);
	II856<= not (Y_23 and II810);
	II860<= not (Y_21 and II873);
	II864<= not (II804 and II873);
	II917<= not (II1047_1 and II1047_2);
	II1004<= not (Y_26 and Y_25);
	II1008<= not (Y_27 and II962);
	II1012<= not (Y_25 and II1025);
	II1016<= not (II956 and II1025);
	II1069<= not (II1199_1 and II1199_2);
	II1156<= not (Y_30 and Y_29);
	II1160<= not (Y_31 and II1114);
	II1164<= not (Y_29 and II1177);
	II1168<= not (II1108 and II1177);
	II1226<= not (X and Y_1);
	II1228<= not (Y_3 and II1259);
	II1229<= not (Y_4 and II1230);
	II1253<= not (II1223 and II1259);
	II1262<= not (X and II1221);
	II1288<= not (Y_7 and II1321);
	II1289<= not (Y_8 and II1290);
	II1316<= not (II1283 and II1321);
	II1324<= not (II1281 and II1329);
	II1328<= not (II1219_1 and II1280);
	II1356<= not (Y_11 and II1389);
	II1357<= not (Y_12 and II1358);
	II1384<= not (II1351 and II1389);
	II1392<= not (II1349 and II1397);
	II1396<= not (II1219_2 and II1348);
	II1424<= not (Y_15 and II1457);
	II1425<= not (Y_16 and II1426);
	II1452<= not (II1419 and II1457);
	II1460<= not (II1417 and II1465);
	II1464<= not (II1219_3 and II1416);
	II1492<= not (Y_19 and II1525);
	II1493<= not (Y_20 and II1494);
	II1520<= not (II1487 and II1525);
	II1528<= not (II1485 and II1533);
	II1532<= not (II1219_4 and II1484);
	II1560<= not (Y_23 and II1593);
	II1561<= not (Y_24 and II1562);
	II1588<= not (II1555 and II1593);
	II1596<= not (II1553 and II1601);
	II1600<= not (II1219_5 and II1552);
	II1628<= not (Y_27 and II1661);
	II1629<= not (Y_28 and II1630);
	II1656<= not (II1623 and II1661);
	II1664<= not (II1621 and II1669);
	II1668<= not (II1219_6 and II1620);
	II1694<= not (Y_30 and II1726);
	II1698<= not (II1726 and II1690);
	II1729<= not (II1688 and II1219_7);
	II1821<= not (P_1 and C_1);
	II1833<= not (P_4 and C_4);
	II1841<= not (P_6 and C_6);
	II1865<= not (P_12 and C_12);
	II1885<= not (P_17 and C_17);
	II1901<= not (P_21 and C_21);
	II1905<= not (P_22 and C_22);
	II1995<= not (II1986 and II1990 and II1982 and II1885);
	II1997<= not (II1950 and II1833 and II1821 and II1905);
	II2001<= not (II1865 and II1841 and II1978 and II1901);
	Z<= not (II2002 and II2008 and II1996 and II1976);
	II135_1<=II43 or II104;
	II135_2<=Y_2 or II100;
	II287_1<=II195 or II256;
	II287_2<=Y_6 or II252;
	II439_1<=II347 or II408;
	II439_2<=Y_10 or II404;
	II591_1<=II499 or II560;
	II591_2<=Y_14 or II556;
	II743_1<=II651 or II712;
	II743_2<=Y_18 or II708;
	II895_1<=II803 or II864;
	II895_2<=Y_22 or II860;
	II1047_1<=II955 or II1016;
	II1047_2<=Y_26 or II1012;
	II1199_1<=II1107 or II1168;
	II1199_2<=Y_30 or II1164;
	II1_1<= not (II41 or II96);
	II1_2<= not (II193 or II248);
	II1_3<= not (II345 or II400);
	II1_4<= not (II497 or II552);
	II1_5<= not (II649 or II704);
	II1_6<= not (II801 or II856);
	II1_7<= not (II953 or II1008);
	II46<= not (II127_1 or II127_2);
	II47<= not (II131_1 or II131_2);
	II109<= not (II43 or II100);
	II113<= not (CLEAR or II40);
	II198<= not (II279_1 or II279_2);
	II199<= not (II283_1 or II283_2);
	II261<= not (II195 or II252);
	II265<= not (CLEAR or II192);
	II350<= not (II431_1 or II431_2);
	II351<= not (II435_1 or II435_2);
	II413<= not (II347 or II404);
	II417<= not (CLEAR or II344);
	II502<= not (II583_1 or II583_2);
	II503<= not (II587_1 or II587_2);
	II565<= not (II499 or II556);
	II569<= not (CLEAR or II496);
	II654<= not (II735_1 or II735_2);
	II655<= not (II739_1 or II739_2);
	II717<= not (II651 or II708);
	II721<= not (CLEAR or II648);
	II806<= not (II887_1 or II887_2);
	II807<= not (II891_1 or II891_2);
	II869<= not (II803 or II860);
	II873<= not (CLEAR or II800);
	II958<= not (II1039_1 or II1039_2);
	II959<= not (II1043_1 or II1043_2);
	II1021<= not (II955 or II1012);
	II1025<= not (CLEAR or II952);
	II1110<= not (II1191_1 or II1191_2);
	II1111<= not (II1195_1 or II1195_2);
	II1173<= not (II1107 or II1164);
	II1177<= not (CLEAR or II1104);
	II1259<= not (Y_2 or II1262);
	II1321<= not (Y_6 or II1324);
	II1389<= not (Y_10 or II1392);
	II1457<= not (Y_14 or II1460);
	II1525<= not (Y_18 or II1528);
	II1593<= not (Y_22 or II1596);
	II1661<= not (Y_26 or II1664);
	II1726<= not (II1729 or Y_29);
	II1948<= not (II2017_1 or II2017_2);
	II1950<= not (II2021_1 or II2021_2);
	II1952<= not (II2025_1 or II2025_2);
	II1956<= not (II1951 or II2029_1);
	II1964<= not (II2032_1 or II2032_2 or II2032_3);
	II1966<= not (II1955 or II2037_1);
	II1972<= not (II1947 or II2040_1);
	II1974<= not (II2043_1 or II2043_2);
	II1976<= not (II2047_1 or II2047_2 or II1963);
	II1978<= not (II2051_1 or II2051_2 or II1971);
	II1982<= not (II2055_1 or II2055_2 or II1965);
	II1986<= not (II2059_1 or II2059_2);
	II1990<= not (II2063_1 or II2063_2 or II1973);
	II2008<= not (II2070_1 or II2070_2 or II1997);
	P_2<= not (II1222 or II1262);
	P_5<= not (II1281 or II1328);
	P_6<= not (II1282 or II1324);
	P_9<= not (II1349 or II1396);
	P_10<= not (II1350 or II1392);
	P_13<= not (II1417 or II1464);
	P_14<= not (II1418 or II1460);
	P_17<= not (II1485 or II1532);
	P_18<= not (II1486 or II1528);
	P_21<= not (II1553 or II1600);
	P_22<= not (II1554 or II1596);
	P_25<= not (II1621 or II1668);
	P_26<= not (II1622 or II1664);
	P_29<= not (II1689 or II1729);
	P_31<= not (II1691 or II1698);
	P_32<= not (Y_31 or II1698 or II1692);
	W<= not (II1105 or II1160);
end RTL;
