-- File created by Bench2VHDL
-- Name: s38417
-- File: bench/s38417.bench
-- Timestamp: 2019-05-21T22:08:28.326284
--
-- Original File
-- =============
--	# s38417
--	# 28 inputs
--	# 106 outputs
--	# 1636 D-type flipflops
--	# 13470 inverters
--	# 8709 gates (4154 ANDs + 2050 NANDs + 226 ORs + 2279 NORs)
--	
--	INPUT(g51)
--	INPUT(g563)
--	INPUT(g1249)
--	INPUT(g1943)
--	INPUT(g2637)
--	INPUT(g3212)
--	INPUT(g3213)
--	INPUT(g3214)
--	INPUT(g3215)
--	INPUT(g3216)
--	INPUT(g3217)
--	INPUT(g3218)
--	INPUT(g3219)
--	INPUT(g3220)
--	INPUT(g3221)
--	INPUT(g3222)
--	INPUT(g3223)
--	INPUT(g3224)
--	INPUT(g3225)
--	INPUT(g3226)
--	INPUT(g3227)
--	INPUT(g3228)
--	INPUT(g3229)
--	INPUT(g3230)
--	INPUT(g3231)
--	INPUT(g3232)
--	INPUT(g3233)
--	INPUT(g3234)
--	
--	OUTPUT(g3993)
--	OUTPUT(g4088)
--	OUTPUT(g4090)
--	OUTPUT(g4200)
--	OUTPUT(g4321)
--	OUTPUT(g4323)
--	OUTPUT(g4450)
--	OUTPUT(g4590)
--	OUTPUT(g5388)
--	OUTPUT(g5437)
--	OUTPUT(g5472)
--	OUTPUT(g5511)
--	OUTPUT(g5549)
--	OUTPUT(g5555)
--	OUTPUT(g5595)
--	OUTPUT(g5612)
--	OUTPUT(g5629)
--	OUTPUT(g5637)
--	OUTPUT(g5648)
--	OUTPUT(g5657)
--	OUTPUT(g5686)
--	OUTPUT(g5695)
--	OUTPUT(g5738)
--	OUTPUT(g5747)
--	OUTPUT(g5796)
--	OUTPUT(g6225)
--	OUTPUT(g6231)
--	OUTPUT(g6313)
--	OUTPUT(g6368)
--	OUTPUT(g6442)
--	OUTPUT(g6447)
--	OUTPUT(g6485)
--	OUTPUT(g6518)
--	OUTPUT(g6573)
--	OUTPUT(g6642)
--	OUTPUT(g6677)
--	OUTPUT(g6712)
--	OUTPUT(g6750)
--	OUTPUT(g6782)
--	OUTPUT(g6837)
--	OUTPUT(g6895)
--	OUTPUT(g6911)
--	OUTPUT(g6944)
--	OUTPUT(g6979)
--	OUTPUT(g7014)
--	OUTPUT(g7052)
--	OUTPUT(g7084)
--	OUTPUT(g7161)
--	OUTPUT(g7194)
--	OUTPUT(g7229)
--	OUTPUT(g7264)
--	OUTPUT(g7302)
--	OUTPUT(g7334)
--	OUTPUT(g7357)
--	OUTPUT(g7390)
--	OUTPUT(g7425)
--	OUTPUT(g7487)
--	OUTPUT(g7519)
--	OUTPUT(g7909)
--	OUTPUT(g7956)
--	OUTPUT(g7961)
--	OUTPUT(g8007)
--	OUTPUT(g8012)
--	OUTPUT(g8021)
--	OUTPUT(g8023)
--	OUTPUT(g8030)
--	OUTPUT(g8082)
--	OUTPUT(g8087)
--	OUTPUT(g8096)
--	OUTPUT(g8106)
--	OUTPUT(g8167)
--	OUTPUT(g8175)
--	OUTPUT(g8249)
--	OUTPUT(g8251)
--	OUTPUT(g8258)
--	OUTPUT(g8259)
--	OUTPUT(g8260)
--	OUTPUT(g8261)
--	OUTPUT(g8262)
--	OUTPUT(g8263)
--	OUTPUT(g8264)
--	OUTPUT(g8265)
--	OUTPUT(g8266)
--	OUTPUT(g8267)
--	OUTPUT(g8268)
--	OUTPUT(g8269)
--	OUTPUT(g8270)
--	OUTPUT(g8271)
--	OUTPUT(g8272)
--	OUTPUT(g8273)
--	OUTPUT(g8274)
--	OUTPUT(g8275)
--	OUTPUT(g16297)
--	OUTPUT(g16355)
--	OUTPUT(g16399)
--	OUTPUT(g16437)
--	OUTPUT(g16496)
--	OUTPUT(g24734)
--	OUTPUT(g25420)
--	OUTPUT(g25435)
--	OUTPUT(g25442)
--	OUTPUT(g25489)
--	OUTPUT(g26104)
--	OUTPUT(g26135)
--	OUTPUT(g26149)
--	OUTPUT(g27380)
--	
--	g2814 = DFF(g16475)
--	g2817 = DFF(g20571)
--	g2933 = DFF(g20588)
--	g2950 = DFF(g21951)
--	g2883 = DFF(g23315)
--	g2888 = DFF(g24423)
--	g2896 = DFF(g25175)
--	g2892 = DFF(g26019)
--	g2903 = DFF(g26747)
--	g2900 = DFF(g27237)
--	g2908 = DFF(g27715)
--	g2912 = DFF(g24424)
--	g2917 = DFF(g25174)
--	g2924 = DFF(g26020)
--	g2920 = DFF(g26746)
--	g2984 = DFF(g19061)
--	g2985 = DFF(g19060)
--	g2930 = DFF(g19062)
--	g2929 = DFF(g2930)
--	g2879 = DFF(g16494)
--	g2934 = DFF(g16476)
--	g2935 = DFF(g16477)
--	g2938 = DFF(g16478)
--	g2941 = DFF(g16479)
--	g2944 = DFF(g16480)
--	g2947 = DFF(g16481)
--	g2953 = DFF(g16482)
--	g2956 = DFF(g16483)
--	g2959 = DFF(g16484)
--	g2962 = DFF(g16485)
--	g2963 = DFF(g16486)
--	g2966 = DFF(g16487)
--	g2969 = DFF(g16488)
--	g2972 = DFF(g16489)
--	g2975 = DFF(g16490)
--	g2978 = DFF(g16491)
--	g2981 = DFF(g16492)
--	g2874 = DFF(g16493)
--	g1506 = DFF(g20572)
--	g1501 = DFF(g20573)
--	g1496 = DFF(g20574)
--	g1491 = DFF(g20575)
--	g1486 = DFF(g20576)
--	g1481 = DFF(g20577)
--	g1476 = DFF(g20578)
--	g1471 = DFF(g20579)
--	g2877 = DFF(g23313)
--	g2861 = DFF(g21960)
--	g813 = DFF(g2861)
--	g2864 = DFF(g21961)
--	g809 = DFF(g2864)
--	g2867 = DFF(g21962)
--	g805 = DFF(g2867)
--	g2870 = DFF(g21963)
--	g801 = DFF(g2870)
--	g2818 = DFF(g21947)
--	g797 = DFF(g2818)
--	g2821 = DFF(g21948)
--	g793 = DFF(g2821)
--	g2824 = DFF(g21949)
--	g789 = DFF(g2824)
--	g2827 = DFF(g21950)
--	g785 = DFF(g2827)
--	g2830 = DFF(g23312)
--	g2873 = DFF(g2830)
--	g2833 = DFF(g21952)
--	g125 = DFF(g2833)
--	g2836 = DFF(g21953)
--	g121 = DFF(g2836)
--	g2839 = DFF(g21954)
--	g117 = DFF(g2839)
--	g2842 = DFF(g21955)
--	g113 = DFF(g2842)
--	g2845 = DFF(g21956)
--	g109 = DFF(g2845)
--	g2848 = DFF(g21957)
--	g105 = DFF(g2848)
--	g2851 = DFF(g21958)
--	g101 = DFF(g2851)
--	g2854 = DFF(g21959)
--	g97 = DFF(g2854)
--	g2858 = DFF(g23316)
--	g2857 = DFF(g2858)
--	g2200 = DFF(g20587)
--	g2195 = DFF(g20585)
--	g2190 = DFF(g20586)
--	g2185 = DFF(g20584)
--	g2180 = DFF(g20583)
--	g2175 = DFF(g20582)
--	g2170 = DFF(g20581)
--	g2165 = DFF(g20580)
--	g2878 = DFF(g23314)
--	g3129 = DFF(g13475)
--	g3117 = DFF(g3129)
--	g3109 = DFF(g3117)
--	g3210 = DFF(g20630)
--	g3211 = DFF(g20631)
--	g3084 = DFF(g20632)
--	g3085 = DFF(g20609)
--	g3086 = DFF(g20610)
--	g3087 = DFF(g20611)
--	g3091 = DFF(g20612)
--	g3092 = DFF(g20613)
--	g3093 = DFF(g20614)
--	g3094 = DFF(g20615)
--	g3095 = DFF(g20616)
--	g3096 = DFF(g20617)
--	g3097 = DFF(g26751)
--	g3098 = DFF(g26752)
--	g3099 = DFF(g26753)
--	g3100 = DFF(g29163)
--	g3101 = DFF(g29164)
--	g3102 = DFF(g29165)
--	g3103 = DFF(g30120)
--	g3104 = DFF(g30121)
--	g3105 = DFF(g30122)
--	g3106 = DFF(g30941)
--	g3107 = DFF(g30942)
--	g3108 = DFF(g30943)
--	g3155 = DFF(g20618)
--	g3158 = DFF(g20619)
--	g3161 = DFF(g20620)
--	g3164 = DFF(g20621)
--	g3167 = DFF(g20622)
--	g3170 = DFF(g20623)
--	g3173 = DFF(g20624)
--	g3176 = DFF(g20625)
--	g3179 = DFF(g20626)
--	g3182 = DFF(g20627)
--	g3185 = DFF(g20628)
--	g3088 = DFF(g20629)
--	g3191 = DFF(g27717)
--	g3194 = DFF(g28316)
--	g3197 = DFF(g28317)
--	g3198 = DFF(g28318)
--	g3201 = DFF(g28704)
--	g3204 = DFF(g28705)
--	g3207 = DFF(g28706)
--	g3188 = DFF(g29463)
--	g3133 = DFF(g29656)
--	g3132 = DFF(g28698)
--	g3128 = DFF(g29166)
--	g3127 = DFF(g28697)
--	g3126 = DFF(g28315)
--	g3125 = DFF(g28696)
--	g3124 = DFF(g28314)
--	g3123 = DFF(g28313)
--	g3120 = DFF(g28695)
--	g3114 = DFF(g28694)
--	g3113 = DFF(g28693)
--	g3112 = DFF(g28312)
--	g3110 = DFF(g28311)
--	g3111 = DFF(g28310)
--	g3139 = DFF(g29461)
--	g3136 = DFF(g28701)
--	g3134 = DFF(g28700)
--	g3135 = DFF(g28699)
--	g3151 = DFF(g29462)
--	g3142 = DFF(g28703)
--	g3147 = DFF(g28702)
--	g185 = DFF(g29657)
--	g138 = DFF(g13405)
--	g135 = DFF(g138)
--	g165 = DFF(g135)
--	g130 = DFF(g24259)
--	g131 = DFF(g24260)
--	g129 = DFF(g24261)
--	g133 = DFF(g24262)
--	g134 = DFF(g24263)
--	g132 = DFF(g24264)
--	g142 = DFF(g24265)
--	g143 = DFF(g24266)
--	g141 = DFF(g24267)
--	g145 = DFF(g24268)
--	g146 = DFF(g24269)
--	g144 = DFF(g24270)
--	g148 = DFF(g24271)
--	g149 = DFF(g24272)
--	g147 = DFF(g24273)
--	g151 = DFF(g24274)
--	g152 = DFF(g24275)
--	g150 = DFF(g24276)
--	g154 = DFF(g24277)
--	g155 = DFF(g24278)
--	g153 = DFF(g24279)
--	g157 = DFF(g24280)
--	g158 = DFF(g24281)
--	g156 = DFF(g24282)
--	g160 = DFF(g24283)
--	g161 = DFF(g24284)
--	g159 = DFF(g24285)
--	g163 = DFF(g24286)
--	g164 = DFF(g24287)
--	g162 = DFF(g24288)
--	g169 = DFF(g26679)
--	g170 = DFF(g26680)
--	g168 = DFF(g26681)
--	g172 = DFF(g26682)
--	g173 = DFF(g26683)
--	g171 = DFF(g26684)
--	g175 = DFF(g26685)
--	g176 = DFF(g26686)
--	g174 = DFF(g26687)
--	g178 = DFF(g26688)
--	g179 = DFF(g26689)
--	g177 = DFF(g26690)
--	g186 = DFF(g30506)
--	g189 = DFF(g30507)
--	g192 = DFF(g30508)
--	g231 = DFF(g30842)
--	g234 = DFF(g30843)
--	g237 = DFF(g30844)
--	g195 = DFF(g30836)
--	g198 = DFF(g30837)
--	g201 = DFF(g30838)
--	g240 = DFF(g30845)
--	g243 = DFF(g30846)
--	g246 = DFF(g30847)
--	g204 = DFF(g30509)
--	g207 = DFF(g30510)
--	g210 = DFF(g30511)
--	g249 = DFF(g30515)
--	g252 = DFF(g30516)
--	g255 = DFF(g30517)
--	g213 = DFF(g30512)
--	g216 = DFF(g30513)
--	g219 = DFF(g30514)
--	g258 = DFF(g30518)
--	g261 = DFF(g30519)
--	g264 = DFF(g30520)
--	g222 = DFF(g30839)
--	g225 = DFF(g30840)
--	g228 = DFF(g30841)
--	g267 = DFF(g30848)
--	g270 = DFF(g30849)
--	g273 = DFF(g30850)
--	g92 = DFF(g25983)
--	g88 = DFF(g26678)
--	g83 = DFF(g27189)
--	g79 = DFF(g27683)
--	g74 = DFF(g28206)
--	g70 = DFF(g28673)
--	g65 = DFF(g29131)
--	g61 = DFF(g29413)
--	g56 = DFF(g29627)
--	g52 = DFF(g29794)
--	g180 = DFF(g20555)
--	g182 = DFF(g180)
--	g181 = DFF(g182)
--	g276 = DFF(g13406)
--	g405 = DFF(g276)
--	g401 = DFF(g405)
--	g309 = DFF(g11496)
--	g354 = DFF(g28207)
--	g343 = DFF(g28208)
--	g346 = DFF(g28209)
--	g369 = DFF(g28210)
--	g358 = DFF(g28211)
--	g361 = DFF(g28212)
--	g384 = DFF(g28213)
--	g373 = DFF(g28214)
--	g376 = DFF(g28215)
--	g398 = DFF(g28216)
--	g388 = DFF(g28217)
--	g391 = DFF(g28218)
--	g408 = DFF(g29414)
--	g411 = DFF(g29415)
--	g414 = DFF(g29416)
--	g417 = DFF(g29631)
--	g420 = DFF(g29632)
--	g423 = DFF(g29633)
--	g427 = DFF(g29417)
--	g428 = DFF(g29418)
--	g426 = DFF(g29419)
--	g429 = DFF(g27684)
--	g432 = DFF(g27685)
--	g435 = DFF(g27686)
--	g438 = DFF(g27687)
--	g441 = DFF(g27688)
--	g444 = DFF(g27689)
--	g448 = DFF(g28674)
--	g449 = DFF(g28675)
--	g447 = DFF(g28676)
--	g312 = DFF(g29795)
--	g313 = DFF(g29796)
--	g314 = DFF(g29797)
--	g315 = DFF(g30851)
--	g316 = DFF(g30852)
--	g317 = DFF(g30853)
--	g318 = DFF(g30710)
--	g319 = DFF(g30711)
--	g320 = DFF(g30712)
--	g322 = DFF(g29628)
--	g323 = DFF(g29629)
--	g321 = DFF(g29630)
--	g403 = DFF(g27191)
--	g404 = DFF(g27192)
--	g402 = DFF(g27193)
--	g450 = DFF(g11509)
--	g451 = DFF(g450)
--	g452 = DFF(g11510)
--	g453 = DFF(g452)
--	g454 = DFF(g11511)
--	g279 = DFF(g454)
--	g280 = DFF(g11491)
--	g281 = DFF(g280)
--	g282 = DFF(g11492)
--	g283 = DFF(g282)
--	g284 = DFF(g11493)
--	g285 = DFF(g284)
--	g286 = DFF(g11494)
--	g287 = DFF(g286)
--	g288 = DFF(g11495)
--	g289 = DFF(g288)
--	g290 = DFF(g13407)
--	g291 = DFF(g290)
--	g299 = DFF(g19012)
--	g305 = DFF(g23148)
--	g308 = DFF(g23149)
--	g297 = DFF(g23150)
--	g296 = DFF(g23151)
--	g295 = DFF(g23152)
--	g294 = DFF(g23153)
--	g304 = DFF(g19016)
--	g303 = DFF(g19015)
--	g302 = DFF(g19014)
--	g301 = DFF(g19013)
--	g300 = DFF(g25130)
--	g298 = DFF(g27190)
--	g342 = DFF(g11497)
--	g349 = DFF(g342)
--	g350 = DFF(g11498)
--	g351 = DFF(g350)
--	g352 = DFF(g11499)
--	g353 = DFF(g352)
--	g357 = DFF(g11500)
--	g364 = DFF(g357)
--	g365 = DFF(g11501)
--	g366 = DFF(g365)
--	g367 = DFF(g11502)
--	g368 = DFF(g367)
--	g372 = DFF(g11503)
--	g379 = DFF(g372)
--	g380 = DFF(g11504)
--	g381 = DFF(g380)
--	g382 = DFF(g11505)
--	g383 = DFF(g382)
--	g387 = DFF(g11506)
--	g394 = DFF(g387)
--	g395 = DFF(g11507)
--	g396 = DFF(g395)
--	g397 = DFF(g11508)
--	g324 = DFF(g397)
--	g325 = DFF(g13408)
--	g331 = DFF(g325)
--	g337 = DFF(g331)
--	g545 = DFF(g13419)
--	g551 = DFF(g545)
--	g550 = DFF(g551)
--	g554 = DFF(g23160)
--	g557 = DFF(g20556)
--	g510 = DFF(g20557)
--	g513 = DFF(g16467)
--	g523 = DFF(g513)
--	g524 = DFF(g523)
--	g564 = DFF(g11512)
--	g569 = DFF(g564)
--	g570 = DFF(g11515)
--	g571 = DFF(g570)
--	g572 = DFF(g11516)
--	g573 = DFF(g572)
--	g574 = DFF(g11517)
--	g565 = DFF(g574)
--	g566 = DFF(g11513)
--	g567 = DFF(g566)
--	g568 = DFF(g11514)
--	g489 = DFF(g568)
--	g474 = DFF(g13409)
--	g481 = DFF(g474)
--	g485 = DFF(g481)
--	g486 = DFF(g24292)
--	g487 = DFF(g24293)
--	g488 = DFF(g24294)
--	g455 = DFF(g25139)
--	g458 = DFF(g25131)
--	g461 = DFF(g25132)
--	g477 = DFF(g25136)
--	g478 = DFF(g25137)
--	g479 = DFF(g25138)
--	g480 = DFF(g24289)
--	g484 = DFF(g24290)
--	g464 = DFF(g24291)
--	g465 = DFF(g25133)
--	g468 = DFF(g25134)
--	g471 = DFF(g25135)
--	g528 = DFF(g16468)
--	g535 = DFF(g528)
--	g542 = DFF(g535)
--	g543 = DFF(g19021)
--	g544 = DFF(g543)
--	g548 = DFF(g23159)
--	g549 = DFF(g19022)
--	g499 = DFF(g549)
--	g558 = DFF(g19023)
--	g559 = DFF(g558)
--	g576 = DFF(g28219)
--	g577 = DFF(g28220)
--	g575 = DFF(g28221)
--	g579 = DFF(g28222)
--	g580 = DFF(g28223)
--	g578 = DFF(g28224)
--	g582 = DFF(g28225)
--	g583 = DFF(g28226)
--	g581 = DFF(g28227)
--	g585 = DFF(g28228)
--	g586 = DFF(g28229)
--	g584 = DFF(g28230)
--	g587 = DFF(g25985)
--	g590 = DFF(g25986)
--	g593 = DFF(g25987)
--	g596 = DFF(g25988)
--	g599 = DFF(g25989)
--	g602 = DFF(g25990)
--	g614 = DFF(g29135)
--	g617 = DFF(g29136)
--	g620 = DFF(g29137)
--	g605 = DFF(g29132)
--	g608 = DFF(g29133)
--	g611 = DFF(g29134)
--	g490 = DFF(g27194)
--	g493 = DFF(g27195)
--	g496 = DFF(g27196)
--	g506 = DFF(g8284)
--	g507 = DFF(g24295)
--	g508 = DFF(g19017)
--	g509 = DFF(g19018)
--	g514 = DFF(g19019)
--	g515 = DFF(g19020)
--	g516 = DFF(g23158)
--	g517 = DFF(g23157)
--	g518 = DFF(g23156)
--	g519 = DFF(g23155)
--	g520 = DFF(g23154)
--	g525 = DFF(g520)
--	g529 = DFF(g13410)
--	g530 = DFF(g13411)
--	g531 = DFF(g13412)
--	g532 = DFF(g13413)
--	g533 = DFF(g13414)
--	g534 = DFF(g13415)
--	g536 = DFF(g13416)
--	g537 = DFF(g13417)
--	g538 = DFF(g25984)
--	g541 = DFF(g13418)
--	g623 = DFF(g13420)
--	g626 = DFF(g623)
--	g629 = DFF(g626)
--	g630 = DFF(g20558)
--	g659 = DFF(g21943)
--	g640 = DFF(g23161)
--	g633 = DFF(g24296)
--	g653 = DFF(g25140)
--	g646 = DFF(g25991)
--	g660 = DFF(g26691)
--	g672 = DFF(g27197)
--	g666 = DFF(g27690)
--	g679 = DFF(g28231)
--	g686 = DFF(g28677)
--	g692 = DFF(g29138)
--	g699 = DFF(g23162)
--	g700 = DFF(g23163)
--	g698 = DFF(g23164)
--	g702 = DFF(g23165)
--	g703 = DFF(g23166)
--	g701 = DFF(g23167)
--	g705 = DFF(g23168)
--	g706 = DFF(g23169)
--	g704 = DFF(g23170)
--	g708 = DFF(g23171)
--	g709 = DFF(g23172)
--	g707 = DFF(g23173)
--	g711 = DFF(g23174)
--	g712 = DFF(g23175)
--	g710 = DFF(g23176)
--	g714 = DFF(g23177)
--	g715 = DFF(g23178)
--	g713 = DFF(g23179)
--	g717 = DFF(g23180)
--	g718 = DFF(g23181)
--	g716 = DFF(g23182)
--	g720 = DFF(g23183)
--	g721 = DFF(g23184)
--	g719 = DFF(g23185)
--	g723 = DFF(g23186)
--	g724 = DFF(g23187)
--	g722 = DFF(g23188)
--	g726 = DFF(g23189)
--	g727 = DFF(g23190)
--	g725 = DFF(g23191)
--	g729 = DFF(g23192)
--	g730 = DFF(g23193)
--	g728 = DFF(g23194)
--	g732 = DFF(g23195)
--	g733 = DFF(g23196)
--	g731 = DFF(g23197)
--	g735 = DFF(g26692)
--	g736 = DFF(g26693)
--	g734 = DFF(g26694)
--	g738 = DFF(g24297)
--	g739 = DFF(g24298)
--	g737 = DFF(g24299)
--	g826 = DFF(g13421)
--	g823 = DFF(g826)
--	g853 = DFF(g823)
--	g818 = DFF(g24300)
--	g819 = DFF(g24301)
--	g817 = DFF(g24302)
--	g821 = DFF(g24303)
--	g822 = DFF(g24304)
--	g820 = DFF(g24305)
--	g830 = DFF(g24306)
--	g831 = DFF(g24307)
--	g829 = DFF(g24308)
--	g833 = DFF(g24309)
--	g834 = DFF(g24310)
--	g832 = DFF(g24311)
--	g836 = DFF(g24312)
--	g837 = DFF(g24313)
--	g835 = DFF(g24314)
--	g839 = DFF(g24315)
--	g840 = DFF(g24316)
--	g838 = DFF(g24317)
--	g842 = DFF(g24318)
--	g843 = DFF(g24319)
--	g841 = DFF(g24320)
--	g845 = DFF(g24321)
--	g846 = DFF(g24322)
--	g844 = DFF(g24323)
--	g848 = DFF(g24324)
--	g849 = DFF(g24325)
--	g847 = DFF(g24326)
--	g851 = DFF(g24327)
--	g852 = DFF(g24328)
--	g850 = DFF(g24329)
--	g857 = DFF(g26696)
--	g858 = DFF(g26697)
--	g856 = DFF(g26698)
--	g860 = DFF(g26699)
--	g861 = DFF(g26700)
--	g859 = DFF(g26701)
--	g863 = DFF(g26702)
--	g864 = DFF(g26703)
--	g862 = DFF(g26704)
--	g866 = DFF(g26705)
--	g867 = DFF(g26706)
--	g865 = DFF(g26707)
--	g873 = DFF(g30521)
--	g876 = DFF(g30522)
--	g879 = DFF(g30523)
--	g918 = DFF(g30860)
--	g921 = DFF(g30861)
--	g924 = DFF(g30862)
--	g882 = DFF(g30854)
--	g885 = DFF(g30855)
--	g888 = DFF(g30856)
--	g927 = DFF(g30863)
--	g930 = DFF(g30864)
--	g933 = DFF(g30865)
--	g891 = DFF(g30524)
--	g894 = DFF(g30525)
--	g897 = DFF(g30526)
--	g936 = DFF(g30530)
--	g939 = DFF(g30531)
--	g942 = DFF(g30532)
--	g900 = DFF(g30527)
--	g903 = DFF(g30528)
--	g906 = DFF(g30529)
--	g945 = DFF(g30533)
--	g948 = DFF(g30534)
--	g951 = DFF(g30535)
--	g909 = DFF(g30857)
--	g912 = DFF(g30858)
--	g915 = DFF(g30859)
--	g954 = DFF(g30866)
--	g957 = DFF(g30867)
--	g960 = DFF(g30868)
--	g780 = DFF(g25992)
--	g776 = DFF(g26695)
--	g771 = DFF(g27198)
--	g767 = DFF(g27691)
--	g762 = DFF(g28232)
--	g758 = DFF(g28678)
--	g753 = DFF(g29139)
--	g749 = DFF(g29420)
--	g744 = DFF(g29634)
--	g740 = DFF(g29798)
--	g868 = DFF(g20559)
--	g870 = DFF(g868)
--	g869 = DFF(g870)
--	g963 = DFF(g13422)
--	g1092 = DFF(g963)
--	g1088 = DFF(g1092)
--	g996 = DFF(g11523)
--	g1041 = DFF(g28233)
--	g1030 = DFF(g28234)
--	g1033 = DFF(g28235)
--	g1056 = DFF(g28236)
--	g1045 = DFF(g28237)
--	g1048 = DFF(g28238)
--	g1071 = DFF(g28239)
--	g1060 = DFF(g28240)
--	g1063 = DFF(g28241)
--	g1085 = DFF(g28242)
--	g1075 = DFF(g28243)
--	g1078 = DFF(g28244)
--	g1095 = DFF(g29421)
--	g1098 = DFF(g29422)
--	g1101 = DFF(g29423)
--	g1104 = DFF(g29638)
--	g1107 = DFF(g29639)
--	g1110 = DFF(g29640)
--	g1114 = DFF(g29424)
--	g1115 = DFF(g29425)
--	g1113 = DFF(g29426)
--	g1116 = DFF(g27692)
--	g1119 = DFF(g27693)
--	g1122 = DFF(g27694)
--	g1125 = DFF(g27695)
--	g1128 = DFF(g27696)
--	g1131 = DFF(g27697)
--	g1135 = DFF(g28679)
--	g1136 = DFF(g28680)
--	g1134 = DFF(g28681)
--	g999 = DFF(g29799)
--	g1000 = DFF(g29800)
--	g1001 = DFF(g29801)
--	g1002 = DFF(g30869)
--	g1003 = DFF(g30870)
--	g1004 = DFF(g30871)
--	g1005 = DFF(g30713)
--	g1006 = DFF(g30714)
--	g1007 = DFF(g30715)
--	g1009 = DFF(g29635)
--	g1010 = DFF(g29636)
--	g1008 = DFF(g29637)
--	g1090 = DFF(g27206)
--	g1091 = DFF(g27207)
--	g1089 = DFF(g27208)
--	g1137 = DFF(g11536)
--	g1138 = DFF(g1137)
--	g1139 = DFF(g11537)
--	g1140 = DFF(g1139)
--	g1141 = DFF(g11538)
--	g966 = DFF(g1141)
--	g967 = DFF(g11518)
--	g968 = DFF(g967)
--	g969 = DFF(g11519)
--	g970 = DFF(g969)
--	g971 = DFF(g11520)
--	g972 = DFF(g971)
--	g973 = DFF(g11521)
--	g974 = DFF(g973)
--	g975 = DFF(g11522)
--	g976 = DFF(g975)
--	g977 = DFF(g13423)
--	g978 = DFF(g977)
--	g986 = DFF(g19024)
--	g992 = DFF(g27200)
--	g995 = DFF(g27201)
--	g984 = DFF(g27202)
--	g983 = DFF(g27203)
--	g982 = DFF(g27204)
--	g981 = DFF(g27205)
--	g991 = DFF(g19028)
--	g990 = DFF(g19027)
--	g989 = DFF(g19026)
--	g988 = DFF(g19025)
--	g987 = DFF(g25141)
--	g985 = DFF(g27199)
--	g1029 = DFF(g11524)
--	g1036 = DFF(g1029)
--	g1037 = DFF(g11525)
--	g1038 = DFF(g1037)
--	g1039 = DFF(g11526)
--	g1040 = DFF(g1039)
--	g1044 = DFF(g11527)
--	g1051 = DFF(g1044)
--	g1052 = DFF(g11528)
--	g1053 = DFF(g1052)
--	g1054 = DFF(g11529)
--	g1055 = DFF(g1054)
--	g1059 = DFF(g11530)
--	g1066 = DFF(g1059)
--	g1067 = DFF(g11531)
--	g1068 = DFF(g1067)
--	g1069 = DFF(g11532)
--	g1070 = DFF(g1069)
--	g1074 = DFF(g11533)
--	g1081 = DFF(g1074)
--	g1082 = DFF(g11534)
--	g1083 = DFF(g1082)
--	g1084 = DFF(g11535)
--	g1011 = DFF(g1084)
--	g1012 = DFF(g13424)
--	g1018 = DFF(g1012)
--	g1024 = DFF(g1018)
--	g1231 = DFF(g13435)
--	g1237 = DFF(g1231)
--	g1236 = DFF(g1237)
--	g1240 = DFF(g23198)
--	g1243 = DFF(g20560)
--	g1196 = DFF(g20561)
--	g1199 = DFF(g16469)
--	g1209 = DFF(g1199)
--	g1210 = DFF(g1209)
--	g1250 = DFF(g11539)
--	g1255 = DFF(g1250)
--	g1256 = DFF(g11542)
--	g1257 = DFF(g1256)
--	g1258 = DFF(g11543)
--	g1259 = DFF(g1258)
--	g1260 = DFF(g11544)
--	g1251 = DFF(g1260)
--	g1252 = DFF(g11540)
--	g1253 = DFF(g1252)
--	g1254 = DFF(g11541)
--	g1176 = DFF(g1254)
--	g1161 = DFF(g13425)
--	g1168 = DFF(g1161)
--	g1172 = DFF(g1168)
--	g1173 = DFF(g24333)
--	g1174 = DFF(g24334)
--	g1175 = DFF(g24335)
--	g1142 = DFF(g25150)
--	g1145 = DFF(g25142)
--	g1148 = DFF(g25143)
--	g1164 = DFF(g25147)
--	g1165 = DFF(g25148)
--	g1166 = DFF(g25149)
--	g1167 = DFF(g24330)
--	g1171 = DFF(g24331)
--	g1151 = DFF(g24332)
--	g1152 = DFF(g25144)
--	g1155 = DFF(g25145)
--	g1158 = DFF(g25146)
--	g1214 = DFF(g16470)
--	g1221 = DFF(g1214)
--	g1228 = DFF(g1221)
--	g1229 = DFF(g19033)
--	g1230 = DFF(g1229)
--	g1234 = DFF(g27217)
--	g1235 = DFF(g19034)
--	g1186 = DFF(g1235)
--	g1244 = DFF(g19035)
--	g1245 = DFF(g1244)
--	g1262 = DFF(g28245)
--	g1263 = DFF(g28246)
--	g1261 = DFF(g28247)
--	g1265 = DFF(g28248)
--	g1266 = DFF(g28249)
--	g1264 = DFF(g28250)
--	g1268 = DFF(g28251)
--	g1269 = DFF(g28252)
--	g1267 = DFF(g28253)
--	g1271 = DFF(g28254)
--	g1272 = DFF(g28255)
--	g1270 = DFF(g28256)
--	g1273 = DFF(g25994)
--	g1276 = DFF(g25995)
--	g1279 = DFF(g25996)
--	g1282 = DFF(g25997)
--	g1285 = DFF(g25998)
--	g1288 = DFF(g25999)
--	g1300 = DFF(g29143)
--	g1303 = DFF(g29144)
--	g1306 = DFF(g29145)
--	g1291 = DFF(g29140)
--	g1294 = DFF(g29141)
--	g1297 = DFF(g29142)
--	g1177 = DFF(g27209)
--	g1180 = DFF(g27210)
--	g1183 = DFF(g27211)
--	g1192 = DFF(g8293)
--	g1193 = DFF(g24336)
--	g1194 = DFF(g19029)
--	g1195 = DFF(g19030)
--	g1200 = DFF(g19031)
--	g1201 = DFF(g19032)
--	g1202 = DFF(g27216)
--	g1203 = DFF(g27215)
--	g1204 = DFF(g27214)
--	g1205 = DFF(g27213)
--	g1206 = DFF(g27212)
--	g1211 = DFF(g1206)
--	g1215 = DFF(g13426)
--	g1216 = DFF(g13427)
--	g1217 = DFF(g13428)
--	g1218 = DFF(g13429)
--	g1219 = DFF(g13430)
--	g1220 = DFF(g13431)
--	g1222 = DFF(g13432)
--	g1223 = DFF(g13433)
--	g1224 = DFF(g25993)
--	g1227 = DFF(g13434)
--	g1309 = DFF(g13436)
--	g1312 = DFF(g1309)
--	g1315 = DFF(g1312)
--	g1316 = DFF(g20562)
--	g1345 = DFF(g21944)
--	g1326 = DFF(g23199)
--	g1319 = DFF(g24337)
--	g1339 = DFF(g25151)
--	g1332 = DFF(g26000)
--	g1346 = DFF(g26708)
--	g1358 = DFF(g27218)
--	g1352 = DFF(g27698)
--	g1365 = DFF(g28257)
--	g1372 = DFF(g28682)
--	g1378 = DFF(g29146)
--	g1385 = DFF(g23200)
--	g1386 = DFF(g23201)
--	g1384 = DFF(g23202)
--	g1388 = DFF(g23203)
--	g1389 = DFF(g23204)
--	g1387 = DFF(g23205)
--	g1391 = DFF(g23206)
--	g1392 = DFF(g23207)
--	g1390 = DFF(g23208)
--	g1394 = DFF(g23209)
--	g1395 = DFF(g23210)
--	g1393 = DFF(g23211)
--	g1397 = DFF(g23212)
--	g1398 = DFF(g23213)
--	g1396 = DFF(g23214)
--	g1400 = DFF(g23215)
--	g1401 = DFF(g23216)
--	g1399 = DFF(g23217)
--	g1403 = DFF(g23218)
--	g1404 = DFF(g23219)
--	g1402 = DFF(g23220)
--	g1406 = DFF(g23221)
--	g1407 = DFF(g23222)
--	g1405 = DFF(g23223)
--	g1409 = DFF(g23224)
--	g1410 = DFF(g23225)
--	g1408 = DFF(g23226)
--	g1412 = DFF(g23227)
--	g1413 = DFF(g23228)
--	g1411 = DFF(g23229)
--	g1415 = DFF(g23230)
--	g1416 = DFF(g23231)
--	g1414 = DFF(g23232)
--	g1418 = DFF(g23233)
--	g1419 = DFF(g23234)
--	g1417 = DFF(g23235)
--	g1421 = DFF(g26709)
--	g1422 = DFF(g26710)
--	g1420 = DFF(g26711)
--	g1424 = DFF(g24338)
--	g1425 = DFF(g24339)
--	g1423 = DFF(g24340)
--	g1520 = DFF(g13437)
--	g1517 = DFF(g1520)
--	g1547 = DFF(g1517)
--	g1512 = DFF(g24341)
--	g1513 = DFF(g24342)
--	g1511 = DFF(g24343)
--	g1515 = DFF(g24344)
--	g1516 = DFF(g24345)
--	g1514 = DFF(g24346)
--	g1524 = DFF(g24347)
--	g1525 = DFF(g24348)
--	g1523 = DFF(g24349)
--	g1527 = DFF(g24350)
--	g1528 = DFF(g24351)
--	g1526 = DFF(g24352)
--	g1530 = DFF(g24353)
--	g1531 = DFF(g24354)
--	g1529 = DFF(g24355)
--	g1533 = DFF(g24356)
--	g1534 = DFF(g24357)
--	g1532 = DFF(g24358)
--	g1536 = DFF(g24359)
--	g1537 = DFF(g24360)
--	g1535 = DFF(g24361)
--	g1539 = DFF(g24362)
--	g1540 = DFF(g24363)
--	g1538 = DFF(g24364)
--	g1542 = DFF(g24365)
--	g1543 = DFF(g24366)
--	g1541 = DFF(g24367)
--	g1545 = DFF(g24368)
--	g1546 = DFF(g24369)
--	g1544 = DFF(g24370)
--	g1551 = DFF(g26713)
--	g1552 = DFF(g26714)
--	g1550 = DFF(g26715)
--	g1554 = DFF(g26716)
--	g1555 = DFF(g26717)
--	g1553 = DFF(g26718)
--	g1557 = DFF(g26719)
--	g1558 = DFF(g26720)
--	g1556 = DFF(g26721)
--	g1560 = DFF(g26722)
--	g1561 = DFF(g26723)
--	g1559 = DFF(g26724)
--	g1567 = DFF(g30536)
--	g1570 = DFF(g30537)
--	g1573 = DFF(g30538)
--	g1612 = DFF(g30878)
--	g1615 = DFF(g30879)
--	g1618 = DFF(g30880)
--	g1576 = DFF(g30872)
--	g1579 = DFF(g30873)
--	g1582 = DFF(g30874)
--	g1621 = DFF(g30881)
--	g1624 = DFF(g30882)
--	g1627 = DFF(g30883)
--	g1585 = DFF(g30539)
--	g1588 = DFF(g30540)
--	g1591 = DFF(g30541)
--	g1630 = DFF(g30545)
--	g1633 = DFF(g30546)
--	g1636 = DFF(g30547)
--	g1594 = DFF(g30542)
--	g1597 = DFF(g30543)
--	g1600 = DFF(g30544)
--	g1639 = DFF(g30548)
--	g1642 = DFF(g30549)
--	g1645 = DFF(g30550)
--	g1603 = DFF(g30875)
--	g1606 = DFF(g30876)
--	g1609 = DFF(g30877)
--	g1648 = DFF(g30884)
--	g1651 = DFF(g30885)
--	g1654 = DFF(g30886)
--	g1466 = DFF(g26001)
--	g1462 = DFF(g26712)
--	g1457 = DFF(g27219)
--	g1453 = DFF(g27699)
--	g1448 = DFF(g28258)
--	g1444 = DFF(g28683)
--	g1439 = DFF(g29147)
--	g1435 = DFF(g29427)
--	g1430 = DFF(g29641)
--	g1426 = DFF(g29802)
--	g1562 = DFF(g20563)
--	g1564 = DFF(g1562)
--	g1563 = DFF(g1564)
--	g1657 = DFF(g13438)
--	g1786 = DFF(g1657)
--	g1782 = DFF(g1786)
--	g1690 = DFF(g11550)
--	g1735 = DFF(g28259)
--	g1724 = DFF(g28260)
--	g1727 = DFF(g28261)
--	g1750 = DFF(g28262)
--	g1739 = DFF(g28263)
--	g1742 = DFF(g28264)
--	g1765 = DFF(g28265)
--	g1754 = DFF(g28266)
--	g1757 = DFF(g28267)
--	g1779 = DFF(g28268)
--	g1769 = DFF(g28269)
--	g1772 = DFF(g28270)
--	g1789 = DFF(g29434)
--	g1792 = DFF(g29435)
--	g1795 = DFF(g29436)
--	g1798 = DFF(g29645)
--	g1801 = DFF(g29646)
--	g1804 = DFF(g29647)
--	g1808 = DFF(g29437)
--	g1809 = DFF(g29438)
--	g1807 = DFF(g29439)
--	g1810 = DFF(g27700)
--	g1813 = DFF(g27701)
--	g1816 = DFF(g27702)
--	g1819 = DFF(g27703)
--	g1822 = DFF(g27704)
--	g1825 = DFF(g27705)
--	g1829 = DFF(g28684)
--	g1830 = DFF(g28685)
--	g1828 = DFF(g28686)
--	g1693 = DFF(g29803)
--	g1694 = DFF(g29804)
--	g1695 = DFF(g29805)
--	g1696 = DFF(g30887)
--	g1697 = DFF(g30888)
--	g1698 = DFF(g30889)
--	g1699 = DFF(g30716)
--	g1700 = DFF(g30717)
--	g1701 = DFF(g30718)
--	g1703 = DFF(g29642)
--	g1704 = DFF(g29643)
--	g1702 = DFF(g29644)
--	g1784 = DFF(g27221)
--	g1785 = DFF(g27222)
--	g1783 = DFF(g27223)
--	g1831 = DFF(g11563)
--	g1832 = DFF(g1831)
--	g1833 = DFF(g11564)
--	g1834 = DFF(g1833)
--	g1835 = DFF(g11565)
--	g1660 = DFF(g1835)
--	g1661 = DFF(g11545)
--	g1662 = DFF(g1661)
--	g1663 = DFF(g11546)
--	g1664 = DFF(g1663)
--	g1665 = DFF(g11547)
--	g1666 = DFF(g1665)
--	g1667 = DFF(g11548)
--	g1668 = DFF(g1667)
--	g1669 = DFF(g11549)
--	g1670 = DFF(g1669)
--	g1671 = DFF(g13439)
--	g1672 = DFF(g1671)
--	g1680 = DFF(g19036)
--	g1686 = DFF(g29428)
--	g1689 = DFF(g29429)
--	g1678 = DFF(g29430)
--	g1677 = DFF(g29431)
--	g1676 = DFF(g29432)
--	g1675 = DFF(g29433)
--	g1685 = DFF(g19040)
--	g1684 = DFF(g19039)
--	g1683 = DFF(g19038)
--	g1682 = DFF(g19037)
--	g1681 = DFF(g25152)
--	g1679 = DFF(g27220)
--	g1723 = DFF(g11551)
--	g1730 = DFF(g1723)
--	g1731 = DFF(g11552)
--	g1732 = DFF(g1731)
--	g1733 = DFF(g11553)
--	g1734 = DFF(g1733)
--	g1738 = DFF(g11554)
--	g1745 = DFF(g1738)
--	g1746 = DFF(g11555)
--	g1747 = DFF(g1746)
--	g1748 = DFF(g11556)
--	g1749 = DFF(g1748)
--	g1753 = DFF(g11557)
--	g1760 = DFF(g1753)
--	g1761 = DFF(g11558)
--	g1762 = DFF(g1761)
--	g1763 = DFF(g11559)
--	g1764 = DFF(g1763)
--	g1768 = DFF(g11560)
--	g1775 = DFF(g1768)
--	g1776 = DFF(g11561)
--	g1777 = DFF(g1776)
--	g1778 = DFF(g11562)
--	g1705 = DFF(g1778)
--	g1706 = DFF(g13440)
--	g1712 = DFF(g1706)
--	g1718 = DFF(g1712)
--	g1925 = DFF(g13451)
--	g1931 = DFF(g1925)
--	g1930 = DFF(g1931)
--	g1934 = DFF(g23236)
--	g1937 = DFF(g20564)
--	g1890 = DFF(g20565)
--	g1893 = DFF(g16471)
--	g1903 = DFF(g1893)
--	g1904 = DFF(g1903)
--	g1944 = DFF(g11566)
--	g1949 = DFF(g1944)
--	g1950 = DFF(g11569)
--	g1951 = DFF(g1950)
--	g1952 = DFF(g11570)
--	g1953 = DFF(g1952)
--	g1954 = DFF(g11571)
--	g1945 = DFF(g1954)
--	g1946 = DFF(g11567)
--	g1947 = DFF(g1946)
--	g1948 = DFF(g11568)
--	g1870 = DFF(g1948)
--	g1855 = DFF(g13441)
--	g1862 = DFF(g1855)
--	g1866 = DFF(g1862)
--	g1867 = DFF(g24374)
--	g1868 = DFF(g24375)
--	g1869 = DFF(g24376)
--	g1836 = DFF(g25161)
--	g1839 = DFF(g25153)
--	g1842 = DFF(g25154)
--	g1858 = DFF(g25158)
--	g1859 = DFF(g25159)
--	g1860 = DFF(g25160)
--	g1861 = DFF(g24371)
--	g1865 = DFF(g24372)
--	g1845 = DFF(g24373)
--	g1846 = DFF(g25155)
--	g1849 = DFF(g25156)
--	g1852 = DFF(g25157)
--	g1908 = DFF(g16472)
--	g1915 = DFF(g1908)
--	g1922 = DFF(g1915)
--	g1923 = DFF(g19045)
--	g1924 = DFF(g1923)
--	g1928 = DFF(g29445)
--	g1929 = DFF(g19046)
--	g1880 = DFF(g1929)
--	g1938 = DFF(g19047)
--	g1939 = DFF(g1938)
--	g1956 = DFF(g28271)
--	g1957 = DFF(g28272)
--	g1955 = DFF(g28273)
--	g1959 = DFF(g28274)
--	g1960 = DFF(g28275)
--	g1958 = DFF(g28276)
--	g1962 = DFF(g28277)
--	g1963 = DFF(g28278)
--	g1961 = DFF(g28279)
--	g1965 = DFF(g28280)
--	g1966 = DFF(g28281)
--	g1964 = DFF(g28282)
--	g1967 = DFF(g26003)
--	g1970 = DFF(g26004)
--	g1973 = DFF(g26005)
--	g1976 = DFF(g26006)
--	g1979 = DFF(g26007)
--	g1982 = DFF(g26008)
--	g1994 = DFF(g29151)
--	g1997 = DFF(g29152)
--	g2000 = DFF(g29153)
--	g1985 = DFF(g29148)
--	g1988 = DFF(g29149)
--	g1991 = DFF(g29150)
--	g1871 = DFF(g27224)
--	g1874 = DFF(g27225)
--	g1877 = DFF(g27226)
--	g1886 = DFF(g8302)
--	g1887 = DFF(g24377)
--	g1888 = DFF(g19041)
--	g1889 = DFF(g19042)
--	g1894 = DFF(g19043)
--	g1895 = DFF(g19044)
--	g1896 = DFF(g29444)
--	g1897 = DFF(g29443)
--	g1898 = DFF(g29442)
--	g1899 = DFF(g29441)
--	g1900 = DFF(g29440)
--	g1905 = DFF(g1900)
--	g1909 = DFF(g13442)
--	g1910 = DFF(g13443)
--	g1911 = DFF(g13444)
--	g1912 = DFF(g13445)
--	g1913 = DFF(g13446)
--	g1914 = DFF(g13447)
--	g1916 = DFF(g13448)
--	g1917 = DFF(g13449)
--	g1918 = DFF(g26002)
--	g1921 = DFF(g13450)
--	g2003 = DFF(g13452)
--	g2006 = DFF(g2003)
--	g2009 = DFF(g2006)
--	g2010 = DFF(g20566)
--	g2039 = DFF(g21945)
--	g2020 = DFF(g23237)
--	g2013 = DFF(g24378)
--	g2033 = DFF(g25162)
--	g2026 = DFF(g26009)
--	g2040 = DFF(g26725)
--	g2052 = DFF(g27227)
--	g2046 = DFF(g27706)
--	g2059 = DFF(g28283)
--	g2066 = DFF(g28687)
--	g2072 = DFF(g29154)
--	g2079 = DFF(g23238)
--	g2080 = DFF(g23239)
--	g2078 = DFF(g23240)
--	g2082 = DFF(g23241)
--	g2083 = DFF(g23242)
--	g2081 = DFF(g23243)
--	g2085 = DFF(g23244)
--	g2086 = DFF(g23245)
--	g2084 = DFF(g23246)
--	g2088 = DFF(g23247)
--	g2089 = DFF(g23248)
--	g2087 = DFF(g23249)
--	g2091 = DFF(g23250)
--	g2092 = DFF(g23251)
--	g2090 = DFF(g23252)
--	g2094 = DFF(g23253)
--	g2095 = DFF(g23254)
--	g2093 = DFF(g23255)
--	g2097 = DFF(g23256)
--	g2098 = DFF(g23257)
--	g2096 = DFF(g23258)
--	g2100 = DFF(g23259)
--	g2101 = DFF(g23260)
--	g2099 = DFF(g23261)
--	g2103 = DFF(g23262)
--	g2104 = DFF(g23263)
--	g2102 = DFF(g23264)
--	g2106 = DFF(g23265)
--	g2107 = DFF(g23266)
--	g2105 = DFF(g23267)
--	g2109 = DFF(g23268)
--	g2110 = DFF(g23269)
--	g2108 = DFF(g23270)
--	g2112 = DFF(g23271)
--	g2113 = DFF(g23272)
--	g2111 = DFF(g23273)
--	g2115 = DFF(g26726)
--	g2116 = DFF(g26727)
--	g2114 = DFF(g26728)
--	g2118 = DFF(g24379)
--	g2119 = DFF(g24380)
--	g2117 = DFF(g24381)
--	g2214 = DFF(g13453)
--	g2211 = DFF(g2214)
--	g2241 = DFF(g2211)
--	g2206 = DFF(g24382)
--	g2207 = DFF(g24383)
--	g2205 = DFF(g24384)
--	g2209 = DFF(g24385)
--	g2210 = DFF(g24386)
--	g2208 = DFF(g24387)
--	g2218 = DFF(g24388)
--	g2219 = DFF(g24389)
--	g2217 = DFF(g24390)
--	g2221 = DFF(g24391)
--	g2222 = DFF(g24392)
--	g2220 = DFF(g24393)
--	g2224 = DFF(g24394)
--	g2225 = DFF(g24395)
--	g2223 = DFF(g24396)
--	g2227 = DFF(g24397)
--	g2228 = DFF(g24398)
--	g2226 = DFF(g24399)
--	g2230 = DFF(g24400)
--	g2231 = DFF(g24401)
--	g2229 = DFF(g24402)
--	g2233 = DFF(g24403)
--	g2234 = DFF(g24404)
--	g2232 = DFF(g24405)
--	g2236 = DFF(g24406)
--	g2237 = DFF(g24407)
--	g2235 = DFF(g24408)
--	g2239 = DFF(g24409)
--	g2240 = DFF(g24410)
--	g2238 = DFF(g24411)
--	g2245 = DFF(g26730)
--	g2246 = DFF(g26731)
--	g2244 = DFF(g26732)
--	g2248 = DFF(g26733)
--	g2249 = DFF(g26734)
--	g2247 = DFF(g26735)
--	g2251 = DFF(g26736)
--	g2252 = DFF(g26737)
--	g2250 = DFF(g26738)
--	g2254 = DFF(g26739)
--	g2255 = DFF(g26740)
--	g2253 = DFF(g26741)
--	g2261 = DFF(g30551)
--	g2264 = DFF(g30552)
--	g2267 = DFF(g30553)
--	g2306 = DFF(g30896)
--	g2309 = DFF(g30897)
--	g2312 = DFF(g30898)
--	g2270 = DFF(g30890)
--	g2273 = DFF(g30891)
--	g2276 = DFF(g30892)
--	g2315 = DFF(g30899)
--	g2318 = DFF(g30900)
--	g2321 = DFF(g30901)
--	g2279 = DFF(g30554)
--	g2282 = DFF(g30555)
--	g2285 = DFF(g30556)
--	g2324 = DFF(g30560)
--	g2327 = DFF(g30561)
--	g2330 = DFF(g30562)
--	g2288 = DFF(g30557)
--	g2291 = DFF(g30558)
--	g2294 = DFF(g30559)
--	g2333 = DFF(g30563)
--	g2336 = DFF(g30564)
--	g2339 = DFF(g30565)
--	g2297 = DFF(g30893)
--	g2300 = DFF(g30894)
--	g2303 = DFF(g30895)
--	g2342 = DFF(g30902)
--	g2345 = DFF(g30903)
--	g2348 = DFF(g30904)
--	g2160 = DFF(g26010)
--	g2156 = DFF(g26729)
--	g2151 = DFF(g27228)
--	g2147 = DFF(g27707)
--	g2142 = DFF(g28284)
--	g2138 = DFF(g28688)
--	g2133 = DFF(g29155)
--	g2129 = DFF(g29446)
--	g2124 = DFF(g29648)
--	g2120 = DFF(g29806)
--	g2256 = DFF(g20567)
--	g2258 = DFF(g2256)
--	g2257 = DFF(g2258)
--	g2351 = DFF(g13454)
--	g2480 = DFF(g2351)
--	g2476 = DFF(g2480)
--	g2384 = DFF(g11577)
--	g2429 = DFF(g28285)
--	g2418 = DFF(g28286)
--	g2421 = DFF(g28287)
--	g2444 = DFF(g28288)
--	g2433 = DFF(g28289)
--	g2436 = DFF(g28290)
--	g2459 = DFF(g28291)
--	g2448 = DFF(g28292)
--	g2451 = DFF(g28293)
--	g2473 = DFF(g28294)
--	g2463 = DFF(g28295)
--	g2466 = DFF(g28296)
--	g2483 = DFF(g29447)
--	g2486 = DFF(g29448)
--	g2489 = DFF(g29449)
--	g2492 = DFF(g29652)
--	g2495 = DFF(g29653)
--	g2498 = DFF(g29654)
--	g2502 = DFF(g29450)
--	g2503 = DFF(g29451)
--	g2501 = DFF(g29452)
--	g2504 = DFF(g27708)
--	g2507 = DFF(g27709)
--	g2510 = DFF(g27710)
--	g2513 = DFF(g27711)
--	g2516 = DFF(g27712)
--	g2519 = DFF(g27713)
--	g2523 = DFF(g28689)
--	g2524 = DFF(g28690)
--	g2522 = DFF(g28691)
--	g2387 = DFF(g29807)
--	g2388 = DFF(g29808)
--	g2389 = DFF(g29809)
--	g2390 = DFF(g30905)
--	g2391 = DFF(g30906)
--	g2392 = DFF(g30907)
--	g2393 = DFF(g30719)
--	g2394 = DFF(g30720)
--	g2395 = DFF(g30721)
--	g2397 = DFF(g29649)
--	g2398 = DFF(g29650)
--	g2396 = DFF(g29651)
--	g2478 = DFF(g27230)
--	g2479 = DFF(g27231)
--	g2477 = DFF(g27232)
--	g2525 = DFF(g11590)
--	g2526 = DFF(g2525)
--	g2527 = DFF(g11591)
--	g2528 = DFF(g2527)
--	g2529 = DFF(g11592)
--	g2354 = DFF(g2529)
--	g2355 = DFF(g11572)
--	g2356 = DFF(g2355)
--	g2357 = DFF(g11573)
--	g2358 = DFF(g2357)
--	g2359 = DFF(g11574)
--	g2360 = DFF(g2359)
--	g2361 = DFF(g11575)
--	g2362 = DFF(g2361)
--	g2363 = DFF(g11576)
--	g2364 = DFF(g2363)
--	g2365 = DFF(g13455)
--	g2366 = DFF(g2365)
--	g2374 = DFF(g19048)
--	g2380 = DFF(g30314)
--	g2383 = DFF(g30315)
--	g2372 = DFF(g30316)
--	g2371 = DFF(g30317)
--	g2370 = DFF(g30318)
--	g2369 = DFF(g30319)
--	g2379 = DFF(g19052)
--	g2378 = DFF(g19051)
--	g2377 = DFF(g19050)
--	g2376 = DFF(g19049)
--	g2375 = DFF(g25163)
--	g2373 = DFF(g27229)
--	g2417 = DFF(g11578)
--	g2424 = DFF(g2417)
--	g2425 = DFF(g11579)
--	g2426 = DFF(g2425)
--	g2427 = DFF(g11580)
--	g2428 = DFF(g2427)
--	g2432 = DFF(g11581)
--	g2439 = DFF(g2432)
--	g2440 = DFF(g11582)
--	g2441 = DFF(g2440)
--	g2442 = DFF(g11583)
--	g2443 = DFF(g2442)
--	g2447 = DFF(g11584)
--	g2454 = DFF(g2447)
--	g2455 = DFF(g11585)
--	g2456 = DFF(g2455)
--	g2457 = DFF(g11586)
--	g2458 = DFF(g2457)
--	g2462 = DFF(g11587)
--	g2469 = DFF(g2462)
--	g2470 = DFF(g11588)
--	g2471 = DFF(g2470)
--	g2472 = DFF(g11589)
--	g2399 = DFF(g2472)
--	g2400 = DFF(g13456)
--	g2406 = DFF(g2400)
--	g2412 = DFF(g2406)
--	g2619 = DFF(g13467)
--	g2625 = DFF(g2619)
--	g2624 = DFF(g2625)
--	g2628 = DFF(g23274)
--	g2631 = DFF(g20568)
--	g2584 = DFF(g20569)
--	g2587 = DFF(g16473)
--	g2597 = DFF(g2587)
--	g2598 = DFF(g2597)
--	g2638 = DFF(g11593)
--	g2643 = DFF(g2638)
--	g2644 = DFF(g11596)
--	g2645 = DFF(g2644)
--	g2646 = DFF(g11597)
--	g2647 = DFF(g2646)
--	g2648 = DFF(g11598)
--	g2639 = DFF(g2648)
--	g2640 = DFF(g11594)
--	g2641 = DFF(g2640)
--	g2642 = DFF(g11595)
--	g2564 = DFF(g2642)
--	g2549 = DFF(g13457)
--	g2556 = DFF(g2549)
--	g2560 = DFF(g2556)
--	g2561 = DFF(g24415)
--	g2562 = DFF(g24416)
--	g2563 = DFF(g24417)
--	g2530 = DFF(g25172)
--	g2533 = DFF(g25164)
--	g2536 = DFF(g25165)
--	g2552 = DFF(g25169)
--	g2553 = DFF(g25170)
--	g2554 = DFF(g25171)
--	g2555 = DFF(g24412)
--	g2559 = DFF(g24413)
--	g2539 = DFF(g24414)
--	g2540 = DFF(g25166)
--	g2543 = DFF(g25167)
--	g2546 = DFF(g25168)
--	g2602 = DFF(g16474)
--	g2609 = DFF(g2602)
--	g2616 = DFF(g2609)
--	g2617 = DFF(g19057)
--	g2618 = DFF(g2617)
--	g2622 = DFF(g30325)
--	g2623 = DFF(g19058)
--	g2574 = DFF(g2623)
--	g2632 = DFF(g19059)
--	g2633 = DFF(g2632)
--	g2650 = DFF(g28297)
--	g2651 = DFF(g28298)
--	g2649 = DFF(g28299)
--	g2653 = DFF(g28300)
--	g2654 = DFF(g28301)
--	g2652 = DFF(g28302)
--	g2656 = DFF(g28303)
--	g2657 = DFF(g28304)
--	g2655 = DFF(g28305)
--	g2659 = DFF(g28306)
--	g2660 = DFF(g28307)
--	g2658 = DFF(g28308)
--	g2661 = DFF(g26012)
--	g2664 = DFF(g26013)
--	g2667 = DFF(g26014)
--	g2670 = DFF(g26015)
--	g2673 = DFF(g26016)
--	g2676 = DFF(g26017)
--	g2688 = DFF(g29159)
--	g2691 = DFF(g29160)
--	g2694 = DFF(g29161)
--	g2679 = DFF(g29156)
--	g2682 = DFF(g29157)
--	g2685 = DFF(g29158)
--	g2565 = DFF(g27233)
--	g2568 = DFF(g27234)
--	g2571 = DFF(g27235)
--	g2580 = DFF(g8311)
--	g2581 = DFF(g24418)
--	g2582 = DFF(g19053)
--	g2583 = DFF(g19054)
--	g2588 = DFF(g19055)
--	g2589 = DFF(g19056)
--	g2590 = DFF(g30324)
--	g2591 = DFF(g30323)
--	g2592 = DFF(g30322)
--	g2593 = DFF(g30321)
--	g2594 = DFF(g30320)
--	g2599 = DFF(g2594)
--	g2603 = DFF(g13458)
--	g2604 = DFF(g13459)
--	g2605 = DFF(g13460)
--	g2606 = DFF(g13461)
--	g2607 = DFF(g13462)
--	g2608 = DFF(g13463)
--	g2610 = DFF(g13464)
--	g2611 = DFF(g13465)
--	g2612 = DFF(g26011)
--	g2615 = DFF(g13466)
--	g2697 = DFF(g13468)
--	g2700 = DFF(g2697)
--	g2703 = DFF(g2700)
--	g2704 = DFF(g20570)
--	g2733 = DFF(g21946)
--	g2714 = DFF(g23275)
--	g2707 = DFF(g24419)
--	g2727 = DFF(g25173)
--	g2720 = DFF(g26018)
--	g2734 = DFF(g26742)
--	g2746 = DFF(g27236)
--	g2740 = DFF(g27714)
--	g2753 = DFF(g28309)
--	g2760 = DFF(g28692)
--	g2766 = DFF(g29162)
--	g2773 = DFF(g23276)
--	g2774 = DFF(g23277)
--	g2772 = DFF(g23278)
--	g2776 = DFF(g23279)
--	g2777 = DFF(g23280)
--	g2775 = DFF(g23281)
--	g2779 = DFF(g23282)
--	g2780 = DFF(g23283)
--	g2778 = DFF(g23284)
--	g2782 = DFF(g23285)
--	g2783 = DFF(g23286)
--	g2781 = DFF(g23287)
--	g2785 = DFF(g23288)
--	g2786 = DFF(g23289)
--	g2784 = DFF(g23290)
--	g2788 = DFF(g23291)
--	g2789 = DFF(g23292)
--	g2787 = DFF(g23293)
--	g2791 = DFF(g23294)
--	g2792 = DFF(g23295)
--	g2790 = DFF(g23296)
--	g2794 = DFF(g23297)
--	g2795 = DFF(g23298)
--	g2793 = DFF(g23299)
--	g2797 = DFF(g23300)
--	g2798 = DFF(g23301)
--	g2796 = DFF(g23302)
--	g2800 = DFF(g23303)
--	g2801 = DFF(g23304)
--	g2799 = DFF(g23305)
--	g2803 = DFF(g23306)
--	g2804 = DFF(g23307)
--	g2802 = DFF(g23308)
--	g2806 = DFF(g23309)
--	g2807 = DFF(g23310)
--	g2805 = DFF(g23311)
--	g2809 = DFF(g26743)
--	g2810 = DFF(g26744)
--	g2808 = DFF(g26745)
--	g2812 = DFF(g24420)
--	g2813 = DFF(g24421)
--	g2811 = DFF(g24422)
--	g3054 = DFF(g23317)
--	g3079 = DFF(g23318)
--	g3080 = DFF(g21965)
--	g3043 = DFF(g29453)
--	g3044 = DFF(g29454)
--	g3045 = DFF(g29455)
--	g3046 = DFF(g29456)
--	g3047 = DFF(g29457)
--	g3048 = DFF(g29458)
--	g3049 = DFF(g29459)
--	g3050 = DFF(g29460)
--	g3051 = DFF(g29655)
--	g3052 = DFF(g29972)
--	g3053 = DFF(g29973)
--	g3055 = DFF(g29974)
--	g3056 = DFF(g29975)
--	g3057 = DFF(g29976)
--	g3058 = DFF(g29977)
--	g3059 = DFF(g29978)
--	g3060 = DFF(g29979)
--	g3061 = DFF(g30119)
--	g3062 = DFF(g30908)
--	g3063 = DFF(g30909)
--	g3064 = DFF(g30910)
--	g3065 = DFF(g30911)
--	g3066 = DFF(g30912)
--	g3067 = DFF(g30913)
--	g3068 = DFF(g30914)
--	g3069 = DFF(g30915)
--	g3070 = DFF(g30940)
--	g3071 = DFF(g30980)
--	g3072 = DFF(g30981)
--	g3073 = DFF(g30982)
--	g3074 = DFF(g30983)
--	g3075 = DFF(g30984)
--	g3076 = DFF(g30985)
--	g3077 = DFF(g30986)
--	g3078 = DFF(g30987)
--	g2997 = DFF(g30989)
--	g2993 = DFF(g26748)
--	g2998 = DFF(g27238)
--	g3006 = DFF(g25177)
--	g3002 = DFF(g26021)
--	g3013 = DFF(g26750)
--	g3010 = DFF(g27239)
--	g3024 = DFF(g27716)
--	g3018 = DFF(g24425)
--	g3028 = DFF(g25176)
--	g3036 = DFF(g26022)
--	g3032 = DFF(g26749)
--	g3040 = DFF(g16497)
--	g2986 = DFF(g3040)
--	g2987 = DFF(g16495)
--	g48 = DFF(g20595)
--	g45 = DFF(g20596)
--	g42 = DFF(g20597)
--	g39 = DFF(g20598)
--	g27 = DFF(g20599)
--	g30 = DFF(g20600)
--	g33 = DFF(g20601)
--	g36 = DFF(g20602)
--	g3083 = DFF(g20603)
--	g26 = DFF(g20604)
--	g2992 = DFF(g21966)
--	g23 = DFF(g20605)
--	g20 = DFF(g20606)
--	g17 = DFF(g20607)
--	g11 = DFF(g20608)
--	g14 = DFF(g20589)
--	g5 = DFF(g20590)
--	g8 = DFF(g20591)
--	g2 = DFF(g20592)
--	g2990 = DFF(g20593)
--	g2991 = DFF(g21964)
--	g1 = DFF(g20594)
--	
--	I13089 = NOT(g563)
--	g562 = NOT(I13089)
--	I13092 = NOT(g1249)
--	g1248 = NOT(I13092)
--	I13095 = NOT(g1943)
--	g1942 = NOT(I13095)
--	I13098 = NOT(g2637)
--	g2636 = NOT(I13098)
--	I13101 = NOT(g1)
--	g3235 = NOT(I13101)
--	I13104 = NOT(g2)
--	g3236 = NOT(I13104)
--	I13107 = NOT(g5)
--	g3237 = NOT(I13107)
--	I13110 = NOT(g8)
--	g3238 = NOT(I13110)
--	I13113 = NOT(g11)
--	g3239 = NOT(I13113)
--	I13116 = NOT(g14)
--	g3240 = NOT(I13116)
--	I13119 = NOT(g17)
--	g3241 = NOT(I13119)
--	I13122 = NOT(g20)
--	g3242 = NOT(I13122)
--	I13125 = NOT(g23)
--	g3243 = NOT(I13125)
--	I13128 = NOT(g26)
--	g3244 = NOT(I13128)
--	I13131 = NOT(g27)
--	g3245 = NOT(I13131)
--	I13134 = NOT(g30)
--	g3246 = NOT(I13134)
--	I13137 = NOT(g33)
--	g3247 = NOT(I13137)
--	I13140 = NOT(g36)
--	g3248 = NOT(I13140)
--	I13143 = NOT(g39)
--	g3249 = NOT(I13143)
--	I13146 = NOT(g42)
--	g3250 = NOT(I13146)
--	I13149 = NOT(g45)
--	g3251 = NOT(I13149)
--	I13152 = NOT(g48)
--	g3252 = NOT(I13152)
--	I13155 = NOT(g51)
--	g3253 = NOT(I13155)
--	I13158 = NOT(g165)
--	g3254 = NOT(I13158)
--	I13161 = NOT(g308)
--	g3304 = NOT(I13161)
--	g3305 = NOT(g305)
--	I13165 = NOT(g401)
--	g3306 = NOT(I13165)
--	g3337 = NOT(g309)
--	I13169 = NOT(g550)
--	g3338 = NOT(I13169)
--	g3365 = NOT(g499)
--	I13173 = NOT(g629)
--	g3366 = NOT(I13173)
--	I13176 = NOT(g630)
--	g3398 = NOT(I13176)
--	I13179 = NOT(g853)
--	g3410 = NOT(I13179)
--	I13182 = NOT(g995)
--	g3460 = NOT(I13182)
--	g3461 = NOT(g992)
--	I13186 = NOT(g1088)
--	g3462 = NOT(I13186)
--	g3493 = NOT(g996)
--	I13190 = NOT(g1236)
--	g3494 = NOT(I13190)
--	g3521 = NOT(g1186)
--	I13194 = NOT(g1315)
--	g3522 = NOT(I13194)
--	I13197 = NOT(g1316)
--	g3554 = NOT(I13197)
--	I13200 = NOT(g1547)
--	g3566 = NOT(I13200)
--	I13203 = NOT(g1689)
--	g3616 = NOT(I13203)
--	g3617 = NOT(g1686)
--	I13207 = NOT(g1782)
--	g3618 = NOT(I13207)
--	g3649 = NOT(g1690)
--	I13211 = NOT(g1930)
--	g3650 = NOT(I13211)
--	g3677 = NOT(g1880)
--	I13215 = NOT(g2009)
--	g3678 = NOT(I13215)
--	I13218 = NOT(g2010)
--	g3710 = NOT(I13218)
--	I13221 = NOT(g2241)
--	g3722 = NOT(I13221)
--	I13224 = NOT(g2383)
--	g3772 = NOT(I13224)
--	g3773 = NOT(g2380)
--	I13228 = NOT(g2476)
--	g3774 = NOT(I13228)
--	g3805 = NOT(g2384)
--	I13232 = NOT(g2624)
--	g3806 = NOT(I13232)
--	g3833 = NOT(g2574)
--	I13236 = NOT(g2703)
--	g3834 = NOT(I13236)
--	I13239 = NOT(g2704)
--	g3866 = NOT(I13239)
--	I13242 = NOT(g2879)
--	g3878 = NOT(I13242)
--	g3897 = NOT(g2950)
--	I13246 = NOT(g2987)
--	g3900 = NOT(I13246)
--	g3919 = NOT(g3080)
--	g3922 = NOT(g150)
--	g3925 = NOT(g155)
--	g3928 = NOT(g157)
--	g3931 = NOT(g171)
--	g3934 = NOT(g176)
--	g3937 = NOT(g178)
--	g3940 = NOT(g408)
--	g3941 = NOT(g455)
--	g3942 = NOT(g699)
--	g3945 = NOT(g726)
--	g3948 = NOT(g835)
--	g3951 = NOT(g840)
--	g3954 = NOT(g842)
--	g3957 = NOT(g856)
--	g3960 = NOT(g861)
--	g3963 = NOT(g863)
--	g3966 = NOT(g1526)
--	g3969 = NOT(g1531)
--	g3972 = NOT(g1533)
--	g3975 = NOT(g1552)
--	g3978 = NOT(g1554)
--	g3981 = NOT(g2217)
--	g3984 = NOT(g2222)
--	g3987 = NOT(g2224)
--	g3990 = NOT(g2245)
--	I13275 = NOT(g2848)
--	g3993 = NOT(I13275)
--	g3994 = NOT(g2848)
--	g3995 = NOT(g3064)
--	g3996 = NOT(g3073)
--	g3997 = NOT(g45)
--	g3998 = NOT(g23)
--	g3999 = NOT(g3204)
--	g4000 = NOT(g153)
--	g4003 = NOT(g158)
--	g4006 = NOT(g160)
--	g4009 = NOT(g174)
--	g4012 = NOT(g179)
--	g4015 = NOT(g411)
--	g4016 = NOT(g417)
--	g4017 = NOT(g427)
--	g4020 = NOT(g700)
--	g4023 = NOT(g702)
--	g4026 = NOT(g727)
--	g4029 = NOT(g838)
--	g4032 = NOT(g843)
--	g4035 = NOT(g845)
--	g4038 = NOT(g859)
--	g4041 = NOT(g864)
--	g4044 = NOT(g866)
--	g4047 = NOT(g1095)
--	g4048 = NOT(g1142)
--	g4049 = NOT(g1385)
--	g4052 = NOT(g1412)
--	g4055 = NOT(g1529)
--	g4058 = NOT(g1534)
--	g4061 = NOT(g1536)
--	g4064 = NOT(g1550)
--	g4067 = NOT(g1555)
--	g4070 = NOT(g1557)
--	g4073 = NOT(g2220)
--	g4076 = NOT(g2225)
--	g4079 = NOT(g2227)
--	g4082 = NOT(g2246)
--	g4085 = NOT(g2248)
--	I13316 = NOT(g2836)
--	g4088 = NOT(I13316)
--	g4089 = NOT(g2836)
--	I13320 = NOT(g2864)
--	g4090 = NOT(I13320)
--	g4091 = NOT(g2864)
--	g4092 = NOT(g3074)
--	g4093 = NOT(g33)
--	g4094 = NOT(g3207)
--	g4095 = NOT(g130)
--	g4098 = NOT(g156)
--	g4101 = NOT(g161)
--	g4104 = NOT(g163)
--	g4107 = NOT(g177)
--	g4110 = NOT(g414)
--	g4111 = NOT(g420)
--	g4112 = NOT(g428)
--	g4115 = NOT(g698)
--	g4118 = NOT(g703)
--	g4121 = NOT(g705)
--	g4124 = NOT(g725)
--	g4127 = NOT(g841)
--	g4130 = NOT(g846)
--	g4133 = NOT(g848)
--	g4136 = NOT(g862)
--	g4139 = NOT(g867)
--	g4142 = NOT(g1098)
--	g4143 = NOT(g1104)
--	g4144 = NOT(g1114)
--	g4147 = NOT(g1386)
--	g4150 = NOT(g1388)
--	g4153 = NOT(g1413)
--	g4156 = NOT(g1532)
--	g4159 = NOT(g1537)
--	g4162 = NOT(g1539)
--	g4165 = NOT(g1553)
--	g4168 = NOT(g1558)
--	g4171 = NOT(g1560)
--	g4174 = NOT(g1789)
--	g4175 = NOT(g1836)
--	g4176 = NOT(g2079)
--	g4179 = NOT(g2106)
--	g4182 = NOT(g2223)
--	g4185 = NOT(g2228)
--	g4188 = NOT(g2230)
--	g4191 = NOT(g2244)
--	g4194 = NOT(g2249)
--	g4197 = NOT(g2251)
--	I13366 = NOT(g2851)
--	g4200 = NOT(I13366)
--	g4201 = NOT(g2851)
--	g4202 = NOT(g42)
--	g4203 = NOT(g20)
--	g4204 = NOT(g3188)
--	g4205 = NOT(g131)
--	g4208 = NOT(g133)
--	g4211 = NOT(g159)
--	g4214 = NOT(g164)
--	g4217 = NOT(g354)
--	g4220 = NOT(g423)
--	g4221 = NOT(g426)
--	g4224 = NOT(g429)
--	g4225 = NOT(g701)
--	g4228 = NOT(g706)
--	g4231 = NOT(g708)
--	g4234 = NOT(g818)
--	g4237 = NOT(g844)
--	g4240 = NOT(g849)
--	g4243 = NOT(g851)
--	g4246 = NOT(g865)
--	g4249 = NOT(g1101)
--	g4250 = NOT(g1107)
--	g4251 = NOT(g1115)
--	g4254 = NOT(g1384)
--	g4257 = NOT(g1389)
--	g4260 = NOT(g1391)
--	g4263 = NOT(g1411)
--	g4266 = NOT(g1535)
--	g4269 = NOT(g1540)
--	g4272 = NOT(g1542)
--	g4275 = NOT(g1556)
--	g4278 = NOT(g1561)
--	g4281 = NOT(g1792)
--	g4282 = NOT(g1798)
--	g4283 = NOT(g1808)
--	g4286 = NOT(g2080)
--	g4289 = NOT(g2082)
--	g4292 = NOT(g2107)
--	g4295 = NOT(g2226)
--	g4298 = NOT(g2231)
--	g4301 = NOT(g2233)
--	g4304 = NOT(g2247)
--	g4307 = NOT(g2252)
--	g4310 = NOT(g2254)
--	g4313 = NOT(g2483)
--	g4314 = NOT(g2530)
--	g4315 = NOT(g2773)
--	g4318 = NOT(g2800)
--	I13417 = NOT(g2839)
--	g4321 = NOT(I13417)
--	g4322 = NOT(g2839)
--	I13421 = NOT(g2867)
--	g4323 = NOT(I13421)
--	g4324 = NOT(g2867)
--	g4325 = NOT(g36)
--	g4326 = NOT(g181)
--	g4329 = NOT(g129)
--	g4332 = NOT(g134)
--	g4335 = NOT(g162)
--	I13430 = NOT(g101)
--	g4338 = NOT(I13430)
--	I13433 = NOT(g105)
--	g4339 = NOT(I13433)
--	g4340 = NOT(g343)
--	g4343 = NOT(g369)
--	g4346 = NOT(g432)
--	g4347 = NOT(g438)
--	g4348 = NOT(g704)
--	g4351 = NOT(g709)
--	g4354 = NOT(g711)
--	g4357 = NOT(g729)
--	g4360 = NOT(g819)
--	g4363 = NOT(g821)
--	g4366 = NOT(g847)
--	g4369 = NOT(g852)
--	g4372 = NOT(g1041)
--	g4375 = NOT(g1110)
--	g4376 = NOT(g1113)
--	g4379 = NOT(g1116)
--	g4380 = NOT(g1387)
--	g4383 = NOT(g1392)
--	g4386 = NOT(g1394)
--	g4389 = NOT(g1512)
--	g4392 = NOT(g1538)
--	g4395 = NOT(g1543)
--	g4398 = NOT(g1545)
--	g4401 = NOT(g1559)
--	g4404 = NOT(g1795)
--	g4405 = NOT(g1801)
--	g4406 = NOT(g1809)
--	g4409 = NOT(g2078)
--	g4412 = NOT(g2083)
--	g4415 = NOT(g2085)
--	g4418 = NOT(g2105)
--	g4421 = NOT(g2229)
--	g4424 = NOT(g2234)
--	g4427 = NOT(g2236)
--	g4430 = NOT(g2250)
--	g4433 = NOT(g2255)
--	g4436 = NOT(g2486)
--	g4437 = NOT(g2492)
--	g4438 = NOT(g2502)
--	g4441 = NOT(g2774)
--	g4444 = NOT(g2776)
--	g4447 = NOT(g2801)
--	I13478 = NOT(g2854)
--	g4450 = NOT(I13478)
--	g4451 = NOT(g2854)
--	g4452 = NOT(g17)
--	g4453 = NOT(g132)
--	g4456 = NOT(g309)
--	g4465 = NOT(g346)
--	g4468 = NOT(g358)
--	g4471 = NOT(g384)
--	g4474 = NOT(g435)
--	g4475 = NOT(g441)
--	g4476 = NOT(g576)
--	g4479 = NOT(g587)
--	g4480 = NOT(g707)
--	g4483 = NOT(g712)
--	g4486 = NOT(g714)
--	g4489 = NOT(g730)
--	g4492 = NOT(g732)
--	g4495 = NOT(g869)
--	g4498 = NOT(g817)
--	g4501 = NOT(g822)
--	g4504 = NOT(g850)
--	I13501 = NOT(g789)
--	g4507 = NOT(I13501)
--	I13504 = NOT(g793)
--	g4508 = NOT(I13504)
--	g4509 = NOT(g1030)
--	g4512 = NOT(g1056)
--	g4515 = NOT(g1119)
--	g4516 = NOT(g1125)
--	g4517 = NOT(g1390)
--	g4520 = NOT(g1395)
--	g4523 = NOT(g1397)
--	g4526 = NOT(g1415)
--	g4529 = NOT(g1513)
--	g4532 = NOT(g1515)
--	g4535 = NOT(g1541)
--	g4538 = NOT(g1546)
--	g4541 = NOT(g1735)
--	g4544 = NOT(g1804)
--	g4545 = NOT(g1807)
--	g4548 = NOT(g1810)
--	g4549 = NOT(g2081)
--	g4552 = NOT(g2086)
--	g4555 = NOT(g2088)
--	g4558 = NOT(g2206)
--	g4561 = NOT(g2232)
--	g4564 = NOT(g2237)
--	g4567 = NOT(g2239)
--	g4570 = NOT(g2253)
--	g4573 = NOT(g2489)
--	g4574 = NOT(g2495)
--	g4575 = NOT(g2503)
--	g4578 = NOT(g2772)
--	g4581 = NOT(g2777)
--	g4584 = NOT(g2779)
--	g4587 = NOT(g2799)
--	I13538 = NOT(g2870)
--	g4590 = NOT(I13538)
--	g4591 = NOT(g2870)
--	g4592 = NOT(g361)
--	g4595 = NOT(g373)
--	g4598 = NOT(g398)
--	g4601 = NOT(g444)
--	g4602 = NOT(g525)
--	g4603 = NOT(g577)
--	g4606 = NOT(g579)
--	g4609 = NOT(g590)
--	g4610 = NOT(g596)
--	g4611 = NOT(g710)
--	g4614 = NOT(g715)
--	g4617 = NOT(g717)
--	g4620 = NOT(g728)
--	g4623 = NOT(g733)
--	g4626 = NOT(g735)
--	g4629 = NOT(g820)
--	g4632 = NOT(g996)
--	g4641 = NOT(g1033)
--	g4644 = NOT(g1045)
--	g4647 = NOT(g1071)
--	g4650 = NOT(g1122)
--	g4651 = NOT(g1128)
--	g4652 = NOT(g1262)
--	g4655 = NOT(g1273)
--	g4656 = NOT(g1393)
--	g4659 = NOT(g1398)
--	g4662 = NOT(g1400)
--	g4665 = NOT(g1416)
--	g4668 = NOT(g1418)
--	g4671 = NOT(g1563)
--	g4674 = NOT(g1511)
--	g4677 = NOT(g1516)
--	g4680 = NOT(g1544)
--	I13575 = NOT(g1476)
--	g4683 = NOT(I13575)
--	I13578 = NOT(g1481)
--	g4684 = NOT(I13578)
--	g4685 = NOT(g1724)
--	g4688 = NOT(g1750)
--	g4691 = NOT(g1813)
--	g4692 = NOT(g1819)
--	g4693 = NOT(g2084)
--	g4696 = NOT(g2089)
--	g4699 = NOT(g2091)
--	g4702 = NOT(g2109)
--	g4705 = NOT(g2207)
--	g4708 = NOT(g2209)
--	g4711 = NOT(g2235)
--	g4714 = NOT(g2240)
--	g4717 = NOT(g2429)
--	g4720 = NOT(g2498)
--	g4721 = NOT(g2501)
--	g4724 = NOT(g2504)
--	g4725 = NOT(g2775)
--	g4728 = NOT(g2780)
--	g4731 = NOT(g2782)
--	g4734 = NOT(g11)
--	I13601 = NOT(g121)
--	g4735 = NOT(I13601)
--	I13604 = NOT(g125)
--	g4736 = NOT(I13604)
--	g4737 = NOT(g376)
--	g4740 = NOT(g388)
--	g4743 = NOT(g575)
--	g4746 = NOT(g580)
--	g4749 = NOT(g582)
--	g4752 = NOT(g593)
--	g4753 = NOT(g599)
--	g4754 = NOT(g713)
--	g4757 = NOT(g718)
--	g4760 = NOT(g720)
--	g4763 = NOT(g731)
--	g4766 = NOT(g736)
--	g4769 = NOT(g1048)
--	g4772 = NOT(g1060)
--	g4775 = NOT(g1085)
--	g4778 = NOT(g1131)
--	g4779 = NOT(g1211)
--	g4780 = NOT(g1263)
--	g4783 = NOT(g1265)
--	g4786 = NOT(g1276)
--	g4787 = NOT(g1282)
--	g4788 = NOT(g1396)
--	g4791 = NOT(g1401)
--	g4794 = NOT(g1403)
--	g4797 = NOT(g1414)
--	g4800 = NOT(g1419)
--	g4803 = NOT(g1421)
--	g4806 = NOT(g1514)
--	g4809 = NOT(g1690)
--	g4818 = NOT(g1727)
--	g4821 = NOT(g1739)
--	g4824 = NOT(g1765)
--	g4827 = NOT(g1816)
--	g4828 = NOT(g1822)
--	g4829 = NOT(g1956)
--	g4832 = NOT(g1967)
--	g4833 = NOT(g2087)
--	g4836 = NOT(g2092)
--	g4839 = NOT(g2094)
--	g4842 = NOT(g2110)
--	g4845 = NOT(g2112)
--	g4848 = NOT(g2257)
--	g4851 = NOT(g2205)
--	g4854 = NOT(g2210)
--	g4857 = NOT(g2238)
--	I13652 = NOT(g2170)
--	g4860 = NOT(I13652)
--	I13655 = NOT(g2175)
--	g4861 = NOT(I13655)
--	g4862 = NOT(g2418)
--	g4865 = NOT(g2444)
--	g4868 = NOT(g2507)
--	g4869 = NOT(g2513)
--	g4870 = NOT(g2778)
--	g4873 = NOT(g2783)
--	g4876 = NOT(g2785)
--	g4879 = NOT(g2803)
--	g4882 = NOT(g391)
--	g4885 = NOT(g448)
--	g4888 = NOT(g578)
--	g4891 = NOT(g583)
--	g4894 = NOT(g585)
--	g4897 = NOT(g602)
--	g4898 = NOT(g605)
--	g4899 = NOT(g716)
--	g4902 = NOT(g721)
--	g4905 = NOT(g723)
--	g4908 = NOT(g734)
--	I13677 = NOT(g809)
--	g4911 = NOT(I13677)
--	I13680 = NOT(g813)
--	g4912 = NOT(I13680)
--	g4913 = NOT(g1063)
--	g4916 = NOT(g1075)
--	g4919 = NOT(g1261)
--	g4922 = NOT(g1266)
--	g4925 = NOT(g1268)
--	g4928 = NOT(g1279)
--	g4929 = NOT(g1285)
--	g4930 = NOT(g1399)
--	g4933 = NOT(g1404)
--	g4936 = NOT(g1406)
--	g4939 = NOT(g1417)
--	g4942 = NOT(g1422)
--	g4945 = NOT(g1742)
--	g4948 = NOT(g1754)
--	g4951 = NOT(g1779)
--	g4954 = NOT(g1825)
--	g4955 = NOT(g1905)
--	g4956 = NOT(g1957)
--	g4959 = NOT(g1959)
--	g4962 = NOT(g1970)
--	g4963 = NOT(g1976)
--	g4964 = NOT(g2090)
--	g4967 = NOT(g2095)
--	g4970 = NOT(g2097)
--	g4973 = NOT(g2108)
--	g4976 = NOT(g2113)
--	g4979 = NOT(g2115)
--	g4982 = NOT(g2208)
--	g4985 = NOT(g2384)
--	g4994 = NOT(g2421)
--	g4997 = NOT(g2433)
--	g5000 = NOT(g2459)
--	g5003 = NOT(g2510)
--	g5004 = NOT(g2516)
--	g5005 = NOT(g2650)
--	g5008 = NOT(g2661)
--	g5009 = NOT(g2781)
--	g5012 = NOT(g2786)
--	g5015 = NOT(g2788)
--	g5018 = NOT(g2804)
--	g5021 = NOT(g2806)
--	g5024 = NOT(g449)
--	g5027 = NOT(g581)
--	g5030 = NOT(g586)
--	g5033 = NOT(g608)
--	g5034 = NOT(g614)
--	g5035 = NOT(g719)
--	g5038 = NOT(g724)
--	g5041 = NOT(g1078)
--	g5044 = NOT(g1135)
--	g5047 = NOT(g1264)
--	g5050 = NOT(g1269)
--	g5053 = NOT(g1271)
--	g5056 = NOT(g1288)
--	g5057 = NOT(g1291)
--	g5058 = NOT(g1402)
--	g5061 = NOT(g1407)
--	g5064 = NOT(g1409)
--	g5067 = NOT(g1420)
--	I13742 = NOT(g1501)
--	g5070 = NOT(I13742)
--	I13745 = NOT(g1506)
--	g5071 = NOT(I13745)
--	g5072 = NOT(g1757)
--	g5075 = NOT(g1769)
--	g5078 = NOT(g1955)
--	g5081 = NOT(g1960)
--	g5084 = NOT(g1962)
--	g5087 = NOT(g1973)
--	g5088 = NOT(g1979)
--	g5089 = NOT(g2093)
--	g5092 = NOT(g2098)
--	g5095 = NOT(g2100)
--	g5098 = NOT(g2111)
--	g5101 = NOT(g2116)
--	g5104 = NOT(g2436)
--	g5107 = NOT(g2448)
--	g5110 = NOT(g2473)
--	g5113 = NOT(g2519)
--	g5114 = NOT(g2599)
--	g5115 = NOT(g2651)
--	g5118 = NOT(g2653)
--	g5121 = NOT(g2664)
--	g5122 = NOT(g2670)
--	g5123 = NOT(g2784)
--	g5126 = NOT(g2789)
--	g5129 = NOT(g2791)
--	g5132 = NOT(g2802)
--	g5135 = NOT(g2807)
--	g5138 = NOT(g2809)
--	I13775 = NOT(g109)
--	g5141 = NOT(I13775)
--	g5142 = NOT(g447)
--	g5145 = NOT(g584)
--	g5148 = NOT(g611)
--	g5149 = NOT(g617)
--	g5150 = NOT(g722)
--	g5153 = NOT(g1136)
--	g5156 = NOT(g1267)
--	g5159 = NOT(g1272)
--	g5162 = NOT(g1294)
--	g5163 = NOT(g1300)
--	g5164 = NOT(g1405)
--	g5167 = NOT(g1410)
--	g5170 = NOT(g1772)
--	g5173 = NOT(g1829)
--	g5176 = NOT(g1958)
--	g5179 = NOT(g1963)
--	g5182 = NOT(g1965)
--	g5185 = NOT(g1982)
--	g5186 = NOT(g1985)
--	g5187 = NOT(g2096)
--	g5190 = NOT(g2101)
--	g5193 = NOT(g2103)
--	g5196 = NOT(g2114)
--	I13801 = NOT(g2195)
--	g5199 = NOT(I13801)
--	I13804 = NOT(g2200)
--	g5200 = NOT(I13804)
--	g5201 = NOT(g2451)
--	g5204 = NOT(g2463)
--	g5207 = NOT(g2649)
--	g5210 = NOT(g2654)
--	g5213 = NOT(g2656)
--	g5216 = NOT(g2667)
--	g5217 = NOT(g2673)
--	g5218 = NOT(g2787)
--	g5221 = NOT(g2792)
--	g5224 = NOT(g2794)
--	g5227 = NOT(g2805)
--	g5230 = NOT(g2810)
--	g5233 = NOT(g620)
--	I13820 = NOT(g797)
--	g5234 = NOT(I13820)
--	g5235 = NOT(g1134)
--	g5238 = NOT(g1270)
--	g5241 = NOT(g1297)
--	g5242 = NOT(g1303)
--	g5243 = NOT(g1408)
--	g5246 = NOT(g1830)
--	g5249 = NOT(g1961)
--	g5252 = NOT(g1966)
--	g5255 = NOT(g1988)
--	g5256 = NOT(g1994)
--	g5257 = NOT(g2099)
--	g5260 = NOT(g2104)
--	g5263 = NOT(g2466)
--	g5266 = NOT(g2523)
--	g5269 = NOT(g2652)
--	g5272 = NOT(g2657)
--	g5275 = NOT(g2659)
--	g5278 = NOT(g2676)
--	g5279 = NOT(g2679)
--	g5280 = NOT(g2790)
--	g5283 = NOT(g2795)
--	g5286 = NOT(g2797)
--	g5289 = NOT(g2808)
--	g5292 = NOT(g2857)
--	g5293 = NOT(g738)
--	g5296 = NOT(g1306)
--	I13849 = NOT(g1486)
--	g5297 = NOT(I13849)
--	g5298 = NOT(g1828)
--	g5301 = NOT(g1964)
--	g5304 = NOT(g1991)
--	g5305 = NOT(g1997)
--	g5306 = NOT(g2102)
--	g5309 = NOT(g2524)
--	g5312 = NOT(g2655)
--	g5315 = NOT(g2660)
--	g5318 = NOT(g2682)
--	g5319 = NOT(g2688)
--	g5320 = NOT(g2793)
--	g5323 = NOT(g2798)
--	g5326 = NOT(g2873)
--	g5327 = NOT(g739)
--	g5330 = NOT(g1424)
--	g5333 = NOT(g2000)
--	I13868 = NOT(g2180)
--	g5334 = NOT(I13868)
--	g5335 = NOT(g2522)
--	g5338 = NOT(g2658)
--	g5341 = NOT(g2685)
--	g5342 = NOT(g2691)
--	g5343 = NOT(g2796)
--	g5346 = NOT(g3106)
--	g5349 = NOT(g2877)
--	g5352 = NOT(g737)
--	g5355 = NOT(g1425)
--	g5358 = NOT(g2118)
--	g5361 = NOT(g2694)
--	g5362 = NOT(g2817)
--	g5363 = NOT(g3107)
--	g5366 = NOT(g2878)
--	g5369 = NOT(g1423)
--	g5372 = NOT(g2119)
--	g5375 = NOT(g2812)
--	g5378 = NOT(g2933)
--	g5379 = NOT(g3108)
--	g5382 = NOT(g2117)
--	g5385 = NOT(g2813)
--	I13892 = NOT(g3040)
--	g5388 = NOT(I13892)
--	g5389 = NOT(g3040)
--	I13896 = NOT(g343)
--	g5390 = NOT(I13896)
--	g5391 = NOT(g2811)
--	g5394 = NOT(g3054)
--	I13901 = NOT(g346)
--	g5395 = NOT(I13901)
--	I13904 = NOT(g358)
--	g5396 = NOT(I13904)
--	I13907 = NOT(g1030)
--	g5397 = NOT(I13907)
--	I13910 = NOT(g361)
--	g5398 = NOT(I13910)
--	I13913 = NOT(g373)
--	g5399 = NOT(I13913)
--	I13916 = NOT(g1033)
--	g5400 = NOT(I13916)
--	I13919 = NOT(g1045)
--	g5401 = NOT(I13919)
--	I13922 = NOT(g1724)
--	g5402 = NOT(I13922)
--	I13925 = NOT(g376)
--	g5403 = NOT(I13925)
--	I13928 = NOT(g388)
--	g5404 = NOT(I13928)
--	I13931 = NOT(g1048)
--	g5405 = NOT(I13931)
--	I13934 = NOT(g1060)
--	g5406 = NOT(I13934)
--	I13937 = NOT(g1727)
--	g5407 = NOT(I13937)
--	I13940 = NOT(g1739)
--	g5408 = NOT(I13940)
--	I13943 = NOT(g2418)
--	g5409 = NOT(I13943)
--	g5410 = NOT(g3079)
--	I13947 = NOT(g391)
--	g5411 = NOT(I13947)
--	I13950 = NOT(g1063)
--	g5412 = NOT(I13950)
--	I13953 = NOT(g1075)
--	g5413 = NOT(I13953)
--	I13956 = NOT(g1742)
--	g5414 = NOT(I13956)
--	I13959 = NOT(g1754)
--	g5415 = NOT(I13959)
--	I13962 = NOT(g2421)
--	g5416 = NOT(I13962)
--	I13965 = NOT(g2433)
--	g5417 = NOT(I13965)
--	I13968 = NOT(g1078)
--	g5418 = NOT(I13968)
--	I13971 = NOT(g1757)
--	g5419 = NOT(I13971)
--	I13974 = NOT(g1769)
--	g5420 = NOT(I13974)
--	I13977 = NOT(g2436)
--	g5421 = NOT(I13977)
--	I13980 = NOT(g2448)
--	g5422 = NOT(I13980)
--	g5423 = NOT(g2879)
--	I13984 = NOT(g1772)
--	g5424 = NOT(I13984)
--	I13987 = NOT(g2451)
--	g5425 = NOT(I13987)
--	I13990 = NOT(g2463)
--	g5426 = NOT(I13990)
--	I13993 = NOT(g2466)
--	g5427 = NOT(I13993)
--	g5428 = NOT(g3210)
--	g5431 = NOT(g3211)
--	g5434 = NOT(g3084)
--	I13999 = NOT(g276)
--	g5437 = NOT(I13999)
--	I14002 = NOT(g276)
--	g5438 = NOT(I14002)
--	g5469 = NOT(g3085)
--	I14006 = NOT(g963)
--	g5472 = NOT(I14006)
--	I14009 = NOT(g963)
--	g5473 = NOT(I14009)
--	g5504 = NOT(g3086)
--	g5507 = NOT(g3155)
--	I14014 = NOT(g499)
--	g5508 = NOT(I14014)
--	I14017 = NOT(g1657)
--	g5511 = NOT(I14017)
--	I14020 = NOT(g1657)
--	g5512 = NOT(I14020)
--	g5543 = NOT(g3087)
--	g5546 = NOT(g3164)
--	g5547 = NOT(g101)
--	g5548 = NOT(g105)
--	I14027 = NOT(g182)
--	g5549 = NOT(I14027)
--	I14030 = NOT(g182)
--	g5550 = NOT(I14030)
--	g5551 = NOT(g514)
--	I14034 = NOT(g1186)
--	g5552 = NOT(I14034)
--	I14037 = NOT(g2351)
--	g5555 = NOT(I14037)
--	I14040 = NOT(g2351)
--	g5556 = NOT(I14040)
--	g5587 = NOT(g3091)
--	g5590 = NOT(g3158)
--	g5591 = NOT(g3173)
--	g5592 = NOT(g515)
--	g5593 = NOT(g789)
--	g5594 = NOT(g793)
--	I14049 = NOT(g870)
--	g5595 = NOT(I14049)
--	I14052 = NOT(g870)
--	g5596 = NOT(I14052)
--	g5597 = NOT(g1200)
--	I14056 = NOT(g1880)
--	g5598 = NOT(I14056)
--	g5601 = NOT(g3092)
--	g5604 = NOT(g3167)
--	g5605 = NOT(g3182)
--	g5606 = NOT(g79)
--	g5609 = NOT(g1201)
--	g5610 = NOT(g1476)
--	g5611 = NOT(g1481)
--	I14066 = NOT(g1564)
--	g5612 = NOT(I14066)
--	I14069 = NOT(g1564)
--	g5613 = NOT(I14069)
--	g5614 = NOT(g1894)
--	I14073 = NOT(g2574)
--	g5615 = NOT(I14073)
--	g5618 = NOT(g3093)
--	g5621 = NOT(g3161)
--	g5622 = NOT(g3176)
--	g5623 = NOT(g70)
--	g5626 = NOT(g121)
--	g5627 = NOT(g125)
--	g5628 = NOT(g300)
--	I14083 = NOT(g325)
--	g5629 = NOT(I14083)
--	g5631 = NOT(g767)
--	g5634 = NOT(g1895)
--	g5635 = NOT(g2170)
--	g5636 = NOT(g2175)
--	I14091 = NOT(g2258)
--	g5637 = NOT(I14091)
--	I14094 = NOT(g2258)
--	g5638 = NOT(I14094)
--	g5639 = NOT(g2588)
--	g5640 = NOT(g3170)
--	g5641 = NOT(g3185)
--	g5642 = NOT(g61)
--	g5645 = NOT(g101)
--	g5646 = NOT(g213)
--	g5647 = NOT(g301)
--	I14104 = NOT(g331)
--	g5648 = NOT(I14104)
--	g5651 = NOT(g758)
--	g5654 = NOT(g809)
--	g5655 = NOT(g813)
--	g5656 = NOT(g987)
--	I14113 = NOT(g1012)
--	g5657 = NOT(I14113)
--	g5659 = NOT(g1453)
--	g5662 = NOT(g2589)
--	g5663 = NOT(g3179)
--	g5664 = NOT(g65)
--	g5665 = NOT(g105)
--	g5666 = NOT(g216)
--	g5667 = NOT(g222)
--	g5668 = NOT(g299)
--	g5675 = NOT(g302)
--	g5679 = NOT(g506)
--	g5680 = NOT(g749)
--	g5683 = NOT(g789)
--	g5684 = NOT(g900)
--	g5685 = NOT(g988)
--	I14134 = NOT(g1018)
--	g5686 = NOT(I14134)
--	g5689 = NOT(g1444)
--	g5692 = NOT(g1501)
--	g5693 = NOT(g1506)
--	g5694 = NOT(g1681)
--	I14143 = NOT(g1706)
--	g5695 = NOT(I14143)
--	g5697 = NOT(g2147)
--	g5700 = NOT(g3088)
--	I14149 = NOT(g3231)
--	g5701 = NOT(I14149)
--	g5702 = NOT(g56)
--	g5703 = NOT(g109)
--	g5704 = NOT(g219)
--	g5705 = NOT(g225)
--	g5706 = NOT(g231)
--	g5707 = NOT(g109)
--	g5708 = NOT(g303)
--	g5712 = NOT(g305)
--	I14163 = NOT(g113)
--	g5713 = NOT(I14163)
--	g5714 = NOT(g507)
--	g5715 = NOT(g541)
--	g5716 = NOT(g753)
--	g5717 = NOT(g793)
--	g5718 = NOT(g903)
--	g5719 = NOT(g909)
--	g5720 = NOT(g986)
--	g5727 = NOT(g989)
--	g5731 = NOT(g1192)
--	g5732 = NOT(g1435)
--	g5735 = NOT(g1476)
--	g5736 = NOT(g1594)
--	g5737 = NOT(g1682)
--	I14182 = NOT(g1712)
--	g5738 = NOT(I14182)
--	g5741 = NOT(g2138)
--	g5744 = NOT(g2195)
--	g5745 = NOT(g2200)
--	g5746 = NOT(g2375)
--	I14191 = NOT(g2400)
--	g5747 = NOT(I14191)
--	I14195 = NOT(g3212)
--	g5749 = NOT(I14195)
--	g5750 = NOT(g92)
--	g5751 = NOT(g52)
--	g5752 = NOT(g113)
--	g5753 = NOT(g228)
--	g5754 = NOT(g234)
--	g5755 = NOT(g240)
--	g5756 = NOT(g304)
--	g5759 = NOT(g508)
--	g5760 = NOT(g744)
--	g5761 = NOT(g797)
--	g5762 = NOT(g906)
--	g5763 = NOT(g912)
--	g5764 = NOT(g918)
--	g5765 = NOT(g797)
--	g5766 = NOT(g990)
--	g5770 = NOT(g992)
--	I14219 = NOT(g801)
--	g5771 = NOT(I14219)
--	g5772 = NOT(g1193)
--	g5773 = NOT(g1227)
--	g5774 = NOT(g1439)
--	g5775 = NOT(g1481)
--	g5776 = NOT(g1597)
--	g5777 = NOT(g1603)
--	g5778 = NOT(g1680)
--	g5785 = NOT(g1683)
--	g5789 = NOT(g1886)
--	g5790 = NOT(g2129)
--	g5793 = NOT(g2170)
--	g5794 = NOT(g2288)
--	g5795 = NOT(g2376)
--	I14238 = NOT(g2406)
--	g5796 = NOT(I14238)
--	I14243 = NOT(g3221)
--	g5799 = NOT(I14243)
--	I14246 = NOT(g3227)
--	g5800 = NOT(I14246)
--	I14249 = NOT(g3216)
--	g5801 = NOT(I14249)
--	g5802 = NOT(g83)
--	g5803 = NOT(g117)
--	g5804 = NOT(g237)
--	g5805 = NOT(g243)
--	g5806 = NOT(g249)
--	g5808 = NOT(g509)
--	g5809 = NOT(g780)
--	g5810 = NOT(g740)
--	g5811 = NOT(g801)
--	g5812 = NOT(g915)
--	g5813 = NOT(g921)
--	g5814 = NOT(g927)
--	g5815 = NOT(g991)
--	g5818 = NOT(g1194)
--	g5819 = NOT(g1430)
--	g5820 = NOT(g1486)
--	g5821 = NOT(g1600)
--	g5822 = NOT(g1606)
--	g5823 = NOT(g1612)
--	g5824 = NOT(g1486)
--	g5825 = NOT(g1684)
--	g5829 = NOT(g1686)
--	I14280 = NOT(g1491)
--	g5830 = NOT(I14280)
--	g5831 = NOT(g1887)
--	g5832 = NOT(g1921)
--	g5833 = NOT(g2133)
--	g5834 = NOT(g2175)
--	g5835 = NOT(g2291)
--	g5836 = NOT(g2297)
--	g5837 = NOT(g2374)
--	g5844 = NOT(g2377)
--	g5848 = NOT(g2580)
--	I14295 = NOT(g3228)
--	g5849 = NOT(I14295)
--	I14298 = NOT(g3217)
--	g5850 = NOT(I14298)
--	g5851 = NOT(g74)
--	g5852 = NOT(g121)
--	g5853 = NOT(g246)
--	g5854 = NOT(g252)
--	g5855 = NOT(g258)
--	I14306 = NOT(g97)
--	g5856 = NOT(I14306)
--	g5857 = NOT(g538)
--	g5858 = NOT(g771)
--	g5859 = NOT(g805)
--	g5860 = NOT(g924)
--	g5861 = NOT(g930)
--	g5862 = NOT(g936)
--	g5864 = NOT(g1195)
--	g5865 = NOT(g1466)
--	g5866 = NOT(g1426)
--	g5867 = NOT(g1491)
--	g5868 = NOT(g1609)
--	g5869 = NOT(g1615)
--	g5870 = NOT(g1621)
--	g5871 = NOT(g1685)
--	g5874 = NOT(g1888)
--	g5875 = NOT(g2124)
--	g5876 = NOT(g2180)
--	g5877 = NOT(g2294)
--	g5878 = NOT(g2300)
--	g5879 = NOT(g2306)
--	g5880 = NOT(g2180)
--	g5881 = NOT(g2378)
--	g5885 = NOT(g2380)
--	I14338 = NOT(g2185)
--	g5886 = NOT(I14338)
--	g5887 = NOT(g2581)
--	g5888 = NOT(g2615)
--	I14343 = NOT(g3219)
--	g5889 = NOT(I14343)
--	g5890 = NOT(g88)
--	g5893 = NOT(g125)
--	g5894 = NOT(g186)
--	g5895 = NOT(g255)
--	g5896 = NOT(g261)
--	g5897 = NOT(g267)
--	g5898 = NOT(g762)
--	g5899 = NOT(g809)
--	g5900 = NOT(g933)
--	g5901 = NOT(g939)
--	g5902 = NOT(g945)
--	I14357 = NOT(g785)
--	g5903 = NOT(I14357)
--	g5904 = NOT(g1224)
--	g5905 = NOT(g1457)
--	g5906 = NOT(g1496)
--	g5907 = NOT(g1618)
--	g5908 = NOT(g1624)
--	g5909 = NOT(g1630)
--	g5911 = NOT(g1889)
--	g5912 = NOT(g2160)
--	g5913 = NOT(g2120)
--	g5914 = NOT(g2185)
--	g5915 = NOT(g2303)
--	g5916 = NOT(g2309)
--	g5917 = NOT(g2315)
--	g5918 = NOT(g2379)
--	g5921 = NOT(g2582)
--	I14378 = NOT(g3234)
--	g5922 = NOT(I14378)
--	I14381 = NOT(g3223)
--	g5923 = NOT(I14381)
--	I14384 = NOT(g3218)
--	g5924 = NOT(I14384)
--	g5925 = NOT(g189)
--	g5926 = NOT(g195)
--	g5927 = NOT(g264)
--	g5928 = NOT(g270)
--	g5929 = NOT(g776)
--	g5932 = NOT(g813)
--	g5933 = NOT(g873)
--	g5934 = NOT(g942)
--	g5935 = NOT(g948)
--	g5936 = NOT(g954)
--	g5937 = NOT(g1448)
--	g5938 = NOT(g1501)
--	g5939 = NOT(g1627)
--	g5940 = NOT(g1633)
--	g5941 = NOT(g1639)
--	I14402 = NOT(g1471)
--	g5942 = NOT(I14402)
--	g5943 = NOT(g1918)
--	g5944 = NOT(g2151)
--	g5945 = NOT(g2190)
--	g5946 = NOT(g2312)
--	g5947 = NOT(g2318)
--	g5948 = NOT(g2324)
--	g5950 = NOT(g2583)
--	I14413 = NOT(g3233)
--	g5951 = NOT(I14413)
--	I14416 = NOT(g3222)
--	g5952 = NOT(I14416)
--	g5953 = NOT(g97)
--	g5954 = NOT(g192)
--	g5955 = NOT(g198)
--	g5956 = NOT(g204)
--	g5957 = NOT(g273)
--	I14424 = NOT(g117)
--	g5958 = NOT(I14424)
--	g5959 = NOT(g876)
--	g5960 = NOT(g882)
--	g5961 = NOT(g951)
--	g5962 = NOT(g957)
--	g5963 = NOT(g1462)
--	g5966 = NOT(g1506)
--	g5967 = NOT(g1567)
--	g5968 = NOT(g1636)
--	g5969 = NOT(g1642)
--	g5970 = NOT(g1648)
--	g5971 = NOT(g2142)
--	g5972 = NOT(g2195)
--	g5973 = NOT(g2321)
--	g5974 = NOT(g2327)
--	g5975 = NOT(g2333)
--	I14442 = NOT(g2165)
--	g5976 = NOT(I14442)
--	g5977 = NOT(g2612)
--	I14446 = NOT(g3230)
--	g5978 = NOT(I14446)
--	I14449 = NOT(g3224)
--	g5979 = NOT(I14449)
--	g5980 = NOT(g201)
--	g5981 = NOT(g207)
--	g5982 = NOT(g785)
--	g5983 = NOT(g879)
--	g5984 = NOT(g885)
--	g5985 = NOT(g891)
--	g5986 = NOT(g960)
--	I14459 = NOT(g805)
--	g5987 = NOT(I14459)
--	g5988 = NOT(g1570)
--	g5989 = NOT(g1576)
--	g5990 = NOT(g1645)
--	g5991 = NOT(g1651)
--	g5992 = NOT(g2156)
--	g5995 = NOT(g2200)
--	g5996 = NOT(g2261)
--	g5997 = NOT(g2330)
--	g5998 = NOT(g2336)
--	g5999 = NOT(g2342)
--	I14472 = NOT(g3080)
--	g6000 = NOT(I14472)
--	I14475 = NOT(g3225)
--	g6014 = NOT(I14475)
--	I14478 = NOT(g3213)
--	g6015 = NOT(I14478)
--	g6016 = NOT(g210)
--	g6017 = NOT(g888)
--	g6018 = NOT(g894)
--	g6019 = NOT(g1471)
--	g6020 = NOT(g1573)
--	g6021 = NOT(g1579)
--	g6022 = NOT(g1585)
--	g6023 = NOT(g1654)
--	I14489 = NOT(g1496)
--	g6024 = NOT(I14489)
--	g6025 = NOT(g2264)
--	g6026 = NOT(g2270)
--	g6027 = NOT(g2339)
--	g6028 = NOT(g2345)
--	I14496 = NOT(g3226)
--	g6029 = NOT(I14496)
--	I14499 = NOT(g3214)
--	g6030 = NOT(I14499)
--	I14502 = NOT(g471)
--	g6031 = NOT(I14502)
--	g6032 = NOT(g897)
--	g6033 = NOT(g1582)
--	g6034 = NOT(g1588)
--	g6035 = NOT(g2165)
--	g6036 = NOT(g2267)
--	g6037 = NOT(g2273)
--	g6038 = NOT(g2279)
--	g6039 = NOT(g2348)
--	I14513 = NOT(g2190)
--	g6040 = NOT(I14513)
--	I14516 = NOT(g3215)
--	g6041 = NOT(I14516)
--	I14519 = NOT(g1158)
--	g6042 = NOT(I14519)
--	g6043 = NOT(g1591)
--	g6044 = NOT(g2276)
--	g6045 = NOT(g2282)
--	I14525 = NOT(g1852)
--	g6046 = NOT(I14525)
--	g6047 = NOT(g2285)
--	I14529 = NOT(g3142)
--	g6048 = NOT(I14529)
--	I14532 = NOT(g354)
--	g6051 = NOT(I14532)
--	I14535 = NOT(g2546)
--	g6052 = NOT(I14535)
--	I14538 = NOT(g369)
--	g6053 = NOT(I14538)
--	I14541 = NOT(g455)
--	g6054 = NOT(I14541)
--	I14544 = NOT(g1041)
--	g6055 = NOT(I14544)
--	I14547 = NOT(g384)
--	g6056 = NOT(I14547)
--	I14550 = NOT(g458)
--	g6057 = NOT(I14550)
--	I14553 = NOT(g1056)
--	g6058 = NOT(I14553)
--	I14556 = NOT(g1142)
--	g6059 = NOT(I14556)
--	I14559 = NOT(g1735)
--	g6060 = NOT(I14559)
--	I14562 = NOT(g398)
--	g6061 = NOT(I14562)
--	I14565 = NOT(g461)
--	g6062 = NOT(I14565)
--	I14568 = NOT(g1071)
--	g6063 = NOT(I14568)
--	I14571 = NOT(g1145)
--	g6064 = NOT(I14571)
--	I14574 = NOT(g1750)
--	g6065 = NOT(I14574)
--	I14577 = NOT(g1836)
--	g6066 = NOT(I14577)
--	I14580 = NOT(g2429)
--	g6067 = NOT(I14580)
--	g6068 = NOT(g499)
--	I14584 = NOT(g465)
--	g6079 = NOT(I14584)
--	I14587 = NOT(g1085)
--	g6080 = NOT(I14587)
--	I14590 = NOT(g1148)
--	g6081 = NOT(I14590)
--	I14593 = NOT(g1765)
--	g6082 = NOT(I14593)
--	I14596 = NOT(g1839)
--	g6083 = NOT(I14596)
--	I14599 = NOT(g2444)
--	g6084 = NOT(I14599)
--	I14602 = NOT(g2530)
--	g6085 = NOT(I14602)
--	I14605 = NOT(g468)
--	g6086 = NOT(I14605)
--	g6087 = NOT(g1186)
--	I14609 = NOT(g1152)
--	g6098 = NOT(I14609)
--	I14612 = NOT(g1779)
--	g6099 = NOT(I14612)
--	I14615 = NOT(g1842)
--	g6100 = NOT(I14615)
--	I14618 = NOT(g2459)
--	g6101 = NOT(I14618)
--	I14621 = NOT(g2533)
--	g6102 = NOT(I14621)
--	I14624 = NOT(g1155)
--	g6103 = NOT(I14624)
--	g6104 = NOT(g1880)
--	I14628 = NOT(g1846)
--	g6115 = NOT(I14628)
--	I14631 = NOT(g2473)
--	g6116 = NOT(I14631)
--	I14634 = NOT(g2536)
--	g6117 = NOT(I14634)
--	I14637 = NOT(g1849)
--	g6118 = NOT(I14637)
--	g6119 = NOT(g2574)
--	I14641 = NOT(g2540)
--	g6130 = NOT(I14641)
--	I14644 = NOT(g3142)
--	g6131 = NOT(I14644)
--	I14647 = NOT(g2543)
--	g6134 = NOT(I14647)
--	I14650 = NOT(g525)
--	g6135 = NOT(I14650)
--	g6136 = NOT(g672)
--	I14654 = NOT(g3220)
--	g6139 = NOT(I14654)
--	g6140 = NOT(g524)
--	g6141 = NOT(g554)
--	g6142 = NOT(g679)
--	I14660 = NOT(g1211)
--	g6145 = NOT(I14660)
--	g6146 = NOT(g1358)
--	g6149 = NOT(g3097)
--	I14665 = NOT(g3147)
--	g6153 = NOT(I14665)
--	I14668 = NOT(g3232)
--	g6156 = NOT(I14668)
--	g6157 = NOT(g686)
--	g6161 = NOT(g1210)
--	g6162 = NOT(g1240)
--	g6163 = NOT(g1365)
--	I14675 = NOT(g1905)
--	g6166 = NOT(I14675)
--	g6167 = NOT(g2052)
--	g6170 = NOT(g3098)
--	g6173 = NOT(g557)
--	g6177 = NOT(g633)
--	g6180 = NOT(g692)
--	g6183 = NOT(g291)
--	g6184 = NOT(g1372)
--	g6188 = NOT(g1904)
--	g6189 = NOT(g1934)
--	g6190 = NOT(g2059)
--	I14688 = NOT(g2599)
--	g6193 = NOT(I14688)
--	g6194 = NOT(g2746)
--	g6197 = NOT(g3099)
--	g6200 = NOT(g542)
--	g6201 = NOT(g646)
--	g6204 = NOT(g289)
--	g6205 = NOT(g1243)
--	g6209 = NOT(g1319)
--	g6212 = NOT(g1378)
--	g6215 = NOT(g978)
--	g6216 = NOT(g2066)
--	g6220 = NOT(g2598)
--	g6221 = NOT(g2628)
--	g6222 = NOT(g2753)
--	I14704 = NOT(g2818)
--	g6225 = NOT(I14704)
--	g6226 = NOT(g2818)
--	g6227 = NOT(g3100)
--	I14709 = NOT(g3229)
--	g6230 = NOT(I14709)
--	I14712 = NOT(g138)
--	g6231 = NOT(I14712)
--	I14715 = NOT(g138)
--	g6232 = NOT(I14715)
--	g6281 = NOT(g510)
--	g6284 = NOT(g640)
--	g6288 = NOT(g287)
--	g6289 = NOT(g1228)
--	g6290 = NOT(g1332)
--	g6293 = NOT(g976)
--	g6294 = NOT(g1937)
--	g6298 = NOT(g2013)
--	g6301 = NOT(g2072)
--	g6304 = NOT(g1672)
--	g6305 = NOT(g2760)
--	g6309 = NOT(g14)
--	g6310 = NOT(g3101)
--	I14731 = NOT(g135)
--	g6313 = NOT(I14731)
--	I14734 = NOT(g135)
--	g6314 = NOT(I14734)
--	g6363 = NOT(g653)
--	g6367 = NOT(g285)
--	I14739 = NOT(g826)
--	g6368 = NOT(I14739)
--	I14742 = NOT(g826)
--	g6369 = NOT(I14742)
--	g6418 = NOT(g1196)
--	g6421 = NOT(g1326)
--	g6425 = NOT(g974)
--	g6426 = NOT(g1922)
--	g6427 = NOT(g2026)
--	g6430 = NOT(g1670)
--	g6431 = NOT(g2631)
--	g6435 = NOT(g2707)
--	g6438 = NOT(g2766)
--	g6441 = NOT(g2366)
--	I14755 = NOT(g2821)
--	g6442 = NOT(I14755)
--	g6443 = NOT(g2821)
--	g6444 = NOT(g3102)
--	I14760 = NOT(g405)
--	g6447 = NOT(I14760)
--	I14763 = NOT(g405)
--	g6448 = NOT(I14763)
--	I14766 = NOT(g545)
--	g6485 = NOT(I14766)
--	I14769 = NOT(g545)
--	g6486 = NOT(I14769)
--	g6512 = NOT(g544)
--	g6513 = NOT(g660)
--	g6517 = NOT(g283)
--	I14775 = NOT(g823)
--	g6518 = NOT(I14775)
--	I14778 = NOT(g823)
--	g6519 = NOT(I14778)
--	g6568 = NOT(g1339)
--	g6572 = NOT(g972)
--	I14783 = NOT(g1520)
--	g6573 = NOT(I14783)
--	I14786 = NOT(g1520)
--	g6574 = NOT(I14786)
--	g6623 = NOT(g1890)
--	g6626 = NOT(g2020)
--	g6630 = NOT(g1668)
--	g6631 = NOT(g2616)
--	g6632 = NOT(g2720)
--	g6635 = NOT(g2364)
--	g6636 = NOT(g1491)
--	g6637 = NOT(g5)
--	g6638 = NOT(g3103)
--	g6641 = NOT(g113)
--	I14799 = NOT(g551)
--	g6642 = NOT(I14799)
--	I14802 = NOT(g551)
--	g6643 = NOT(I14802)
--	g6672 = NOT(g464)
--	g6675 = NOT(g458)
--	g6676 = NOT(g559)
--	I14808 = NOT(g623)
--	g6677 = NOT(I14808)
--	I14811 = NOT(g623)
--	g6678 = NOT(I14811)
--	g6707 = NOT(g666)
--	g6711 = NOT(g281)
--	I14816 = NOT(g1092)
--	g6712 = NOT(I14816)
--	I14819 = NOT(g1092)
--	g6713 = NOT(I14819)
--	I14822 = NOT(g1231)
--	g6750 = NOT(I14822)
--	I14825 = NOT(g1231)
--	g6751 = NOT(I14825)
--	g6776 = NOT(g1230)
--	g6777 = NOT(g1346)
--	g6781 = NOT(g970)
--	I14831 = NOT(g1517)
--	g6782 = NOT(I14831)
--	I14834 = NOT(g1517)
--	g6783 = NOT(I14834)
--	g6832 = NOT(g2033)
--	g6836 = NOT(g1666)
--	I14839 = NOT(g2214)
--	g6837 = NOT(I14839)
--	I14842 = NOT(g2214)
--	g6838 = NOT(I14842)
--	g6887 = NOT(g2584)
--	g6890 = NOT(g2714)
--	g6894 = NOT(g2362)
--	I14848 = NOT(g2824)
--	g6895 = NOT(I14848)
--	g6896 = NOT(g2824)
--	g6897 = NOT(g1486)
--	g6898 = NOT(g2993)
--	g6901 = NOT(g3006)
--	g6905 = NOT(g3104)
--	g6908 = NOT(g484)
--	I14857 = NOT(g626)
--	g6911 = NOT(I14857)
--	I14860 = NOT(g626)
--	g6912 = NOT(I14860)
--	g6942 = NOT(g279)
--	g6943 = NOT(g801)
--	I14865 = NOT(g1237)
--	g6944 = NOT(I14865)
--	I14868 = NOT(g1237)
--	g6945 = NOT(I14868)
--	g6974 = NOT(g1151)
--	g6977 = NOT(g1145)
--	g6978 = NOT(g1245)
--	I14874 = NOT(g1309)
--	g6979 = NOT(I14874)
--	I14877 = NOT(g1309)
--	g6980 = NOT(I14877)
--	g7009 = NOT(g1352)
--	g7013 = NOT(g968)
--	I14882 = NOT(g1786)
--	g7014 = NOT(I14882)
--	I14885 = NOT(g1786)
--	g7015 = NOT(I14885)
--	I14888 = NOT(g1925)
--	g7052 = NOT(I14888)
--	I14891 = NOT(g1925)
--	g7053 = NOT(I14891)
--	g7078 = NOT(g1924)
--	g7079 = NOT(g2040)
--	g7083 = NOT(g1664)
--	I14897 = NOT(g2211)
--	g7084 = NOT(I14897)
--	I14900 = NOT(g2211)
--	g7085 = NOT(I14900)
--	g7134 = NOT(g2727)
--	g7138 = NOT(g2360)
--	g7139 = NOT(g1481)
--	g7140 = NOT(g2170)
--	g7141 = NOT(g2195)
--	g7142 = NOT(g8)
--	g7143 = NOT(g2998)
--	g7146 = NOT(g3013)
--	g7149 = NOT(g3105)
--	g7152 = NOT(g3136)
--	g7153 = NOT(g480)
--	g7156 = NOT(g461)
--	g7157 = NOT(g453)
--	g7158 = NOT(g1171)
--	I14917 = NOT(g1312)
--	g7161 = NOT(I14917)
--	I14920 = NOT(g1312)
--	g7162 = NOT(I14920)
--	g7192 = NOT(g966)
--	g7193 = NOT(g1491)
--	I14925 = NOT(g1931)
--	g7194 = NOT(I14925)
--	I14928 = NOT(g1931)
--	g7195 = NOT(I14928)
--	g7224 = NOT(g1845)
--	g7227 = NOT(g1839)
--	g7228 = NOT(g1939)
--	I14934 = NOT(g2003)
--	g7229 = NOT(I14934)
--	I14937 = NOT(g2003)
--	g7230 = NOT(I14937)
--	g7259 = NOT(g2046)
--	g7263 = NOT(g1662)
--	I14942 = NOT(g2480)
--	g7264 = NOT(I14942)
--	I14945 = NOT(g2480)
--	g7265 = NOT(I14945)
--	I14948 = NOT(g2619)
--	g7302 = NOT(I14948)
--	I14951 = NOT(g2619)
--	g7303 = NOT(I14951)
--	g7328 = NOT(g2618)
--	g7329 = NOT(g2734)
--	g7333 = NOT(g2358)
--	I14957 = NOT(g2827)
--	g7334 = NOT(I14957)
--	g7335 = NOT(g2827)
--	g7336 = NOT(g1476)
--	g7337 = NOT(g2190)
--	g7338 = NOT(g3002)
--	g7342 = NOT(g3024)
--	g7345 = NOT(g3139)
--	g7346 = NOT(g97)
--	g7347 = NOT(g490)
--	g7348 = NOT(g451)
--	g7349 = NOT(g1167)
--	g7352 = NOT(g1148)
--	g7353 = NOT(g1140)
--	g7354 = NOT(g1865)
--	I14973 = NOT(g2006)
--	g7357 = NOT(I14973)
--	I14976 = NOT(g2006)
--	g7358 = NOT(I14976)
--	g7388 = NOT(g1660)
--	g7389 = NOT(g2185)
--	I14981 = NOT(g2625)
--	g7390 = NOT(I14981)
--	I14984 = NOT(g2625)
--	g7391 = NOT(I14984)
--	g7420 = NOT(g2539)
--	g7423 = NOT(g2533)
--	g7424 = NOT(g2633)
--	I14990 = NOT(g2697)
--	g7425 = NOT(I14990)
--	I14993 = NOT(g2697)
--	g7426 = NOT(I14993)
--	g7455 = NOT(g2740)
--	g7459 = NOT(g2356)
--	g7460 = NOT(g1471)
--	g7461 = NOT(g2175)
--	g7462 = NOT(g2912)
--	g7465 = NOT(g2)
--	g7466 = NOT(g3010)
--	g7471 = NOT(g3036)
--	g7475 = NOT(g493)
--	g7476 = NOT(g785)
--	g7477 = NOT(g1177)
--	g7478 = NOT(g1138)
--	g7479 = NOT(g1861)
--	g7482 = NOT(g1842)
--	g7483 = NOT(g1834)
--	g7484 = NOT(g2559)
--	I15012 = NOT(g2700)
--	g7487 = NOT(I15012)
--	I15015 = NOT(g2700)
--	g7488 = NOT(I15015)
--	g7518 = NOT(g2354)
--	I15019 = NOT(g2830)
--	g7519 = NOT(I15019)
--	g7520 = NOT(g2830)
--	g7521 = NOT(g2200)
--	g7522 = NOT(g2917)
--	g7527 = NOT(g3018)
--	g7529 = NOT(g465)
--	g7530 = NOT(g496)
--	g7531 = NOT(g1180)
--	g7532 = NOT(g1471)
--	g7533 = NOT(g1871)
--	g7534 = NOT(g1832)
--	g7535 = NOT(g2555)
--	g7538 = NOT(g2536)
--	g7539 = NOT(g2528)
--	g7540 = NOT(g1506)
--	g7541 = NOT(g2180)
--	g7542 = NOT(g2883)
--	g7545 = NOT(g2920)
--	g7548 = NOT(g2990)
--	g7549 = NOT(g3028)
--	g7553 = NOT(g3114)
--	g7554 = NOT(g117)
--	g7555 = NOT(g1152)
--	g7556 = NOT(g1183)
--	g7557 = NOT(g1874)
--	g7558 = NOT(g2165)
--	g7559 = NOT(g2565)
--	g7560 = NOT(g2526)
--	g7561 = NOT(g1501)
--	g7562 = NOT(g2888)
--	g7566 = NOT(g2896)
--	g7570 = NOT(g3032)
--	g7573 = NOT(g3120)
--	g7574 = NOT(g3128)
--	g7576 = NOT(g468)
--	g7577 = NOT(g805)
--	g7578 = NOT(g1846)
--	g7579 = NOT(g1877)
--	g7580 = NOT(g2568)
--	g7581 = NOT(g1496)
--	g7582 = NOT(g2185)
--	g7583 = NOT(g2892)
--	g7587 = NOT(g2903)
--	g7590 = NOT(g1155)
--	g7591 = NOT(g1496)
--	g7592 = NOT(g2540)
--	g7593 = NOT(g2571)
--	g7594 = NOT(g2165)
--	g7595 = NOT(g2900)
--	g7600 = NOT(g2908)
--	g7603 = NOT(g3133)
--	g7604 = NOT(g471)
--	g7605 = NOT(g1849)
--	g7606 = NOT(g2190)
--	g7607 = NOT(g2924)
--	g7610 = NOT(g312)
--	g7613 = NOT(g1158)
--	g7614 = NOT(g2543)
--	g7615 = NOT(g3123)
--	g7616 = NOT(g313)
--	g7619 = NOT(g999)
--	g7622 = NOT(g1852)
--	g7623 = NOT(g314)
--	g7626 = NOT(g315)
--	g7629 = NOT(g403)
--	g7632 = NOT(g1000)
--	g7635 = NOT(g1693)
--	g7638 = NOT(g2546)
--	g7639 = NOT(g3094)
--	g7642 = NOT(g3125)
--	g7643 = NOT(g316)
--	g7646 = NOT(g318)
--	g7649 = NOT(g404)
--	g7652 = NOT(g1001)
--	g7655 = NOT(g1002)
--	g7658 = NOT(g1090)
--	g7661 = NOT(g1694)
--	g7664 = NOT(g2387)
--	g7667 = NOT(g3095)
--	g7670 = NOT(g317)
--	g7673 = NOT(g319)
--	g7676 = NOT(g402)
--	g7679 = NOT(g1003)
--	g7682 = NOT(g1005)
--	g7685 = NOT(g1091)
--	g7688 = NOT(g1695)
--	g7691 = NOT(g1696)
--	g7694 = NOT(g1784)
--	g7697 = NOT(g2388)
--	g7700 = NOT(g3096)
--	g7703 = NOT(g320)
--	g7706 = NOT(g1004)
--	g7709 = NOT(g1006)
--	g7712 = NOT(g1089)
--	g7715 = NOT(g1697)
--	g7718 = NOT(g1699)
--	g7721 = NOT(g1785)
--	g7724 = NOT(g2389)
--	g7727 = NOT(g2390)
--	g7730 = NOT(g2478)
--	g7733 = NOT(g1007)
--	g7736 = NOT(g1698)
--	g7739 = NOT(g1700)
--	g7742 = NOT(g1783)
--	g7745 = NOT(g2391)
--	g7748 = NOT(g2393)
--	g7751 = NOT(g2479)
--	g7754 = NOT(g322)
--	g7757 = NOT(g1701)
--	g7760 = NOT(g2392)
--	g7763 = NOT(g2394)
--	g7766 = NOT(g2477)
--	g7769 = NOT(g323)
--	g7772 = NOT(g659)
--	g7776 = NOT(g1009)
--	g7779 = NOT(g2395)
--	g7782 = NOT(g321)
--	g7785 = NOT(g1010)
--	g7788 = NOT(g1345)
--	g7792 = NOT(g1703)
--	g7796 = NOT(g1008)
--	g7799 = NOT(g1704)
--	g7802 = NOT(g2039)
--	g7806 = NOT(g2397)
--	g7809 = NOT(g1702)
--	g7812 = NOT(g2398)
--	g7815 = NOT(g2733)
--	g7819 = NOT(g479)
--	g7822 = NOT(g510)
--	g7823 = NOT(g2396)
--	g7826 = NOT(g2987)
--	g7827 = NOT(g478)
--	g7830 = NOT(g1166)
--	g7833 = NOT(g1196)
--	g7834 = NOT(g2953)
--	g7837 = NOT(g3044)
--	g7838 = NOT(g477)
--	g7841 = NOT(g630)
--	g7842 = NOT(g1165)
--	g7845 = NOT(g1860)
--	g7848 = NOT(g1890)
--	g7849 = NOT(g2956)
--	g7852 = NOT(g2981)
--	g7856 = NOT(g3045)
--	g7857 = NOT(g3055)
--	g7858 = NOT(g1164)
--	g7861 = NOT(g1316)
--	g7862 = NOT(g1859)
--	g7865 = NOT(g2554)
--	g7868 = NOT(g2584)
--	g7869 = NOT(g2959)
--	g7872 = NOT(g2874)
--	g7877 = NOT(g3046)
--	g7878 = NOT(g3056)
--	g7879 = NOT(g3065)
--	g7880 = NOT(g3201)
--	g7888 = NOT(g1858)
--	g7891 = NOT(g2010)
--	g7892 = NOT(g2553)
--	g7897 = NOT(g3047)
--	g7898 = NOT(g3057)
--	g7899 = NOT(g3066)
--	g7900 = NOT(g3075)
--	I15222 = NOT(g3151)
--	g7901 = NOT(I15222)
--	g7906 = NOT(g488)
--	I15226 = NOT(g474)
--	g7909 = NOT(I15226)
--	g7910 = NOT(g474)
--	I15230 = NOT(g499)
--	g7911 = NOT(I15230)
--	g7912 = NOT(g2552)
--	g7915 = NOT(g2704)
--	g7916 = NOT(g2935)
--	g7919 = NOT(g2963)
--	g7924 = NOT(g3048)
--	g7925 = NOT(g3058)
--	g7926 = NOT(g3067)
--	g7927 = NOT(g3076)
--	g7928 = NOT(g3204)
--	I15256 = NOT(g2950)
--	g7936 = NOT(I15256)
--	g7949 = NOT(g165)
--	g7950 = NOT(g142)
--	g7953 = NOT(g487)
--	I15262 = NOT(g481)
--	g7956 = NOT(I15262)
--	g7957 = NOT(g481)
--	g7958 = NOT(g1175)
--	I15267 = NOT(g1161)
--	g7961 = NOT(I15267)
--	g7962 = NOT(g1161)
--	I15271 = NOT(g1186)
--	g7963 = NOT(I15271)
--	g7964 = NOT(g2938)
--	g7967 = NOT(g2966)
--	g7971 = NOT(g3049)
--	g7972 = NOT(g3059)
--	g7973 = NOT(g3068)
--	g7974 = NOT(g3077)
--	g7975 = NOT(g39)
--	I15288 = NOT(g3109)
--	g7976 = NOT(I15288)
--	g7989 = NOT(g3191)
--	g7990 = NOT(g143)
--	g7993 = NOT(g145)
--	g7996 = NOT(g486)
--	g7999 = NOT(g485)
--	g8000 = NOT(g853)
--	g8001 = NOT(g830)
--	g8004 = NOT(g1174)
--	I15299 = NOT(g1168)
--	g8007 = NOT(I15299)
--	g8008 = NOT(g1168)
--	g8009 = NOT(g1869)
--	I15304 = NOT(g1855)
--	g8012 = NOT(I15304)
--	g8013 = NOT(g1855)
--	I15308 = NOT(g1880)
--	g8014 = NOT(I15308)
--	g8015 = NOT(g2941)
--	g8018 = NOT(g2969)
--	I15313 = NOT(g2930)
--	g8021 = NOT(I15313)
--	g8022 = NOT(g2930)
--	I15317 = NOT(g2842)
--	g8023 = NOT(I15317)
--	g8024 = NOT(g2842)
--	g8025 = NOT(g3050)
--	g8026 = NOT(g3060)
--	g8027 = NOT(g3069)
--	g8028 = NOT(g3078)
--	g8029 = NOT(g3083)
--	I15326 = NOT(g3117)
--	g8030 = NOT(I15326)
--	I15329 = NOT(g3117)
--	g8031 = NOT(I15329)
--	g8044 = NOT(g3194)
--	g8045 = NOT(g3207)
--	g8053 = NOT(g141)
--	g8056 = NOT(g146)
--	g8059 = NOT(g148)
--	g8062 = NOT(g169)
--	g8065 = NOT(g831)
--	g8068 = NOT(g833)
--	g8071 = NOT(g1173)
--	g8074 = NOT(g1172)
--	g8075 = NOT(g1547)
--	g8076 = NOT(g1524)
--	g8079 = NOT(g1868)
--	I15345 = NOT(g1862)
--	g8082 = NOT(I15345)
--	g8083 = NOT(g1862)
--	g8084 = NOT(g2563)
--	I15350 = NOT(g2549)
--	g8087 = NOT(I15350)
--	g8088 = NOT(g2549)
--	I15354 = NOT(g2574)
--	g8089 = NOT(I15354)
--	g8090 = NOT(g2944)
--	g8093 = NOT(g2972)
--	I15359 = NOT(g2858)
--	g8096 = NOT(I15359)
--	g8097 = NOT(g2858)
--	g8098 = NOT(g3051)
--	g8099 = NOT(g3061)
--	g8100 = NOT(g3070)
--	g8101 = NOT(g2997)
--	g8102 = NOT(g27)
--	g8103 = NOT(g185)
--	I15369 = NOT(g3129)
--	g8106 = NOT(I15369)
--	I15372 = NOT(g3129)
--	g8107 = NOT(I15372)
--	g8120 = NOT(g3197)
--	g8123 = NOT(g144)
--	g8126 = NOT(g149)
--	g8129 = NOT(g151)
--	g8132 = NOT(g170)
--	g8135 = NOT(g172)
--	g8138 = NOT(g829)
--	g8141 = NOT(g834)
--	g8144 = NOT(g836)
--	g8147 = NOT(g857)
--	g8150 = NOT(g1525)
--	g8153 = NOT(g1527)
--	g8156 = NOT(g1867)
--	g8159 = NOT(g1866)
--	g8160 = NOT(g2241)
--	g8161 = NOT(g2218)
--	g8164 = NOT(g2562)
--	I15392 = NOT(g2556)
--	g8167 = NOT(I15392)
--	g8168 = NOT(g2556)
--	g8169 = NOT(g2947)
--	g8172 = NOT(g2975)
--	I15398 = NOT(g2845)
--	g8175 = NOT(I15398)
--	g8176 = NOT(g2845)
--	g8177 = NOT(g3043)
--	g8178 = NOT(g3052)
--	g8179 = NOT(g3062)
--	g8180 = NOT(g3071)
--	g8181 = NOT(g48)
--	g8182 = NOT(g3198)
--	g8183 = NOT(g3188)
--	g8191 = NOT(g147)
--	g8194 = NOT(g152)
--	g8197 = NOT(g154)
--	g8200 = NOT(g168)
--	g8203 = NOT(g173)
--	g8206 = NOT(g175)
--	g8209 = NOT(g832)
--	g8212 = NOT(g837)
--	g8215 = NOT(g839)
--	g8218 = NOT(g858)
--	g8221 = NOT(g860)
--	g8224 = NOT(g1523)
--	g8227 = NOT(g1528)
--	g8230 = NOT(g1530)
--	g8233 = NOT(g1551)
--	g8236 = NOT(g2219)
--	g8239 = NOT(g2221)
--	g8242 = NOT(g2561)
--	g8245 = NOT(g2560)
--	g8246 = NOT(g2978)
--	I15429 = NOT(g2833)
--	g8249 = NOT(I15429)
--	g8250 = NOT(g2833)
--	I15433 = NOT(g2861)
--	g8251 = NOT(I15433)
--	g8252 = NOT(g2861)
--	g8253 = NOT(g3053)
--	g8254 = NOT(g3063)
--	g8255 = NOT(g3072)
--	g8256 = NOT(g30)
--	g8257 = NOT(g3201)
--	I15442 = NOT(g3235)
--	g8258 = NOT(I15442)
--	I15445 = NOT(g3236)
--	g8259 = NOT(I15445)
--	I15448 = NOT(g3237)
--	g8260 = NOT(I15448)
--	I15451 = NOT(g3238)
--	g8261 = NOT(I15451)
--	I15454 = NOT(g3239)
--	g8262 = NOT(I15454)
--	I15457 = NOT(g3240)
--	g8263 = NOT(I15457)
--	I15460 = NOT(g3241)
--	g8264 = NOT(I15460)
--	I15463 = NOT(g3242)
--	g8265 = NOT(I15463)
--	I15466 = NOT(g3243)
--	g8266 = NOT(I15466)
--	I15469 = NOT(g3244)
--	g8267 = NOT(I15469)
--	I15472 = NOT(g3245)
--	g8268 = NOT(I15472)
--	I15475 = NOT(g3246)
--	g8269 = NOT(I15475)
--	I15478 = NOT(g3247)
--	g8270 = NOT(I15478)
--	I15481 = NOT(g3248)
--	g8271 = NOT(I15481)
--	I15484 = NOT(g3249)
--	g8272 = NOT(I15484)
--	I15487 = NOT(g3250)
--	g8273 = NOT(I15487)
--	I15490 = NOT(g3251)
--	g8274 = NOT(I15490)
--	I15493 = NOT(g3252)
--	g8275 = NOT(I15493)
--	g8276 = NOT(g3253)
--	g8277 = NOT(g3305)
--	g8278 = NOT(g3337)
--	I15499 = NOT(g7911)
--	g8284 = NOT(I15499)
--	g8285 = NOT(g3365)
--	g8286 = NOT(g3461)
--	g8287 = NOT(g3493)
--	I15505 = NOT(g7963)
--	g8293 = NOT(I15505)
--	g8294 = NOT(g3521)
--	g8295 = NOT(g3617)
--	g8296 = NOT(g3649)
--	I15511 = NOT(g8014)
--	g8302 = NOT(I15511)
--	g8303 = NOT(g3677)
--	g8304 = NOT(g3773)
--	g8305 = NOT(g3805)
--	I15517 = NOT(g8089)
--	g8311 = NOT(I15517)
--	g8312 = NOT(g3833)
--	g8313 = NOT(g3897)
--	g8317 = NOT(g3919)
--	I15523 = NOT(g3254)
--	g8321 = NOT(I15523)
--	I15526 = NOT(g6314)
--	g8324 = NOT(I15526)
--	I15532 = NOT(g3410)
--	g8330 = NOT(I15532)
--	I15535 = NOT(g6519)
--	g8333 = NOT(I15535)
--	I15538 = NOT(g6369)
--	g8336 = NOT(I15538)
--	I15543 = NOT(g3410)
--	g8341 = NOT(I15543)
--	I15546 = NOT(g6783)
--	g8344 = NOT(I15546)
--	I15549 = NOT(g6574)
--	g8347 = NOT(I15549)
--	I15553 = NOT(g3566)
--	g8351 = NOT(I15553)
--	I15556 = NOT(g6783)
--	g8354 = NOT(I15556)
--	I15559 = NOT(g7015)
--	g8357 = NOT(I15559)
--	I15562 = NOT(g5778)
--	g8360 = NOT(I15562)
--	I15565 = NOT(g6838)
--	g8363 = NOT(I15565)
--	I15568 = NOT(g3722)
--	g8366 = NOT(I15568)
--	I15571 = NOT(g7085)
--	g8369 = NOT(I15571)
--	I15574 = NOT(g6838)
--	g8372 = NOT(I15574)
--	I15577 = NOT(g7265)
--	g8375 = NOT(I15577)
--	I15580 = NOT(g5837)
--	g8378 = NOT(I15580)
--	I15584 = NOT(g3254)
--	g8382 = NOT(I15584)
--	I15590 = NOT(g3410)
--	g8388 = NOT(I15590)
--	I15593 = NOT(g6519)
--	g8391 = NOT(I15593)
--	I15599 = NOT(g3566)
--	g8397 = NOT(I15599)
--	I15602 = NOT(g6783)
--	g8400 = NOT(I15602)
--	I15605 = NOT(g6574)
--	g8403 = NOT(I15605)
--	I15610 = NOT(g3566)
--	g8408 = NOT(I15610)
--	I15613 = NOT(g7085)
--	g8411 = NOT(I15613)
--	I15616 = NOT(g6838)
--	g8414 = NOT(I15616)
--	I15620 = NOT(g3722)
--	g8418 = NOT(I15620)
--	I15623 = NOT(g7085)
--	g8421 = NOT(I15623)
--	I15626 = NOT(g7265)
--	g8424 = NOT(I15626)
--	I15629 = NOT(g5837)
--	g8427 = NOT(I15629)
--	I15636 = NOT(g3410)
--	g8434 = NOT(I15636)
--	I15642 = NOT(g3566)
--	g8440 = NOT(I15642)
--	I15645 = NOT(g6783)
--	g8443 = NOT(I15645)
--	I15651 = NOT(g3722)
--	g8449 = NOT(I15651)
--	I15654 = NOT(g7085)
--	g8452 = NOT(I15654)
--	I15657 = NOT(g6838)
--	g8455 = NOT(I15657)
--	I15662 = NOT(g3722)
--	g8460 = NOT(I15662)
--	I15671 = NOT(g3566)
--	g8469 = NOT(I15671)
--	I15677 = NOT(g3722)
--	g8475 = NOT(I15677)
--	I15680 = NOT(g7085)
--	g8478 = NOT(I15680)
--	I15696 = NOT(g3722)
--	g8494 = NOT(I15696)
--	g8514 = NOT(g6139)
--	g8530 = NOT(g6156)
--	g8568 = NOT(g6230)
--	I15771 = NOT(g6000)
--	g8569 = NOT(I15771)
--	I15779 = NOT(g6000)
--	g8575 = NOT(I15779)
--	I15784 = NOT(g6000)
--	g8578 = NOT(I15784)
--	I15787 = NOT(g6000)
--	g8579 = NOT(I15787)
--	g8580 = NOT(g6281)
--	g8587 = NOT(g6418)
--	g8594 = NOT(g6623)
--	I15794 = NOT(g3338)
--	g8602 = NOT(I15794)
--	g8605 = NOT(g6887)
--	I15800 = NOT(g3494)
--	g8614 = NOT(I15800)
--	I15803 = NOT(g8107)
--	g8617 = NOT(I15803)
--	I15806 = NOT(g5550)
--	g8620 = NOT(I15806)
--	I15810 = NOT(g3338)
--	g8622 = NOT(I15810)
--	I15815 = NOT(g3650)
--	g8627 = NOT(I15815)
--	I15818 = NOT(g5596)
--	g8630 = NOT(I15818)
--	I15822 = NOT(g3494)
--	g8632 = NOT(I15822)
--	I15827 = NOT(g3806)
--	g8637 = NOT(I15827)
--	I15830 = NOT(g8031)
--	g8640 = NOT(I15830)
--	I15833 = NOT(g3338)
--	g8643 = NOT(I15833)
--	I15836 = NOT(g3366)
--	g8646 = NOT(I15836)
--	I15839 = NOT(g5613)
--	g8649 = NOT(I15839)
--	I15843 = NOT(g3650)
--	g8651 = NOT(I15843)
--	I15847 = NOT(g3878)
--	g8655 = NOT(I15847)
--	I15850 = NOT(g5627)
--	g8658 = NOT(I15850)
--	I15853 = NOT(g3494)
--	g8659 = NOT(I15853)
--	I15856 = NOT(g3522)
--	g8662 = NOT(I15856)
--	I15859 = NOT(g5638)
--	g8665 = NOT(I15859)
--	I15863 = NOT(g3806)
--	g8667 = NOT(I15863)
--	I15866 = NOT(g3878)
--	g8670 = NOT(I15866)
--	I15869 = NOT(g7976)
--	g8673 = NOT(I15869)
--	I15873 = NOT(g5655)
--	g8677 = NOT(I15873)
--	I15876 = NOT(g3650)
--	g8678 = NOT(I15876)
--	I15879 = NOT(g3678)
--	g8681 = NOT(I15879)
--	I15882 = NOT(g3878)
--	g8684 = NOT(I15882)
--	I15887 = NOT(g5693)
--	g8689 = NOT(I15887)
--	I15890 = NOT(g3806)
--	g8690 = NOT(I15890)
--	I15893 = NOT(g3834)
--	g8693 = NOT(I15893)
--	I15896 = NOT(g3878)
--	g8696 = NOT(I15896)
--	I15899 = NOT(g5626)
--	g8699 = NOT(I15899)
--	I15902 = NOT(g6486)
--	g8700 = NOT(I15902)
--	I15909 = NOT(g5745)
--	g8707 = NOT(I15909)
--	I15912 = NOT(g3878)
--	g8708 = NOT(I15912)
--	I15915 = NOT(g3878)
--	g8711 = NOT(I15915)
--	I15918 = NOT(g6643)
--	g8714 = NOT(I15918)
--	I15922 = NOT(g5654)
--	g8718 = NOT(I15922)
--	I15925 = NOT(g6751)
--	g8719 = NOT(I15925)
--	I15932 = NOT(g5423)
--	g8726 = NOT(I15932)
--	I15935 = NOT(g3878)
--	g8745 = NOT(I15935)
--	I15938 = NOT(g3338)
--	g8748 = NOT(I15938)
--	I15942 = NOT(g6945)
--	g8752 = NOT(I15942)
--	I15946 = NOT(g5692)
--	g8756 = NOT(I15946)
--	I15949 = NOT(g7053)
--	g8757 = NOT(I15949)
--	I15955 = NOT(g3878)
--	g8763 = NOT(I15955)
--	I15958 = NOT(g3878)
--	g8766 = NOT(I15958)
--	I15961 = NOT(g6051)
--	g8769 = NOT(I15961)
--	I15964 = NOT(g7554)
--	g8770 = NOT(I15964)
--	I15967 = NOT(g3494)
--	g8771 = NOT(I15967)
--	I15971 = NOT(g7195)
--	g8775 = NOT(I15971)
--	I15975 = NOT(g5744)
--	g8779 = NOT(I15975)
--	I15978 = NOT(g7303)
--	g8780 = NOT(I15978)
--	I15983 = NOT(g3878)
--	g8785 = NOT(I15983)
--	I15986 = NOT(g3878)
--	g8788 = NOT(I15986)
--	I15989 = NOT(g6053)
--	g8791 = NOT(I15989)
--	I15992 = NOT(g6055)
--	g8792 = NOT(I15992)
--	I15995 = NOT(g7577)
--	g8793 = NOT(I15995)
--	I15998 = NOT(g3650)
--	g8794 = NOT(I15998)
--	I16002 = NOT(g7391)
--	g8798 = NOT(I16002)
--	I16006 = NOT(g3878)
--	g8802 = NOT(I16006)
--	I16009 = NOT(g3878)
--	g8805 = NOT(I16009)
--	I16012 = NOT(g5390)
--	g8808 = NOT(I16012)
--	I16015 = NOT(g6056)
--	g8809 = NOT(I16015)
--	I16018 = NOT(g6058)
--	g8810 = NOT(I16018)
--	I16021 = NOT(g6060)
--	g8811 = NOT(I16021)
--	I16024 = NOT(g7591)
--	g8812 = NOT(I16024)
--	I16027 = NOT(g3806)
--	g8813 = NOT(I16027)
--	I16031 = NOT(g3878)
--	g8817 = NOT(I16031)
--	I16034 = NOT(g5396)
--	g8820 = NOT(I16034)
--	I16037 = NOT(g6061)
--	g8821 = NOT(I16037)
--	g8822 = NOT(g4602)
--	I16041 = NOT(g6486)
--	g8823 = NOT(I16041)
--	I16044 = NOT(g5397)
--	g8824 = NOT(I16044)
--	I16047 = NOT(g6063)
--	g8825 = NOT(I16047)
--	I16050 = NOT(g6065)
--	g8826 = NOT(I16050)
--	I16053 = NOT(g6067)
--	g8827 = NOT(I16053)
--	I16056 = NOT(g7606)
--	g8828 = NOT(I16056)
--	I16059 = NOT(g3878)
--	g8829 = NOT(I16059)
--	I16062 = NOT(g3900)
--	g8832 = NOT(I16062)
--	I16065 = NOT(g7936)
--	g8835 = NOT(I16065)
--	I16068 = NOT(g5438)
--	g8836 = NOT(I16068)
--	I16071 = NOT(g5395)
--	g8839 = NOT(I16071)
--	I16074 = NOT(g5399)
--	g8840 = NOT(I16074)
--	I16079 = NOT(g6086)
--	g8843 = NOT(I16079)
--	I16082 = NOT(g5401)
--	g8844 = NOT(I16082)
--	I16085 = NOT(g6080)
--	g8845 = NOT(I16085)
--	g8846 = NOT(g4779)
--	I16089 = NOT(g6751)
--	g8847 = NOT(I16089)
--	I16092 = NOT(g5402)
--	g8850 = NOT(I16092)
--	I16095 = NOT(g6082)
--	g8851 = NOT(I16095)
--	I16098 = NOT(g6084)
--	g8852 = NOT(I16098)
--	I16101 = NOT(g3878)
--	g8853 = NOT(I16101)
--	I16104 = NOT(g6448)
--	g8856 = NOT(I16104)
--	I16107 = NOT(g5398)
--	g8859 = NOT(I16107)
--	I16110 = NOT(g5404)
--	g8860 = NOT(I16110)
--	I16114 = NOT(g7936)
--	g8862 = NOT(I16114)
--	I16117 = NOT(g5473)
--	g8863 = NOT(I16117)
--	I16120 = NOT(g5400)
--	g8866 = NOT(I16120)
--	I16123 = NOT(g5406)
--	g8867 = NOT(I16123)
--	I16128 = NOT(g6103)
--	g8870 = NOT(I16128)
--	I16131 = NOT(g5408)
--	g8871 = NOT(I16131)
--	I16134 = NOT(g6099)
--	g8872 = NOT(I16134)
--	g8873 = NOT(g4955)
--	I16138 = NOT(g7053)
--	g8874 = NOT(I16138)
--	I16141 = NOT(g5409)
--	g8877 = NOT(I16141)
--	I16144 = NOT(g6101)
--	g8878 = NOT(I16144)
--	I16147 = NOT(g3878)
--	g8879 = NOT(I16147)
--	I16150 = NOT(g3900)
--	g8882 = NOT(I16150)
--	I16153 = NOT(g3306)
--	g8885 = NOT(I16153)
--	I16156 = NOT(g5438)
--	g8888 = NOT(I16156)
--	I16159 = NOT(g5403)
--	g8891 = NOT(I16159)
--	I16163 = NOT(g6031)
--	g8893 = NOT(I16163)
--	I16166 = NOT(g6713)
--	g8894 = NOT(I16166)
--	I16169 = NOT(g5405)
--	g8897 = NOT(I16169)
--	I16172 = NOT(g5413)
--	g8898 = NOT(I16172)
--	I16176 = NOT(g7936)
--	g8900 = NOT(I16176)
--	I16179 = NOT(g5512)
--	g8901 = NOT(I16179)
--	I16182 = NOT(g5407)
--	g8904 = NOT(I16182)
--	I16185 = NOT(g5415)
--	g8905 = NOT(I16185)
--	I16190 = NOT(g6118)
--	g8908 = NOT(I16190)
--	I16193 = NOT(g5417)
--	g8909 = NOT(I16193)
--	I16196 = NOT(g6116)
--	g8910 = NOT(I16196)
--	g8911 = NOT(g5114)
--	I16200 = NOT(g7303)
--	g8912 = NOT(I16200)
--	I16203 = NOT(g3878)
--	g8915 = NOT(I16203)
--	I16206 = NOT(g6448)
--	g8918 = NOT(I16206)
--	I16209 = NOT(g5438)
--	g8921 = NOT(I16209)
--	I16212 = NOT(g5411)
--	g8924 = NOT(I16212)
--	I16215 = NOT(g3462)
--	g8925 = NOT(I16215)
--	I16218 = NOT(g5473)
--	g8928 = NOT(I16218)
--	I16221 = NOT(g5412)
--	g8931 = NOT(I16221)
--	I16225 = NOT(g6042)
--	g8933 = NOT(I16225)
--	I16228 = NOT(g7015)
--	g8934 = NOT(I16228)
--	I16231 = NOT(g5414)
--	g8937 = NOT(I16231)
--	I16234 = NOT(g5420)
--	g8938 = NOT(I16234)
--	I16238 = NOT(g7936)
--	g8940 = NOT(I16238)
--	I16241 = NOT(g5556)
--	g8941 = NOT(I16241)
--	I16244 = NOT(g5416)
--	g8944 = NOT(I16244)
--	I16247 = NOT(g5422)
--	g8945 = NOT(I16247)
--	I16252 = NOT(g6134)
--	g8948 = NOT(I16252)
--	I16255 = NOT(g3900)
--	g8949 = NOT(I16255)
--	I16258 = NOT(g3306)
--	g8952 = NOT(I16258)
--	I16261 = NOT(g6448)
--	g8955 = NOT(I16261)
--	I16264 = NOT(g6713)
--	g8958 = NOT(I16264)
--	I16267 = NOT(g5473)
--	g8961 = NOT(I16267)
--	I16270 = NOT(g5418)
--	g8964 = NOT(I16270)
--	I16273 = NOT(g3618)
--	g8965 = NOT(I16273)
--	I16276 = NOT(g5512)
--	g8968 = NOT(I16276)
--	I16279 = NOT(g5419)
--	g8971 = NOT(I16279)
--	I16283 = NOT(g6046)
--	g8973 = NOT(I16283)
--	I16286 = NOT(g7265)
--	g8974 = NOT(I16286)
--	I16289 = NOT(g5421)
--	g8977 = NOT(I16289)
--	I16292 = NOT(g5426)
--	g8978 = NOT(I16292)
--	I16296 = NOT(g3306)
--	g8980 = NOT(I16296)
--	g8983 = NOT(g6486)
--	I16300 = NOT(g3462)
--	g8984 = NOT(I16300)
--	I16303 = NOT(g6713)
--	g8987 = NOT(I16303)
--	I16306 = NOT(g7015)
--	g8990 = NOT(I16306)
--	I16309 = NOT(g5512)
--	g8993 = NOT(I16309)
--	I16312 = NOT(g5424)
--	g8996 = NOT(I16312)
--	I16315 = NOT(g3774)
--	g8997 = NOT(I16315)
--	I16318 = NOT(g5556)
--	g9000 = NOT(I16318)
--	I16321 = NOT(g5425)
--	g9003 = NOT(I16321)
--	I16325 = NOT(g6052)
--	g9005 = NOT(I16325)
--	I16328 = NOT(g3900)
--	g9006 = NOT(I16328)
--	I16332 = NOT(g3462)
--	g9010 = NOT(I16332)
--	I16335 = NOT(g3618)
--	g9013 = NOT(I16335)
--	I16338 = NOT(g7015)
--	g9016 = NOT(I16338)
--	I16341 = NOT(g7265)
--	g9019 = NOT(I16341)
--	I16344 = NOT(g5556)
--	g9022 = NOT(I16344)
--	I16347 = NOT(g5427)
--	g9025 = NOT(I16347)
--	g9027 = NOT(g5679)
--	I16354 = NOT(g3618)
--	g9035 = NOT(I16354)
--	I16357 = NOT(g3774)
--	g9038 = NOT(I16357)
--	I16360 = NOT(g7265)
--	g9041 = NOT(I16360)
--	I16363 = NOT(g3900)
--	g9044 = NOT(I16363)
--	g9050 = NOT(g5731)
--	I16372 = NOT(g3774)
--	g9058 = NOT(I16372)
--	g9067 = NOT(g5789)
--	g9084 = NOT(g5848)
--	I16432 = NOT(g3366)
--	g9128 = NOT(I16432)
--	I16438 = NOT(g3522)
--	g9134 = NOT(I16438)
--	I16444 = NOT(g3678)
--	g9140 = NOT(I16444)
--	I16450 = NOT(g3834)
--	g9146 = NOT(I16450)
--	I16453 = NOT(g7936)
--	g9149 = NOT(I16453)
--	g9150 = NOT(g5893)
--	I16457 = NOT(g7936)
--	g9159 = NOT(I16457)
--	g9160 = NOT(g6170)
--	g9161 = NOT(g5852)
--	I16462 = NOT(g5438)
--	g9170 = NOT(I16462)
--	I16465 = NOT(g6000)
--	g9173 = NOT(I16465)
--	g9174 = NOT(g5932)
--	I16469 = NOT(g7936)
--	g9183 = NOT(I16469)
--	I16472 = NOT(g7901)
--	g9184 = NOT(I16472)
--	g9187 = NOT(g5803)
--	I16476 = NOT(g6448)
--	g9196 = NOT(I16476)
--	I16479 = NOT(g5438)
--	g9199 = NOT(I16479)
--	I16482 = NOT(g6000)
--	g9202 = NOT(I16482)
--	g9203 = NOT(g5899)
--	I16486 = NOT(g5473)
--	g9212 = NOT(I16486)
--	I16489 = NOT(g6000)
--	g9215 = NOT(I16489)
--	g9216 = NOT(g5966)
--	I16493 = NOT(g7936)
--	g9225 = NOT(I16493)
--	g9226 = NOT(g5434)
--	g9227 = NOT(g5587)
--	g9228 = NOT(g7667)
--	I16499 = NOT(g7901)
--	g9229 = NOT(I16499)
--	g9232 = NOT(g5752)
--	I16504 = NOT(g3306)
--	g9242 = NOT(I16504)
--	I16507 = NOT(g6448)
--	g9245 = NOT(I16507)
--	g9248 = NOT(g5859)
--	I16511 = NOT(g6713)
--	g9257 = NOT(I16511)
--	I16514 = NOT(g5473)
--	g9260 = NOT(I16514)
--	I16517 = NOT(g6000)
--	g9263 = NOT(I16517)
--	g9264 = NOT(g5938)
--	I16521 = NOT(g5512)
--	g9273 = NOT(I16521)
--	I16524 = NOT(g6000)
--	g9276 = NOT(I16524)
--	g9277 = NOT(g5995)
--	g9286 = NOT(g6197)
--	g9287 = NOT(g6638)
--	g9288 = NOT(g5363)
--	g9289 = NOT(g5379)
--	I16532 = NOT(g7901)
--	g9290 = NOT(I16532)
--	g9293 = NOT(g5703)
--	I16538 = NOT(g3306)
--	g9303 = NOT(I16538)
--	I16541 = NOT(g5438)
--	g9306 = NOT(I16541)
--	I16544 = NOT(g6054)
--	g9309 = NOT(I16544)
--	g9310 = NOT(g5811)
--	I16549 = NOT(g3462)
--	g9320 = NOT(I16549)
--	I16552 = NOT(g6713)
--	g9323 = NOT(I16552)
--	g9326 = NOT(g5906)
--	I16556 = NOT(g7015)
--	g9335 = NOT(I16556)
--	I16559 = NOT(g5512)
--	g9338 = NOT(I16559)
--	I16562 = NOT(g6000)
--	g9341 = NOT(I16562)
--	g9342 = NOT(g5972)
--	I16566 = NOT(g5556)
--	g9351 = NOT(I16566)
--	I16569 = NOT(g6000)
--	g9354 = NOT(I16569)
--	g9355 = NOT(g7639)
--	g9356 = NOT(g5665)
--	I16578 = NOT(g6448)
--	g9368 = NOT(I16578)
--	I16581 = NOT(g5438)
--	g9371 = NOT(I16581)
--	g9374 = NOT(g5761)
--	I16587 = NOT(g3462)
--	g9384 = NOT(I16587)
--	I16590 = NOT(g5473)
--	g9387 = NOT(I16590)
--	I16593 = NOT(g6059)
--	g9390 = NOT(I16593)
--	g9391 = NOT(g5867)
--	I16598 = NOT(g3618)
--	g9401 = NOT(I16598)
--	I16601 = NOT(g7015)
--	g9404 = NOT(I16601)
--	g9407 = NOT(g5945)
--	I16605 = NOT(g7265)
--	g9416 = NOT(I16605)
--	I16608 = NOT(g5556)
--	g9419 = NOT(I16608)
--	I16611 = NOT(g6000)
--	g9422 = NOT(I16611)
--	g9423 = NOT(g5428)
--	g9424 = NOT(g5469)
--	g9425 = NOT(g5346)
--	g9426 = NOT(g5543)
--	g9427 = NOT(g5645)
--	I16624 = NOT(g3306)
--	g9443 = NOT(I16624)
--	I16627 = NOT(g6448)
--	g9446 = NOT(I16627)
--	I16630 = NOT(g6057)
--	g9449 = NOT(I16630)
--	I16633 = NOT(g6486)
--	g9450 = NOT(I16633)
--	g9453 = NOT(g5717)
--	I16641 = NOT(g6713)
--	g9465 = NOT(I16641)
--	I16644 = NOT(g5473)
--	g9468 = NOT(I16644)
--	g9471 = NOT(g5820)
--	I16650 = NOT(g3618)
--	g9481 = NOT(I16650)
--	I16653 = NOT(g5512)
--	g9484 = NOT(I16653)
--	I16656 = NOT(g6066)
--	g9487 = NOT(I16656)
--	g9488 = NOT(g5914)
--	I16661 = NOT(g3774)
--	g9498 = NOT(I16661)
--	I16664 = NOT(g7265)
--	g9501 = NOT(I16664)
--	g9504 = NOT(g6149)
--	g9505 = NOT(g6227)
--	g9506 = NOT(g6444)
--	g9507 = NOT(g5953)
--	I16677 = NOT(g3306)
--	g9524 = NOT(I16677)
--	g9527 = NOT(g5508)
--	I16681 = NOT(g6643)
--	g9528 = NOT(I16681)
--	I16684 = NOT(g6486)
--	g9531 = NOT(I16684)
--	g9569 = NOT(g5683)
--	I16694 = NOT(g3462)
--	g9585 = NOT(I16694)
--	I16697 = NOT(g6713)
--	g9588 = NOT(I16697)
--	I16700 = NOT(g6064)
--	g9591 = NOT(I16700)
--	I16703 = NOT(g6751)
--	g9592 = NOT(I16703)
--	g9595 = NOT(g5775)
--	I16711 = NOT(g7015)
--	g9607 = NOT(I16711)
--	I16714 = NOT(g5512)
--	g9610 = NOT(I16714)
--	g9613 = NOT(g5876)
--	I16720 = NOT(g3774)
--	g9623 = NOT(I16720)
--	I16723 = NOT(g5556)
--	g9626 = NOT(I16723)
--	I16726 = NOT(g6085)
--	g9629 = NOT(I16726)
--	I16741 = NOT(g6062)
--	g9640 = NOT(I16741)
--	I16744 = NOT(g3338)
--	g9641 = NOT(I16744)
--	I16747 = NOT(g6643)
--	g9644 = NOT(I16747)
--	g9649 = NOT(g5982)
--	I16759 = NOT(g3462)
--	g9666 = NOT(I16759)
--	g9669 = NOT(g5552)
--	I16763 = NOT(g6945)
--	g9670 = NOT(I16763)
--	I16766 = NOT(g6751)
--	g9673 = NOT(I16766)
--	g9711 = NOT(g5735)
--	I16776 = NOT(g3618)
--	g9727 = NOT(I16776)
--	I16779 = NOT(g7015)
--	g9730 = NOT(I16779)
--	I16782 = NOT(g6083)
--	g9733 = NOT(I16782)
--	I16785 = NOT(g7053)
--	g9734 = NOT(I16785)
--	g9737 = NOT(g5834)
--	I16793 = NOT(g7265)
--	g9749 = NOT(I16793)
--	I16796 = NOT(g5556)
--	g9752 = NOT(I16796)
--	g9755 = NOT(g5431)
--	g9756 = NOT(g5504)
--	g9757 = NOT(g5601)
--	g9758 = NOT(g5618)
--	I16811 = NOT(g3338)
--	g9767 = NOT(I16811)
--	I16814 = NOT(g6486)
--	g9770 = NOT(I16814)
--	I16832 = NOT(g6081)
--	g9786 = NOT(I16832)
--	I16835 = NOT(g3494)
--	g9787 = NOT(I16835)
--	I16838 = NOT(g6945)
--	g9790 = NOT(I16838)
--	g9795 = NOT(g6019)
--	I16850 = NOT(g3618)
--	g9812 = NOT(I16850)
--	g9815 = NOT(g5598)
--	I16854 = NOT(g7195)
--	g9816 = NOT(I16854)
--	I16857 = NOT(g7053)
--	g9819 = NOT(I16857)
--	g9857 = NOT(g5793)
--	I16867 = NOT(g3774)
--	g9873 = NOT(I16867)
--	I16870 = NOT(g7265)
--	g9876 = NOT(I16870)
--	I16873 = NOT(g6102)
--	g9879 = NOT(I16873)
--	I16876 = NOT(g7303)
--	g9880 = NOT(I16876)
--	g9884 = NOT(g6310)
--	g9885 = NOT(g6905)
--	g9886 = NOT(g7149)
--	I16897 = NOT(g6643)
--	g9895 = NOT(I16897)
--	I16900 = NOT(g6486)
--	g9898 = NOT(I16900)
--	I16915 = NOT(g3494)
--	g9913 = NOT(I16915)
--	I16918 = NOT(g6751)
--	g9916 = NOT(I16918)
--	I16936 = NOT(g6100)
--	g9932 = NOT(I16936)
--	I16939 = NOT(g3650)
--	g9933 = NOT(I16939)
--	I16942 = NOT(g7195)
--	g9936 = NOT(I16942)
--	g9941 = NOT(g6035)
--	I16954 = NOT(g3774)
--	g9958 = NOT(I16954)
--	g9961 = NOT(g5615)
--	I16958 = NOT(g7391)
--	g9962 = NOT(I16958)
--	I16961 = NOT(g7303)
--	g9965 = NOT(I16961)
--	I16972 = NOT(g3900)
--	g10004 = NOT(I16972)
--	g10015 = NOT(g5292)
--	I16984 = NOT(g7936)
--	g10016 = NOT(I16984)
--	I16987 = NOT(g6079)
--	g10017 = NOT(I16987)
--	I16990 = NOT(g3338)
--	g10018 = NOT(I16990)
--	I16993 = NOT(g6643)
--	g10021 = NOT(I16993)
--	I17009 = NOT(g6945)
--	g10049 = NOT(I17009)
--	I17012 = NOT(g6751)
--	g10052 = NOT(I17012)
--	I17027 = NOT(g3650)
--	g10067 = NOT(I17027)
--	I17030 = NOT(g7053)
--	g10070 = NOT(I17030)
--	I17048 = NOT(g6117)
--	g10086 = NOT(I17048)
--	I17051 = NOT(g3806)
--	g10087 = NOT(I17051)
--	I17054 = NOT(g7391)
--	g10090 = NOT(I17054)
--	I17066 = NOT(g3900)
--	g10096 = NOT(I17066)
--	g10099 = NOT(g7700)
--	I17070 = NOT(g7528)
--	g10100 = NOT(I17070)
--	I17081 = NOT(g3338)
--	g10109 = NOT(I17081)
--	g10124 = NOT(g5326)
--	I17097 = NOT(g7936)
--	g10125 = NOT(I17097)
--	I17100 = NOT(g6098)
--	g10126 = NOT(I17100)
--	I17103 = NOT(g3494)
--	g10127 = NOT(I17103)
--	I17106 = NOT(g6945)
--	g10130 = NOT(I17106)
--	I17122 = NOT(g7195)
--	g10158 = NOT(I17122)
--	I17125 = NOT(g7053)
--	g10161 = NOT(I17125)
--	I17140 = NOT(g3806)
--	g10176 = NOT(I17140)
--	I17143 = NOT(g7303)
--	g10179 = NOT(I17143)
--	I17159 = NOT(g3900)
--	g10189 = NOT(I17159)
--	I17184 = NOT(g3494)
--	g10214 = NOT(I17184)
--	g10229 = NOT(g5349)
--	I17200 = NOT(g7936)
--	g10230 = NOT(I17200)
--	I17203 = NOT(g6115)
--	g10231 = NOT(I17203)
--	I17206 = NOT(g3650)
--	g10232 = NOT(I17206)
--	I17209 = NOT(g7195)
--	g10235 = NOT(I17209)
--	I17225 = NOT(g7391)
--	g10263 = NOT(I17225)
--	I17228 = NOT(g7303)
--	g10266 = NOT(I17228)
--	I17235 = NOT(g3900)
--	g10273 = NOT(I17235)
--	I17238 = NOT(g3900)
--	g10276 = NOT(I17238)
--	I17278 = NOT(g3650)
--	g10316 = NOT(I17278)
--	g10331 = NOT(g5366)
--	I17294 = NOT(g7936)
--	g10332 = NOT(I17294)
--	I17297 = NOT(g6130)
--	g10333 = NOT(I17297)
--	I17300 = NOT(g3806)
--	g10334 = NOT(I17300)
--	I17303 = NOT(g7391)
--	g10337 = NOT(I17303)
--	I17311 = NOT(g3900)
--	g10357 = NOT(I17311)
--	I17363 = NOT(g3806)
--	g10409 = NOT(I17363)
--	I17370 = NOT(g3900)
--	g10416 = NOT(I17370)
--	I17373 = NOT(g3900)
--	g10419 = NOT(I17373)
--	g10424 = NOT(g7910)
--	g10481 = NOT(g7826)
--	I17433 = NOT(g3900)
--	g10482 = NOT(I17433)
--	g10486 = NOT(g7957)
--	g10500 = NOT(g7962)
--	I17483 = NOT(g3900)
--	g10542 = NOT(I17483)
--	I17486 = NOT(g3900)
--	g10545 = NOT(I17486)
--	g10549 = NOT(g7999)
--	g10560 = NOT(g8008)
--	g10574 = NOT(g8013)
--	I17527 = NOT(g3900)
--	g10601 = NOT(I17527)
--	g10606 = NOT(g8074)
--	g10617 = NOT(g8083)
--	g10631 = NOT(g8088)
--	I17557 = NOT(g3900)
--	g10646 = NOT(I17557)
--	g10653 = NOT(g8159)
--	g10664 = NOT(g8168)
--	g10683 = NOT(g8245)
--	g10694 = NOT(g4326)
--	g10714 = NOT(g4495)
--	g10730 = NOT(g6173)
--	g10735 = NOT(g4671)
--	g10749 = NOT(g6205)
--	g10754 = NOT(g4848)
--	g10765 = NOT(g6048)
--	g10766 = NOT(g6676)
--	g10767 = NOT(g6294)
--	g10772 = NOT(g6978)
--	g10773 = NOT(g6431)
--	I17627 = NOT(g7575)
--	g10779 = NOT(I17627)
--	g10783 = NOT(g7228)
--	I17632 = NOT(g6183)
--	g10787 = NOT(I17632)
--	g10788 = NOT(g7424)
--	I17637 = NOT(g6204)
--	g10792 = NOT(I17637)
--	I17641 = NOT(g6215)
--	g10796 = NOT(I17641)
--	I17645 = NOT(g6288)
--	g10800 = NOT(I17645)
--	I17649 = NOT(g6293)
--	g10804 = NOT(I17649)
--	I17653 = NOT(g6304)
--	g10808 = NOT(I17653)
--	g10809 = NOT(g5701)
--	I17658 = NOT(g6367)
--	g10813 = NOT(I17658)
--	I17662 = NOT(g6425)
--	g10817 = NOT(I17662)
--	I17666 = NOT(g6430)
--	g10821 = NOT(I17666)
--	I17670 = NOT(g6441)
--	g10825 = NOT(I17670)
--	I17673 = NOT(g8107)
--	g10826 = NOT(I17673)
--	g10829 = NOT(g5749)
--	I17677 = NOT(g6517)
--	g10830 = NOT(I17677)
--	I17681 = NOT(g6572)
--	g10834 = NOT(I17681)
--	I17685 = NOT(g6630)
--	g10838 = NOT(I17685)
--	I17689 = NOT(g6635)
--	g10842 = NOT(I17689)
--	I17692 = NOT(g8107)
--	g10843 = NOT(I17692)
--	g10846 = NOT(g5799)
--	g10847 = NOT(g5800)
--	g10848 = NOT(g5801)
--	I17698 = NOT(g6711)
--	g10849 = NOT(I17698)
--	I17701 = NOT(g6781)
--	g10850 = NOT(I17701)
--	I17705 = NOT(g6836)
--	g10854 = NOT(I17705)
--	I17709 = NOT(g6894)
--	g10858 = NOT(I17709)
--	I17712 = NOT(g8031)
--	g10859 = NOT(I17712)
--	I17715 = NOT(g8107)
--	g10862 = NOT(I17715)
--	g10865 = NOT(g6131)
--	g10866 = NOT(g5849)
--	g10867 = NOT(g5850)
--	I17721 = NOT(g6641)
--	g10868 = NOT(I17721)
--	I17724 = NOT(g6942)
--	g10869 = NOT(I17724)
--	I17727 = NOT(g7013)
--	g10870 = NOT(I17727)
--	I17730 = NOT(g7083)
--	g10871 = NOT(I17730)
--	I17734 = NOT(g7138)
--	g10875 = NOT(I17734)
--	I17737 = NOT(g6000)
--	g10876 = NOT(I17737)
--	I17740 = NOT(g8031)
--	g10877 = NOT(I17740)
--	I17743 = NOT(g8107)
--	g10880 = NOT(I17743)
--	I17746 = NOT(g8107)
--	g10883 = NOT(I17746)
--	g10886 = NOT(g5889)
--	I17750 = NOT(g7157)
--	g10887 = NOT(I17750)
--	I17753 = NOT(g6943)
--	g10888 = NOT(I17753)
--	I17756 = NOT(g7192)
--	g10889 = NOT(I17756)
--	I17759 = NOT(g7263)
--	g10890 = NOT(I17759)
--	I17762 = NOT(g7333)
--	g10891 = NOT(I17762)
--	I17765 = NOT(g7976)
--	g10892 = NOT(I17765)
--	I17768 = NOT(g8031)
--	g10895 = NOT(I17768)
--	I17771 = NOT(g8107)
--	g10898 = NOT(I17771)
--	I17774 = NOT(g8107)
--	g10901 = NOT(I17774)
--	g10904 = NOT(g5922)
--	g10905 = NOT(g5923)
--	g10906 = NOT(g5924)
--	I17780 = NOT(g7348)
--	g10907 = NOT(I17780)
--	I17783 = NOT(g7353)
--	g10908 = NOT(I17783)
--	I17786 = NOT(g7193)
--	g10909 = NOT(I17786)
--	I17789 = NOT(g7388)
--	g10910 = NOT(I17789)
--	I17792 = NOT(g7459)
--	g10911 = NOT(I17792)
--	I17795 = NOT(g7976)
--	g10912 = NOT(I17795)
--	I17798 = NOT(g8031)
--	g10915 = NOT(I17798)
--	I17801 = NOT(g8107)
--	g10918 = NOT(I17801)
--	I17804 = NOT(g8031)
--	g10921 = NOT(I17804)
--	I17807 = NOT(g8107)
--	g10924 = NOT(I17807)
--	g10927 = NOT(g6153)
--	g10928 = NOT(g5951)
--	g10929 = NOT(g5952)
--	I17813 = NOT(g5707)
--	g10930 = NOT(I17813)
--	I17816 = NOT(g7346)
--	g10931 = NOT(I17816)
--	I17819 = NOT(g6448)
--	g10932 = NOT(I17819)
--	I17822 = NOT(g7478)
--	g10933 = NOT(I17822)
--	I17825 = NOT(g7483)
--	g10934 = NOT(I17825)
--	I17828 = NOT(g7389)
--	g10935 = NOT(I17828)
--	I17831 = NOT(g7518)
--	g10936 = NOT(I17831)
--	I17834 = NOT(g7976)
--	g10937 = NOT(I17834)
--	I17837 = NOT(g8031)
--	g10940 = NOT(I17837)
--	I17840 = NOT(g8107)
--	g10943 = NOT(I17840)
--	I17843 = NOT(g8031)
--	g10946 = NOT(I17843)
--	I17846 = NOT(g8107)
--	g10949 = NOT(I17846)
--	I17849 = NOT(g8103)
--	g10952 = NOT(I17849)
--	g10961 = NOT(g5978)
--	g10962 = NOT(g5979)
--	I17854 = NOT(g6232)
--	g10963 = NOT(I17854)
--	I17857 = NOT(g6448)
--	g10966 = NOT(I17857)
--	I17860 = NOT(g5765)
--	g10967 = NOT(I17860)
--	I17863 = NOT(g7476)
--	g10968 = NOT(I17863)
--	I17866 = NOT(g6713)
--	g10969 = NOT(I17866)
--	I17869 = NOT(g7534)
--	g10972 = NOT(I17869)
--	I17872 = NOT(g7539)
--	g10973 = NOT(I17872)
--	I17875 = NOT(g7976)
--	g10974 = NOT(I17875)
--	I17878 = NOT(g8031)
--	g10977 = NOT(I17878)
--	I17881 = NOT(g7976)
--	g10980 = NOT(I17881)
--	I17884 = NOT(g8031)
--	g10983 = NOT(I17884)
--	g10986 = NOT(g6014)
--	g10987 = NOT(g6015)
--	I17889 = NOT(g6314)
--	g10988 = NOT(I17889)
--	I17892 = NOT(g6232)
--	g10991 = NOT(I17892)
--	I17895 = NOT(g6448)
--	g10994 = NOT(I17895)
--	I17898 = NOT(g6643)
--	g10995 = NOT(I17898)
--	I17901 = NOT(g6369)
--	g10996 = NOT(I17901)
--	I17904 = NOT(g6713)
--	g10999 = NOT(I17904)
--	I17907 = NOT(g5824)
--	g11002 = NOT(I17907)
--	I17910 = NOT(g7532)
--	g11003 = NOT(I17910)
--	I17913 = NOT(g7015)
--	g11004 = NOT(I17913)
--	I17916 = NOT(g7560)
--	g11007 = NOT(I17916)
--	I17919 = NOT(g7976)
--	g11008 = NOT(I17919)
--	I17922 = NOT(g8031)
--	g11011 = NOT(I17922)
--	I17925 = NOT(g7976)
--	g11014 = NOT(I17925)
--	I17928 = NOT(g8031)
--	g11017 = NOT(I17928)
--	g11020 = NOT(g6029)
--	g11021 = NOT(g6030)
--	I17933 = NOT(g3254)
--	g11022 = NOT(I17933)
--	I17936 = NOT(g6314)
--	g11025 = NOT(I17936)
--	I17939 = NOT(g6232)
--	g11028 = NOT(I17939)
--	I17942 = NOT(g5548)
--	g11031 = NOT(I17942)
--	I17945 = NOT(g5668)
--	g11032 = NOT(I17945)
--	I17948 = NOT(g6643)
--	g11035 = NOT(I17948)
--	I17951 = NOT(g6519)
--	g11036 = NOT(I17951)
--	I17954 = NOT(g6369)
--	g11039 = NOT(I17954)
--	I17957 = NOT(g6713)
--	g11042 = NOT(I17957)
--	I17960 = NOT(g6945)
--	g11045 = NOT(I17960)
--	I17963 = NOT(g6574)
--	g11048 = NOT(I17963)
--	I17966 = NOT(g7015)
--	g11051 = NOT(I17966)
--	I17969 = NOT(g5880)
--	g11054 = NOT(I17969)
--	I17972 = NOT(g7558)
--	g11055 = NOT(I17972)
--	I17975 = NOT(g7265)
--	g11056 = NOT(I17975)
--	I17978 = NOT(g7795)
--	g11059 = NOT(I17978)
--	I17981 = NOT(g7976)
--	g11063 = NOT(I17981)
--	I17984 = NOT(g7976)
--	g11066 = NOT(I17984)
--	g11069 = NOT(g8257)
--	g11078 = NOT(g6041)
--	I17989 = NOT(g3254)
--	g11079 = NOT(I17989)
--	I17992 = NOT(g6314)
--	g11082 = NOT(I17992)
--	I17995 = NOT(g6232)
--	g11085 = NOT(I17995)
--	I17998 = NOT(g5668)
--	g11088 = NOT(I17998)
--	I18001 = NOT(g6643)
--	g11091 = NOT(I18001)
--	I18004 = NOT(g3410)
--	g11092 = NOT(I18004)
--	I18007 = NOT(g6519)
--	g11095 = NOT(I18007)
--	I18010 = NOT(g6369)
--	g11098 = NOT(I18010)
--	I18013 = NOT(g5594)
--	g11101 = NOT(I18013)
--	I18016 = NOT(g5720)
--	g11102 = NOT(I18016)
--	I18019 = NOT(g6945)
--	g11105 = NOT(I18019)
--	I18022 = NOT(g6783)
--	g11108 = NOT(I18022)
--	I18025 = NOT(g6574)
--	g11111 = NOT(I18025)
--	I18028 = NOT(g7015)
--	g11114 = NOT(I18028)
--	I18031 = NOT(g7195)
--	g11117 = NOT(I18031)
--	I18034 = NOT(g6838)
--	g11120 = NOT(I18034)
--	I18037 = NOT(g7265)
--	g11123 = NOT(I18037)
--	I18040 = NOT(g7976)
--	g11126 = NOT(I18040)
--	I18043 = NOT(g7976)
--	g11129 = NOT(I18043)
--	I18046 = NOT(g3254)
--	g11132 = NOT(I18046)
--	I18049 = NOT(g6314)
--	g11135 = NOT(I18049)
--	I18052 = NOT(g6232)
--	g11138 = NOT(I18052)
--	I18055 = NOT(g5668)
--	g11141 = NOT(I18055)
--	I18058 = NOT(g6643)
--	g11144 = NOT(I18058)
--	I18061 = NOT(g3410)
--	g11145 = NOT(I18061)
--	I18064 = NOT(g6519)
--	g11148 = NOT(I18064)
--	I18067 = NOT(g6369)
--	g11151 = NOT(I18067)
--	I18070 = NOT(g5720)
--	g11154 = NOT(I18070)
--	I18073 = NOT(g6945)
--	g11157 = NOT(I18073)
--	I18076 = NOT(g3566)
--	g11160 = NOT(I18076)
--	I18079 = NOT(g6783)
--	g11163 = NOT(I18079)
--	I18082 = NOT(g6574)
--	g11166 = NOT(I18082)
--	I18085 = NOT(g5611)
--	g11169 = NOT(I18085)
--	I18088 = NOT(g5778)
--	g11170 = NOT(I18088)
--	I18091 = NOT(g7195)
--	g11173 = NOT(I18091)
--	I18094 = NOT(g7085)
--	g11176 = NOT(I18094)
--	I18097 = NOT(g6838)
--	g11179 = NOT(I18097)
--	I18100 = NOT(g7265)
--	g11182 = NOT(I18100)
--	I18103 = NOT(g7391)
--	g11185 = NOT(I18103)
--	g11190 = NOT(g3999)
--	I18121 = NOT(g3254)
--	g11199 = NOT(I18121)
--	I18124 = NOT(g6314)
--	g11202 = NOT(I18124)
--	I18127 = NOT(g6232)
--	g11205 = NOT(I18127)
--	I18130 = NOT(g5547)
--	g11208 = NOT(I18130)
--	I18133 = NOT(g6448)
--	g11209 = NOT(I18133)
--	I18136 = NOT(g5668)
--	g11210 = NOT(I18136)
--	I18139 = NOT(g6643)
--	g11213 = NOT(I18139)
--	I18142 = NOT(g3410)
--	g11216 = NOT(I18142)
--	I18145 = NOT(g6519)
--	g11219 = NOT(I18145)
--	I18148 = NOT(g6369)
--	g11222 = NOT(I18148)
--	I18151 = NOT(g5720)
--	g11225 = NOT(I18151)
--	I18154 = NOT(g6945)
--	g11228 = NOT(I18154)
--	I18157 = NOT(g3566)
--	g11231 = NOT(I18157)
--	I18160 = NOT(g6783)
--	g11234 = NOT(I18160)
--	I18163 = NOT(g6574)
--	g11237 = NOT(I18163)
--	I18166 = NOT(g5778)
--	g11240 = NOT(I18166)
--	I18169 = NOT(g7195)
--	g11243 = NOT(I18169)
--	I18172 = NOT(g3722)
--	g11246 = NOT(I18172)
--	I18175 = NOT(g7085)
--	g11249 = NOT(I18175)
--	I18178 = NOT(g6838)
--	g11252 = NOT(I18178)
--	I18181 = NOT(g5636)
--	g11255 = NOT(I18181)
--	I18184 = NOT(g5837)
--	g11256 = NOT(I18184)
--	I18187 = NOT(g7391)
--	g11259 = NOT(I18187)
--	I18211 = NOT(g6232)
--	g11265 = NOT(I18211)
--	I18214 = NOT(g3254)
--	g11268 = NOT(I18214)
--	I18217 = NOT(g6314)
--	g11271 = NOT(I18217)
--	I18220 = NOT(g6232)
--	g11274 = NOT(I18220)
--	I18223 = NOT(g6448)
--	g11277 = NOT(I18223)
--	I18226 = NOT(g5668)
--	g11278 = NOT(I18226)
--	I18229 = NOT(g3410)
--	g11281 = NOT(I18229)
--	I18232 = NOT(g6519)
--	g11284 = NOT(I18232)
--	I18235 = NOT(g6369)
--	g11287 = NOT(I18235)
--	I18238 = NOT(g5593)
--	g11290 = NOT(I18238)
--	I18241 = NOT(g6713)
--	g11291 = NOT(I18241)
--	I18244 = NOT(g5720)
--	g11294 = NOT(I18244)
--	I18247 = NOT(g6945)
--	g11297 = NOT(I18247)
--	I18250 = NOT(g3566)
--	g11300 = NOT(I18250)
--	I18253 = NOT(g6783)
--	g11303 = NOT(I18253)
--	I18256 = NOT(g6574)
--	g11306 = NOT(I18256)
--	I18259 = NOT(g5778)
--	g11309 = NOT(I18259)
--	I18262 = NOT(g7195)
--	g11312 = NOT(I18262)
--	I18265 = NOT(g3722)
--	g11315 = NOT(I18265)
--	I18268 = NOT(g7085)
--	g11318 = NOT(I18268)
--	I18271 = NOT(g6838)
--	g11321 = NOT(I18271)
--	I18274 = NOT(g5837)
--	g11324 = NOT(I18274)
--	I18277 = NOT(g7391)
--	g11327 = NOT(I18277)
--	g11332 = NOT(g4094)
--	I18295 = NOT(g6314)
--	g11341 = NOT(I18295)
--	I18298 = NOT(g6232)
--	g11344 = NOT(I18298)
--	I18302 = NOT(g3254)
--	g11348 = NOT(I18302)
--	I18305 = NOT(g6314)
--	g11351 = NOT(I18305)
--	I18308 = NOT(g6448)
--	g11354 = NOT(I18308)
--	I18311 = NOT(g5668)
--	g11355 = NOT(I18311)
--	I18314 = NOT(g6369)
--	g11358 = NOT(I18314)
--	I18317 = NOT(g3410)
--	g11361 = NOT(I18317)
--	I18320 = NOT(g6519)
--	g11364 = NOT(I18320)
--	I18323 = NOT(g6369)
--	g11367 = NOT(I18323)
--	I18326 = NOT(g6713)
--	g11370 = NOT(I18326)
--	I18329 = NOT(g5720)
--	g11373 = NOT(I18329)
--	I18332 = NOT(g3566)
--	g11376 = NOT(I18332)
--	I18335 = NOT(g6783)
--	g11379 = NOT(I18335)
--	I18338 = NOT(g6574)
--	g11382 = NOT(I18338)
--	I18341 = NOT(g5610)
--	g11385 = NOT(I18341)
--	I18344 = NOT(g7015)
--	g11386 = NOT(I18344)
--	I18347 = NOT(g5778)
--	g11389 = NOT(I18347)
--	I18350 = NOT(g7195)
--	g11392 = NOT(I18350)
--	I18353 = NOT(g3722)
--	g11395 = NOT(I18353)
--	I18356 = NOT(g7085)
--	g11398 = NOT(I18356)
--	I18359 = NOT(g6838)
--	g11401 = NOT(I18359)
--	I18362 = NOT(g5837)
--	g11404 = NOT(I18362)
--	I18365 = NOT(g7391)
--	g11407 = NOT(I18365)
--	I18375 = NOT(g3254)
--	g11411 = NOT(I18375)
--	I18378 = NOT(g6314)
--	g11414 = NOT(I18378)
--	I18381 = NOT(g6232)
--	g11417 = NOT(I18381)
--	I18386 = NOT(g3254)
--	g11422 = NOT(I18386)
--	I18389 = NOT(g6519)
--	g11425 = NOT(I18389)
--	I18392 = NOT(g6369)
--	g11428 = NOT(I18392)
--	I18396 = NOT(g3410)
--	g11432 = NOT(I18396)
--	I18399 = NOT(g6519)
--	g11435 = NOT(I18399)
--	I18402 = NOT(g6713)
--	g11438 = NOT(I18402)
--	I18405 = NOT(g5720)
--	g11441 = NOT(I18405)
--	I18408 = NOT(g6574)
--	g11444 = NOT(I18408)
--	I18411 = NOT(g3566)
--	g11447 = NOT(I18411)
--	I18414 = NOT(g6783)
--	g11450 = NOT(I18414)
--	I18417 = NOT(g6574)
--	g11453 = NOT(I18417)
--	I18420 = NOT(g7015)
--	g11456 = NOT(I18420)
--	I18423 = NOT(g5778)
--	g11459 = NOT(I18423)
--	I18426 = NOT(g3722)
--	g11462 = NOT(I18426)
--	I18429 = NOT(g7085)
--	g11465 = NOT(I18429)
--	I18432 = NOT(g6838)
--	g11468 = NOT(I18432)
--	I18435 = NOT(g5635)
--	g11471 = NOT(I18435)
--	I18438 = NOT(g7265)
--	g11472 = NOT(I18438)
--	I18441 = NOT(g5837)
--	g11475 = NOT(I18441)
--	I18444 = NOT(g7391)
--	g11478 = NOT(I18444)
--	g11481 = NOT(g4204)
--	g11490 = NOT(g8276)
--	I18449 = NOT(g10868)
--	g11491 = NOT(I18449)
--	I18452 = NOT(g10930)
--	g11492 = NOT(I18452)
--	I18455 = NOT(g11031)
--	g11493 = NOT(I18455)
--	I18458 = NOT(g11208)
--	g11494 = NOT(I18458)
--	I18461 = NOT(g10931)
--	g11495 = NOT(I18461)
--	I18464 = NOT(g8620)
--	g11496 = NOT(I18464)
--	I18467 = NOT(g8769)
--	g11497 = NOT(I18467)
--	I18470 = NOT(g8808)
--	g11498 = NOT(I18470)
--	I18473 = NOT(g8839)
--	g11499 = NOT(I18473)
--	I18476 = NOT(g8791)
--	g11500 = NOT(I18476)
--	I18479 = NOT(g8820)
--	g11501 = NOT(I18479)
--	I18482 = NOT(g8859)
--	g11502 = NOT(I18482)
--	I18485 = NOT(g8809)
--	g11503 = NOT(I18485)
--	I18488 = NOT(g8840)
--	g11504 = NOT(I18488)
--	I18491 = NOT(g8891)
--	g11505 = NOT(I18491)
--	I18494 = NOT(g8821)
--	g11506 = NOT(I18494)
--	I18497 = NOT(g8860)
--	g11507 = NOT(I18497)
--	I18500 = NOT(g8924)
--	g11508 = NOT(I18500)
--	I18503 = NOT(g8658)
--	g11509 = NOT(I18503)
--	I18506 = NOT(g8699)
--	g11510 = NOT(I18506)
--	I18509 = NOT(g8770)
--	g11511 = NOT(I18509)
--	I18512 = NOT(g9309)
--	g11512 = NOT(I18512)
--	I18515 = NOT(g8843)
--	g11513 = NOT(I18515)
--	I18518 = NOT(g8893)
--	g11514 = NOT(I18518)
--	I18521 = NOT(g9449)
--	g11515 = NOT(I18521)
--	I18524 = NOT(g9640)
--	g11516 = NOT(I18524)
--	I18527 = NOT(g10017)
--	g11517 = NOT(I18527)
--	I18530 = NOT(g10888)
--	g11518 = NOT(I18530)
--	I18533 = NOT(g10967)
--	g11519 = NOT(I18533)
--	I18536 = NOT(g11101)
--	g11520 = NOT(I18536)
--	I18539 = NOT(g11290)
--	g11521 = NOT(I18539)
--	I18542 = NOT(g10968)
--	g11522 = NOT(I18542)
--	I18545 = NOT(g8630)
--	g11523 = NOT(I18545)
--	I18548 = NOT(g8792)
--	g11524 = NOT(I18548)
--	I18551 = NOT(g8824)
--	g11525 = NOT(I18551)
--	I18554 = NOT(g8866)
--	g11526 = NOT(I18554)
--	I18557 = NOT(g8810)
--	g11527 = NOT(I18557)
--	I18560 = NOT(g8844)
--	g11528 = NOT(I18560)
--	I18563 = NOT(g8897)
--	g11529 = NOT(I18563)
--	I18566 = NOT(g8825)
--	g11530 = NOT(I18566)
--	I18569 = NOT(g8867)
--	g11531 = NOT(I18569)
--	I18572 = NOT(g8931)
--	g11532 = NOT(I18572)
--	I18575 = NOT(g8845)
--	g11533 = NOT(I18575)
--	I18578 = NOT(g8898)
--	g11534 = NOT(I18578)
--	I18581 = NOT(g8964)
--	g11535 = NOT(I18581)
--	I18584 = NOT(g8677)
--	g11536 = NOT(I18584)
--	I18587 = NOT(g8718)
--	g11537 = NOT(I18587)
--	I18590 = NOT(g8793)
--	g11538 = NOT(I18590)
--	I18593 = NOT(g9390)
--	g11539 = NOT(I18593)
--	I18596 = NOT(g8870)
--	g11540 = NOT(I18596)
--	I18599 = NOT(g8933)
--	g11541 = NOT(I18599)
--	I18602 = NOT(g9591)
--	g11542 = NOT(I18602)
--	I18605 = NOT(g9786)
--	g11543 = NOT(I18605)
--	I18608 = NOT(g10126)
--	g11544 = NOT(I18608)
--	I18611 = NOT(g10909)
--	g11545 = NOT(I18611)
--	I18614 = NOT(g11002)
--	g11546 = NOT(I18614)
--	I18617 = NOT(g11169)
--	g11547 = NOT(I18617)
--	I18620 = NOT(g11385)
--	g11548 = NOT(I18620)
--	I18623 = NOT(g11003)
--	g11549 = NOT(I18623)
--	I18626 = NOT(g8649)
--	g11550 = NOT(I18626)
--	I18629 = NOT(g8811)
--	g11551 = NOT(I18629)
--	I18632 = NOT(g8850)
--	g11552 = NOT(I18632)
--	I18635 = NOT(g8904)
--	g11553 = NOT(I18635)
--	I18638 = NOT(g8826)
--	g11554 = NOT(I18638)
--	I18641 = NOT(g8871)
--	g11555 = NOT(I18641)
--	I18644 = NOT(g8937)
--	g11556 = NOT(I18644)
--	I18647 = NOT(g8851)
--	g11557 = NOT(I18647)
--	I18650 = NOT(g8905)
--	g11558 = NOT(I18650)
--	I18653 = NOT(g8971)
--	g11559 = NOT(I18653)
--	I18656 = NOT(g8872)
--	g11560 = NOT(I18656)
--	I18659 = NOT(g8938)
--	g11561 = NOT(I18659)
--	I18662 = NOT(g8996)
--	g11562 = NOT(I18662)
--	I18665 = NOT(g8689)
--	g11563 = NOT(I18665)
--	I18668 = NOT(g8756)
--	g11564 = NOT(I18668)
--	I18671 = NOT(g8812)
--	g11565 = NOT(I18671)
--	I18674 = NOT(g9487)
--	g11566 = NOT(I18674)
--	I18677 = NOT(g8908)
--	g11567 = NOT(I18677)
--	I18680 = NOT(g8973)
--	g11568 = NOT(I18680)
--	I18683 = NOT(g9733)
--	g11569 = NOT(I18683)
--	I18686 = NOT(g9932)
--	g11570 = NOT(I18686)
--	I18689 = NOT(g10231)
--	g11571 = NOT(I18689)
--	I18692 = NOT(g10935)
--	g11572 = NOT(I18692)
--	I18695 = NOT(g11054)
--	g11573 = NOT(I18695)
--	I18698 = NOT(g11255)
--	g11574 = NOT(I18698)
--	I18701 = NOT(g11471)
--	g11575 = NOT(I18701)
--	I18704 = NOT(g11055)
--	g11576 = NOT(I18704)
--	I18707 = NOT(g8665)
--	g11577 = NOT(I18707)
--	I18710 = NOT(g8827)
--	g11578 = NOT(I18710)
--	I18713 = NOT(g8877)
--	g11579 = NOT(I18713)
--	I18716 = NOT(g8944)
--	g11580 = NOT(I18716)
--	I18719 = NOT(g8852)
--	g11581 = NOT(I18719)
--	I18722 = NOT(g8909)
--	g11582 = NOT(I18722)
--	I18725 = NOT(g8977)
--	g11583 = NOT(I18725)
--	I18728 = NOT(g8878)
--	g11584 = NOT(I18728)
--	I18731 = NOT(g8945)
--	g11585 = NOT(I18731)
--	I18734 = NOT(g9003)
--	g11586 = NOT(I18734)
--	I18737 = NOT(g8910)
--	g11587 = NOT(I18737)
--	I18740 = NOT(g8978)
--	g11588 = NOT(I18740)
--	I18743 = NOT(g9025)
--	g11589 = NOT(I18743)
--	I18746 = NOT(g8707)
--	g11590 = NOT(I18746)
--	I18749 = NOT(g8779)
--	g11591 = NOT(I18749)
--	I18752 = NOT(g8828)
--	g11592 = NOT(I18752)
--	I18755 = NOT(g9629)
--	g11593 = NOT(I18755)
--	I18758 = NOT(g8948)
--	g11594 = NOT(I18758)
--	I18761 = NOT(g9005)
--	g11595 = NOT(I18761)
--	I18764 = NOT(g9879)
--	g11596 = NOT(I18764)
--	I18767 = NOT(g10086)
--	g11597 = NOT(I18767)
--	I18770 = NOT(g10333)
--	g11598 = NOT(I18770)
--	I18773 = NOT(g10830)
--	g11599 = NOT(I18773)
--	I18777 = NOT(g9050)
--	g11603 = NOT(I18777)
--	I18780 = NOT(g10870)
--	g11606 = NOT(I18780)
--	I18784 = NOT(g9067)
--	g11608 = NOT(I18784)
--	I18787 = NOT(g10910)
--	g11611 = NOT(I18787)
--	I18791 = NOT(g9084)
--	g11613 = NOT(I18791)
--	I18794 = NOT(g10973)
--	g11616 = NOT(I18794)
--	g11620 = NOT(g10601)
--	g11623 = NOT(g10961)
--	I18810 = NOT(g10813)
--	g11628 = NOT(I18810)
--	I18813 = NOT(g10850)
--	g11629 = NOT(I18813)
--	I18817 = NOT(g9067)
--	g11633 = NOT(I18817)
--	I18820 = NOT(g10890)
--	g11636 = NOT(I18820)
--	I18824 = NOT(g9084)
--	g11638 = NOT(I18824)
--	I18827 = NOT(g10936)
--	g11641 = NOT(I18827)
--	g11642 = NOT(g10646)
--	I18835 = NOT(g10834)
--	g11651 = NOT(I18835)
--	I18838 = NOT(g10871)
--	g11652 = NOT(I18838)
--	I18842 = NOT(g9084)
--	g11656 = NOT(I18842)
--	I18845 = NOT(g10911)
--	g11659 = NOT(I18845)
--	I18854 = NOT(g10854)
--	g11670 = NOT(I18854)
--	I18857 = NOT(g10891)
--	g11671 = NOT(I18857)
--	I18866 = NOT(g10875)
--	g11682 = NOT(I18866)
--	g11706 = NOT(g10928)
--	g11732 = NOT(g10826)
--	g11734 = NOT(g10843)
--	g11735 = NOT(g10859)
--	g11736 = NOT(g10862)
--	g11737 = NOT(g10809)
--	g11740 = NOT(g10877)
--	g11741 = NOT(g10880)
--	g11742 = NOT(g10883)
--	g11743 = NOT(g8530)
--	g11745 = NOT(g10892)
--	g11746 = NOT(g10895)
--	g11747 = NOT(g10898)
--	g11748 = NOT(g10901)
--	I18929 = NOT(g10711)
--	g11749 = NOT(I18929)
--	g11758 = NOT(g8514)
--	g11761 = NOT(g10912)
--	g11762 = NOT(g10915)
--	g11763 = NOT(g10918)
--	g11764 = NOT(g10921)
--	g11765 = NOT(g10924)
--	g11766 = NOT(g10886)
--	I18943 = NOT(g9149)
--	g11769 = NOT(I18943)
--	g11770 = NOT(g10932)
--	g11774 = NOT(g10937)
--	g11775 = NOT(g10940)
--	g11776 = NOT(g10943)
--	g11777 = NOT(g10946)
--	g11778 = NOT(g10949)
--	g11779 = NOT(g10906)
--	g11782 = NOT(g10963)
--	g11783 = NOT(g10966)
--	I18962 = NOT(g9159)
--	g11786 = NOT(I18962)
--	g11787 = NOT(g10969)
--	I18969 = NOT(g8726)
--	g11791 = NOT(I18969)
--	g11794 = NOT(g10974)
--	g11795 = NOT(g10977)
--	g11796 = NOT(g10980)
--	g11797 = NOT(g10983)
--	g11798 = NOT(g10867)
--	g11801 = NOT(g10988)
--	g11802 = NOT(g10991)
--	g11803 = NOT(g10994)
--	g11804 = NOT(g10995)
--	g11808 = NOT(g10996)
--	g11809 = NOT(g10999)
--	I18990 = NOT(g9183)
--	g11812 = NOT(I18990)
--	g11813 = NOT(g11004)
--	g11817 = NOT(g11008)
--	g11818 = NOT(g11011)
--	g11819 = NOT(g11014)
--	g11820 = NOT(g11017)
--	g11821 = NOT(g10848)
--	g11824 = NOT(g11022)
--	g11825 = NOT(g11025)
--	g11826 = NOT(g11028)
--	g11827 = NOT(g11032)
--	g11829 = NOT(g11035)
--	g11834 = NOT(g11036)
--	g11835 = NOT(g11039)
--	g11836 = NOT(g11042)
--	g11837 = NOT(g11045)
--	g11841 = NOT(g11048)
--	g11842 = NOT(g11051)
--	I19025 = NOT(g9225)
--	g11845 = NOT(I19025)
--	g11846 = NOT(g11056)
--	I19030 = NOT(g8726)
--	g11848 = NOT(I19030)
--	g11852 = NOT(g11063)
--	g11853 = NOT(g11066)
--	g11854 = NOT(g11078)
--	g11856 = NOT(g11079)
--	g11857 = NOT(g11082)
--	g11858 = NOT(g11085)
--	g11859 = NOT(g11088)
--	g11862 = NOT(g11091)
--	g11866 = NOT(g11092)
--	g11867 = NOT(g11095)
--	g11868 = NOT(g11098)
--	g11869 = NOT(g11102)
--	g11871 = NOT(g11105)
--	g11876 = NOT(g11108)
--	g11877 = NOT(g11111)
--	g11878 = NOT(g11114)
--	g11879 = NOT(g11117)
--	g11883 = NOT(g11120)
--	g11884 = NOT(g11123)
--	g11886 = NOT(g11126)
--	g11887 = NOT(g11129)
--	g11888 = NOT(g11021)
--	g11891 = NOT(g11132)
--	g11892 = NOT(g11135)
--	g11893 = NOT(g11138)
--	g11894 = NOT(g11141)
--	g11895 = NOT(g11144)
--	g11898 = NOT(g11145)
--	g11899 = NOT(g11148)
--	g11900 = NOT(g11151)
--	g11901 = NOT(g11154)
--	g11904 = NOT(g11157)
--	g11908 = NOT(g11160)
--	g11909 = NOT(g11163)
--	g11910 = NOT(g11166)
--	g11911 = NOT(g11170)
--	g11913 = NOT(g11173)
--	g11918 = NOT(g11176)
--	g11919 = NOT(g11179)
--	g11920 = NOT(g11182)
--	g11921 = NOT(g11185)
--	I19105 = NOT(g8726)
--	g11923 = NOT(I19105)
--	g11927 = NOT(g10987)
--	g11929 = NOT(g11199)
--	g11930 = NOT(g11202)
--	g11931 = NOT(g11205)
--	g11932 = NOT(g11209)
--	g11933 = NOT(g11210)
--	g11936 = NOT(g11213)
--	I19119 = NOT(g9202)
--	g11937 = NOT(I19119)
--	g11941 = NOT(g11216)
--	g11942 = NOT(g11219)
--	g11943 = NOT(g11222)
--	g11944 = NOT(g11225)
--	g11945 = NOT(g11228)
--	g11948 = NOT(g11231)
--	g11949 = NOT(g11234)
--	g11950 = NOT(g11237)
--	g11951 = NOT(g11240)
--	g11954 = NOT(g11243)
--	g11958 = NOT(g11246)
--	g11959 = NOT(g11249)
--	g11960 = NOT(g11252)
--	g11961 = NOT(g11256)
--	g11963 = NOT(g11259)
--	g11968 = NOT(g11265)
--	g11969 = NOT(g11268)
--	g11970 = NOT(g11271)
--	g11971 = NOT(g11274)
--	g11972 = NOT(g11277)
--	g11973 = NOT(g11278)
--	I19160 = NOT(g10549)
--	g11976 = NOT(I19160)
--	g11982 = NOT(g11281)
--	g11983 = NOT(g11284)
--	g11984 = NOT(g11287)
--	g11985 = NOT(g11291)
--	g11986 = NOT(g11294)
--	g11989 = NOT(g11297)
--	I19174 = NOT(g9263)
--	g11990 = NOT(I19174)
--	g11994 = NOT(g11300)
--	g11995 = NOT(g11303)
--	g11996 = NOT(g11306)
--	g11997 = NOT(g11309)
--	g11998 = NOT(g11312)
--	g12001 = NOT(g11315)
--	g12002 = NOT(g11318)
--	g12003 = NOT(g11321)
--	g12004 = NOT(g11324)
--	g12007 = NOT(g11327)
--	I19195 = NOT(g8726)
--	g12009 = NOT(I19195)
--	g12013 = NOT(g10772)
--	g12017 = NOT(g10100)
--	g12020 = NOT(g11341)
--	g12021 = NOT(g11344)
--	g12022 = NOT(g11348)
--	g12023 = NOT(g11351)
--	g12024 = NOT(g11354)
--	g12025 = NOT(g11355)
--	I19208 = NOT(g10424)
--	g12027 = NOT(I19208)
--	I19211 = NOT(g10486)
--	g12030 = NOT(I19211)
--	g12037 = NOT(g11358)
--	g12038 = NOT(g11361)
--	g12039 = NOT(g11364)
--	g12040 = NOT(g11367)
--	g12041 = NOT(g11370)
--	g12042 = NOT(g11373)
--	I19226 = NOT(g10606)
--	g12045 = NOT(I19226)
--	g12051 = NOT(g11376)
--	g12052 = NOT(g11379)
--	g12053 = NOT(g11382)
--	g12054 = NOT(g11386)
--	g12055 = NOT(g11389)
--	g12058 = NOT(g11392)
--	I19240 = NOT(g9341)
--	g12059 = NOT(I19240)
--	g12063 = NOT(g11395)
--	g12064 = NOT(g11398)
--	g12065 = NOT(g11401)
--	g12066 = NOT(g11404)
--	g12067 = NOT(g11407)
--	g12071 = NOT(g10783)
--	g12075 = NOT(g11411)
--	g12076 = NOT(g11414)
--	g12077 = NOT(g11417)
--	g12078 = NOT(g11422)
--	g12084 = NOT(g11425)
--	g12085 = NOT(g11428)
--	g12086 = NOT(g11432)
--	g12087 = NOT(g11435)
--	g12088 = NOT(g11438)
--	g12089 = NOT(g11441)
--	I19271 = NOT(g10500)
--	g12091 = NOT(I19271)
--	I19274 = NOT(g10560)
--	g12094 = NOT(I19274)
--	g12101 = NOT(g11444)
--	g12102 = NOT(g11447)
--	g12103 = NOT(g11450)
--	g12104 = NOT(g11453)
--	g12105 = NOT(g11456)
--	g12106 = NOT(g11459)
--	I19289 = NOT(g10653)
--	g12109 = NOT(I19289)
--	g12115 = NOT(g11462)
--	g12116 = NOT(g11465)
--	g12117 = NOT(g11468)
--	g12118 = NOT(g11472)
--	g12119 = NOT(g11475)
--	g12122 = NOT(g11478)
--	I19303 = NOT(g9422)
--	g12123 = NOT(I19303)
--	I19307 = NOT(g8726)
--	g12125 = NOT(I19307)
--	g12130 = NOT(g10788)
--	g12134 = NOT(g8321)
--	g12135 = NOT(g8324)
--	I19315 = NOT(g10424)
--	g12136 = NOT(I19315)
--	I19318 = NOT(g10486)
--	g12139 = NOT(I19318)
--	I19321 = NOT(g10549)
--	g12142 = NOT(I19321)
--	g12147 = NOT(g8330)
--	g12148 = NOT(g8333)
--	g12149 = NOT(g8336)
--	g12150 = NOT(g8341)
--	g12156 = NOT(g8344)
--	g12157 = NOT(g8347)
--	g12158 = NOT(g8351)
--	g12159 = NOT(g8354)
--	g12160 = NOT(g8357)
--	g12161 = NOT(g8360)
--	I19342 = NOT(g10574)
--	g12163 = NOT(I19342)
--	I19345 = NOT(g10617)
--	g12166 = NOT(I19345)
--	g12173 = NOT(g8363)
--	g12174 = NOT(g8366)
--	g12175 = NOT(g8369)
--	g12176 = NOT(g8372)
--	g12177 = NOT(g8375)
--	g12178 = NOT(g8378)
--	I19360 = NOT(g10683)
--	g12181 = NOT(I19360)
--	g12187 = NOT(g8285)
--	g12191 = NOT(g8382)
--	g12196 = NOT(g8388)
--	g12197 = NOT(g8391)
--	I19374 = NOT(g10500)
--	g12198 = NOT(I19374)
--	I19377 = NOT(g10560)
--	g12201 = NOT(I19377)
--	I19380 = NOT(g10606)
--	g12204 = NOT(I19380)
--	g12209 = NOT(g8397)
--	g12210 = NOT(g8400)
--	g12211 = NOT(g8403)
--	g12212 = NOT(g8408)
--	g12218 = NOT(g8411)
--	g12219 = NOT(g8414)
--	g12220 = NOT(g8418)
--	g12221 = NOT(g8421)
--	g12222 = NOT(g8424)
--	g12223 = NOT(g8427)
--	I19401 = NOT(g10631)
--	g12225 = NOT(I19401)
--	I19404 = NOT(g10664)
--	g12228 = NOT(I19404)
--	g12235 = NOT(g8294)
--	I19412 = NOT(g10486)
--	g12239 = NOT(I19412)
--	I19415 = NOT(g10549)
--	g12242 = NOT(I19415)
--	g12246 = NOT(g8434)
--	g12251 = NOT(g8440)
--	g12252 = NOT(g8443)
--	I19426 = NOT(g10574)
--	g12253 = NOT(I19426)
--	I19429 = NOT(g10617)
--	g12256 = NOT(I19429)
--	I19432 = NOT(g10653)
--	g12259 = NOT(I19432)
--	g12264 = NOT(g8449)
--	g12265 = NOT(g8452)
--	g12266 = NOT(g8455)
--	g12267 = NOT(g8460)
--	g12275 = NOT(g8303)
--	I19449 = NOT(g10424)
--	g12279 = NOT(I19449)
--	I19452 = NOT(g10560)
--	g12282 = NOT(I19452)
--	I19455 = NOT(g10606)
--	g12285 = NOT(I19455)
--	g12289 = NOT(g8469)
--	g12294 = NOT(g8475)
--	g12295 = NOT(g8478)
--	I19466 = NOT(g10631)
--	g12296 = NOT(I19466)
--	I19469 = NOT(g10664)
--	g12299 = NOT(I19469)
--	I19472 = NOT(g10683)
--	g12302 = NOT(I19472)
--	g12308 = NOT(g8312)
--	I19479 = NOT(g10549)
--	g12312 = NOT(I19479)
--	I19482 = NOT(g10500)
--	g12315 = NOT(I19482)
--	I19485 = NOT(g10617)
--	g12318 = NOT(I19485)
--	I19488 = NOT(g10653)
--	g12321 = NOT(I19488)
--	g12325 = NOT(g8494)
--	g12332 = NOT(g10829)
--	I19500 = NOT(g10424)
--	g12333 = NOT(I19500)
--	I19503 = NOT(g10486)
--	g12336 = NOT(I19503)
--	I19507 = NOT(g10606)
--	g12340 = NOT(I19507)
--	I19510 = NOT(g10574)
--	g12343 = NOT(I19510)
--	I19513 = NOT(g10664)
--	g12346 = NOT(I19513)
--	I19516 = NOT(g10683)
--	g12349 = NOT(I19516)
--	g12354 = NOT(g8381)
--	g12362 = NOT(g10866)
--	I19523 = NOT(g10500)
--	g12363 = NOT(I19523)
--	I19526 = NOT(g10560)
--	g12366 = NOT(I19526)
--	I19530 = NOT(g10653)
--	g12370 = NOT(I19530)
--	I19533 = NOT(g10631)
--	g12373 = NOT(I19533)
--	g12378 = NOT(g10847)
--	I19539 = NOT(g10549)
--	g12379 = NOT(I19539)
--	I19542 = NOT(g10574)
--	g12382 = NOT(I19542)
--	I19545 = NOT(g10617)
--	g12385 = NOT(I19545)
--	I19549 = NOT(g10683)
--	g12389 = NOT(I19549)
--	I19552 = NOT(g8430)
--	g12392 = NOT(I19552)
--	g12408 = NOT(g11020)
--	I19557 = NOT(g10606)
--	g12409 = NOT(I19557)
--	I19560 = NOT(g10631)
--	g12412 = NOT(I19560)
--	I19563 = NOT(g10664)
--	g12415 = NOT(I19563)
--	g12420 = NOT(g10986)
--	I19569 = NOT(g10653)
--	g12421 = NOT(I19569)
--	g12424 = NOT(g10962)
--	I19573 = NOT(g8835)
--	g12425 = NOT(I19573)
--	I19576 = NOT(g10683)
--	g12426 = NOT(I19576)
--	g12430 = NOT(g10905)
--	I19582 = NOT(g8862)
--	g12432 = NOT(I19582)
--	g12434 = NOT(g10929)
--	I19587 = NOT(g9173)
--	g12435 = NOT(I19587)
--	I19591 = NOT(g8900)
--	g12437 = NOT(I19591)
--	g12438 = NOT(g10846)
--	I19595 = NOT(g10810)
--	g12439 = NOT(I19595)
--	I19598 = NOT(g9215)
--	g12440 = NOT(I19598)
--	I19602 = NOT(g8940)
--	g12442 = NOT(I19602)
--	I19605 = NOT(g10797)
--	g12443 = NOT(I19605)
--	I19608 = NOT(g10831)
--	g12444 = NOT(I19608)
--	I19611 = NOT(g9276)
--	g12445 = NOT(I19611)
--	I19615 = NOT(g10789)
--	g12447 = NOT(I19615)
--	I19618 = NOT(g10814)
--	g12448 = NOT(I19618)
--	I19621 = NOT(g10851)
--	g12449 = NOT(I19621)
--	I19624 = NOT(g9354)
--	g12450 = NOT(I19624)
--	I19628 = NOT(g10784)
--	g12452 = NOT(I19628)
--	I19631 = NOT(g10801)
--	g12453 = NOT(I19631)
--	I19634 = NOT(g10835)
--	g12454 = NOT(I19634)
--	I19637 = NOT(g10872)
--	g12455 = NOT(I19637)
--	g12456 = NOT(g8602)
--	I19642 = NOT(g10793)
--	g12460 = NOT(I19642)
--	I19645 = NOT(g10818)
--	g12461 = NOT(I19645)
--	I19648 = NOT(g10855)
--	g12462 = NOT(I19648)
--	g12463 = NOT(g10730)
--	g12466 = NOT(g8614)
--	I19654 = NOT(g10805)
--	g12470 = NOT(I19654)
--	I19657 = NOT(g10839)
--	g12471 = NOT(I19657)
--	g12472 = NOT(g8617)
--	g12473 = NOT(g8580)
--	g12476 = NOT(g8622)
--	g12478 = NOT(g10749)
--	g12481 = NOT(g8627)
--	I19667 = NOT(g10822)
--	g12485 = NOT(I19667)
--	g12490 = NOT(g8587)
--	g12493 = NOT(g8632)
--	g12495 = NOT(g10767)
--	g12498 = NOT(g8637)
--	g12502 = NOT(g8640)
--	g12504 = NOT(g8643)
--	g12505 = NOT(g8646)
--	g12510 = NOT(g8594)
--	g12513 = NOT(g8651)
--	g12515 = NOT(g10773)
--	g12518 = NOT(g8655)
--	I19689 = NOT(g10016)
--	g12519 = NOT(I19689)
--	g12521 = NOT(g8659)
--	g12522 = NOT(g8662)
--	g12527 = NOT(g8605)
--	g12530 = NOT(g8667)
--	g12532 = NOT(g8670)
--	g12533 = NOT(g8673)
--	I19702 = NOT(g10125)
--	g12534 = NOT(I19702)
--	g12536 = NOT(g8678)
--	g12537 = NOT(g8681)
--	g12542 = NOT(g8684)
--	I19711 = NOT(g10230)
--	g12543 = NOT(I19711)
--	g12545 = NOT(g8690)
--	g12546 = NOT(g8693)
--	g12547 = NOT(g8696)
--	I19718 = NOT(g8726)
--	g12548 = NOT(I19718)
--	g12551 = NOT(g8700)
--	I19722 = NOT(g10332)
--	g12552 = NOT(I19722)
--	g12553 = NOT(g8708)
--	g12554 = NOT(g8711)
--	I19727 = NOT(g8726)
--	g12555 = NOT(I19727)
--	g12558 = NOT(g8714)
--	g12559 = NOT(g8719)
--	g12560 = NOT(g8745)
--	I19733 = NOT(g8726)
--	g12561 = NOT(I19733)
--	I19736 = NOT(g9184)
--	g12564 = NOT(I19736)
--	I19739 = NOT(g10694)
--	g12565 = NOT(I19739)
--	g12596 = NOT(g8748)
--	g12597 = NOT(g8752)
--	g12598 = NOT(g8757)
--	g12599 = NOT(g8763)
--	g12600 = NOT(g8766)
--	I19747 = NOT(g8726)
--	g12601 = NOT(I19747)
--	I19750 = NOT(g8726)
--	g12604 = NOT(I19750)
--	I19753 = NOT(g9229)
--	g12607 = NOT(I19753)
--	I19756 = NOT(g10424)
--	g12608 = NOT(I19756)
--	I19759 = NOT(g10714)
--	g12611 = NOT(I19759)
--	g12642 = NOT(g8771)
--	g12643 = NOT(g8775)
--	g12644 = NOT(g8780)
--	g12645 = NOT(g8785)
--	g12646 = NOT(g8788)
--	I19767 = NOT(g8726)
--	g12647 = NOT(I19767)
--	I19771 = NOT(g10038)
--	g12651 = NOT(I19771)
--	I19774 = NOT(g10500)
--	g12654 = NOT(I19774)
--	I19777 = NOT(g10735)
--	g12657 = NOT(I19777)
--	g12688 = NOT(g8794)
--	g12689 = NOT(g8798)
--	g12690 = NOT(g8802)
--	g12691 = NOT(g8805)
--	I19784 = NOT(g8726)
--	g12692 = NOT(I19784)
--	I19787 = NOT(g8726)
--	g12695 = NOT(I19787)
--	I19791 = NOT(g10486)
--	g12699 = NOT(I19791)
--	I19794 = NOT(g10676)
--	g12702 = NOT(I19794)
--	I19797 = NOT(g10147)
--	g12705 = NOT(I19797)
--	I19800 = NOT(g10574)
--	g12708 = NOT(I19800)
--	I19803 = NOT(g10754)
--	g12711 = NOT(I19803)
--	g12742 = NOT(g8813)
--	g12743 = NOT(g8817)
--	I19808 = NOT(g8726)
--	g12744 = NOT(I19808)
--	g12748 = NOT(g8823)
--	I19813 = NOT(g10649)
--	g12749 = NOT(I19813)
--	I19816 = NOT(g10703)
--	g12752 = NOT(I19816)
--	I19820 = NOT(g10560)
--	g12756 = NOT(I19820)
--	I19823 = NOT(g10705)
--	g12759 = NOT(I19823)
--	I19826 = NOT(g10252)
--	g12762 = NOT(I19826)
--	I19829 = NOT(g10631)
--	g12765 = NOT(I19829)
--	g12768 = NOT(g8829)
--	I19833 = NOT(g8726)
--	g12769 = NOT(I19833)
--	I19836 = NOT(g8726)
--	g12772 = NOT(I19836)
--	g12775 = NOT(g8832)
--	g12776 = NOT(g10766)
--	g12782 = NOT(g8836)
--	I19844 = NOT(g8533)
--	g12783 = NOT(I19844)
--	I19847 = NOT(g10677)
--	g12786 = NOT(I19847)
--	g12790 = NOT(g8847)
--	I19852 = NOT(g10679)
--	g12791 = NOT(I19852)
--	I19855 = NOT(g10723)
--	g12794 = NOT(I19855)
--	I19859 = NOT(g10617)
--	g12798 = NOT(I19859)
--	I19862 = NOT(g10725)
--	g12801 = NOT(I19862)
--	I19865 = NOT(g10354)
--	g12804 = NOT(I19865)
--	g12807 = NOT(g8853)
--	I19869 = NOT(g8726)
--	g12808 = NOT(I19869)
--	I19872 = NOT(g8317)
--	g12811 = NOT(I19872)
--	g12815 = NOT(g8856)
--	I19877 = NOT(g8547)
--	g12816 = NOT(I19877)
--	g12821 = NOT(g8863)
--	I19883 = NOT(g8550)
--	g12822 = NOT(I19883)
--	I19886 = NOT(g10706)
--	g12825 = NOT(I19886)
--	g12829 = NOT(g8874)
--	I19891 = NOT(g10708)
--	g12830 = NOT(I19891)
--	I19894 = NOT(g10744)
--	g12833 = NOT(I19894)
--	I19898 = NOT(g10664)
--	g12837 = NOT(I19898)
--	I19901 = NOT(g10746)
--	g12840 = NOT(I19901)
--	g12843 = NOT(g8879)
--	I19905 = NOT(g8726)
--	g12844 = NOT(I19905)
--	g12847 = NOT(g8882)
--	g12848 = NOT(g11059)
--	g12850 = NOT(g8885)
--	g12851 = NOT(g8888)
--	g12853 = NOT(g8894)
--	I19915 = NOT(g8560)
--	g12854 = NOT(I19915)
--	g12859 = NOT(g8901)
--	I19921 = NOT(g8563)
--	g12860 = NOT(I19921)
--	I19924 = NOT(g10726)
--	g12863 = NOT(I19924)
--	g12867 = NOT(g8912)
--	I19929 = NOT(g10728)
--	g12868 = NOT(I19929)
--	I19932 = NOT(g10763)
--	g12871 = NOT(I19932)
--	g12874 = NOT(g8915)
--	g12875 = NOT(g10779)
--	g12881 = NOT(g8918)
--	g12882 = NOT(g8921)
--	g12891 = NOT(g8925)
--	g12892 = NOT(g8928)
--	g12894 = NOT(g8934)
--	I19952 = NOT(g8571)
--	g12895 = NOT(I19952)
--	g12900 = NOT(g8941)
--	I19958 = NOT(g8574)
--	g12901 = NOT(I19958)
--	I19961 = NOT(g10747)
--	g12904 = NOT(I19961)
--	g12907 = NOT(g8949)
--	g12909 = NOT(g10904)
--	g12914 = NOT(g8952)
--	g12915 = NOT(g8955)
--	g12921 = NOT(g8958)
--	g12922 = NOT(g8961)
--	g12931 = NOT(g8965)
--	g12932 = NOT(g8968)
--	g12934 = NOT(g8974)
--	I19986 = NOT(g8577)
--	g12935 = NOT(I19986)
--	g12940 = NOT(g8980)
--	g12943 = NOT(g8984)
--	g12944 = NOT(g8987)
--	g12950 = NOT(g8990)
--	g12951 = NOT(g8993)
--	g12960 = NOT(g8997)
--	g12961 = NOT(g9000)
--	I20009 = NOT(g8313)
--	g12962 = NOT(I20009)
--	g12965 = NOT(g9006)
--	g12969 = NOT(g9010)
--	g12972 = NOT(g9013)
--	g12973 = NOT(g9016)
--	g12979 = NOT(g9019)
--	g12980 = NOT(g9022)
--	g12993 = NOT(g9035)
--	g12996 = NOT(g9038)
--	g12997 = NOT(g9041)
--	g12998 = NOT(g9044)
--	g13003 = NOT(g9058)
--	I20062 = NOT(g10480)
--	g13011 = NOT(I20062)
--	g13025 = NOT(g10810)
--	g13033 = NOT(g10797)
--	g13036 = NOT(g10831)
--	g13043 = NOT(g10789)
--	g13046 = NOT(g10814)
--	g13049 = NOT(g10851)
--	g13057 = NOT(g10784)
--	g13060 = NOT(g10801)
--	g13063 = NOT(g10835)
--	g13066 = NOT(g10872)
--	I20117 = NOT(g10876)
--	g13070 = NOT(I20117)
--	g13073 = NOT(g10793)
--	g13076 = NOT(g10818)
--	g13079 = NOT(g10855)
--	g13092 = NOT(g10805)
--	g13095 = NOT(g10839)
--	g13101 = NOT(g9128)
--	g13107 = NOT(g10822)
--	g13117 = NOT(g9134)
--	g13130 = NOT(g9140)
--	g13141 = NOT(g9146)
--	g13148 = NOT(g9170)
--	g13151 = NOT(g9184)
--	g13152 = NOT(g9196)
--	g13153 = NOT(g9199)
--	g13154 = NOT(g9212)
--	g13157 = NOT(g9229)
--	g13158 = NOT(g9242)
--	g13159 = NOT(g9245)
--	g13161 = NOT(g9257)
--	g13162 = NOT(g9260)
--	g13163 = NOT(g9273)
--	g13166 = NOT(g9290)
--	g13167 = NOT(g9303)
--	g13168 = NOT(g9306)
--	g13169 = NOT(g9320)
--	g13170 = NOT(g9323)
--	g13172 = NOT(g9335)
--	g13173 = NOT(g9338)
--	g13174 = NOT(g9351)
--	g13176 = NOT(g9368)
--	g13177 = NOT(g9371)
--	g13178 = NOT(g9384)
--	g13179 = NOT(g9387)
--	g13180 = NOT(g9401)
--	g13181 = NOT(g9404)
--	g13183 = NOT(g9416)
--	g13184 = NOT(g9419)
--	g13185 = NOT(g9443)
--	g13186 = NOT(g9446)
--	g13187 = NOT(g9450)
--	g13188 = NOT(g9465)
--	g13189 = NOT(g9468)
--	g13190 = NOT(g9481)
--	g13191 = NOT(g9484)
--	g13192 = NOT(g9498)
--	g13193 = NOT(g9501)
--	g13195 = NOT(g9524)
--	g13196 = NOT(g9528)
--	g13197 = NOT(g9531)
--	g13198 = NOT(g9585)
--	g13199 = NOT(g9588)
--	g13200 = NOT(g9592)
--	g13201 = NOT(g9607)
--	g13202 = NOT(g9610)
--	g13203 = NOT(g9623)
--	g13204 = NOT(g9626)
--	g13205 = NOT(g9641)
--	g13206 = NOT(g9644)
--	g13207 = NOT(g9666)
--	g13208 = NOT(g9670)
--	g13209 = NOT(g9673)
--	g13210 = NOT(g9727)
--	g13211 = NOT(g9730)
--	g13212 = NOT(g9734)
--	g13213 = NOT(g9749)
--	g13214 = NOT(g9752)
--	I20264 = NOT(g9027)
--	g13215 = NOT(I20264)
--	g13218 = NOT(g9767)
--	g13219 = NOT(g9770)
--	g13220 = NOT(g9787)
--	g13221 = NOT(g9790)
--	g13222 = NOT(g9812)
--	g13223 = NOT(g9816)
--	g13224 = NOT(g9819)
--	g13225 = NOT(g9873)
--	g13226 = NOT(g9876)
--	g13227 = NOT(g9880)
--	I20278 = NOT(g9027)
--	g13229 = NOT(I20278)
--	g13232 = NOT(g9895)
--	g13233 = NOT(g9898)
--	I20283 = NOT(g9050)
--	g13234 = NOT(I20283)
--	g13237 = NOT(g9913)
--	g13238 = NOT(g9916)
--	g13239 = NOT(g9933)
--	g13240 = NOT(g9936)
--	g13241 = NOT(g9958)
--	g13242 = NOT(g9962)
--	g13243 = NOT(g9965)
--	g13244 = NOT(g10004)
--	I20295 = NOT(g10015)
--	g13246 = NOT(I20295)
--	I20299 = NOT(g10800)
--	g13248 = NOT(I20299)
--	g13249 = NOT(g10018)
--	g13250 = NOT(g10021)
--	I20305 = NOT(g9050)
--	g13252 = NOT(I20305)
--	g13255 = NOT(g10049)
--	g13256 = NOT(g10052)
--	I20310 = NOT(g9067)
--	g13257 = NOT(I20310)
--	g13260 = NOT(g10067)
--	g13261 = NOT(g10070)
--	g13262 = NOT(g10087)
--	g13263 = NOT(g10090)
--	g13264 = NOT(g10096)
--	g13265 = NOT(g8568)
--	I20320 = NOT(g10792)
--	g13267 = NOT(I20320)
--	g13268 = NOT(g10109)
--	I20324 = NOT(g10124)
--	g13269 = NOT(I20324)
--	I20328 = NOT(g10817)
--	g13271 = NOT(I20328)
--	g13272 = NOT(g10127)
--	g13273 = NOT(g10130)
--	I20334 = NOT(g9067)
--	g13275 = NOT(I20334)
--	g13278 = NOT(g10158)
--	g13279 = NOT(g10161)
--	I20339 = NOT(g9084)
--	g13280 = NOT(I20339)
--	g13283 = NOT(g10176)
--	g13284 = NOT(g10179)
--	g13285 = NOT(g10189)
--	I20347 = NOT(g10787)
--	g13290 = NOT(I20347)
--	I20351 = NOT(g10804)
--	g13292 = NOT(I20351)
--	g13293 = NOT(g10214)
--	I20355 = NOT(g10229)
--	g13294 = NOT(I20355)
--	I20359 = NOT(g10838)
--	g13296 = NOT(I20359)
--	g13297 = NOT(g10232)
--	g13298 = NOT(g10235)
--	I20365 = NOT(g9084)
--	g13300 = NOT(I20365)
--	g13303 = NOT(g10263)
--	g13304 = NOT(g10266)
--	g13308 = NOT(g10273)
--	g13309 = NOT(g10276)
--	I20376 = NOT(g8569)
--	g13317 = NOT(I20376)
--	I20379 = NOT(g11213)
--	g13318 = NOT(I20379)
--	I20382 = NOT(g10907)
--	g13319 = NOT(I20382)
--	I20386 = NOT(g10796)
--	g13321 = NOT(I20386)
--	I20390 = NOT(g10821)
--	g13323 = NOT(I20390)
--	g13324 = NOT(g10316)
--	I20394 = NOT(g10331)
--	g13325 = NOT(I20394)
--	I20398 = NOT(g10858)
--	g13327 = NOT(I20398)
--	g13328 = NOT(g10334)
--	g13329 = NOT(g10337)
--	g13330 = NOT(g10357)
--	I20407 = NOT(g9027)
--	g13336 = NOT(I20407)
--	I20410 = NOT(g10887)
--	g13339 = NOT(I20410)
--	I20414 = NOT(g8575)
--	g13341 = NOT(I20414)
--	I20417 = NOT(g10933)
--	g13342 = NOT(I20417)
--	I20421 = NOT(g10808)
--	g13344 = NOT(I20421)
--	I20425 = NOT(g10842)
--	g13346 = NOT(I20425)
--	g13347 = NOT(g10409)
--	g13351 = NOT(g10416)
--	g13352 = NOT(g10419)
--	I20441 = NOT(g9027)
--	g13356 = NOT(I20441)
--	I20444 = NOT(g10869)
--	g13359 = NOT(I20444)
--	I20448 = NOT(g9050)
--	g13361 = NOT(I20448)
--	I20451 = NOT(g10908)
--	g13364 = NOT(I20451)
--	I20455 = NOT(g8578)
--	g13366 = NOT(I20455)
--	I20458 = NOT(g10972)
--	g13367 = NOT(I20458)
--	I20462 = NOT(g10825)
--	g13369 = NOT(I20462)
--	g13373 = NOT(g10482)
--	I20476 = NOT(g9027)
--	g13381 = NOT(I20476)
--	I20479 = NOT(g10849)
--	g13384 = NOT(I20479)
--	I20483 = NOT(g9050)
--	g13386 = NOT(I20483)
--	I20486 = NOT(g10889)
--	g13389 = NOT(I20486)
--	I20490 = NOT(g9067)
--	g13391 = NOT(I20490)
--	I20493 = NOT(g10934)
--	g13394 = NOT(I20493)
--	I20497 = NOT(g8579)
--	g13396 = NOT(I20497)
--	I20500 = NOT(g11007)
--	g13397 = NOT(I20500)
--	g13398 = NOT(g10542)
--	g13400 = NOT(g10545)
--	I20514 = NOT(g11769)
--	g13405 = NOT(I20514)
--	I20517 = NOT(g12425)
--	g13406 = NOT(I20517)
--	I20520 = NOT(g13246)
--	g13407 = NOT(I20520)
--	I20523 = NOT(g13317)
--	g13408 = NOT(I20523)
--	I20526 = NOT(g12519)
--	g13409 = NOT(I20526)
--	I20529 = NOT(g13319)
--	g13410 = NOT(I20529)
--	I20532 = NOT(g13339)
--	g13411 = NOT(I20532)
--	I20535 = NOT(g13359)
--	g13412 = NOT(I20535)
--	I20538 = NOT(g13384)
--	g13413 = NOT(I20538)
--	I20541 = NOT(g11599)
--	g13414 = NOT(I20541)
--	I20544 = NOT(g11628)
--	g13415 = NOT(I20544)
--	I20547 = NOT(g13248)
--	g13416 = NOT(I20547)
--	I20550 = NOT(g13267)
--	g13417 = NOT(I20550)
--	I20553 = NOT(g13290)
--	g13418 = NOT(I20553)
--	I20556 = NOT(g12435)
--	g13419 = NOT(I20556)
--	I20559 = NOT(g11937)
--	g13420 = NOT(I20559)
--	I20562 = NOT(g11786)
--	g13421 = NOT(I20562)
--	I20565 = NOT(g12432)
--	g13422 = NOT(I20565)
--	I20568 = NOT(g13269)
--	g13423 = NOT(I20568)
--	I20571 = NOT(g13341)
--	g13424 = NOT(I20571)
--	I20574 = NOT(g12534)
--	g13425 = NOT(I20574)
--	I20577 = NOT(g13342)
--	g13426 = NOT(I20577)
--	I20580 = NOT(g13364)
--	g13427 = NOT(I20580)
--	I20583 = NOT(g13389)
--	g13428 = NOT(I20583)
--	I20586 = NOT(g11606)
--	g13429 = NOT(I20586)
--	I20589 = NOT(g11629)
--	g13430 = NOT(I20589)
--	I20592 = NOT(g11651)
--	g13431 = NOT(I20592)
--	I20595 = NOT(g13271)
--	g13432 = NOT(I20595)
--	I20598 = NOT(g13292)
--	g13433 = NOT(I20598)
--	I20601 = NOT(g13321)
--	g13434 = NOT(I20601)
--	I20604 = NOT(g12440)
--	g13435 = NOT(I20604)
--	I20607 = NOT(g11990)
--	g13436 = NOT(I20607)
--	I20610 = NOT(g11812)
--	g13437 = NOT(I20610)
--	I20613 = NOT(g12437)
--	g13438 = NOT(I20613)
--	I20616 = NOT(g13294)
--	g13439 = NOT(I20616)
--	I20619 = NOT(g13366)
--	g13440 = NOT(I20619)
--	I20622 = NOT(g12543)
--	g13441 = NOT(I20622)
--	I20625 = NOT(g13367)
--	g13442 = NOT(I20625)
--	I20628 = NOT(g13394)
--	g13443 = NOT(I20628)
--	I20631 = NOT(g11611)
--	g13444 = NOT(I20631)
--	I20634 = NOT(g11636)
--	g13445 = NOT(I20634)
--	I20637 = NOT(g11652)
--	g13446 = NOT(I20637)
--	I20640 = NOT(g11670)
--	g13447 = NOT(I20640)
--	I20643 = NOT(g13296)
--	g13448 = NOT(I20643)
--	I20646 = NOT(g13323)
--	g13449 = NOT(I20646)
--	I20649 = NOT(g13344)
--	g13450 = NOT(I20649)
--	I20652 = NOT(g12445)
--	g13451 = NOT(I20652)
--	I20655 = NOT(g12059)
--	g13452 = NOT(I20655)
--	I20658 = NOT(g11845)
--	g13453 = NOT(I20658)
--	I20661 = NOT(g12442)
--	g13454 = NOT(I20661)
--	I20664 = NOT(g13325)
--	g13455 = NOT(I20664)
--	I20667 = NOT(g13396)
--	g13456 = NOT(I20667)
--	I20670 = NOT(g12552)
--	g13457 = NOT(I20670)
--	I20673 = NOT(g13397)
--	g13458 = NOT(I20673)
--	I20676 = NOT(g11616)
--	g13459 = NOT(I20676)
--	I20679 = NOT(g11641)
--	g13460 = NOT(I20679)
--	I20682 = NOT(g11659)
--	g13461 = NOT(I20682)
--	I20685 = NOT(g11671)
--	g13462 = NOT(I20685)
--	I20688 = NOT(g11682)
--	g13463 = NOT(I20688)
--	I20691 = NOT(g13327)
--	g13464 = NOT(I20691)
--	I20694 = NOT(g13346)
--	g13465 = NOT(I20694)
--	I20697 = NOT(g13369)
--	g13466 = NOT(I20697)
--	I20700 = NOT(g12450)
--	g13467 = NOT(I20700)
--	I20703 = NOT(g12123)
--	g13468 = NOT(I20703)
--	I20706 = NOT(g11490)
--	g13469 = NOT(I20706)
--	I20709 = NOT(g13070)
--	g13475 = NOT(I20709)
--	g13519 = NOT(g13228)
--	g13530 = NOT(g13251)
--	g13541 = NOT(g13274)
--	g13552 = NOT(g13299)
--	g13565 = NOT(g12192)
--	g13568 = NOT(g11627)
--	I20791 = NOT(g13149)
--	g13571 = NOT(I20791)
--	I20794 = NOT(g13111)
--	g13572 = NOT(I20794)
--	g13573 = NOT(g12247)
--	g13576 = NOT(g11650)
--	I20799 = NOT(g13155)
--	g13579 = NOT(I20799)
--	I20802 = NOT(g13160)
--	g13580 = NOT(I20802)
--	I20805 = NOT(g13124)
--	g13581 = NOT(I20805)
--	g13582 = NOT(g12290)
--	g13585 = NOT(g11669)
--	I20810 = NOT(g13164)
--	g13588 = NOT(I20810)
--	I20813 = NOT(g13265)
--	g13589 = NOT(I20813)
--	I20816 = NOT(g12487)
--	g13598 = NOT(I20816)
--	I20820 = NOT(g13171)
--	g13600 = NOT(I20820)
--	I20823 = NOT(g13135)
--	g13601 = NOT(I20823)
--	g13602 = NOT(g12326)
--	g13605 = NOT(g11681)
--	I20828 = NOT(g13175)
--	g13608 = NOT(I20828)
--	I20832 = NOT(g12507)
--	g13610 = NOT(I20832)
--	I20836 = NOT(g13182)
--	g13612 = NOT(I20836)
--	I20839 = NOT(g13143)
--	g13613 = NOT(I20839)
--	g13614 = NOT(g11690)
--	I20844 = NOT(g12524)
--	g13620 = NOT(I20844)
--	I20848 = NOT(g13194)
--	g13622 = NOT(I20848)
--	I20852 = NOT(g12457)
--	g13624 = NOT(I20852)
--	g13626 = NOT(g11697)
--	I20858 = NOT(g12539)
--	g13632 = NOT(I20858)
--	I20863 = NOT(g12467)
--	g13635 = NOT(I20863)
--	g13637 = NOT(g11703)
--	g13644 = NOT(g13215)
--	I20873 = NOT(g12482)
--	g13647 = NOT(I20873)
--	g13649 = NOT(g11711)
--	g13657 = NOT(g12452)
--	g13669 = NOT(g13229)
--	g13670 = NOT(g13234)
--	I20886 = NOT(g12499)
--	g13673 = NOT(I20886)
--	g13677 = NOT(g12447)
--	g13687 = NOT(g12460)
--	g13699 = NOT(g13252)
--	g13700 = NOT(g13257)
--	g13706 = NOT(g12443)
--	g13714 = NOT(g12453)
--	g13724 = NOT(g12470)
--	g13736 = NOT(g13275)
--	g13737 = NOT(g13280)
--	I20909 = NOT(g13055)
--	g13741 = NOT(I20909)
--	g13750 = NOT(g12439)
--	g13756 = NOT(g12448)
--	g13764 = NOT(g12461)
--	g13774 = NOT(g12485)
--	g13786 = NOT(g13300)
--	g13791 = NOT(g12444)
--	g13797 = NOT(g12454)
--	g13805 = NOT(g12471)
--	g13817 = NOT(g13336)
--	g13819 = NOT(g12449)
--	g13825 = NOT(g12462)
--	g13836 = NOT(g13356)
--	g13838 = NOT(g13361)
--	g13840 = NOT(g12455)
--	g13848 = NOT(g11744)
--	g13849 = NOT(g13381)
--	g13850 = NOT(g13386)
--	g13852 = NOT(g13391)
--	g13856 = NOT(g11759)
--	g13857 = NOT(g11760)
--	g13858 = NOT(g11603)
--	g13859 = NOT(g11608)
--	g13861 = NOT(g11613)
--	I20959 = NOT(g11713)
--	g13863 = NOT(I20959)
--	g13864 = NOT(g11767)
--	g13866 = NOT(g11772)
--	g13867 = NOT(g11773)
--	g13868 = NOT(g11633)
--	g13869 = NOT(g11638)
--	g13872 = NOT(g11780)
--	g13873 = NOT(g12698)
--	g13879 = NOT(g11784)
--	g13881 = NOT(g11789)
--	g13882 = NOT(g11790)
--	g13883 = NOT(g11656)
--	g13885 = NOT(g11799)
--	g13886 = NOT(g12747)
--	g13894 = NOT(g11806)
--	g13895 = NOT(g12755)
--	g13901 = NOT(g11810)
--	g13903 = NOT(g11815)
--	g13906 = NOT(g11822)
--	g13907 = NOT(g12781)
--	g13918 = NOT(g11830)
--	g13922 = NOT(g11831)
--	g13926 = NOT(g11832)
--	g13927 = NOT(g12789)
--	g13935 = NOT(g11839)
--	g13936 = NOT(g12797)
--	g13942 = NOT(g11843)
--	g13945 = NOT(g11855)
--	g13946 = NOT(g12814)
--	I21012 = NOT(g12503)
--	g13954 = NOT(I21012)
--	g13958 = NOT(g11863)
--	g13962 = NOT(g11864)
--	g13963 = NOT(g12820)
--	g13974 = NOT(g11872)
--	g13978 = NOT(g11873)
--	g13982 = NOT(g11874)
--	g13983 = NOT(g12828)
--	g13991 = NOT(g11881)
--	g13992 = NOT(g12836)
--	g13999 = NOT(g11889)
--	g14000 = NOT(g11890)
--	g14001 = NOT(g12849)
--	I21037 = NOT(g12486)
--	g14008 = NOT(I21037)
--	g14011 = NOT(g11896)
--	g14015 = NOT(g11897)
--	g14016 = NOT(g12852)
--	I21045 = NOT(g12520)
--	g14024 = NOT(I21045)
--	g14028 = NOT(g11905)
--	g14032 = NOT(g11906)
--	g14033 = NOT(g12858)
--	g14044 = NOT(g11914)
--	g14048 = NOT(g11915)
--	g14052 = NOT(g11916)
--	g14053 = NOT(g12866)
--	g14061 = NOT(g11928)
--	g14062 = NOT(g12880)
--	I21064 = NOT(g13147)
--	g14068 = NOT(I21064)
--	g14071 = NOT(g11934)
--	g14079 = NOT(g11935)
--	g14086 = NOT(g11938)
--	g14090 = NOT(g11939)
--	g14091 = NOT(g11940)
--	g14092 = NOT(g12890)
--	I21075 = NOT(g12506)
--	g14099 = NOT(I21075)
--	g14102 = NOT(g11946)
--	g14106 = NOT(g11947)
--	g14107 = NOT(g12893)
--	I21083 = NOT(g12535)
--	g14115 = NOT(I21083)
--	g14119 = NOT(g11955)
--	g14123 = NOT(g11956)
--	g14124 = NOT(g12899)
--	g14135 = NOT(g11964)
--	g14139 = NOT(g11965)
--	I21096 = NOT(g11749)
--	g14144 = NOT(I21096)
--	g14148 = NOT(g12912)
--	g14153 = NOT(g12913)
--	g14158 = NOT(g11974)
--	g14165 = NOT(g11975)
--	g14171 = NOT(g11979)
--	g14175 = NOT(g11980)
--	g14176 = NOT(g11981)
--	g14177 = NOT(g12920)
--	I21108 = NOT(g13150)
--	g14183 = NOT(I21108)
--	g14186 = NOT(g11987)
--	g14194 = NOT(g11988)
--	g14201 = NOT(g11991)
--	g14205 = NOT(g11992)
--	g14206 = NOT(g11993)
--	g14207 = NOT(g12930)
--	I21119 = NOT(g12523)
--	g14214 = NOT(I21119)
--	g14217 = NOT(g11999)
--	g14221 = NOT(g12000)
--	g14222 = NOT(g12933)
--	I21127 = NOT(g12544)
--	g14230 = NOT(I21127)
--	g14234 = NOT(g12008)
--	g14238 = NOT(g12939)
--	g14244 = NOT(g12026)
--	g14249 = NOT(g12034)
--	g14252 = NOT(g12035)
--	g14256 = NOT(g12036)
--	I21137 = NOT(g11749)
--	g14259 = NOT(I21137)
--	g14263 = NOT(g12941)
--	g14268 = NOT(g12942)
--	g14273 = NOT(g12043)
--	g14280 = NOT(g12044)
--	g14286 = NOT(g12048)
--	g14290 = NOT(g12049)
--	g14291 = NOT(g12050)
--	g14292 = NOT(g12949)
--	I21149 = NOT(g13156)
--	g14298 = NOT(I21149)
--	g14301 = NOT(g12056)
--	g14309 = NOT(g12057)
--	g14316 = NOT(g12060)
--	g14320 = NOT(g12061)
--	g14321 = NOT(g12062)
--	g14322 = NOT(g12959)
--	I21160 = NOT(g12538)
--	g14329 = NOT(I21160)
--	g14332 = NOT(g12068)
--	I21165 = NOT(g13110)
--	g14337 = NOT(I21165)
--	g14342 = NOT(g12967)
--	g14347 = NOT(g12079)
--	g14352 = NOT(g12081)
--	g14355 = NOT(g12082)
--	g14359 = NOT(g12083)
--	g14360 = NOT(g12968)
--	g14366 = NOT(g12090)
--	g14371 = NOT(g12098)
--	g14374 = NOT(g12099)
--	g14378 = NOT(g12100)
--	I21178 = NOT(g11749)
--	g14381 = NOT(I21178)
--	g14385 = NOT(g12970)
--	g14390 = NOT(g12971)
--	g14395 = NOT(g12107)
--	g14402 = NOT(g12108)
--	g14408 = NOT(g12112)
--	g14412 = NOT(g12113)
--	g14413 = NOT(g12114)
--	g14414 = NOT(g12978)
--	I21190 = NOT(g13165)
--	g14420 = NOT(I21190)
--	g14423 = NOT(g12120)
--	g14431 = NOT(g12121)
--	g14438 = NOT(g12124)
--	g14442 = NOT(g11768)
--	g14450 = NOT(g12146)
--	g14454 = NOT(g12991)
--	g14459 = NOT(g12151)
--	g14464 = NOT(g12153)
--	g14467 = NOT(g12154)
--	g14471 = NOT(g12155)
--	g14472 = NOT(g12992)
--	g14478 = NOT(g12162)
--	g14483 = NOT(g12170)
--	g14486 = NOT(g12171)
--	g14490 = NOT(g12172)
--	I21208 = NOT(g11749)
--	g14493 = NOT(I21208)
--	g14497 = NOT(g12994)
--	g14502 = NOT(g12995)
--	g14507 = NOT(g12179)
--	g14514 = NOT(g12180)
--	g14520 = NOT(g12184)
--	g14524 = NOT(g12185)
--	g14525 = NOT(g12195)
--	g14529 = NOT(g11785)
--	g14537 = NOT(g12208)
--	g14541 = NOT(g13001)
--	g14546 = NOT(g12213)
--	g14551 = NOT(g12215)
--	g14554 = NOT(g12216)
--	g14558 = NOT(g12217)
--	g14559 = NOT(g13002)
--	g14565 = NOT(g12224)
--	g14570 = NOT(g12232)
--	g14573 = NOT(g12233)
--	g14577 = NOT(g12234)
--	g14580 = NOT(g12250)
--	g14584 = NOT(g11811)
--	g14592 = NOT(g12263)
--	g14596 = NOT(g13022)
--	g14601 = NOT(g12268)
--	g14606 = NOT(g12270)
--	g14609 = NOT(g12271)
--	g14613 = NOT(g12272)
--	g14614 = NOT(g12293)
--	g14618 = NOT(g11844)
--	g14626 = NOT(g12306)
--	I21241 = NOT(g13378)
--	g14630 = NOT(I21241)
--	g14637 = NOT(g12329)
--	g14641 = NOT(g11823)
--	I21246 = NOT(g11624)
--	g14642 = NOT(I21246)
--	I21249 = NOT(g11600)
--	g14650 = NOT(I21249)
--	I21252 = NOT(g11644)
--	g14657 = NOT(I21252)
--	g14668 = NOT(g11865)
--	I21256 = NOT(g11647)
--	g14669 = NOT(I21256)
--	I21259 = NOT(g11630)
--	g14677 = NOT(I21259)
--	I21262 = NOT(g11713)
--	g14684 = NOT(I21262)
--	g14685 = NOT(g12245)
--	I21267 = NOT(g11663)
--	g14691 = NOT(I21267)
--	g14702 = NOT(g11907)
--	I21271 = NOT(g11666)
--	g14703 = NOT(I21271)
--	I21274 = NOT(g11653)
--	g14711 = NOT(I21274)
--	I21277 = NOT(g12430)
--	g14718 = NOT(I21277)
--	g14719 = NOT(g12288)
--	I21282 = NOT(g11675)
--	g14725 = NOT(I21282)
--	g14736 = NOT(g11957)
--	I21286 = NOT(g11678)
--	g14737 = NOT(I21286)
--	I21289 = NOT(g12434)
--	g14745 = NOT(I21289)
--	I21292 = NOT(g11888)
--	g14746 = NOT(I21292)
--	g14747 = NOT(g12324)
--	I21297 = NOT(g11687)
--	g14753 = NOT(I21297)
--	g14764 = NOT(g11791)
--	I21301 = NOT(g12438)
--	g14765 = NOT(I21301)
--	I21304 = NOT(g11927)
--	g14766 = NOT(I21304)
--	g14768 = NOT(g12352)
--	I21310 = NOT(g12332)
--	g14774 = NOT(I21310)
--	I21313 = NOT(g11743)
--	g14775 = NOT(I21313)
--	g14776 = NOT(g12033)
--	g14794 = NOT(g11848)
--	I21318 = NOT(g12362)
--	g14795 = NOT(I21318)
--	I21321 = NOT(g11758)
--	g14796 = NOT(I21321)
--	g14797 = NOT(g12080)
--	g14811 = NOT(g12097)
--	I21326 = NOT(g12378)
--	g14829 = NOT(I21326)
--	I21329 = NOT(g11766)
--	g14830 = NOT(I21329)
--	g14831 = NOT(g11828)
--	g14837 = NOT(g12145)
--	g14849 = NOT(g12152)
--	g14863 = NOT(g12169)
--	g14881 = NOT(g11923)
--	I21337 = NOT(g12408)
--	g14882 = NOT(I21337)
--	I21340 = NOT(g11779)
--	g14883 = NOT(I21340)
--	g14885 = NOT(g11860)
--	g14895 = NOT(g12193)
--	g14904 = NOT(g11870)
--	g14910 = NOT(g12207)
--	g14922 = NOT(g12214)
--	g14936 = NOT(g12231)
--	I21351 = NOT(g12420)
--	g14954 = NOT(I21351)
--	I21354 = NOT(g11798)
--	g14955 = NOT(I21354)
--	g14959 = NOT(g11976)
--	I21361 = NOT(g13026)
--	g14960 = NOT(I21361)
--	I21364 = NOT(g13028)
--	g14963 = NOT(I21364)
--	g14966 = NOT(g11902)
--	g14976 = NOT(g12248)
--	g14985 = NOT(g11912)
--	g14991 = NOT(g12262)
--	g15003 = NOT(g12269)
--	g15017 = NOT(g12009)
--	I21374 = NOT(g12424)
--	g15018 = NOT(I21374)
--	I21377 = NOT(g11821)
--	g15019 = NOT(I21377)
--	I21381 = NOT(g13157)
--	g15021 = NOT(I21381)
--	g15022 = NOT(g11781)
--	g15032 = NOT(g12027)
--	g15033 = NOT(g12030)
--	I21389 = NOT(g12883)
--	g15034 = NOT(I21389)
--	I21392 = NOT(g13020)
--	g15037 = NOT(I21392)
--	I21395 = NOT(g13034)
--	g15040 = NOT(I21395)
--	I21398 = NOT(g13021)
--	g15043 = NOT(I21398)
--	g15048 = NOT(g12045)
--	I21404 = NOT(g13037)
--	g15049 = NOT(I21404)
--	I21407 = NOT(g13039)
--	g15052 = NOT(I21407)
--	g15055 = NOT(g11952)
--	g15065 = NOT(g12291)
--	g15074 = NOT(g11962)
--	g15080 = NOT(g12305)
--	I21415 = NOT(g11854)
--	g15092 = NOT(I21415)
--	I21420 = NOT(g13166)
--	g15095 = NOT(I21420)
--	g15096 = NOT(g11800)
--	I21426 = NOT(g11661)
--	g15106 = NOT(I21426)
--	I21429 = NOT(g13027)
--	g15109 = NOT(I21429)
--	I21432 = NOT(g13044)
--	g15112 = NOT(I21432)
--	I21435 = NOT(g11662)
--	g15115 = NOT(I21435)
--	g15118 = NOT(g11807)
--	g15128 = NOT(g12091)
--	g15129 = NOT(g12094)
--	I21443 = NOT(g12923)
--	g15130 = NOT(I21443)
--	I21446 = NOT(g13029)
--	g15133 = NOT(I21446)
--	I21449 = NOT(g13047)
--	g15136 = NOT(I21449)
--	I21452 = NOT(g13030)
--	g15139 = NOT(I21452)
--	g15144 = NOT(g12109)
--	I21458 = NOT(g13050)
--	g15145 = NOT(I21458)
--	I21461 = NOT(g13052)
--	g15148 = NOT(I21461)
--	g15151 = NOT(g12005)
--	g15161 = NOT(g12327)
--	g15170 = NOT(g12125)
--	g15174 = NOT(g12136)
--	g15175 = NOT(g12139)
--	g15176 = NOT(g12142)
--	g15177 = NOT(g12339)
--	I21476 = NOT(g11672)
--	g15179 = NOT(I21476)
--	I21479 = NOT(g13035)
--	g15182 = NOT(I21479)
--	I21482 = NOT(g13058)
--	g15185 = NOT(I21482)
--	g15188 = NOT(g11833)
--	I21488 = NOT(g11673)
--	g15198 = NOT(I21488)
--	I21491 = NOT(g13038)
--	g15201 = NOT(I21491)
--	I21494 = NOT(g13061)
--	g15204 = NOT(I21494)
--	I21497 = NOT(g11674)
--	g15207 = NOT(I21497)
--	g15210 = NOT(g11840)
--	g15220 = NOT(g12163)
--	g15221 = NOT(g12166)
--	I21505 = NOT(g12952)
--	g15222 = NOT(I21505)
--	I21508 = NOT(g13040)
--	g15225 = NOT(I21508)
--	I21511 = NOT(g13064)
--	g15228 = NOT(I21511)
--	I21514 = NOT(g13041)
--	g15231 = NOT(I21514)
--	g15236 = NOT(g12181)
--	I21520 = NOT(g13067)
--	g15237 = NOT(I21520)
--	I21523 = NOT(g13069)
--	g15240 = NOT(I21523)
--	I21531 = NOT(g11683)
--	g15248 = NOT(I21531)
--	I21534 = NOT(g13045)
--	g15251 = NOT(I21534)
--	I21537 = NOT(g13071)
--	g15254 = NOT(I21537)
--	g15260 = NOT(g12198)
--	g15261 = NOT(g12201)
--	g15262 = NOT(g12204)
--	g15263 = NOT(g12369)
--	I21548 = NOT(g11684)
--	g15265 = NOT(I21548)
--	I21551 = NOT(g13048)
--	g15268 = NOT(I21551)
--	I21554 = NOT(g13074)
--	g15271 = NOT(I21554)
--	g15274 = NOT(g11875)
--	I21560 = NOT(g11685)
--	g15284 = NOT(I21560)
--	I21563 = NOT(g13051)
--	g15287 = NOT(I21563)
--	I21566 = NOT(g13077)
--	g15290 = NOT(I21566)
--	I21569 = NOT(g11686)
--	g15293 = NOT(I21569)
--	g15296 = NOT(g11882)
--	g15306 = NOT(g12225)
--	g15307 = NOT(g12228)
--	I21577 = NOT(g12981)
--	g15308 = NOT(I21577)
--	I21580 = NOT(g13053)
--	g15311 = NOT(I21580)
--	I21583 = NOT(g13080)
--	g15314 = NOT(I21583)
--	I21586 = NOT(g13054)
--	g15317 = NOT(I21586)
--	g15322 = NOT(g12239)
--	g15323 = NOT(g12242)
--	I21595 = NOT(g11691)
--	g15326 = NOT(I21595)
--	I21598 = NOT(g13059)
--	g15329 = NOT(I21598)
--	I21601 = NOT(g13087)
--	g15332 = NOT(I21601)
--	I21609 = NOT(g11692)
--	g15340 = NOT(I21609)
--	I21612 = NOT(g13062)
--	g15343 = NOT(I21612)
--	I21615 = NOT(g13090)
--	g15346 = NOT(I21615)
--	g15352 = NOT(g12253)
--	g15353 = NOT(g12256)
--	g15354 = NOT(g12259)
--	g15355 = NOT(g12388)
--	I21626 = NOT(g11693)
--	g15357 = NOT(I21626)
--	I21629 = NOT(g13065)
--	g15360 = NOT(I21629)
--	I21632 = NOT(g13093)
--	g15363 = NOT(I21632)
--	g15366 = NOT(g11917)
--	I21638 = NOT(g11694)
--	g15376 = NOT(I21638)
--	I21641 = NOT(g13068)
--	g15379 = NOT(I21641)
--	I21644 = NOT(g13096)
--	g15382 = NOT(I21644)
--	I21647 = NOT(g11695)
--	g15385 = NOT(I21647)
--	g15390 = NOT(g12279)
--	I21655 = NOT(g11696)
--	g15393 = NOT(I21655)
--	I21658 = NOT(g13072)
--	g15396 = NOT(I21658)
--	I21661 = NOT(g13098)
--	g15399 = NOT(I21661)
--	I21666 = NOT(g13100)
--	g15404 = NOT(I21666)
--	g15408 = NOT(g12282)
--	g15409 = NOT(g12285)
--	I21674 = NOT(g11698)
--	g15412 = NOT(I21674)
--	I21677 = NOT(g13075)
--	g15415 = NOT(I21677)
--	I21680 = NOT(g13102)
--	g15418 = NOT(I21680)
--	I21688 = NOT(g11699)
--	g15426 = NOT(I21688)
--	I21691 = NOT(g13078)
--	g15429 = NOT(I21691)
--	I21694 = NOT(g13105)
--	g15432 = NOT(I21694)
--	g15438 = NOT(g12296)
--	g15439 = NOT(g12299)
--	g15440 = NOT(g12302)
--	g15441 = NOT(g12418)
--	I21705 = NOT(g11700)
--	g15443 = NOT(I21705)
--	I21708 = NOT(g13081)
--	g15446 = NOT(I21708)
--	I21711 = NOT(g13108)
--	g15449 = NOT(I21711)
--	g15458 = NOT(g12312)
--	I21720 = NOT(g11701)
--	g15461 = NOT(I21720)
--	I21723 = NOT(g13088)
--	g15464 = NOT(I21723)
--	I21726 = NOT(g13112)
--	g15467 = NOT(I21726)
--	I21730 = NOT(g13089)
--	g15471 = NOT(I21730)
--	g15474 = NOT(g12315)
--	I21736 = NOT(g11702)
--	g15477 = NOT(I21736)
--	I21739 = NOT(g13091)
--	g15480 = NOT(I21739)
--	I21742 = NOT(g13114)
--	g15483 = NOT(I21742)
--	I21747 = NOT(g13116)
--	g15488 = NOT(I21747)
--	g15492 = NOT(g12318)
--	g15493 = NOT(g12321)
--	I21755 = NOT(g11704)
--	g15496 = NOT(I21755)
--	I21758 = NOT(g13094)
--	g15499 = NOT(I21758)
--	I21761 = NOT(g13118)
--	g15502 = NOT(I21761)
--	I21769 = NOT(g11705)
--	g15510 = NOT(I21769)
--	I21772 = NOT(g13097)
--	g15513 = NOT(I21772)
--	I21775 = NOT(g13121)
--	g15516 = NOT(I21775)
--	I21780 = NOT(g13305)
--	g15521 = NOT(I21780)
--	g15524 = NOT(g12333)
--	g15525 = NOT(g12336)
--	I21787 = NOT(g11707)
--	g15528 = NOT(I21787)
--	I21790 = NOT(g13099)
--	g15531 = NOT(I21790)
--	I21793 = NOT(g13123)
--	g15534 = NOT(I21793)
--	I21796 = NOT(g11708)
--	g15537 = NOT(I21796)
--	g15544 = NOT(g12340)
--	I21803 = NOT(g11709)
--	g15547 = NOT(I21803)
--	I21806 = NOT(g13103)
--	g15550 = NOT(I21806)
--	I21809 = NOT(g13125)
--	g15553 = NOT(I21809)
--	I21813 = NOT(g13104)
--	g15557 = NOT(I21813)
--	g15560 = NOT(g12343)
--	I21819 = NOT(g11710)
--	g15563 = NOT(I21819)
--	I21822 = NOT(g13106)
--	g15566 = NOT(I21822)
--	I21825 = NOT(g13127)
--	g15569 = NOT(I21825)
--	I21830 = NOT(g13129)
--	g15574 = NOT(I21830)
--	g15578 = NOT(g12346)
--	g15579 = NOT(g12349)
--	I21838 = NOT(g11712)
--	g15582 = NOT(I21838)
--	I21841 = NOT(g13109)
--	g15585 = NOT(I21841)
--	I21844 = NOT(g13131)
--	g15588 = NOT(I21844)
--	I21852 = NOT(g11716)
--	g15596 = NOT(I21852)
--	I21855 = NOT(g13113)
--	g15599 = NOT(I21855)
--	g15602 = NOT(g12363)
--	g15603 = NOT(g12366)
--	I21862 = NOT(g11717)
--	g15606 = NOT(I21862)
--	I21865 = NOT(g13115)
--	g15609 = NOT(I21865)
--	I21868 = NOT(g13134)
--	g15612 = NOT(I21868)
--	I21871 = NOT(g11718)
--	g15615 = NOT(I21871)
--	g15622 = NOT(g12370)
--	I21878 = NOT(g11719)
--	g15625 = NOT(I21878)
--	I21881 = NOT(g13119)
--	g15628 = NOT(I21881)
--	I21884 = NOT(g13136)
--	g15631 = NOT(I21884)
--	I21888 = NOT(g13120)
--	g15635 = NOT(I21888)
--	g15638 = NOT(g12373)
--	I21894 = NOT(g11720)
--	g15641 = NOT(I21894)
--	I21897 = NOT(g13122)
--	g15644 = NOT(I21897)
--	I21900 = NOT(g13138)
--	g15647 = NOT(I21900)
--	I21905 = NOT(g13140)
--	g15652 = NOT(I21905)
--	I21908 = NOT(g13082)
--	g15655 = NOT(I21908)
--	g15659 = NOT(g11706)
--	g15665 = NOT(g12379)
--	I21918 = NOT(g11721)
--	g15667 = NOT(I21918)
--	I21923 = NOT(g11722)
--	g15672 = NOT(I21923)
--	I21926 = NOT(g13126)
--	g15675 = NOT(I21926)
--	g15678 = NOT(g12382)
--	g15679 = NOT(g12385)
--	I21933 = NOT(g11723)
--	g15682 = NOT(I21933)
--	I21936 = NOT(g13128)
--	g15685 = NOT(I21936)
--	I21939 = NOT(g13142)
--	g15688 = NOT(I21939)
--	I21942 = NOT(g11724)
--	g15691 = NOT(I21942)
--	g15698 = NOT(g12389)
--	I21949 = NOT(g11725)
--	g15701 = NOT(I21949)
--	I21952 = NOT(g13132)
--	g15704 = NOT(I21952)
--	I21955 = NOT(g13144)
--	g15707 = NOT(I21955)
--	I21959 = NOT(g13133)
--	g15711 = NOT(I21959)
--	I21962 = NOT(g13004)
--	g15714 = NOT(I21962)
--	g15722 = NOT(g13011)
--	g15724 = NOT(g12409)
--	I21974 = NOT(g11726)
--	g15726 = NOT(I21974)
--	I21979 = NOT(g11727)
--	g15731 = NOT(I21979)
--	I21982 = NOT(g13137)
--	g15734 = NOT(I21982)
--	g15737 = NOT(g12412)
--	g15738 = NOT(g12415)
--	I21989 = NOT(g11728)
--	g15741 = NOT(I21989)
--	I21992 = NOT(g13139)
--	g15744 = NOT(I21992)
--	I21995 = NOT(g13146)
--	g15747 = NOT(I21995)
--	I21998 = NOT(g11729)
--	g15750 = NOT(I21998)
--	g15762 = NOT(g13011)
--	g15764 = NOT(g12421)
--	I22014 = NOT(g11730)
--	g15766 = NOT(I22014)
--	I22019 = NOT(g11731)
--	g15771 = NOT(I22019)
--	I22022 = NOT(g13145)
--	g15774 = NOT(I22022)
--	I22025 = NOT(g11617)
--	g15777 = NOT(I22025)
--	g15790 = NOT(g13011)
--	g15792 = NOT(g12426)
--	I22044 = NOT(g11733)
--	g15794 = NOT(I22044)
--	g15800 = NOT(g12909)
--	g15813 = NOT(g13011)
--	g15859 = NOT(g13378)
--	I22120 = NOT(g12909)
--	g15876 = NOT(I22120)
--	g15880 = NOT(g11624)
--	g15890 = NOT(g11600)
--	g15904 = NOT(g11644)
--	g15913 = NOT(g11647)
--	g15923 = NOT(g11630)
--	g15933 = NOT(g11663)
--	g15942 = NOT(g11666)
--	g15952 = NOT(g11653)
--	g15962 = NOT(g11675)
--	g15971 = NOT(g11678)
--	g15981 = NOT(g11687)
--	I22163 = NOT(g12433)
--	g15989 = NOT(I22163)
--	g15991 = NOT(g12548)
--	g15994 = NOT(g12555)
--	g15997 = NOT(g12561)
--	g16001 = NOT(g12601)
--	g16002 = NOT(g12604)
--	g16005 = NOT(g12608)
--	g16007 = NOT(g12647)
--	g16011 = NOT(g12651)
--	g16012 = NOT(g12654)
--	g16013 = NOT(g12692)
--	g16014 = NOT(g12695)
--	g16023 = NOT(g12699)
--	g16024 = NOT(g12702)
--	g16025 = NOT(g12705)
--	g16026 = NOT(g12708)
--	g16027 = NOT(g12744)
--	g16034 = NOT(g12749)
--	g16035 = NOT(g12752)
--	g16039 = NOT(g12756)
--	g16040 = NOT(g12759)
--	g16041 = NOT(g12762)
--	g16042 = NOT(g12765)
--	g16043 = NOT(g12769)
--	g16044 = NOT(g12772)
--	g16054 = NOT(g12783)
--	g16055 = NOT(g12786)
--	g16056 = NOT(g12791)
--	g16057 = NOT(g12794)
--	g16061 = NOT(g12798)
--	g16062 = NOT(g12801)
--	g16063 = NOT(g12804)
--	g16064 = NOT(g12808)
--	g16065 = NOT(g12811)
--	g16075 = NOT(g11861)
--	g16088 = NOT(g12816)
--	g16090 = NOT(g12822)
--	g16091 = NOT(g12825)
--	g16092 = NOT(g12830)
--	g16093 = NOT(g12833)
--	g16097 = NOT(g12837)
--	g16098 = NOT(g12840)
--	g16099 = NOT(g12844)
--	g16113 = NOT(g11903)
--	g16126 = NOT(g12854)
--	g16128 = NOT(g12860)
--	g16129 = NOT(g12863)
--	g16130 = NOT(g12868)
--	g16131 = NOT(g12871)
--	g16142 = NOT(g13057)
--	g16154 = NOT(g12194)
--	g16164 = NOT(g11953)
--	g16177 = NOT(g12895)
--	g16179 = NOT(g12901)
--	g16180 = NOT(g12904)
--	g16189 = NOT(g13043)
--	g16201 = NOT(g13073)
--	g16213 = NOT(g12249)
--	g16223 = NOT(g12006)
--	g16236 = NOT(g12935)
--	g16243 = NOT(g13033)
--	g16254 = NOT(g13060)
--	g16266 = NOT(g13092)
--	g16278 = NOT(g12292)
--	g16287 = NOT(g12962)
--	g16293 = NOT(g13025)
--	I22382 = NOT(g520)
--	g16297 = NOT(I22382)
--	g16302 = NOT(g13046)
--	g16313 = NOT(g13076)
--	g16325 = NOT(g13107)
--	g16337 = NOT(g12328)
--	g16351 = NOT(g13036)
--	I22414 = NOT(g1206)
--	g16355 = NOT(I22414)
--	g16360 = NOT(g13063)
--	g16371 = NOT(g13095)
--	g16395 = NOT(g13049)
--	I22444 = NOT(g1900)
--	g16399 = NOT(I22444)
--	g16404 = NOT(g13079)
--	g16433 = NOT(g13066)
--	I22475 = NOT(g2594)
--	g16437 = NOT(I22475)
--	g16466 = NOT(g12017)
--	I22503 = NOT(g13598)
--	g16467 = NOT(I22503)
--	I22506 = NOT(g13624)
--	g16468 = NOT(I22506)
--	I22509 = NOT(g13610)
--	g16469 = NOT(I22509)
--	I22512 = NOT(g13635)
--	g16470 = NOT(I22512)
--	I22515 = NOT(g13620)
--	g16471 = NOT(I22515)
--	I22518 = NOT(g13647)
--	g16472 = NOT(I22518)
--	I22521 = NOT(g13632)
--	g16473 = NOT(I22521)
--	I22524 = NOT(g13673)
--	g16474 = NOT(I22524)
--	I22527 = NOT(g13469)
--	g16475 = NOT(I22527)
--	I22530 = NOT(g14774)
--	g16476 = NOT(I22530)
--	I22533 = NOT(g14795)
--	g16477 = NOT(I22533)
--	I22536 = NOT(g14829)
--	g16478 = NOT(I22536)
--	I22539 = NOT(g14882)
--	g16479 = NOT(I22539)
--	I22542 = NOT(g14954)
--	g16480 = NOT(I22542)
--	I22545 = NOT(g15018)
--	g16481 = NOT(I22545)
--	I22548 = NOT(g14718)
--	g16482 = NOT(I22548)
--	I22551 = NOT(g14745)
--	g16483 = NOT(I22551)
--	I22554 = NOT(g14765)
--	g16484 = NOT(I22554)
--	I22557 = NOT(g14775)
--	g16485 = NOT(I22557)
--	I22560 = NOT(g14796)
--	g16486 = NOT(I22560)
--	I22563 = NOT(g14830)
--	g16487 = NOT(I22563)
--	I22566 = NOT(g14883)
--	g16488 = NOT(I22566)
--	I22569 = NOT(g14955)
--	g16489 = NOT(I22569)
--	I22572 = NOT(g15019)
--	g16490 = NOT(I22572)
--	I22575 = NOT(g15092)
--	g16491 = NOT(I22575)
--	I22578 = NOT(g14746)
--	g16492 = NOT(I22578)
--	I22581 = NOT(g14766)
--	g16493 = NOT(I22581)
--	I22584 = NOT(g15989)
--	g16494 = NOT(I22584)
--	I22587 = NOT(g14684)
--	g16495 = NOT(I22587)
--	I22590 = NOT(g13863)
--	g16496 = NOT(I22590)
--	I22593 = NOT(g15876)
--	g16497 = NOT(I22593)
--	g16501 = NOT(g14158)
--	I22599 = NOT(g14966)
--	g16506 = NOT(I22599)
--	g16507 = NOT(g14186)
--	I22604 = NOT(g15080)
--	g16514 = NOT(I22604)
--	g16515 = NOT(g14244)
--	g16523 = NOT(g14273)
--	I22611 = NOT(g15055)
--	g16528 = NOT(I22611)
--	g16529 = NOT(g14301)
--	I22618 = NOT(g14630)
--	g16540 = NOT(I22618)
--	g16543 = NOT(g14347)
--	g16546 = NOT(g14366)
--	g16554 = NOT(g14395)
--	I22626 = NOT(g15151)
--	g16559 = NOT(I22626)
--	g16560 = NOT(g14423)
--	I22640 = NOT(g14650)
--	g16572 = NOT(I22640)
--	g16575 = NOT(g14459)
--	g16578 = NOT(g14478)
--	g16586 = NOT(g14507)
--	I22651 = NOT(g14677)
--	g16596 = NOT(I22651)
--	g16599 = NOT(g14546)
--	g16602 = NOT(g14565)
--	I22657 = NOT(g14657)
--	g16608 = NOT(I22657)
--	I22663 = NOT(g14711)
--	g16616 = NOT(I22663)
--	g16619 = NOT(g14601)
--	I22667 = NOT(g14642)
--	g16622 = NOT(I22667)
--	I22671 = NOT(g14691)
--	g16626 = NOT(I22671)
--	I22676 = NOT(g14630)
--	g16633 = NOT(I22676)
--	I22679 = NOT(g14669)
--	g16636 = NOT(I22679)
--	I22683 = NOT(g14725)
--	g16640 = NOT(I22683)
--	I22687 = NOT(g14650)
--	g16644 = NOT(I22687)
--	I22690 = NOT(g14703)
--	g16647 = NOT(I22690)
--	I22694 = NOT(g14753)
--	g16651 = NOT(I22694)
--	I22699 = NOT(g14677)
--	g16656 = NOT(I22699)
--	I22702 = NOT(g14737)
--	g16659 = NOT(I22702)
--	g16665 = NOT(g14776)
--	I22715 = NOT(g14711)
--	g16673 = NOT(I22715)
--	I22718 = NOT(g14657)
--	g16676 = NOT(I22718)
--	g16682 = NOT(g14797)
--	g16686 = NOT(g14811)
--	I22726 = NOT(g14642)
--	g16694 = NOT(I22726)
--	g16697 = NOT(g14837)
--	I22730 = NOT(g14691)
--	g16702 = NOT(I22730)
--	g16708 = NOT(g14849)
--	g16712 = NOT(g14863)
--	I22737 = NOT(g14630)
--	g16719 = NOT(I22737)
--	g16722 = NOT(g14895)
--	I22741 = NOT(g14669)
--	g16725 = NOT(I22741)
--	g16728 = NOT(g14910)
--	I22745 = NOT(g14725)
--	g16733 = NOT(I22745)
--	g16739 = NOT(g14922)
--	g16743 = NOT(g14936)
--	g16749 = NOT(g15782)
--	I22752 = NOT(g14657)
--	g16758 = NOT(I22752)
--	I22755 = NOT(g14650)
--	g16761 = NOT(I22755)
--	g16764 = NOT(g14976)
--	I22759 = NOT(g14703)
--	g16767 = NOT(I22759)
--	g16770 = NOT(g14991)
--	I22763 = NOT(g14753)
--	g16775 = NOT(I22763)
--	g16781 = NOT(g15003)
--	I22768 = NOT(g14691)
--	g16785 = NOT(I22768)
--	I22771 = NOT(g14677)
--	g16788 = NOT(I22771)
--	g16791 = NOT(g15065)
--	I22775 = NOT(g14737)
--	g16794 = NOT(I22775)
--	g16797 = NOT(g15080)
--	g16804 = NOT(g15803)
--	g16809 = NOT(g15842)
--	I22783 = NOT(g13572)
--	g16813 = NOT(I22783)
--	I22786 = NOT(g14725)
--	g16814 = NOT(I22786)
--	I22789 = NOT(g14711)
--	g16817 = NOT(I22789)
--	g16820 = NOT(g15161)
--	g16825 = NOT(g15855)
--	I22797 = NOT(g14165)
--	g16830 = NOT(I22797)
--	I22800 = NOT(g13581)
--	g16831 = NOT(I22800)
--	I22803 = NOT(g14753)
--	g16832 = NOT(I22803)
--	g16836 = NOT(g15818)
--	g16840 = NOT(g15878)
--	I22810 = NOT(g14280)
--	g16842 = NOT(I22810)
--	I22813 = NOT(g13601)
--	g16843 = NOT(I22813)
--	g16846 = NOT(g15903)
--	I22820 = NOT(g14402)
--	g16848 = NOT(I22820)
--	I22823 = NOT(g13613)
--	g16849 = NOT(I22823)
--	I22828 = NOT(g14514)
--	g16852 = NOT(I22828)
--	I22836 = NOT(g13571)
--	g16858 = NOT(I22836)
--	I22842 = NOT(g13580)
--	g16862 = NOT(I22842)
--	I22845 = NOT(g13579)
--	g16863 = NOT(I22845)
--	g16867 = NOT(g13589)
--	I22852 = NOT(g13600)
--	g16877 = NOT(I22852)
--	I22855 = NOT(g13588)
--	g16878 = NOT(I22855)
--	I22860 = NOT(g14885)
--	g16881 = NOT(I22860)
--	g16884 = NOT(g13589)
--	g16895 = NOT(g13589)
--	I22866 = NOT(g13612)
--	g16905 = NOT(I22866)
--	I22869 = NOT(g13608)
--	g16906 = NOT(I22869)
--	I22875 = NOT(g14966)
--	g16910 = NOT(I22875)
--	g16913 = NOT(g13589)
--	g16924 = NOT(g13589)
--	I22881 = NOT(g13622)
--	g16934 = NOT(I22881)
--	I22893 = NOT(g15055)
--	g16940 = NOT(I22893)
--	g16943 = NOT(g13589)
--	g16954 = NOT(g13589)
--	I22912 = NOT(g15151)
--	g16971 = NOT(I22912)
--	g16974 = NOT(g13589)
--	g17029 = NOT(g14685)
--	g17057 = NOT(g13519)
--	g17063 = NOT(g14719)
--	g17092 = NOT(g13530)
--	g17098 = NOT(g14747)
--	g17130 = NOT(g13541)
--	g17136 = NOT(g14768)
--	g17157 = NOT(g13552)
--	I23253 = NOT(g13741)
--	g17189 = NOT(I23253)
--	I23274 = NOT(g13741)
--	g17200 = NOT(I23274)
--	g17203 = NOT(g13568)
--	I23287 = NOT(g13741)
--	g17207 = NOT(I23287)
--	g17208 = NOT(g13576)
--	I23292 = NOT(g13741)
--	g17212 = NOT(I23292)
--	g17214 = NOT(g13585)
--	g17217 = NOT(g13605)
--	I23309 = NOT(g16132)
--	g17227 = NOT(I23309)
--	I23314 = NOT(g15720)
--	g17230 = NOT(I23314)
--	I23317 = NOT(g16181)
--	g17233 = NOT(I23317)
--	I23323 = NOT(g15664)
--	g17237 = NOT(I23323)
--	I23326 = NOT(g15758)
--	g17240 = NOT(I23326)
--	I23329 = NOT(g15760)
--	g17243 = NOT(I23329)
--	I23335 = NOT(g16412)
--	g17249 = NOT(I23335)
--	I23338 = NOT(g15721)
--	g17252 = NOT(I23338)
--	I23341 = NOT(g15784)
--	g17255 = NOT(I23341)
--	g17258 = NOT(g16053)
--	I23345 = NOT(g15723)
--	g17259 = NOT(I23345)
--	I23348 = NOT(g15786)
--	g17262 = NOT(I23348)
--	I23351 = NOT(g15788)
--	g17265 = NOT(I23351)
--	I23358 = NOT(g16442)
--	g17272 = NOT(I23358)
--	I23361 = NOT(g15759)
--	g17275 = NOT(I23361)
--	I23364 = NOT(g15805)
--	g17278 = NOT(I23364)
--	g17281 = NOT(g16081)
--	I23368 = NOT(g16446)
--	g17282 = NOT(I23368)
--	I23371 = NOT(g15761)
--	g17285 = NOT(I23371)
--	I23374 = NOT(g15807)
--	g17288 = NOT(I23374)
--	I23377 = NOT(g15763)
--	g17291 = NOT(I23377)
--	I23380 = NOT(g15809)
--	g17294 = NOT(I23380)
--	I23383 = NOT(g15811)
--	g17297 = NOT(I23383)
--	I23386 = NOT(g13469)
--	g17300 = NOT(I23386)
--	I23392 = NOT(g13476)
--	g17304 = NOT(I23392)
--	I23395 = NOT(g15785)
--	g17307 = NOT(I23395)
--	I23398 = NOT(g15820)
--	g17310 = NOT(I23398)
--	g17313 = NOT(g16109)
--	g17314 = NOT(g16110)
--	I23403 = NOT(g13478)
--	g17315 = NOT(I23403)
--	I23406 = NOT(g15787)
--	g17318 = NOT(I23406)
--	I23409 = NOT(g15822)
--	g17321 = NOT(I23409)
--	I23412 = NOT(g13482)
--	g17324 = NOT(I23412)
--	I23415 = NOT(g15789)
--	g17327 = NOT(I23415)
--	I23418 = NOT(g15824)
--	g17330 = NOT(I23418)
--	I23421 = NOT(g15791)
--	g17333 = NOT(I23421)
--	I23424 = NOT(g15826)
--	g17336 = NOT(I23424)
--	I23430 = NOT(g13494)
--	g17342 = NOT(I23430)
--	I23433 = NOT(g15806)
--	g17345 = NOT(I23433)
--	I23436 = NOT(g15832)
--	g17348 = NOT(I23436)
--	g17351 = NOT(g16152)
--	I23442 = NOT(g13495)
--	g17354 = NOT(I23442)
--	I23445 = NOT(g15808)
--	g17357 = NOT(I23445)
--	I23448 = NOT(g15834)
--	g17360 = NOT(I23448)
--	I23451 = NOT(g13497)
--	g17363 = NOT(I23451)
--	I23454 = NOT(g15810)
--	g17366 = NOT(I23454)
--	I23457 = NOT(g15836)
--	g17369 = NOT(I23457)
--	I23460 = NOT(g13501)
--	g17372 = NOT(I23460)
--	I23463 = NOT(g15812)
--	g17375 = NOT(I23463)
--	I23466 = NOT(g15838)
--	g17378 = NOT(I23466)
--	I23472 = NOT(g13510)
--	g17384 = NOT(I23472)
--	I23475 = NOT(g15821)
--	g17387 = NOT(I23475)
--	I23478 = NOT(g15844)
--	g17390 = NOT(I23478)
--	g17394 = NOT(g16197)
--	I23487 = NOT(g13511)
--	g17399 = NOT(I23487)
--	I23490 = NOT(g15823)
--	g17402 = NOT(I23490)
--	I23493 = NOT(g15846)
--	g17405 = NOT(I23493)
--	I23498 = NOT(g13512)
--	g17410 = NOT(I23498)
--	I23501 = NOT(g15825)
--	g17413 = NOT(I23501)
--	I23504 = NOT(g15848)
--	g17416 = NOT(I23504)
--	I23507 = NOT(g13514)
--	g17419 = NOT(I23507)
--	I23510 = NOT(g15827)
--	g17422 = NOT(I23510)
--	I23513 = NOT(g15850)
--	g17425 = NOT(I23513)
--	I23518 = NOT(g15856)
--	g17430 = NOT(I23518)
--	I23521 = NOT(g13518)
--	g17433 = NOT(I23521)
--	I23524 = NOT(g15833)
--	g17436 = NOT(I23524)
--	I23527 = NOT(g15858)
--	g17439 = NOT(I23527)
--	I23530 = NOT(g14885)
--	g17442 = NOT(I23530)
--	g17445 = NOT(g16250)
--	I23539 = NOT(g13524)
--	g17451 = NOT(I23539)
--	I23542 = NOT(g15835)
--	g17454 = NOT(I23542)
--	I23545 = NOT(g15867)
--	g17457 = NOT(I23545)
--	I23553 = NOT(g13525)
--	g17465 = NOT(I23553)
--	I23556 = NOT(g15837)
--	g17468 = NOT(I23556)
--	I23559 = NOT(g15869)
--	g17471 = NOT(I23559)
--	I23564 = NOT(g13526)
--	g17476 = NOT(I23564)
--	I23567 = NOT(g15839)
--	g17479 = NOT(I23567)
--	I23570 = NOT(g15871)
--	g17482 = NOT(I23570)
--	I23575 = NOT(g15843)
--	g17487 = NOT(I23575)
--	I23578 = NOT(g15879)
--	g17490 = NOT(I23578)
--	I23581 = NOT(g13528)
--	g17493 = NOT(I23581)
--	I23584 = NOT(g15845)
--	g17496 = NOT(I23584)
--	g17499 = NOT(g16292)
--	I23588 = NOT(g14885)
--	g17500 = NOT(I23588)
--	I23591 = NOT(g14885)
--	g17503 = NOT(I23591)
--	I23599 = NOT(g15887)
--	g17511 = NOT(I23599)
--	I23602 = NOT(g13529)
--	g17514 = NOT(I23602)
--	I23605 = NOT(g15847)
--	g17517 = NOT(I23605)
--	I23608 = NOT(g15889)
--	g17520 = NOT(I23608)
--	I23611 = NOT(g14966)
--	g17523 = NOT(I23611)
--	I23619 = NOT(g13535)
--	g17531 = NOT(I23619)
--	I23622 = NOT(g15849)
--	g17534 = NOT(I23622)
--	I23625 = NOT(g15898)
--	g17537 = NOT(I23625)
--	I23633 = NOT(g13536)
--	g17545 = NOT(I23633)
--	I23636 = NOT(g15851)
--	g17548 = NOT(I23636)
--	I23639 = NOT(g15900)
--	g17551 = NOT(I23639)
--	I23645 = NOT(g13537)
--	g17557 = NOT(I23645)
--	I23648 = NOT(g15857)
--	g17560 = NOT(I23648)
--	I23651 = NOT(g13538)
--	g17563 = NOT(I23651)
--	g17566 = NOT(g16346)
--	I23655 = NOT(g14831)
--	g17567 = NOT(I23655)
--	I23658 = NOT(g14885)
--	g17570 = NOT(I23658)
--	I23661 = NOT(g16085)
--	g17573 = NOT(I23661)
--	I23667 = NOT(g15866)
--	g17579 = NOT(I23667)
--	I23670 = NOT(g15912)
--	g17582 = NOT(I23670)
--	I23673 = NOT(g13539)
--	g17585 = NOT(I23673)
--	I23676 = NOT(g15868)
--	g17588 = NOT(I23676)
--	I23679 = NOT(g14966)
--	g17591 = NOT(I23679)
--	I23682 = NOT(g14966)
--	g17594 = NOT(I23682)
--	I23689 = NOT(g15920)
--	g17601 = NOT(I23689)
--	I23692 = NOT(g13540)
--	g17604 = NOT(I23692)
--	I23695 = NOT(g15870)
--	g17607 = NOT(I23695)
--	I23698 = NOT(g15922)
--	g17610 = NOT(I23698)
--	I23701 = NOT(g15055)
--	g17613 = NOT(I23701)
--	I23709 = NOT(g13546)
--	g17621 = NOT(I23709)
--	I23712 = NOT(g15872)
--	g17624 = NOT(I23712)
--	I23715 = NOT(g15931)
--	g17627 = NOT(I23715)
--	I23725 = NOT(g13547)
--	g17637 = NOT(I23725)
--	g17640 = NOT(g13873)
--	I23729 = NOT(g14337)
--	g17645 = NOT(I23729)
--	g17648 = NOT(g16384)
--	I23733 = NOT(g14831)
--	g17649 = NOT(I23733)
--	I23739 = NOT(g13548)
--	g17655 = NOT(I23739)
--	I23742 = NOT(g15888)
--	g17658 = NOT(I23742)
--	I23745 = NOT(g13549)
--	g17661 = NOT(I23745)
--	I23748 = NOT(g14904)
--	g17664 = NOT(I23748)
--	I23751 = NOT(g14966)
--	g17667 = NOT(I23751)
--	I23754 = NOT(g16123)
--	g17670 = NOT(I23754)
--	I23760 = NOT(g15897)
--	g17676 = NOT(I23760)
--	I23763 = NOT(g15941)
--	g17679 = NOT(I23763)
--	I23766 = NOT(g13550)
--	g17682 = NOT(I23766)
--	I23769 = NOT(g15899)
--	g17685 = NOT(I23769)
--	I23772 = NOT(g15055)
--	g17688 = NOT(I23772)
--	I23775 = NOT(g15055)
--	g17691 = NOT(I23775)
--	I23782 = NOT(g15949)
--	g17698 = NOT(I23782)
--	I23785 = NOT(g13551)
--	g17701 = NOT(I23785)
--	I23788 = NOT(g15901)
--	g17704 = NOT(I23788)
--	I23791 = NOT(g15951)
--	g17707 = NOT(I23791)
--	I23794 = NOT(g15151)
--	g17710 = NOT(I23794)
--	g17720 = NOT(g15853)
--	g17724 = NOT(g13886)
--	I23817 = NOT(g13557)
--	g17738 = NOT(I23817)
--	g17741 = NOT(g13895)
--	I23821 = NOT(g14337)
--	g17746 = NOT(I23821)
--	I23824 = NOT(g14904)
--	g17749 = NOT(I23824)
--	I23830 = NOT(g13558)
--	g17755 = NOT(I23830)
--	I23833 = NOT(g15921)
--	g17758 = NOT(I23833)
--	I23836 = NOT(g13559)
--	g17761 = NOT(I23836)
--	I23839 = NOT(g14985)
--	g17764 = NOT(I23839)
--	I23842 = NOT(g15055)
--	g17767 = NOT(I23842)
--	I23845 = NOT(g16174)
--	g17770 = NOT(I23845)
--	I23851 = NOT(g15930)
--	g17776 = NOT(I23851)
--	I23854 = NOT(g15970)
--	g17779 = NOT(I23854)
--	I23857 = NOT(g13560)
--	g17782 = NOT(I23857)
--	I23860 = NOT(g15932)
--	g17785 = NOT(I23860)
--	I23863 = NOT(g15151)
--	g17788 = NOT(I23863)
--	I23866 = NOT(g15151)
--	g17791 = NOT(I23866)
--	I23874 = NOT(g15797)
--	g17799 = NOT(I23874)
--	g17802 = NOT(g13907)
--	I23888 = NOT(g14685)
--	g17815 = NOT(I23888)
--	g17825 = NOT(g13927)
--	I23904 = NOT(g13561)
--	g17839 = NOT(I23904)
--	g17842 = NOT(g13936)
--	I23908 = NOT(g14337)
--	g17847 = NOT(I23908)
--	I23911 = NOT(g14985)
--	g17850 = NOT(I23911)
--	I23917 = NOT(g13562)
--	g17856 = NOT(I23917)
--	I23920 = NOT(g15950)
--	g17859 = NOT(I23920)
--	I23923 = NOT(g13563)
--	g17862 = NOT(I23923)
--	I23926 = NOT(g15074)
--	g17865 = NOT(I23926)
--	I23929 = NOT(g15151)
--	g17868 = NOT(I23929)
--	I23932 = NOT(g16233)
--	g17871 = NOT(I23932)
--	g17878 = NOT(g15830)
--	g17882 = NOT(g13946)
--	g17892 = NOT(g13954)
--	g17893 = NOT(g14165)
--	I23954 = NOT(g16154)
--	g17903 = NOT(I23954)
--	g17914 = NOT(g13963)
--	I23976 = NOT(g14719)
--	g17927 = NOT(I23976)
--	g17937 = NOT(g13983)
--	I23992 = NOT(g13564)
--	g17951 = NOT(I23992)
--	g17954 = NOT(g13992)
--	I23996 = NOT(g14337)
--	g17959 = NOT(I23996)
--	I23999 = NOT(g15074)
--	g17962 = NOT(I23999)
--	g17969 = NOT(g15841)
--	g17974 = NOT(g14001)
--	g17984 = NOT(g14008)
--	g17988 = NOT(g14685)
--	g17991 = NOT(g14450)
--	g17993 = NOT(g14016)
--	g18003 = NOT(g14024)
--	g18004 = NOT(g14280)
--	I24049 = NOT(g16213)
--	g18014 = NOT(I24049)
--	g18025 = NOT(g14033)
--	I24071 = NOT(g14747)
--	g18038 = NOT(I24071)
--	g18048 = NOT(g14053)
--	g18063 = NOT(g15660)
--	g18070 = NOT(g15854)
--	g18074 = NOT(g14062)
--	g18084 = NOT(g14068)
--	g18089 = NOT(g14355)
--	g18091 = NOT(g14092)
--	g18101 = NOT(g14099)
--	g18105 = NOT(g14719)
--	g18108 = NOT(g14537)
--	g18110 = NOT(g14107)
--	g18120 = NOT(g14115)
--	g18121 = NOT(g14402)
--	I24144 = NOT(g16278)
--	g18131 = NOT(I24144)
--	g18142 = NOT(g14124)
--	I24166 = NOT(g14768)
--	g18155 = NOT(I24166)
--	I24171 = NOT(g16439)
--	g18166 = NOT(I24171)
--	g18170 = NOT(g15877)
--	g18174 = NOT(g14148)
--	g18179 = NOT(g14153)
--	g18188 = NOT(g14252)
--	g18190 = NOT(g14177)
--	g18200 = NOT(g14183)
--	g18205 = NOT(g14467)
--	g18207 = NOT(g14207)
--	g18217 = NOT(g14214)
--	g18221 = NOT(g14747)
--	g18224 = NOT(g14592)
--	g18226 = NOT(g14222)
--	g18236 = NOT(g14230)
--	g18237 = NOT(g14514)
--	I24247 = NOT(g16337)
--	g18247 = NOT(I24247)
--	I24258 = NOT(g16463)
--	g18258 = NOT(I24258)
--	g18261 = NOT(g15719)
--	g18265 = NOT(g14238)
--	g18275 = NOT(g14171)
--	I24285 = NOT(g15992)
--	g18278 = NOT(I24285)
--	g18281 = NOT(g14263)
--	g18286 = NOT(g14268)
--	g18295 = NOT(g14374)
--	g18297 = NOT(g14292)
--	g18307 = NOT(g14298)
--	g18312 = NOT(g14554)
--	g18314 = NOT(g14322)
--	g18324 = NOT(g14329)
--	g18328 = NOT(g14768)
--	g18331 = NOT(g14626)
--	I24346 = NOT(g15873)
--	g18334 = NOT(I24346)
--	g18337 = NOT(g15757)
--	g18341 = NOT(g14342)
--	g18351 = NOT(g13741)
--	g18353 = NOT(g13918)
--	I24368 = NOT(g15990)
--	g18355 = NOT(I24368)
--	g18358 = NOT(g14360)
--	g18368 = NOT(g14286)
--	I24394 = NOT(g15995)
--	g18371 = NOT(I24394)
--	g18374 = NOT(g14385)
--	g18379 = NOT(g14390)
--	g18388 = NOT(g14486)
--	g18390 = NOT(g14414)
--	g18400 = NOT(g14420)
--	g18405 = NOT(g14609)
--	g18407 = NOT(g15959)
--	g18414 = NOT(g15718)
--	g18415 = NOT(g15783)
--	g18429 = NOT(g14831)
--	I24459 = NOT(g13599)
--	g18432 = NOT(I24459)
--	g18435 = NOT(g14359)
--	g18436 = NOT(g14454)
--	g18446 = NOT(g13741)
--	g18448 = NOT(g13974)
--	I24481 = NOT(g15993)
--	g18450 = NOT(I24481)
--	g18453 = NOT(g14472)
--	g18463 = NOT(g14408)
--	I24507 = NOT(g15999)
--	g18466 = NOT(I24507)
--	g18469 = NOT(g14497)
--	g18474 = NOT(g14502)
--	g18483 = NOT(g14573)
--	g18485 = NOT(g15756)
--	g18486 = NOT(g15804)
--	g18490 = NOT(g13565)
--	g18502 = NOT(g14904)
--	I24560 = NOT(g13611)
--	g18505 = NOT(I24560)
--	g18508 = NOT(g14471)
--	g18509 = NOT(g14541)
--	g18519 = NOT(g13741)
--	g18521 = NOT(g14044)
--	I24582 = NOT(g15996)
--	g18523 = NOT(I24582)
--	g18526 = NOT(g14559)
--	g18536 = NOT(g14520)
--	I24608 = NOT(g16006)
--	g18539 = NOT(I24608)
--	g18543 = NOT(g15819)
--	g18552 = NOT(g16154)
--	g18554 = NOT(g13573)
--	g18566 = NOT(g14985)
--	I24662 = NOT(g13621)
--	g18569 = NOT(I24662)
--	g18572 = NOT(g14558)
--	g18573 = NOT(g14596)
--	g18583 = NOT(g13741)
--	g18585 = NOT(g14135)
--	I24684 = NOT(g16000)
--	g18587 = NOT(I24684)
--	g18593 = NOT(g15831)
--	g18602 = NOT(g16213)
--	g18604 = NOT(g13582)
--	g18616 = NOT(g15074)
--	I24732 = NOT(g13633)
--	g18619 = NOT(I24732)
--	g18622 = NOT(g14613)
--	g18634 = NOT(g16278)
--	g18636 = NOT(g13602)
--	g18643 = NOT(g16337)
--	g18646 = NOT(g16341)
--	g18656 = NOT(g14776)
--	g18670 = NOT(g14797)
--	g18679 = NOT(g14811)
--	g18691 = NOT(g14885)
--	g18692 = NOT(g14837)
--	g18699 = NOT(g14849)
--	g18708 = NOT(g14863)
--	g18720 = NOT(g14895)
--	g18725 = NOT(g13865)
--	g18727 = NOT(g14966)
--	g18728 = NOT(g14910)
--	g18735 = NOT(g14922)
--	g18744 = NOT(g14936)
--	g18756 = NOT(g14960)
--	g18757 = NOT(g14963)
--	g18758 = NOT(g14976)
--	g18764 = NOT(g15055)
--	g18765 = NOT(g14991)
--	g18772 = NOT(g15003)
--	g18783 = NOT(g15034)
--	g18784 = NOT(g15037)
--	g18785 = NOT(g15040)
--	g18786 = NOT(g15043)
--	g18787 = NOT(g15049)
--	g18788 = NOT(g15052)
--	g18789 = NOT(g15065)
--	g18795 = NOT(g15151)
--	g18796 = NOT(g15080)
--	g18805 = NOT(g15106)
--	g18806 = NOT(g15109)
--	g18807 = NOT(g15112)
--	g18808 = NOT(g15115)
--	g18809 = NOT(g15130)
--	g18810 = NOT(g15133)
--	g18811 = NOT(g15136)
--	g18812 = NOT(g15139)
--	g18813 = NOT(g15145)
--	g18814 = NOT(g15148)
--	g18815 = NOT(g15161)
--	g18822 = NOT(g15179)
--	g18823 = NOT(g15182)
--	g18824 = NOT(g15185)
--	g18825 = NOT(g15198)
--	g18826 = NOT(g15201)
--	g18827 = NOT(g15204)
--	g18828 = NOT(g15207)
--	g18829 = NOT(g15222)
--	g18830 = NOT(g15225)
--	g18831 = NOT(g15228)
--	g18832 = NOT(g15231)
--	g18833 = NOT(g15237)
--	g18834 = NOT(g15240)
--	g18838 = NOT(g15248)
--	g18839 = NOT(g15251)
--	g18840 = NOT(g15254)
--	g18841 = NOT(g15265)
--	g18842 = NOT(g15268)
--	g18843 = NOT(g15271)
--	g18844 = NOT(g15284)
--	g18845 = NOT(g15287)
--	g18846 = NOT(g15290)
--	g18847 = NOT(g15293)
--	g18848 = NOT(g15308)
--	g18849 = NOT(g15311)
--	g18850 = NOT(g15314)
--	g18851 = NOT(g15317)
--	g18853 = NOT(g15326)
--	g18854 = NOT(g15329)
--	g18855 = NOT(g15332)
--	g18856 = NOT(g15340)
--	g18857 = NOT(g15343)
--	g18858 = NOT(g15346)
--	g18859 = NOT(g15357)
--	g18860 = NOT(g15360)
--	g18861 = NOT(g15363)
--	g18862 = NOT(g15376)
--	g18863 = NOT(g15379)
--	g18864 = NOT(g15382)
--	g18865 = NOT(g15385)
--	I24894 = NOT(g14797)
--	g18869 = NOT(I24894)
--	g18870 = NOT(g15393)
--	g18871 = NOT(g15396)
--	g18872 = NOT(g15399)
--	g18873 = NOT(g15404)
--	g18874 = NOT(g15412)
--	g18875 = NOT(g15415)
--	g18876 = NOT(g15418)
--	g18877 = NOT(g15426)
--	g18878 = NOT(g15429)
--	g18879 = NOT(g15432)
--	g18880 = NOT(g15443)
--	g18881 = NOT(g15446)
--	g18882 = NOT(g15449)
--	g18884 = NOT(g13469)
--	I24913 = NOT(g15800)
--	g18886 = NOT(I24913)
--	I24916 = NOT(g14776)
--	g18890 = NOT(I24916)
--	g18891 = NOT(g15461)
--	g18892 = NOT(g15464)
--	g18893 = NOT(g15467)
--	g18894 = NOT(g15471)
--	I24923 = NOT(g14849)
--	g18895 = NOT(I24923)
--	g18896 = NOT(g15477)
--	g18897 = NOT(g15480)
--	g18898 = NOT(g15483)
--	g18899 = NOT(g15488)
--	g18900 = NOT(g15496)
--	g18901 = NOT(g15499)
--	g18902 = NOT(g15502)
--	g18903 = NOT(g15510)
--	g18904 = NOT(g15513)
--	g18905 = NOT(g15516)
--	g18908 = NOT(g15521)
--	g18909 = NOT(g15528)
--	g18910 = NOT(g15531)
--	g18911 = NOT(g15534)
--	g18912 = NOT(g15537)
--	I24943 = NOT(g14811)
--	g18913 = NOT(I24943)
--	g18914 = NOT(g15547)
--	g18915 = NOT(g15550)
--	g18916 = NOT(g15553)
--	g18917 = NOT(g15557)
--	I24950 = NOT(g14922)
--	g18918 = NOT(I24950)
--	g18919 = NOT(g15563)
--	g18920 = NOT(g15566)
--	g18921 = NOT(g15569)
--	g18922 = NOT(g15574)
--	g18923 = NOT(g15582)
--	g18924 = NOT(g15585)
--	g18925 = NOT(g15588)
--	g18926 = NOT(g15596)
--	g18927 = NOT(g15599)
--	g18928 = NOT(g15606)
--	g18929 = NOT(g15609)
--	g18930 = NOT(g15612)
--	g18931 = NOT(g15615)
--	I24966 = NOT(g14863)
--	g18932 = NOT(I24966)
--	g18933 = NOT(g15625)
--	g18934 = NOT(g15628)
--	g18935 = NOT(g15631)
--	g18936 = NOT(g15635)
--	I24973 = NOT(g15003)
--	g18937 = NOT(I24973)
--	g18938 = NOT(g15641)
--	g18939 = NOT(g15644)
--	g18940 = NOT(g15647)
--	g18941 = NOT(g15652)
--	g18943 = NOT(g15655)
--	I24982 = NOT(g14347)
--	g18944 = NOT(I24982)
--	g18945 = NOT(g15667)
--	g18946 = NOT(g15672)
--	g18947 = NOT(g15675)
--	g18948 = NOT(g15682)
--	g18949 = NOT(g15685)
--	g18950 = NOT(g15688)
--	g18951 = NOT(g15691)
--	I24992 = NOT(g14936)
--	g18952 = NOT(I24992)
--	g18953 = NOT(g15701)
--	g18954 = NOT(g15704)
--	g18955 = NOT(g15707)
--	g18956 = NOT(g15711)
--	g18958 = NOT(g15714)
--	I25001 = NOT(g14244)
--	g18959 = NOT(I25001)
--	I25004 = NOT(g14459)
--	g18960 = NOT(I25004)
--	g18961 = NOT(g15726)
--	g18962 = NOT(g15731)
--	g18963 = NOT(g15734)
--	g18964 = NOT(g15741)
--	g18965 = NOT(g15744)
--	g18966 = NOT(g15747)
--	g18967 = NOT(g15750)
--	I25015 = NOT(g14158)
--	g18969 = NOT(I25015)
--	I25018 = NOT(g14366)
--	g18970 = NOT(I25018)
--	I25021 = NOT(g14546)
--	g18971 = NOT(I25021)
--	g18972 = NOT(g15766)
--	g18973 = NOT(g15771)
--	g18974 = NOT(g15774)
--	g18976 = NOT(g15777)
--	I25037 = NOT(g14071)
--	g18981 = NOT(I25037)
--	I25041 = NOT(g14895)
--	g18983 = NOT(I25041)
--	I25044 = NOT(g14273)
--	g18984 = NOT(I25044)
--	I25047 = NOT(g14478)
--	g18985 = NOT(I25047)
--	I25050 = NOT(g14601)
--	g18986 = NOT(I25050)
--	g18987 = NOT(g15794)
--	I25054 = NOT(g14837)
--	g18988 = NOT(I25054)
--	I25057 = NOT(g14186)
--	g18989 = NOT(I25057)
--	I25061 = NOT(g14976)
--	g18991 = NOT(I25061)
--	I25064 = NOT(g14395)
--	g18992 = NOT(I25064)
--	I25067 = NOT(g14565)
--	g18993 = NOT(I25067)
--	I25071 = NOT(g14910)
--	g18995 = NOT(I25071)
--	I25074 = NOT(g14301)
--	g18996 = NOT(I25074)
--	I25078 = NOT(g15065)
--	g18998 = NOT(I25078)
--	I25081 = NOT(g14507)
--	g18999 = NOT(I25081)
--	I25084 = NOT(g14885)
--	g19000 = NOT(I25084)
--	g19001 = NOT(g14071)
--	I25089 = NOT(g14991)
--	g19008 = NOT(I25089)
--	I25092 = NOT(g14423)
--	g19009 = NOT(I25092)
--	I25096 = NOT(g15161)
--	g19011 = NOT(I25096)
--	I25099 = NOT(g19000)
--	g19012 = NOT(I25099)
--	I25102 = NOT(g18944)
--	g19013 = NOT(I25102)
--	I25105 = NOT(g18959)
--	g19014 = NOT(I25105)
--	I25108 = NOT(g18969)
--	g19015 = NOT(I25108)
--	I25111 = NOT(g18981)
--	g19016 = NOT(I25111)
--	I25114 = NOT(g18983)
--	g19017 = NOT(I25114)
--	I25117 = NOT(g18988)
--	g19018 = NOT(I25117)
--	I25120 = NOT(g18869)
--	g19019 = NOT(I25120)
--	I25123 = NOT(g18890)
--	g19020 = NOT(I25123)
--	I25126 = NOT(g16858)
--	g19021 = NOT(I25126)
--	I25129 = NOT(g16813)
--	g19022 = NOT(I25129)
--	I25132 = NOT(g16862)
--	g19023 = NOT(I25132)
--	I25135 = NOT(g16506)
--	g19024 = NOT(I25135)
--	I25138 = NOT(g18960)
--	g19025 = NOT(I25138)
--	I25141 = NOT(g18970)
--	g19026 = NOT(I25141)
--	I25144 = NOT(g18984)
--	g19027 = NOT(I25144)
--	I25147 = NOT(g18989)
--	g19028 = NOT(I25147)
--	I25150 = NOT(g18991)
--	g19029 = NOT(I25150)
--	I25153 = NOT(g18995)
--	g19030 = NOT(I25153)
--	I25156 = NOT(g18895)
--	g19031 = NOT(I25156)
--	I25159 = NOT(g18913)
--	g19032 = NOT(I25159)
--	I25162 = NOT(g16863)
--	g19033 = NOT(I25162)
--	I25165 = NOT(g16831)
--	g19034 = NOT(I25165)
--	I25168 = NOT(g16877)
--	g19035 = NOT(I25168)
--	I25171 = NOT(g16528)
--	g19036 = NOT(I25171)
--	I25174 = NOT(g18971)
--	g19037 = NOT(I25174)
--	I25177 = NOT(g18985)
--	g19038 = NOT(I25177)
--	I25180 = NOT(g18992)
--	g19039 = NOT(I25180)
--	I25183 = NOT(g18996)
--	g19040 = NOT(I25183)
--	I25186 = NOT(g18998)
--	g19041 = NOT(I25186)
--	I25189 = NOT(g19008)
--	g19042 = NOT(I25189)
--	I25192 = NOT(g18918)
--	g19043 = NOT(I25192)
--	I25195 = NOT(g18932)
--	g19044 = NOT(I25195)
--	I25198 = NOT(g16878)
--	g19045 = NOT(I25198)
--	I25201 = NOT(g16843)
--	g19046 = NOT(I25201)
--	I25204 = NOT(g16905)
--	g19047 = NOT(I25204)
--	I25207 = NOT(g16559)
--	g19048 = NOT(I25207)
--	I25210 = NOT(g18986)
--	g19049 = NOT(I25210)
--	I25213 = NOT(g18993)
--	g19050 = NOT(I25213)
--	I25216 = NOT(g18999)
--	g19051 = NOT(I25216)
--	I25219 = NOT(g19009)
--	g19052 = NOT(I25219)
--	I25222 = NOT(g19011)
--	g19053 = NOT(I25222)
--	I25225 = NOT(g16514)
--	g19054 = NOT(I25225)
--	I25228 = NOT(g18937)
--	g19055 = NOT(I25228)
--	I25231 = NOT(g18952)
--	g19056 = NOT(I25231)
--	I25234 = NOT(g16906)
--	g19057 = NOT(I25234)
--	I25237 = NOT(g16849)
--	g19058 = NOT(I25237)
--	I25240 = NOT(g16934)
--	g19059 = NOT(I25240)
--	I25243 = NOT(g17227)
--	g19060 = NOT(I25243)
--	I25246 = NOT(g17233)
--	g19061 = NOT(I25246)
--	I25249 = NOT(g17300)
--	g19062 = NOT(I25249)
--	I25253 = NOT(g17124)
--	g19064 = NOT(I25253)
--	g19070 = NOT(g18583)
--	I25258 = NOT(g16974)
--	g19075 = NOT(I25258)
--	g19078 = NOT(g18619)
--	I25264 = NOT(g17151)
--	g19081 = NOT(I25264)
--	I25272 = NOT(g17051)
--	g19091 = NOT(I25272)
--	g19096 = NOT(g18980)
--	I25283 = NOT(g17086)
--	g19098 = NOT(I25283)
--	I25294 = NOT(g17124)
--	g19105 = NOT(I25294)
--	I25303 = NOT(g17151)
--	g19110 = NOT(I25303)
--	I25308 = NOT(g16867)
--	g19113 = NOT(I25308)
--	I25315 = NOT(g16895)
--	g19118 = NOT(I25315)
--	I25320 = NOT(g16924)
--	g19125 = NOT(I25320)
--	I25325 = NOT(g16954)
--	g19132 = NOT(I25325)
--	I25334 = NOT(g17645)
--	g19145 = NOT(I25334)
--	I25338 = NOT(g17746)
--	g19147 = NOT(I25338)
--	I25344 = NOT(g17847)
--	g19151 = NOT(I25344)
--	I25351 = NOT(g17959)
--	g19156 = NOT(I25351)
--	I25355 = NOT(g18669)
--	g19158 = NOT(I25355)
--	I25358 = NOT(g18678)
--	g19159 = NOT(I25358)
--	I25365 = NOT(g18707)
--	g19164 = NOT(I25365)
--	I25371 = NOT(g18719)
--	g19168 = NOT(I25371)
--	I25374 = NOT(g18726)
--	g19169 = NOT(I25374)
--	I25377 = NOT(g18743)
--	g19170 = NOT(I25377)
--	I25383 = NOT(g18755)
--	g19174 = NOT(I25383)
--	I25386 = NOT(g18763)
--	g19175 = NOT(I25386)
--	I25389 = NOT(g18780)
--	g19176 = NOT(I25389)
--	I25395 = NOT(g18782)
--	g19180 = NOT(I25395)
--	I25399 = NOT(g18794)
--	g19182 = NOT(I25399)
--	I25402 = NOT(g18821)
--	g19183 = NOT(I25402)
--	I25406 = NOT(g18804)
--	g19185 = NOT(I25406)
--	I25412 = NOT(g18820)
--	g19189 = NOT(I25412)
--	I25415 = NOT(g18835)
--	g19190 = NOT(I25415)
--	I25423 = NOT(g18852)
--	g19196 = NOT(I25423)
--	I25426 = NOT(g18836)
--	g19197 = NOT(I25426)
--	I25429 = NOT(g18975)
--	g19198 = NOT(I25429)
--	I25432 = NOT(g18837)
--	g19199 = NOT(I25432)
--	I25442 = NOT(g18866)
--	g19207 = NOT(I25442)
--	I25445 = NOT(g18968)
--	g19208 = NOT(I25445)
--	I25456 = NOT(g18883)
--	g19217 = NOT(I25456)
--	I25459 = NOT(g18867)
--	g19218 = NOT(I25459)
--	I25463 = NOT(g18868)
--	g19220 = NOT(I25463)
--	I25474 = NOT(g18885)
--	g19229 = NOT(I25474)
--	I25486 = NOT(g18754)
--	g19237 = NOT(I25486)
--	I25489 = NOT(g18906)
--	g19238 = NOT(I25489)
--	I25492 = NOT(g18907)
--	g19239 = NOT(I25492)
--	I25506 = NOT(g18781)
--	g19247 = NOT(I25506)
--	I25510 = NOT(g18542)
--	g19249 = NOT(I25510)
--	g19251 = NOT(g16540)
--	I25525 = NOT(g18803)
--	g19258 = NOT(I25525)
--	I25528 = NOT(g18942)
--	g19259 = NOT(I25528)
--	g19265 = NOT(g16572)
--	I25557 = NOT(g18957)
--	g19270 = NOT(I25557)
--	I25567 = NOT(g17186)
--	g19272 = NOT(I25567)
--	g19280 = NOT(g16596)
--	g19287 = NOT(g16608)
--	I25612 = NOT(g17197)
--	g19291 = NOT(I25612)
--	g19299 = NOT(g16616)
--	g19301 = NOT(g16622)
--	g19302 = NOT(g17025)
--	g19305 = NOT(g16626)
--	I25660 = NOT(g17204)
--	g19309 = NOT(I25660)
--	g19319 = NOT(g16633)
--	g19322 = NOT(g16636)
--	g19323 = NOT(g17059)
--	g19326 = NOT(g16640)
--	I25717 = NOT(g17209)
--	g19330 = NOT(I25717)
--	I25728 = NOT(g17118)
--	g19335 = NOT(I25728)
--	g19346 = NOT(g16644)
--	g19349 = NOT(g16647)
--	g19350 = NOT(g17094)
--	g19353 = NOT(g16651)
--	I25768 = NOT(g17139)
--	g19358 = NOT(I25768)
--	I25778 = NOT(g17145)
--	g19369 = NOT(I25778)
--	g19380 = NOT(g16656)
--	g19383 = NOT(g16659)
--	g19384 = NOT(g17132)
--	g19387 = NOT(g16567)
--	g19388 = NOT(g17139)
--	I25816 = NOT(g17162)
--	g19390 = NOT(I25816)
--	I25826 = NOT(g17168)
--	g19401 = NOT(I25826)
--	g19412 = NOT(g16673)
--	g19415 = NOT(g16676)
--	g19417 = NOT(g16591)
--	g19418 = NOT(g17162)
--	I25862 = NOT(g17177)
--	g19420 = NOT(I25862)
--	I25872 = NOT(g17183)
--	g19431 = NOT(I25872)
--	g19441 = NOT(g17213)
--	g19444 = NOT(g17985)
--	g19448 = NOT(g16694)
--	g19452 = NOT(g16702)
--	g19454 = NOT(g16611)
--	g19455 = NOT(g17177)
--	I25904 = NOT(g17194)
--	g19457 = NOT(I25904)
--	g19467 = NOT(g16719)
--	g19468 = NOT(g17216)
--	g19471 = NOT(g18102)
--	g19475 = NOT(g16725)
--	g19479 = NOT(g16733)
--	g19481 = NOT(g16629)
--	g19482 = NOT(g17194)
--	g19483 = NOT(g16758)
--	g19484 = NOT(g16867)
--	g19490 = NOT(g16761)
--	g19491 = NOT(g17219)
--	g19494 = NOT(g18218)
--	g19498 = NOT(g16767)
--	g19502 = NOT(g16775)
--	g19504 = NOT(g16785)
--	g19505 = NOT(g16895)
--	g19511 = NOT(g16788)
--	g19512 = NOT(g17221)
--	g19515 = NOT(g18325)
--	g19519 = NOT(g16794)
--	g19523 = NOT(g16814)
--	g19524 = NOT(g16924)
--	g19530 = NOT(g16817)
--	g19533 = NOT(g16832)
--	g19534 = NOT(g16954)
--	I25966 = NOT(g16654)
--	g19543 = NOT(I25966)
--	I25971 = NOT(g16671)
--	g19546 = NOT(I25971)
--	I25977 = NOT(g16692)
--	g19550 = NOT(I25977)
--	I25985 = NOT(g16718)
--	g19556 = NOT(I25985)
--	I25994 = NOT(g16860)
--	g19563 = NOT(I25994)
--	I26006 = NOT(g16866)
--	g19573 = NOT(I26006)
--	g19577 = NOT(g16881)
--	g19578 = NOT(g16884)
--	I26025 = NOT(g16803)
--	g19595 = NOT(I26025)
--	I26028 = NOT(g16566)
--	g19596 = NOT(I26028)
--	g19607 = NOT(g16910)
--	g19608 = NOT(g16913)
--	I26051 = NOT(g16824)
--	g19622 = NOT(I26051)
--	g19640 = NOT(g16940)
--	g19641 = NOT(g16943)
--	I26078 = NOT(g16835)
--	g19652 = NOT(I26078)
--	I26085 = NOT(g18085)
--	g19657 = NOT(I26085)
--	g19680 = NOT(g16971)
--	g19681 = NOT(g16974)
--	I26112 = NOT(g16844)
--	g19689 = NOT(I26112)
--	I26115 = NOT(g16845)
--	g19690 = NOT(I26115)
--	I26123 = NOT(g17503)
--	g19696 = NOT(I26123)
--	I26134 = NOT(g18201)
--	g19705 = NOT(I26134)
--	I26154 = NOT(g16851)
--	g19725 = NOT(I26154)
--	I26171 = NOT(g17594)
--	g19740 = NOT(I26171)
--	I26182 = NOT(g18308)
--	g19749 = NOT(I26182)
--	I26195 = NOT(g16853)
--	g19762 = NOT(I26195)
--	I26198 = NOT(g16854)
--	g19763 = NOT(I26198)
--	I26220 = NOT(g17691)
--	g19783 = NOT(I26220)
--	I26231 = NOT(g18401)
--	g19792 = NOT(I26231)
--	I26237 = NOT(g16857)
--	g19798 = NOT(I26237)
--	I26266 = NOT(g17791)
--	g19825 = NOT(I26266)
--	g19830 = NOT(g18886)
--	I26276 = NOT(g16861)
--	g19838 = NOT(I26276)
--	I26334 = NOT(g18977)
--	g19890 = NOT(I26334)
--	I26337 = NOT(g16880)
--	g19893 = NOT(I26337)
--	I26340 = NOT(g17025)
--	g19894 = NOT(I26340)
--	I26365 = NOT(g18626)
--	g19915 = NOT(I26365)
--	g19918 = NOT(g18646)
--	I26369 = NOT(g17059)
--	g19919 = NOT(I26369)
--	g19933 = NOT(g18548)
--	I26388 = NOT(g17094)
--	g19934 = NOT(I26388)
--	I26401 = NOT(g17012)
--	g19945 = NOT(I26401)
--	g19948 = NOT(g17896)
--	g19950 = NOT(g18598)
--	I26407 = NOT(g17132)
--	g19951 = NOT(I26407)
--	I26413 = NOT(g16643)
--	g19957 = NOT(I26413)
--	I26420 = NOT(g17042)
--	g19972 = NOT(I26420)
--	g19975 = NOT(g18007)
--	g19977 = NOT(g18630)
--	I26426 = NOT(g16536)
--	g19978 = NOT(I26426)
--	I26437 = NOT(g16655)
--	g19987 = NOT(I26437)
--	I26444 = NOT(g17076)
--	g20002 = NOT(I26444)
--	g20005 = NOT(g18124)
--	g20007 = NOT(g18639)
--	I26458 = NOT(g17985)
--	g20016 = NOT(I26458)
--	I26469 = NOT(g16672)
--	g20025 = NOT(I26469)
--	I26476 = NOT(g17111)
--	g20040 = NOT(I26476)
--	g20043 = NOT(g18240)
--	I26481 = NOT(g18590)
--	g20045 = NOT(I26481)
--	I26494 = NOT(g18102)
--	g20058 = NOT(I26494)
--	I26505 = NOT(g16693)
--	g20067 = NOT(I26505)
--	I26512 = NOT(g16802)
--	g20082 = NOT(I26512)
--	g20083 = NOT(g17968)
--	I26535 = NOT(g18218)
--	g20099 = NOT(I26535)
--	I26545 = NOT(g16823)
--	g20105 = NOT(I26545)
--	I26574 = NOT(g18325)
--	g20124 = NOT(I26574)
--	g20127 = NOT(g18623)
--	g20140 = NOT(g16830)
--	g20163 = NOT(g17973)
--	I26612 = NOT(g17645)
--	g20164 = NOT(I26612)
--	g20178 = NOT(g16842)
--	g20193 = NOT(g18691)
--	I26642 = NOT(g17746)
--	g20198 = NOT(I26642)
--	g20212 = NOT(g16848)
--	g20223 = NOT(g18727)
--	I26664 = NOT(g17847)
--	g20228 = NOT(I26664)
--	g20242 = NOT(g16852)
--	g20250 = NOT(g18764)
--	I26679 = NOT(g17959)
--	g20255 = NOT(I26679)
--	g20269 = NOT(g17230)
--	g20273 = NOT(g18795)
--	g20278 = NOT(g17237)
--	g20279 = NOT(g17240)
--	g20281 = NOT(g17243)
--	g20286 = NOT(g17249)
--	g20287 = NOT(g17252)
--	g20288 = NOT(g17255)
--	g20289 = NOT(g17259)
--	g20290 = NOT(g17262)
--	g20292 = NOT(g17265)
--	I26714 = NOT(g17720)
--	g20295 = NOT(I26714)
--	g20296 = NOT(g17272)
--	g20297 = NOT(g17275)
--	g20298 = NOT(g17278)
--	g20302 = NOT(g17282)
--	g20303 = NOT(g17285)
--	g20304 = NOT(g17288)
--	g20305 = NOT(g17291)
--	g20306 = NOT(g17294)
--	g20308 = NOT(g17297)
--	g20311 = NOT(g17304)
--	g20312 = NOT(g17307)
--	g20313 = NOT(g17310)
--	g20315 = NOT(g17315)
--	g20316 = NOT(g17318)
--	g20317 = NOT(g17321)
--	g20321 = NOT(g17324)
--	g20322 = NOT(g17327)
--	g20323 = NOT(g17330)
--	g20324 = NOT(g17333)
--	g20325 = NOT(g17336)
--	g20327 = NOT(g17342)
--	g20328 = NOT(g17345)
--	g20329 = NOT(g17348)
--	g20330 = NOT(g17354)
--	g20331 = NOT(g17357)
--	g20332 = NOT(g17360)
--	g20334 = NOT(g17363)
--	g20335 = NOT(g17366)
--	g20336 = NOT(g17369)
--	g20340 = NOT(g17372)
--	g20341 = NOT(g17375)
--	g20342 = NOT(g17378)
--	g20344 = NOT(g17384)
--	g20345 = NOT(g17387)
--	g20346 = NOT(g17390)
--	g20347 = NOT(g17399)
--	g20348 = NOT(g17402)
--	g20349 = NOT(g17405)
--	g20350 = NOT(g17410)
--	g20351 = NOT(g17413)
--	g20352 = NOT(g17416)
--	g20354 = NOT(g17419)
--	g20355 = NOT(g17422)
--	g20356 = NOT(g17425)
--	I26777 = NOT(g17222)
--	g20360 = NOT(I26777)
--	g20361 = NOT(g17430)
--	g20362 = NOT(g17433)
--	g20363 = NOT(g17436)
--	g20364 = NOT(g17439)
--	g20365 = NOT(g17442)
--	g20366 = NOT(g17451)
--	g20367 = NOT(g17454)
--	g20368 = NOT(g17457)
--	g20369 = NOT(g17465)
--	g20370 = NOT(g17468)
--	g20371 = NOT(g17471)
--	g20372 = NOT(g17476)
--	g20373 = NOT(g17479)
--	g20374 = NOT(g17482)
--	I26796 = NOT(g17224)
--	g20377 = NOT(I26796)
--	g20378 = NOT(g17487)
--	g20379 = NOT(g17490)
--	g20380 = NOT(g17493)
--	g20381 = NOT(g17496)
--	g20382 = NOT(g17500)
--	g20383 = NOT(g17503)
--	g20384 = NOT(g17511)
--	g20385 = NOT(g17514)
--	g20386 = NOT(g17517)
--	g20387 = NOT(g17520)
--	g20388 = NOT(g17523)
--	g20389 = NOT(g17531)
--	g20390 = NOT(g17534)
--	g20391 = NOT(g17537)
--	g20392 = NOT(g17545)
--	g20393 = NOT(g17548)
--	g20394 = NOT(g17551)
--	I26816 = NOT(g17225)
--	g20395 = NOT(I26816)
--	I26819 = NOT(g17226)
--	g20396 = NOT(I26819)
--	g20397 = NOT(g17557)
--	g20398 = NOT(g17560)
--	g20399 = NOT(g17563)
--	g20400 = NOT(g17567)
--	g20401 = NOT(g17570)
--	g20402 = NOT(g17573)
--	g20403 = NOT(g17579)
--	g20404 = NOT(g17582)
--	g20405 = NOT(g17585)
--	g20406 = NOT(g17588)
--	g20407 = NOT(g17591)
--	g20408 = NOT(g17594)
--	g20409 = NOT(g17601)
--	g20410 = NOT(g17604)
--	g20411 = NOT(g17607)
--	g20412 = NOT(g17610)
--	g20413 = NOT(g17613)
--	g20414 = NOT(g17621)
--	g20415 = NOT(g17624)
--	g20416 = NOT(g17627)
--	I26843 = NOT(g17228)
--	g20418 = NOT(I26843)
--	I26846 = NOT(g17229)
--	g20419 = NOT(I26846)
--	g20420 = NOT(g17637)
--	g20421 = NOT(g17649)
--	g20422 = NOT(g17655)
--	g20423 = NOT(g17658)
--	g20424 = NOT(g17661)
--	g20425 = NOT(g17664)
--	g20426 = NOT(g17667)
--	g20427 = NOT(g17670)
--	g20428 = NOT(g17676)
--	g20429 = NOT(g17679)
--	g20430 = NOT(g17682)
--	g20431 = NOT(g17685)
--	g20432 = NOT(g17688)
--	g20433 = NOT(g17691)
--	g20434 = NOT(g17698)
--	g20435 = NOT(g17701)
--	g20436 = NOT(g17704)
--	g20437 = NOT(g17707)
--	g20438 = NOT(g17710)
--	I26868 = NOT(g17234)
--	g20439 = NOT(I26868)
--	I26871 = NOT(g17235)
--	g20440 = NOT(I26871)
--	I26874 = NOT(g17236)
--	g20441 = NOT(I26874)
--	g20442 = NOT(g17738)
--	g20443 = NOT(g17749)
--	g20444 = NOT(g17755)
--	g20445 = NOT(g17758)
--	g20446 = NOT(g17761)
--	g20447 = NOT(g17764)
--	g20448 = NOT(g17767)
--	g20449 = NOT(g17770)
--	g20450 = NOT(g17776)
--	g20451 = NOT(g17779)
--	g20452 = NOT(g17782)
--	g20453 = NOT(g17785)
--	g20454 = NOT(g17788)
--	g20455 = NOT(g17791)
--	g20456 = NOT(g17799)
--	I26892 = NOT(g17246)
--	g20457 = NOT(I26892)
--	I26895 = NOT(g17247)
--	g20458 = NOT(I26895)
--	I26898 = NOT(g17248)
--	g20459 = NOT(I26898)
--	g20461 = NOT(g17839)
--	g20462 = NOT(g17850)
--	g20463 = NOT(g17856)
--	g20464 = NOT(g17859)
--	g20465 = NOT(g17862)
--	g20466 = NOT(g17865)
--	g20467 = NOT(g17868)
--	g20468 = NOT(g17871)
--	I26910 = NOT(g17269)
--	g20469 = NOT(I26910)
--	I26913 = NOT(g17270)
--	g20470 = NOT(I26913)
--	I26916 = NOT(g17271)
--	g20471 = NOT(I26916)
--	g20476 = NOT(g17951)
--	g20477 = NOT(g17962)
--	I26923 = NOT(g17302)
--	g20478 = NOT(I26923)
--	I26926 = NOT(g17303)
--	g20479 = NOT(I26926)
--	I26931 = NOT(g17340)
--	g20484 = NOT(I26931)
--	I26934 = NOT(g17341)
--	g20485 = NOT(I26934)
--	g20490 = NOT(g18166)
--	I26940 = NOT(g17383)
--	g20491 = NOT(I26940)
--	g20496 = NOT(g18258)
--	I26947 = NOT(g17429)
--	g20498 = NOT(I26947)
--	g20500 = NOT(g18278)
--	g20501 = NOT(g18334)
--	g20504 = NOT(g18355)
--	g20505 = NOT(g18371)
--	g20507 = NOT(g18351)
--	I26960 = NOT(g16884)
--	g20513 = NOT(I26960)
--	g20516 = NOT(g18432)
--	g20517 = NOT(g18450)
--	g20518 = NOT(g18466)
--	I26966 = NOT(g17051)
--	g20519 = NOT(I26966)
--	g20526 = NOT(g18446)
--	I26972 = NOT(g16913)
--	g20531 = NOT(I26972)
--	g20534 = NOT(g18505)
--	g20535 = NOT(g18523)
--	g20536 = NOT(g18539)
--	I26980 = NOT(g17086)
--	g20539 = NOT(I26980)
--	g20545 = NOT(g18519)
--	I26985 = NOT(g16943)
--	g20550 = NOT(I26985)
--	g20553 = NOT(g18569)
--	g20554 = NOT(g18587)
--	I26990 = NOT(g19145)
--	g20555 = NOT(I26990)
--	I26993 = NOT(g19159)
--	g20556 = NOT(I26993)
--	I26996 = NOT(g19169)
--	g20557 = NOT(I26996)
--	I26999 = NOT(g19543)
--	g20558 = NOT(I26999)
--	I27002 = NOT(g19147)
--	g20559 = NOT(I27002)
--	I27005 = NOT(g19164)
--	g20560 = NOT(I27005)
--	I27008 = NOT(g19175)
--	g20561 = NOT(I27008)
--	I27011 = NOT(g19546)
--	g20562 = NOT(I27011)
--	I27014 = NOT(g19151)
--	g20563 = NOT(I27014)
--	I27017 = NOT(g19170)
--	g20564 = NOT(I27017)
--	I27020 = NOT(g19182)
--	g20565 = NOT(I27020)
--	I27023 = NOT(g19550)
--	g20566 = NOT(I27023)
--	I27026 = NOT(g19156)
--	g20567 = NOT(I27026)
--	I27029 = NOT(g19176)
--	g20568 = NOT(I27029)
--	I27032 = NOT(g19189)
--	g20569 = NOT(I27032)
--	I27035 = NOT(g19556)
--	g20570 = NOT(I27035)
--	I27038 = NOT(g20082)
--	g20571 = NOT(I27038)
--	I27041 = NOT(g19237)
--	g20572 = NOT(I27041)
--	I27044 = NOT(g19247)
--	g20573 = NOT(I27044)
--	I27047 = NOT(g19258)
--	g20574 = NOT(I27047)
--	I27050 = NOT(g19183)
--	g20575 = NOT(I27050)
--	I27053 = NOT(g19190)
--	g20576 = NOT(I27053)
--	I27056 = NOT(g19196)
--	g20577 = NOT(I27056)
--	I27059 = NOT(g19207)
--	g20578 = NOT(I27059)
--	I27062 = NOT(g19217)
--	g20579 = NOT(I27062)
--	I27065 = NOT(g19270)
--	g20580 = NOT(I27065)
--	I27068 = NOT(g19197)
--	g20581 = NOT(I27068)
--	I27071 = NOT(g19218)
--	g20582 = NOT(I27071)
--	I27074 = NOT(g19238)
--	g20583 = NOT(I27074)
--	I27077 = NOT(g19259)
--	g20584 = NOT(I27077)
--	I27080 = NOT(g19198)
--	g20585 = NOT(I27080)
--	I27083 = NOT(g19208)
--	g20586 = NOT(I27083)
--	I27086 = NOT(g19229)
--	g20587 = NOT(I27086)
--	I27089 = NOT(g20105)
--	g20588 = NOT(I27089)
--	I27092 = NOT(g19174)
--	g20589 = NOT(I27092)
--	I27095 = NOT(g19185)
--	g20590 = NOT(I27095)
--	I27098 = NOT(g19199)
--	g20591 = NOT(I27098)
--	I27101 = NOT(g19220)
--	g20592 = NOT(I27101)
--	I27104 = NOT(g19239)
--	g20593 = NOT(I27104)
--	I27107 = NOT(g19249)
--	g20594 = NOT(I27107)
--	I27110 = NOT(g19622)
--	g20595 = NOT(I27110)
--	I27113 = NOT(g19689)
--	g20596 = NOT(I27113)
--	I27116 = NOT(g19762)
--	g20597 = NOT(I27116)
--	I27119 = NOT(g19563)
--	g20598 = NOT(I27119)
--	I27122 = NOT(g19595)
--	g20599 = NOT(I27122)
--	I27125 = NOT(g19652)
--	g20600 = NOT(I27125)
--	I27128 = NOT(g19725)
--	g20601 = NOT(I27128)
--	I27131 = NOT(g19798)
--	g20602 = NOT(I27131)
--	I27134 = NOT(g19573)
--	g20603 = NOT(I27134)
--	I27137 = NOT(g19596)
--	g20604 = NOT(I27137)
--	I27140 = NOT(g19690)
--	g20605 = NOT(I27140)
--	I27143 = NOT(g19763)
--	g20606 = NOT(I27143)
--	I27146 = NOT(g19838)
--	g20607 = NOT(I27146)
--	I27149 = NOT(g19893)
--	g20608 = NOT(I27149)
--	I27152 = NOT(g20360)
--	g20609 = NOT(I27152)
--	I27155 = NOT(g20395)
--	g20610 = NOT(I27155)
--	I27158 = NOT(g20439)
--	g20611 = NOT(I27158)
--	I27161 = NOT(g20377)
--	g20612 = NOT(I27161)
--	I27164 = NOT(g20418)
--	g20613 = NOT(I27164)
--	I27167 = NOT(g20457)
--	g20614 = NOT(I27167)
--	I27170 = NOT(g20396)
--	g20615 = NOT(I27170)
--	I27173 = NOT(g20440)
--	g20616 = NOT(I27173)
--	I27176 = NOT(g20469)
--	g20617 = NOT(I27176)
--	I27179 = NOT(g20419)
--	g20618 = NOT(I27179)
--	I27182 = NOT(g20458)
--	g20619 = NOT(I27182)
--	I27185 = NOT(g20478)
--	g20620 = NOT(I27185)
--	I27188 = NOT(g20441)
--	g20621 = NOT(I27188)
--	I27191 = NOT(g20470)
--	g20622 = NOT(I27191)
--	I27194 = NOT(g20484)
--	g20623 = NOT(I27194)
--	I27197 = NOT(g20459)
--	g20624 = NOT(I27197)
--	I27200 = NOT(g20479)
--	g20625 = NOT(I27200)
--	I27203 = NOT(g20491)
--	g20626 = NOT(I27203)
--	I27206 = NOT(g20471)
--	g20627 = NOT(I27206)
--	I27209 = NOT(g20485)
--	g20628 = NOT(I27209)
--	I27212 = NOT(g20498)
--	g20629 = NOT(I27212)
--	I27215 = NOT(g19158)
--	g20630 = NOT(I27215)
--	I27218 = NOT(g19168)
--	g20631 = NOT(I27218)
--	I27221 = NOT(g19180)
--	g20632 = NOT(I27221)
--	I27225 = NOT(g19358)
--	g20634 = NOT(I27225)
--	I27228 = NOT(g19390)
--	g20637 = NOT(I27228)
--	I27232 = NOT(g19401)
--	g20641 = NOT(I27232)
--	I27235 = NOT(g19420)
--	g20644 = NOT(I27235)
--	I27240 = NOT(g19335)
--	g20649 = NOT(I27240)
--	I27243 = NOT(g19335)
--	g20652 = NOT(I27243)
--	I27246 = NOT(g19335)
--	g20655 = NOT(I27246)
--	I27250 = NOT(g19390)
--	g20659 = NOT(I27250)
--	I27253 = NOT(g19420)
--	g20662 = NOT(I27253)
--	I27257 = NOT(g19431)
--	g20666 = NOT(I27257)
--	I27260 = NOT(g19457)
--	g20669 = NOT(I27260)
--	I27264 = NOT(g19358)
--	g20673 = NOT(I27264)
--	I27267 = NOT(g19358)
--	g20676 = NOT(I27267)
--	I27270 = NOT(g19335)
--	g20679 = NOT(I27270)
--	I27275 = NOT(g19369)
--	g20684 = NOT(I27275)
--	I27278 = NOT(g19369)
--	g20687 = NOT(I27278)
--	I27281 = NOT(g19369)
--	g20690 = NOT(I27281)
--	I27285 = NOT(g19420)
--	g20694 = NOT(I27285)
--	I27288 = NOT(g19457)
--	g20697 = NOT(I27288)
--	I27293 = NOT(g19335)
--	g20704 = NOT(I27293)
--	I27297 = NOT(g19390)
--	g20708 = NOT(I27297)
--	I27300 = NOT(g19390)
--	g20711 = NOT(I27300)
--	I27303 = NOT(g19369)
--	g20714 = NOT(I27303)
--	I27308 = NOT(g19401)
--	g20719 = NOT(I27308)
--	I27311 = NOT(g19401)
--	g20722 = NOT(I27311)
--	I27314 = NOT(g19401)
--	g20725 = NOT(I27314)
--	I27318 = NOT(g19457)
--	g20729 = NOT(I27318)
--	I27321 = NOT(g19335)
--	g20732 = NOT(I27321)
--	I27324 = NOT(g19358)
--	g20735 = NOT(I27324)
--	I27328 = NOT(g19369)
--	g20739 = NOT(I27328)
--	I27332 = NOT(g19420)
--	g20743 = NOT(I27332)
--	I27335 = NOT(g19420)
--	g20746 = NOT(I27335)
--	I27338 = NOT(g19401)
--	g20749 = NOT(I27338)
--	I27343 = NOT(g19431)
--	g20754 = NOT(I27343)
--	I27346 = NOT(g19431)
--	g20757 = NOT(I27346)
--	I27349 = NOT(g19431)
--	g20760 = NOT(I27349)
--	I27352 = NOT(g19358)
--	g20763 = NOT(I27352)
--	I27355 = NOT(g19335)
--	g20766 = NOT(I27355)
--	I27358 = NOT(g19369)
--	g20769 = NOT(I27358)
--	I27361 = NOT(g19390)
--	g20772 = NOT(I27361)
--	I27365 = NOT(g19401)
--	g20776 = NOT(I27365)
--	I27369 = NOT(g19457)
--	g20780 = NOT(I27369)
--	I27372 = NOT(g19457)
--	g20783 = NOT(I27372)
--	I27375 = NOT(g19431)
--	g20786 = NOT(I27375)
--	I27379 = NOT(g19358)
--	g20790 = NOT(I27379)
--	I27382 = NOT(g19390)
--	g20793 = NOT(I27382)
--	I27385 = NOT(g19369)
--	g20796 = NOT(I27385)
--	I27388 = NOT(g19401)
--	g20799 = NOT(I27388)
--	I27391 = NOT(g19420)
--	g20802 = NOT(I27391)
--	I27395 = NOT(g19431)
--	g20806 = NOT(I27395)
--	I27399 = NOT(g19390)
--	g20810 = NOT(I27399)
--	I27402 = NOT(g19420)
--	g20813 = NOT(I27402)
--	I27405 = NOT(g19401)
--	g20816 = NOT(I27405)
--	I27408 = NOT(g19431)
--	g20819 = NOT(I27408)
--	I27411 = NOT(g19457)
--	g20822 = NOT(I27411)
--	I27416 = NOT(g19420)
--	g20827 = NOT(I27416)
--	I27419 = NOT(g19457)
--	g20830 = NOT(I27419)
--	I27422 = NOT(g19431)
--	g20833 = NOT(I27422)
--	I27426 = NOT(g19457)
--	g20837 = NOT(I27426)
--	g20842 = NOT(g19441)
--	g20850 = NOT(g19468)
--	g20858 = NOT(g19491)
--	g20866 = NOT(g19512)
--	g20885 = NOT(g19865)
--	g20904 = NOT(g19896)
--	g20928 = NOT(g19921)
--	I27488 = NOT(g20310)
--	g20942 = NOT(I27488)
--	I27491 = NOT(g20314)
--	g20943 = NOT(I27491)
--	g20956 = NOT(g19936)
--	I27516 = NOT(g20333)
--	g20971 = NOT(I27516)
--	I27531 = NOT(g20343)
--	g20984 = NOT(I27531)
--	I27534 = NOT(g20083)
--	g20985 = NOT(I27534)
--	I27537 = NOT(g19957)
--	g20986 = NOT(I27537)
--	I27549 = NOT(g20353)
--	g20998 = NOT(I27549)
--	I27565 = NOT(g19987)
--	g21012 = NOT(I27565)
--	I27577 = NOT(g20375)
--	g21024 = NOT(I27577)
--	I27585 = NOT(g20376)
--	g21030 = NOT(I27585)
--	I27593 = NOT(g20025)
--	g21036 = NOT(I27593)
--	g21050 = NOT(g20513)
--	I27614 = NOT(g20067)
--	g21057 = NOT(I27614)
--	I27621 = NOT(g20417)
--	g21064 = NOT(I27621)
--	g21066 = NOT(g20519)
--	g21069 = NOT(g20531)
--	g21076 = NOT(g20539)
--	g21079 = NOT(g20550)
--	I27646 = NOT(g20507)
--	g21087 = NOT(I27646)
--	g21090 = NOT(g19064)
--	g21093 = NOT(g19075)
--	I27658 = NOT(g20526)
--	g21099 = NOT(I27658)
--	g21102 = NOT(g19081)
--	I27667 = NOT(g20507)
--	g21108 = NOT(I27667)
--	I27672 = NOT(g20545)
--	g21113 = NOT(I27672)
--	I27684 = NOT(g20526)
--	g21125 = NOT(I27684)
--	I27689 = NOT(g19070)
--	g21130 = NOT(I27689)
--	I27705 = NOT(g20545)
--	g21144 = NOT(I27705)
--	I27727 = NOT(g19070)
--	g21164 = NOT(I27727)
--	I27749 = NOT(g19954)
--	g21184 = NOT(I27749)
--	g21187 = NOT(g19113)
--	I27766 = NOT(g19984)
--	g21199 = NOT(I27766)
--	g21202 = NOT(g19118)
--	I27779 = NOT(g20022)
--	g21214 = NOT(I27779)
--	g21217 = NOT(g19125)
--	I27785 = NOT(g20064)
--	g21222 = NOT(I27785)
--	g21225 = NOT(g19132)
--	g21241 = NOT(g19945)
--	g21249 = NOT(g19972)
--	g21258 = NOT(g20002)
--	g21266 = NOT(g20040)
--	I27822 = NOT(g19865)
--	g21271 = NOT(I27822)
--	I27827 = NOT(g19896)
--	g21278 = NOT(I27827)
--	I27832 = NOT(g19921)
--	g21285 = NOT(I27832)
--	I27838 = NOT(g19936)
--	g21293 = NOT(I27838)
--	I27868 = NOT(g19144)
--	g21327 = NOT(I27868)
--	I27897 = NOT(g19149)
--	g21358 = NOT(I27897)
--	I27900 = NOT(g19096)
--	g21359 = NOT(I27900)
--	I27917 = NOT(g19153)
--	g21376 = NOT(I27917)
--	I27920 = NOT(g19154)
--	g21377 = NOT(I27920)
--	I27927 = NOT(g19957)
--	g21382 = NOT(I27927)
--	I27942 = NOT(g19157)
--	g21399 = NOT(I27942)
--	g21400 = NOT(g19918)
--	I27949 = NOT(g19957)
--	g21404 = NOT(I27949)
--	I27958 = NOT(g19987)
--	g21415 = NOT(I27958)
--	I27969 = NOT(g19162)
--	g21426 = NOT(I27969)
--	I27972 = NOT(g19163)
--	g21427 = NOT(I27972)
--	I27976 = NOT(g19957)
--	g21429 = NOT(I27976)
--	I27984 = NOT(g19987)
--	g21441 = NOT(I27984)
--	I27992 = NOT(g20025)
--	g21449 = NOT(I27992)
--	I28000 = NOT(g19167)
--	g21457 = NOT(I28000)
--	I28003 = NOT(g19957)
--	g21458 = NOT(I28003)
--	g21461 = NOT(g19957)
--	I28009 = NOT(g20473)
--	g21473 = NOT(I28009)
--	I28013 = NOT(g19987)
--	g21477 = NOT(I28013)
--	I28019 = NOT(g20025)
--	g21483 = NOT(I28019)
--	I28027 = NOT(g20067)
--	g21491 = NOT(I28027)
--	I28031 = NOT(g19172)
--	g21495 = NOT(I28031)
--	I28034 = NOT(g19173)
--	g21496 = NOT(I28034)
--	I28038 = NOT(g19957)
--	g21498 = NOT(I28038)
--	I28043 = NOT(g19987)
--	g21505 = NOT(I28043)
--	g21508 = NOT(g19987)
--	I28047 = NOT(g20481)
--	g21514 = NOT(I28047)
--	I28051 = NOT(g20025)
--	g21518 = NOT(I28051)
--	I28057 = NOT(g20067)
--	g21524 = NOT(I28057)
--	I28061 = NOT(g19178)
--	g21528 = NOT(I28061)
--	g21529 = NOT(g19272)
--	I28065 = NOT(g19957)
--	g21530 = NOT(I28065)
--	I28072 = NOT(g19987)
--	g21537 = NOT(I28072)
--	I28076 = NOT(g20025)
--	g21541 = NOT(I28076)
--	g21544 = NOT(g20025)
--	I28080 = NOT(g20487)
--	g21550 = NOT(I28080)
--	I28084 = NOT(g20067)
--	g21554 = NOT(I28084)
--	I28087 = NOT(g19184)
--	g21557 = NOT(I28087)
--	I28090 = NOT(g20008)
--	g21558 = NOT(I28090)
--	I28093 = NOT(g19957)
--	g21561 = NOT(I28093)
--	g21565 = NOT(g19291)
--	I28100 = NOT(g19987)
--	g21566 = NOT(I28100)
--	I28107 = NOT(g20025)
--	g21573 = NOT(I28107)
--	I28111 = NOT(g20067)
--	g21577 = NOT(I28111)
--	g21580 = NOT(g20067)
--	I28115 = NOT(g20493)
--	g21586 = NOT(I28115)
--	I28119 = NOT(g19957)
--	g21590 = NOT(I28119)
--	I28123 = NOT(g19987)
--	g21594 = NOT(I28123)
--	g21598 = NOT(g19309)
--	I28130 = NOT(g20025)
--	g21599 = NOT(I28130)
--	I28137 = NOT(g20067)
--	g21606 = NOT(I28137)
--	I28143 = NOT(g19957)
--	g21612 = NOT(I28143)
--	I28148 = NOT(g19987)
--	g21619 = NOT(I28148)
--	I28152 = NOT(g20025)
--	g21623 = NOT(I28152)
--	g21627 = NOT(g19330)
--	I28159 = NOT(g20067)
--	g21628 = NOT(I28159)
--	I28169 = NOT(g19987)
--	g21640 = NOT(I28169)
--	I28174 = NOT(g20025)
--	g21647 = NOT(I28174)
--	I28178 = NOT(g20067)
--	g21651 = NOT(I28178)
--	I28184 = NOT(g19103)
--	g21655 = NOT(I28184)
--	g21661 = NOT(g19091)
--	I28201 = NOT(g20025)
--	g21671 = NOT(I28201)
--	I28206 = NOT(g20067)
--	g21678 = NOT(I28206)
--	I28210 = NOT(g20537)
--	g21682 = NOT(I28210)
--	g21690 = NOT(g19098)
--	I28229 = NOT(g20067)
--	g21700 = NOT(I28229)
--	I28235 = NOT(g20153)
--	g21708 = NOT(I28235)
--	g21716 = NOT(g19894)
--	g21726 = NOT(g19105)
--	g21742 = NOT(g19919)
--	g21752 = NOT(g19110)
--	g21766 = NOT(g19934)
--	g21782 = NOT(g19951)
--	I28314 = NOT(g19152)
--	g21795 = NOT(I28314)
--	I28357 = NOT(g20497)
--	g21824 = NOT(I28357)
--	I28360 = NOT(g20163)
--	g21825 = NOT(I28360)
--	g21861 = NOT(g19657)
--	g21867 = NOT(g19705)
--	g21872 = NOT(g19749)
--	g21876 = NOT(g19792)
--	g21883 = NOT(g19890)
--	g21886 = NOT(g19915)
--	g21895 = NOT(g19945)
--	g21902 = NOT(g19978)
--	g21907 = NOT(g19972)
--	I28432 = NOT(g19335)
--	g21914 = NOT(I28432)
--	I28435 = NOT(g19358)
--	g21917 = NOT(I28435)
--	g21921 = NOT(g20002)
--	g21927 = NOT(g20045)
--	I28443 = NOT(g19358)
--	g21928 = NOT(I28443)
--	I28447 = NOT(g19369)
--	g21932 = NOT(I28447)
--	I28450 = NOT(g19390)
--	g21935 = NOT(I28450)
--	g21939 = NOT(g20040)
--	I28455 = NOT(g20943)
--	g21943 = NOT(I28455)
--	I28458 = NOT(g20971)
--	g21944 = NOT(I28458)
--	I28461 = NOT(g20998)
--	g21945 = NOT(I28461)
--	I28464 = NOT(g21024)
--	g21946 = NOT(I28464)
--	I28467 = NOT(g20942)
--	g21947 = NOT(I28467)
--	I28470 = NOT(g20984)
--	g21948 = NOT(I28470)
--	I28473 = NOT(g21030)
--	g21949 = NOT(I28473)
--	I28476 = NOT(g21064)
--	g21950 = NOT(I28476)
--	I28479 = NOT(g21795)
--	g21951 = NOT(I28479)
--	I28482 = NOT(g21376)
--	g21952 = NOT(I28482)
--	I28485 = NOT(g21426)
--	g21953 = NOT(I28485)
--	I28488 = NOT(g21495)
--	g21954 = NOT(I28488)
--	I28491 = NOT(g21327)
--	g21955 = NOT(I28491)
--	I28494 = NOT(g21358)
--	g21956 = NOT(I28494)
--	I28497 = NOT(g21399)
--	g21957 = NOT(I28497)
--	I28500 = NOT(g21457)
--	g21958 = NOT(I28500)
--	I28503 = NOT(g21528)
--	g21959 = NOT(I28503)
--	I28506 = NOT(g21377)
--	g21960 = NOT(I28506)
--	I28509 = NOT(g21427)
--	g21961 = NOT(I28509)
--	I28512 = NOT(g21496)
--	g21962 = NOT(I28512)
--	I28515 = NOT(g21557)
--	g21963 = NOT(I28515)
--	I28518 = NOT(g20985)
--	g21964 = NOT(I28518)
--	I28521 = NOT(g21824)
--	g21965 = NOT(I28521)
--	I28524 = NOT(g21359)
--	g21966 = NOT(I28524)
--	I28527 = NOT(g21407)
--	g21967 = NOT(I28527)
--	I28541 = NOT(g21467)
--	g21982 = NOT(I28541)
--	I28550 = NOT(g21432)
--	g21995 = NOT(I28550)
--	I28557 = NOT(g21407)
--	g22003 = NOT(I28557)
--	I28564 = NOT(g21385)
--	g22014 = NOT(I28564)
--	I28628 = NOT(g21842)
--	g22082 = NOT(I28628)
--	I28649 = NOT(g21843)
--	g22107 = NOT(I28649)
--	I28671 = NOT(g21845)
--	g22133 = NOT(I28671)
--	I28693 = NOT(g21847)
--	g22156 = NOT(I28693)
--	I28712 = NOT(g21851)
--	g22176 = NOT(I28712)
--	g22212 = NOT(g21914)
--	g22213 = NOT(g21917)
--	g22217 = NOT(g21928)
--	I28781 = NOT(g21331)
--	g22219 = NOT(I28781)
--	g22221 = NOT(g21932)
--	g22222 = NOT(g21935)
--	I28789 = NOT(g21878)
--	g22225 = NOT(I28789)
--	I28792 = NOT(g21880)
--	g22226 = NOT(I28792)
--	g22230 = NOT(g20634)
--	I28800 = NOT(g21316)
--	g22232 = NOT(I28800)
--	g22233 = NOT(g20637)
--	g22236 = NOT(g20641)
--	g22237 = NOT(g20644)
--	g22239 = NOT(g20649)
--	g22240 = NOT(g20652)
--	g22241 = NOT(g20655)
--	I28813 = NOT(g21502)
--	g22243 = NOT(I28813)
--	g22246 = NOT(g20659)
--	g22248 = NOT(g20662)
--	g22251 = NOT(g20666)
--	g22252 = NOT(g20669)
--	I28825 = NOT(g21882)
--	g22253 = NOT(I28825)
--	g22256 = NOT(g20673)
--	g22257 = NOT(g20676)
--	g22258 = NOT(g20679)
--	I28833 = NOT(g21470)
--	g22259 = NOT(I28833)
--	g22260 = NOT(g20684)
--	g22261 = NOT(g20687)
--	g22262 = NOT(g20690)
--	g22266 = NOT(g20694)
--	g22268 = NOT(g20697)
--	g22271 = NOT(g20704)
--	g22274 = NOT(g20708)
--	g22275 = NOT(g20711)
--	g22276 = NOT(g20714)
--	g22277 = NOT(g20719)
--	g22278 = NOT(g20722)
--	g22279 = NOT(g20725)
--	g22283 = NOT(g20729)
--	g22286 = NOT(g20732)
--	g22287 = NOT(g20735)
--	g22290 = NOT(g20739)
--	g22293 = NOT(g20743)
--	g22294 = NOT(g20746)
--	g22295 = NOT(g20749)
--	g22296 = NOT(g20754)
--	g22297 = NOT(g20757)
--	g22298 = NOT(g20760)
--	I28876 = NOT(g21238)
--	g22300 = NOT(I28876)
--	g22303 = NOT(g20763)
--	g22304 = NOT(g20766)
--	g22306 = NOT(g20769)
--	g22307 = NOT(g20772)
--	g22310 = NOT(g20776)
--	g22313 = NOT(g20780)
--	g22314 = NOT(g20783)
--	g22315 = NOT(g20786)
--	g22316 = NOT(g21149)
--	g22318 = NOT(g20790)
--	g22319 = NOT(g21228)
--	I28896 = NOT(g21246)
--	g22328 = NOT(I28896)
--	g22331 = NOT(g20793)
--	g22332 = NOT(g20796)
--	g22334 = NOT(g20799)
--	g22335 = NOT(g20802)
--	g22338 = NOT(g20806)
--	g22341 = NOT(g21169)
--	g22343 = NOT(g20810)
--	g22344 = NOT(g21233)
--	I28913 = NOT(g21255)
--	g22353 = NOT(I28913)
--	g22356 = NOT(g20813)
--	g22357 = NOT(g20816)
--	g22359 = NOT(g20819)
--	g22360 = NOT(g20822)
--	g22364 = NOT(g21189)
--	g22366 = NOT(g20827)
--	g22367 = NOT(g21242)
--	I28928 = NOT(g21263)
--	g22376 = NOT(I28928)
--	g22379 = NOT(g20830)
--	g22380 = NOT(g20833)
--	g22384 = NOT(g21204)
--	g22386 = NOT(g20837)
--	g22387 = NOT(g21250)
--	g22401 = NOT(g21533)
--	g22402 = NOT(g21569)
--	g22403 = NOT(g21602)
--	g22404 = NOT(g21631)
--	I28949 = NOT(g21685)
--	g22405 = NOT(I28949)
--	g22408 = NOT(g20986)
--	I28953 = NOT(g21659)
--	g22409 = NOT(I28953)
--	I28956 = NOT(g21714)
--	g22412 = NOT(I28956)
--	I28959 = NOT(g21636)
--	g22415 = NOT(I28959)
--	I28962 = NOT(g21721)
--	g22418 = NOT(I28962)
--	g22421 = NOT(g21012)
--	I28966 = NOT(g20633)
--	g22422 = NOT(I28966)
--	I28969 = NOT(g21686)
--	g22425 = NOT(I28969)
--	I28972 = NOT(g21736)
--	g22428 = NOT(I28972)
--	I28975 = NOT(g21688)
--	g22431 = NOT(I28975)
--	I28978 = NOT(g21740)
--	g22434 = NOT(I28978)
--	I28981 = NOT(g21667)
--	g22437 = NOT(I28981)
--	I28984 = NOT(g21747)
--	g22440 = NOT(I28984)
--	g22443 = NOT(g21036)
--	I28988 = NOT(g20874)
--	g22444 = NOT(I28988)
--	I28991 = NOT(g20648)
--	g22445 = NOT(I28991)
--	I28994 = NOT(g21715)
--	g22448 = NOT(I28994)
--	I28997 = NOT(g21759)
--	g22451 = NOT(I28997)
--	I29001 = NOT(g20658)
--	g22455 = NOT(I29001)
--	I29004 = NOT(g21722)
--	g22458 = NOT(I29004)
--	I29007 = NOT(g21760)
--	g22461 = NOT(I29007)
--	I29010 = NOT(g21724)
--	g22464 = NOT(I29010)
--	I29013 = NOT(g21764)
--	g22467 = NOT(I29013)
--	I29016 = NOT(g21696)
--	g22470 = NOT(I29016)
--	I29019 = NOT(g21771)
--	g22473 = NOT(I29019)
--	g22476 = NOT(g21057)
--	I29023 = NOT(g20672)
--	g22477 = NOT(I29023)
--	I29026 = NOT(g21737)
--	g22480 = NOT(I29026)
--	I29030 = NOT(g20683)
--	g22484 = NOT(I29030)
--	I29033 = NOT(g21741)
--	g22487 = NOT(I29033)
--	I29036 = NOT(g21775)
--	g22490 = NOT(I29036)
--	I29040 = NOT(g20693)
--	g22494 = NOT(I29040)
--	I29043 = NOT(g21748)
--	g22497 = NOT(I29043)
--	I29046 = NOT(g21776)
--	g22500 = NOT(I29046)
--	I29049 = NOT(g21750)
--	g22503 = NOT(I29049)
--	I29052 = NOT(g21780)
--	g22506 = NOT(I29052)
--	I29055 = NOT(g21732)
--	g22509 = NOT(I29055)
--	I29058 = NOT(g20703)
--	g22512 = NOT(I29058)
--	I29064 = NOT(g20875)
--	g22518 = NOT(I29064)
--	I29067 = NOT(g20876)
--	g22519 = NOT(I29067)
--	I29070 = NOT(g20707)
--	g22520 = NOT(I29070)
--	I29073 = NOT(g21761)
--	g22523 = NOT(I29073)
--	I29077 = NOT(g20718)
--	g22527 = NOT(I29077)
--	I29080 = NOT(g21765)
--	g22530 = NOT(I29080)
--	I29083 = NOT(g21790)
--	g22533 = NOT(I29083)
--	I29087 = NOT(g20728)
--	g22537 = NOT(I29087)
--	I29090 = NOT(g21772)
--	g22540 = NOT(I29090)
--	I29093 = NOT(g21791)
--	g22543 = NOT(I29093)
--	g22547 = NOT(g21087)
--	I29098 = NOT(g20879)
--	g22548 = NOT(I29098)
--	I29101 = NOT(g20880)
--	g22549 = NOT(I29101)
--	I29104 = NOT(g20881)
--	g22550 = NOT(I29104)
--	I29107 = NOT(g21435)
--	g22551 = NOT(I29107)
--	I29110 = NOT(g20738)
--	g22552 = NOT(I29110)
--	I29116 = NOT(g20882)
--	g22558 = NOT(I29116)
--	I29119 = NOT(g20883)
--	g22559 = NOT(I29119)
--	I29122 = NOT(g20742)
--	g22560 = NOT(I29122)
--	I29125 = NOT(g21777)
--	g22563 = NOT(I29125)
--	I29129 = NOT(g20753)
--	g22567 = NOT(I29129)
--	I29132 = NOT(g21781)
--	g22570 = NOT(I29132)
--	I29135 = NOT(g21804)
--	g22573 = NOT(I29135)
--	I29142 = NOT(g20682)
--	g22582 = NOT(I29142)
--	I29145 = NOT(g20891)
--	g22583 = NOT(I29145)
--	I29148 = NOT(g20892)
--	g22584 = NOT(I29148)
--	I29151 = NOT(g20893)
--	g22585 = NOT(I29151)
--	I29154 = NOT(g20894)
--	g22586 = NOT(I29154)
--	g22588 = NOT(g21099)
--	I29159 = NOT(g20896)
--	g22589 = NOT(I29159)
--	I29162 = NOT(g20897)
--	g22590 = NOT(I29162)
--	I29165 = NOT(g20898)
--	g22591 = NOT(I29165)
--	I29168 = NOT(g20775)
--	g22592 = NOT(I29168)
--	I29174 = NOT(g20899)
--	g22598 = NOT(I29174)
--	I29177 = NOT(g20900)
--	g22599 = NOT(I29177)
--	I29180 = NOT(g20779)
--	g22600 = NOT(I29180)
--	I29183 = NOT(g21792)
--	g22603 = NOT(I29183)
--	g22609 = NOT(g21108)
--	I29191 = NOT(g20901)
--	g22611 = NOT(I29191)
--	I29194 = NOT(g20902)
--	g22612 = NOT(I29194)
--	I29197 = NOT(g20903)
--	g22613 = NOT(I29197)
--	I29203 = NOT(g20717)
--	g22619 = NOT(I29203)
--	I29206 = NOT(g20910)
--	g22620 = NOT(I29206)
--	I29209 = NOT(g20911)
--	g22621 = NOT(I29209)
--	I29212 = NOT(g20912)
--	g22622 = NOT(I29212)
--	I29215 = NOT(g20913)
--	g22623 = NOT(I29215)
--	g22625 = NOT(g21113)
--	I29220 = NOT(g20915)
--	g22626 = NOT(I29220)
--	I29223 = NOT(g20916)
--	g22627 = NOT(I29223)
--	I29226 = NOT(g20917)
--	g22628 = NOT(I29226)
--	I29229 = NOT(g20805)
--	g22629 = NOT(I29229)
--	I29235 = NOT(g20918)
--	g22635 = NOT(I29235)
--	I29238 = NOT(g20919)
--	g22636 = NOT(I29238)
--	I29243 = NOT(g20921)
--	g22639 = NOT(I29243)
--	I29246 = NOT(g20922)
--	g22640 = NOT(I29246)
--	I29249 = NOT(g20923)
--	g22641 = NOT(I29249)
--	I29252 = NOT(g20924)
--	g22642 = NOT(I29252)
--	g22645 = NOT(g21125)
--	I29259 = NOT(g20925)
--	g22647 = NOT(I29259)
--	I29262 = NOT(g20926)
--	g22648 = NOT(I29262)
--	I29265 = NOT(g20927)
--	g22649 = NOT(I29265)
--	I29271 = NOT(g20752)
--	g22655 = NOT(I29271)
--	I29274 = NOT(g20934)
--	g22656 = NOT(I29274)
--	I29277 = NOT(g20935)
--	g22657 = NOT(I29277)
--	I29280 = NOT(g20936)
--	g22658 = NOT(I29280)
--	I29283 = NOT(g20937)
--	g22659 = NOT(I29283)
--	g22661 = NOT(g21130)
--	I29288 = NOT(g20939)
--	g22662 = NOT(I29288)
--	I29291 = NOT(g20940)
--	g22663 = NOT(I29291)
--	I29294 = NOT(g20941)
--	g22664 = NOT(I29294)
--	I29301 = NOT(g20944)
--	g22669 = NOT(I29301)
--	I29304 = NOT(g20945)
--	g22670 = NOT(I29304)
--	I29307 = NOT(g20946)
--	g22671 = NOT(I29307)
--	I29310 = NOT(g20947)
--	g22672 = NOT(I29310)
--	I29313 = NOT(g20948)
--	g22673 = NOT(I29313)
--	I29317 = NOT(g20949)
--	g22675 = NOT(I29317)
--	I29320 = NOT(g20950)
--	g22676 = NOT(I29320)
--	I29323 = NOT(g20951)
--	g22677 = NOT(I29323)
--	I29326 = NOT(g20952)
--	g22678 = NOT(I29326)
--	g22681 = NOT(g21144)
--	I29333 = NOT(g20953)
--	g22683 = NOT(I29333)
--	I29336 = NOT(g20954)
--	g22684 = NOT(I29336)
--	I29339 = NOT(g20955)
--	g22685 = NOT(I29339)
--	I29345 = NOT(g20789)
--	g22691 = NOT(I29345)
--	I29348 = NOT(g20962)
--	g22692 = NOT(I29348)
--	I29351 = NOT(g20963)
--	g22693 = NOT(I29351)
--	I29354 = NOT(g20964)
--	g22694 = NOT(I29354)
--	I29357 = NOT(g20965)
--	g22695 = NOT(I29357)
--	I29360 = NOT(g21796)
--	g22696 = NOT(I29360)
--	I29366 = NOT(g20966)
--	g22702 = NOT(I29366)
--	I29369 = NOT(g20967)
--	g22703 = NOT(I29369)
--	I29372 = NOT(g20968)
--	g22704 = NOT(I29372)
--	I29375 = NOT(g20969)
--	g22705 = NOT(I29375)
--	I29378 = NOT(g20970)
--	g22706 = NOT(I29378)
--	I29383 = NOT(g20972)
--	g22709 = NOT(I29383)
--	I29386 = NOT(g20973)
--	g22710 = NOT(I29386)
--	I29389 = NOT(g20974)
--	g22711 = NOT(I29389)
--	I29392 = NOT(g20975)
--	g22712 = NOT(I29392)
--	I29395 = NOT(g20976)
--	g22713 = NOT(I29395)
--	I29399 = NOT(g20977)
--	g22715 = NOT(I29399)
--	I29402 = NOT(g20978)
--	g22716 = NOT(I29402)
--	I29405 = NOT(g20979)
--	g22717 = NOT(I29405)
--	I29408 = NOT(g20980)
--	g22718 = NOT(I29408)
--	g22721 = NOT(g21164)
--	I29415 = NOT(g20981)
--	g22723 = NOT(I29415)
--	I29418 = NOT(g20982)
--	g22724 = NOT(I29418)
--	I29421 = NOT(g20983)
--	g22725 = NOT(I29421)
--	I29426 = NOT(g20989)
--	g22728 = NOT(I29426)
--	I29429 = NOT(g20990)
--	g22729 = NOT(I29429)
--	I29432 = NOT(g20991)
--	g22730 = NOT(I29432)
--	I29435 = NOT(g20992)
--	g22731 = NOT(I29435)
--	I29439 = NOT(g20993)
--	g22733 = NOT(I29439)
--	I29442 = NOT(g20994)
--	g22734 = NOT(I29442)
--	I29445 = NOT(g20995)
--	g22735 = NOT(I29445)
--	I29448 = NOT(g20996)
--	g22736 = NOT(I29448)
--	I29451 = NOT(g20997)
--	g22737 = NOT(I29451)
--	I29456 = NOT(g20999)
--	g22740 = NOT(I29456)
--	I29459 = NOT(g21000)
--	g22741 = NOT(I29459)
--	I29462 = NOT(g21001)
--	g22742 = NOT(I29462)
--	I29465 = NOT(g21002)
--	g22743 = NOT(I29465)
--	I29468 = NOT(g21003)
--	g22744 = NOT(I29468)
--	I29472 = NOT(g21004)
--	g22746 = NOT(I29472)
--	I29475 = NOT(g21005)
--	g22747 = NOT(I29475)
--	I29478 = NOT(g21006)
--	g22748 = NOT(I29478)
--	I29481 = NOT(g21007)
--	g22749 = NOT(I29481)
--	I29484 = NOT(g21903)
--	g22750 = NOT(I29484)
--	g22753 = NOT(g21184)
--	I29490 = NOT(g21009)
--	g22756 = NOT(I29490)
--	I29493 = NOT(g21010)
--	g22757 = NOT(I29493)
--	I29496 = NOT(g21011)
--	g22758 = NOT(I29496)
--	I29500 = NOT(g21015)
--	g22760 = NOT(I29500)
--	I29503 = NOT(g21016)
--	g22761 = NOT(I29503)
--	I29506 = NOT(g21017)
--	g22762 = NOT(I29506)
--	I29509 = NOT(g21018)
--	g22763 = NOT(I29509)
--	I29513 = NOT(g21019)
--	g22765 = NOT(I29513)
--	I29516 = NOT(g21020)
--	g22766 = NOT(I29516)
--	I29519 = NOT(g21021)
--	g22767 = NOT(I29519)
--	I29522 = NOT(g21022)
--	g22768 = NOT(I29522)
--	I29525 = NOT(g21023)
--	g22769 = NOT(I29525)
--	I29530 = NOT(g21025)
--	g22772 = NOT(I29530)
--	I29533 = NOT(g21026)
--	g22773 = NOT(I29533)
--	I29536 = NOT(g21027)
--	g22774 = NOT(I29536)
--	I29539 = NOT(g21028)
--	g22775 = NOT(I29539)
--	I29542 = NOT(g21029)
--	g22776 = NOT(I29542)
--	g22777 = NOT(g21796)
--	I29547 = NOT(g21031)
--	g22785 = NOT(I29547)
--	I29550 = NOT(g21032)
--	g22786 = NOT(I29550)
--	g22787 = NOT(g21199)
--	I29556 = NOT(g21033)
--	g22790 = NOT(I29556)
--	I29559 = NOT(g21034)
--	g22791 = NOT(I29559)
--	I29562 = NOT(g21035)
--	g22792 = NOT(I29562)
--	I29566 = NOT(g21039)
--	g22794 = NOT(I29566)
--	I29569 = NOT(g21040)
--	g22795 = NOT(I29569)
--	I29572 = NOT(g21041)
--	g22796 = NOT(I29572)
--	I29575 = NOT(g21042)
--	g22797 = NOT(I29575)
--	I29579 = NOT(g21043)
--	g22799 = NOT(I29579)
--	I29582 = NOT(g21044)
--	g22800 = NOT(I29582)
--	I29585 = NOT(g21045)
--	g22801 = NOT(I29585)
--	I29588 = NOT(g21046)
--	g22802 = NOT(I29588)
--	I29591 = NOT(g21047)
--	g22803 = NOT(I29591)
--	g22805 = NOT(g21894)
--	g22806 = NOT(g21615)
--	I29600 = NOT(g21720)
--	g22812 = NOT(I29600)
--	I29603 = NOT(g21051)
--	g22824 = NOT(I29603)
--	I29606 = NOT(g21364)
--	g22825 = NOT(I29606)
--	I29610 = NOT(g21052)
--	g22827 = NOT(I29610)
--	I29613 = NOT(g21053)
--	g22828 = NOT(I29613)
--	g22829 = NOT(g21214)
--	I29619 = NOT(g21054)
--	g22832 = NOT(I29619)
--	I29622 = NOT(g21055)
--	g22833 = NOT(I29622)
--	I29625 = NOT(g21056)
--	g22834 = NOT(I29625)
--	I29629 = NOT(g21060)
--	g22836 = NOT(I29629)
--	I29632 = NOT(g21061)
--	g22837 = NOT(I29632)
--	I29635 = NOT(g21062)
--	g22838 = NOT(I29635)
--	I29638 = NOT(g21063)
--	g22839 = NOT(I29638)
--	I29641 = NOT(g20825)
--	g22840 = NOT(I29641)
--	g22843 = NOT(g21889)
--	g22847 = NOT(g21643)
--	I29653 = NOT(g21746)
--	g22852 = NOT(I29653)
--	I29656 = NOT(g21070)
--	g22864 = NOT(I29656)
--	I29660 = NOT(g21071)
--	g22866 = NOT(I29660)
--	I29663 = NOT(g21072)
--	g22867 = NOT(I29663)
--	g22868 = NOT(g21222)
--	I29669 = NOT(g21073)
--	g22871 = NOT(I29669)
--	I29672 = NOT(g21074)
--	g22872 = NOT(I29672)
--	I29675 = NOT(g21075)
--	g22873 = NOT(I29675)
--	g22875 = NOT(g21884)
--	g22882 = NOT(g21674)
--	I29687 = NOT(g21770)
--	g22887 = NOT(I29687)
--	I29690 = NOT(g21080)
--	g22899 = NOT(I29690)
--	I29694 = NOT(g21081)
--	g22901 = NOT(I29694)
--	I29697 = NOT(g21082)
--	g22902 = NOT(I29697)
--	I29700 = NOT(g20700)
--	g22903 = NOT(I29700)
--	g22907 = NOT(g21711)
--	g22917 = NOT(g21703)
--	I29712 = NOT(g21786)
--	g22922 = NOT(I29712)
--	I29715 = NOT(g21094)
--	g22934 = NOT(I29715)
--	I29724 = NOT(g21851)
--	g22945 = NOT(I29724)
--	I29727 = NOT(g20877)
--	g22948 = NOT(I29727)
--	g22949 = NOT(g21665)
--	g22954 = NOT(g21739)
--	g22958 = NOT(g21694)
--	g22962 = NOT(g21763)
--	g22966 = NOT(g21730)
--	I29736 = NOT(g20884)
--	g22970 = NOT(I29736)
--	g22971 = NOT(g21779)
--	g22975 = NOT(g21756)
--	I29741 = NOT(g21346)
--	g22979 = NOT(I29741)
--	g22980 = NOT(g21794)
--	g22986 = NOT(g21382)
--	g22988 = NOT(g21404)
--	g22989 = NOT(g21415)
--	g22991 = NOT(g21429)
--	g22995 = NOT(g21441)
--	g22996 = NOT(g21449)
--	g22998 = NOT(g21458)
--	g23001 = NOT(g21473)
--	g23002 = NOT(g21477)
--	g23006 = NOT(g21483)
--	g23007 = NOT(g21491)
--	g23008 = NOT(g21498)
--	g23012 = NOT(g21505)
--	g23015 = NOT(g21514)
--	g23016 = NOT(g21518)
--	g23020 = NOT(g21524)
--	g23021 = NOT(g21530)
--	g23024 = NOT(g21537)
--	g23028 = NOT(g21541)
--	g23031 = NOT(g21550)
--	g23032 = NOT(g21554)
--	g23036 = NOT(g21558)
--	g23037 = NOT(g21561)
--	g23038 = NOT(g21566)
--	g23041 = NOT(g21573)
--	g23045 = NOT(g21577)
--	g23048 = NOT(g21586)
--	g23049 = NOT(g21590)
--	I29797 = NOT(g21432)
--	g23050 = NOT(I29797)
--	I29802 = NOT(g21435)
--	g23055 = NOT(I29802)
--	g23056 = NOT(g21594)
--	g23057 = NOT(g21599)
--	g23060 = NOT(g21606)
--	g23064 = NOT(g21612)
--	I29812 = NOT(g21467)
--	g23065 = NOT(I29812)
--	I29817 = NOT(g21470)
--	g23068 = NOT(I29817)
--	g23069 = NOT(g21619)
--	g23074 = NOT(g21623)
--	g23075 = NOT(g21628)
--	I29827 = NOT(g21502)
--	g23078 = NOT(I29827)
--	g23079 = NOT(g21640)
--	g23082 = NOT(g21647)
--	g23087 = NOT(g21651)
--	g23088 = NOT(g21655)
--	I29841 = NOT(g21316)
--	g23094 = NOT(I29841)
--	g23095 = NOT(g21671)
--	g23098 = NOT(g21678)
--	g23103 = NOT(g21682)
--	I29852 = NOT(g21331)
--	g23105 = NOT(I29852)
--	g23112 = NOT(g21700)
--	g23115 = NOT(g21708)
--	I29863 = NOT(g21346)
--	g23116 = NOT(I29863)
--	I29872 = NOT(g21364)
--	g23125 = NOT(I29872)
--	I29881 = NOT(g21385)
--	g23134 = NOT(I29881)
--	g23140 = NOT(g21825)
--	g23141 = NOT(g21825)
--	g23142 = NOT(g21825)
--	g23143 = NOT(g21825)
--	g23144 = NOT(g21825)
--	g23145 = NOT(g21825)
--	g23146 = NOT(g21825)
--	g23147 = NOT(g21825)
--	I29897 = NOT(g23116)
--	g23148 = NOT(I29897)
--	I29900 = NOT(g23125)
--	g23149 = NOT(I29900)
--	I29903 = NOT(g23134)
--	g23150 = NOT(I29903)
--	I29906 = NOT(g21967)
--	g23151 = NOT(I29906)
--	I29909 = NOT(g23050)
--	g23152 = NOT(I29909)
--	I29912 = NOT(g23065)
--	g23153 = NOT(I29912)
--	I29915 = NOT(g23055)
--	g23154 = NOT(I29915)
--	I29918 = NOT(g23068)
--	g23155 = NOT(I29918)
--	I29921 = NOT(g23078)
--	g23156 = NOT(I29921)
--	I29924 = NOT(g23094)
--	g23157 = NOT(I29924)
--	I29927 = NOT(g23105)
--	g23158 = NOT(I29927)
--	I29930 = NOT(g22176)
--	g23159 = NOT(I29930)
--	I29933 = NOT(g22082)
--	g23160 = NOT(I29933)
--	I29936 = NOT(g22582)
--	g23161 = NOT(I29936)
--	I29939 = NOT(g22518)
--	g23162 = NOT(I29939)
--	I29942 = NOT(g22548)
--	g23163 = NOT(I29942)
--	I29945 = NOT(g22583)
--	g23164 = NOT(I29945)
--	I29948 = NOT(g22549)
--	g23165 = NOT(I29948)
--	I29951 = NOT(g22584)
--	g23166 = NOT(I29951)
--	I29954 = NOT(g22611)
--	g23167 = NOT(I29954)
--	I29957 = NOT(g22585)
--	g23168 = NOT(I29957)
--	I29960 = NOT(g22612)
--	g23169 = NOT(I29960)
--	I29963 = NOT(g22639)
--	g23170 = NOT(I29963)
--	I29966 = NOT(g22613)
--	g23171 = NOT(I29966)
--	I29969 = NOT(g22640)
--	g23172 = NOT(I29969)
--	I29972 = NOT(g22669)
--	g23173 = NOT(I29972)
--	I29975 = NOT(g22641)
--	g23174 = NOT(I29975)
--	I29978 = NOT(g22670)
--	g23175 = NOT(I29978)
--	I29981 = NOT(g22702)
--	g23176 = NOT(I29981)
--	I29984 = NOT(g22671)
--	g23177 = NOT(I29984)
--	I29987 = NOT(g22703)
--	g23178 = NOT(I29987)
--	I29990 = NOT(g22728)
--	g23179 = NOT(I29990)
--	I29993 = NOT(g22704)
--	g23180 = NOT(I29993)
--	I29996 = NOT(g22729)
--	g23181 = NOT(I29996)
--	I29999 = NOT(g22756)
--	g23182 = NOT(I29999)
--	I30002 = NOT(g22730)
--	g23183 = NOT(I30002)
--	I30005 = NOT(g22757)
--	g23184 = NOT(I30005)
--	I30008 = NOT(g22785)
--	g23185 = NOT(I30008)
--	I30011 = NOT(g22758)
--	g23186 = NOT(I30011)
--	I30014 = NOT(g22786)
--	g23187 = NOT(I30014)
--	I30017 = NOT(g22824)
--	g23188 = NOT(I30017)
--	I30020 = NOT(g22519)
--	g23189 = NOT(I30020)
--	I30023 = NOT(g22550)
--	g23190 = NOT(I30023)
--	I30026 = NOT(g22586)
--	g23191 = NOT(I30026)
--	I30029 = NOT(g22642)
--	g23192 = NOT(I30029)
--	I30032 = NOT(g22672)
--	g23193 = NOT(I30032)
--	I30035 = NOT(g22705)
--	g23194 = NOT(I30035)
--	I30038 = NOT(g22673)
--	g23195 = NOT(I30038)
--	I30041 = NOT(g22706)
--	g23196 = NOT(I30041)
--	I30044 = NOT(g22731)
--	g23197 = NOT(I30044)
--	I30047 = NOT(g22107)
--	g23198 = NOT(I30047)
--	I30050 = NOT(g22619)
--	g23199 = NOT(I30050)
--	I30053 = NOT(g22558)
--	g23200 = NOT(I30053)
--	I30056 = NOT(g22589)
--	g23201 = NOT(I30056)
--	I30059 = NOT(g22620)
--	g23202 = NOT(I30059)
--	I30062 = NOT(g22590)
--	g23203 = NOT(I30062)
--	I30065 = NOT(g22621)
--	g23204 = NOT(I30065)
--	I30068 = NOT(g22647)
--	g23205 = NOT(I30068)
--	I30071 = NOT(g22622)
--	g23206 = NOT(I30071)
--	I30074 = NOT(g22648)
--	g23207 = NOT(I30074)
--	I30077 = NOT(g22675)
--	g23208 = NOT(I30077)
--	I30080 = NOT(g22649)
--	g23209 = NOT(I30080)
--	I30083 = NOT(g22676)
--	g23210 = NOT(I30083)
--	I30086 = NOT(g22709)
--	g23211 = NOT(I30086)
--	I30089 = NOT(g22677)
--	g23212 = NOT(I30089)
--	I30092 = NOT(g22710)
--	g23213 = NOT(I30092)
--	I30095 = NOT(g22733)
--	g23214 = NOT(I30095)
--	I30098 = NOT(g22711)
--	g23215 = NOT(I30098)
--	I30101 = NOT(g22734)
--	g23216 = NOT(I30101)
--	I30104 = NOT(g22760)
--	g23217 = NOT(I30104)
--	I30107 = NOT(g22735)
--	g23218 = NOT(I30107)
--	I30110 = NOT(g22761)
--	g23219 = NOT(I30110)
--	I30113 = NOT(g22790)
--	g23220 = NOT(I30113)
--	I30116 = NOT(g22762)
--	g23221 = NOT(I30116)
--	I30119 = NOT(g22791)
--	g23222 = NOT(I30119)
--	I30122 = NOT(g22827)
--	g23223 = NOT(I30122)
--	I30125 = NOT(g22792)
--	g23224 = NOT(I30125)
--	I30128 = NOT(g22828)
--	g23225 = NOT(I30128)
--	I30131 = NOT(g22864)
--	g23226 = NOT(I30131)
--	I30134 = NOT(g22559)
--	g23227 = NOT(I30134)
--	I30137 = NOT(g22591)
--	g23228 = NOT(I30137)
--	I30140 = NOT(g22623)
--	g23229 = NOT(I30140)
--	I30143 = NOT(g22678)
--	g23230 = NOT(I30143)
--	I30146 = NOT(g22712)
--	g23231 = NOT(I30146)
--	I30149 = NOT(g22736)
--	g23232 = NOT(I30149)
--	I30152 = NOT(g22713)
--	g23233 = NOT(I30152)
--	I30155 = NOT(g22737)
--	g23234 = NOT(I30155)
--	I30158 = NOT(g22763)
--	g23235 = NOT(I30158)
--	I30161 = NOT(g22133)
--	g23236 = NOT(I30161)
--	I30164 = NOT(g22655)
--	g23237 = NOT(I30164)
--	I30167 = NOT(g22598)
--	g23238 = NOT(I30167)
--	I30170 = NOT(g22626)
--	g23239 = NOT(I30170)
--	I30173 = NOT(g22656)
--	g23240 = NOT(I30173)
--	I30176 = NOT(g22627)
--	g23241 = NOT(I30176)
--	I30179 = NOT(g22657)
--	g23242 = NOT(I30179)
--	I30182 = NOT(g22683)
--	g23243 = NOT(I30182)
--	I30185 = NOT(g22658)
--	g23244 = NOT(I30185)
--	I30188 = NOT(g22684)
--	g23245 = NOT(I30188)
--	I30191 = NOT(g22715)
--	g23246 = NOT(I30191)
--	I30194 = NOT(g22685)
--	g23247 = NOT(I30194)
--	I30197 = NOT(g22716)
--	g23248 = NOT(I30197)
--	I30200 = NOT(g22740)
--	g23249 = NOT(I30200)
--	I30203 = NOT(g22717)
--	g23250 = NOT(I30203)
--	I30206 = NOT(g22741)
--	g23251 = NOT(I30206)
--	I30209 = NOT(g22765)
--	g23252 = NOT(I30209)
--	I30212 = NOT(g22742)
--	g23253 = NOT(I30212)
--	I30215 = NOT(g22766)
--	g23254 = NOT(I30215)
--	I30218 = NOT(g22794)
--	g23255 = NOT(I30218)
--	I30221 = NOT(g22767)
--	g23256 = NOT(I30221)
--	I30224 = NOT(g22795)
--	g23257 = NOT(I30224)
--	I30227 = NOT(g22832)
--	g23258 = NOT(I30227)
--	I30230 = NOT(g22796)
--	g23259 = NOT(I30230)
--	I30233 = NOT(g22833)
--	g23260 = NOT(I30233)
--	I30236 = NOT(g22866)
--	g23261 = NOT(I30236)
--	I30239 = NOT(g22834)
--	g23262 = NOT(I30239)
--	I30242 = NOT(g22867)
--	g23263 = NOT(I30242)
--	I30245 = NOT(g22899)
--	g23264 = NOT(I30245)
--	I30248 = NOT(g22599)
--	g23265 = NOT(I30248)
--	I30251 = NOT(g22628)
--	g23266 = NOT(I30251)
--	I30254 = NOT(g22659)
--	g23267 = NOT(I30254)
--	I30257 = NOT(g22718)
--	g23268 = NOT(I30257)
--	I30260 = NOT(g22743)
--	g23269 = NOT(I30260)
--	I30263 = NOT(g22768)
--	g23270 = NOT(I30263)
--	I30266 = NOT(g22744)
--	g23271 = NOT(I30266)
--	I30269 = NOT(g22769)
--	g23272 = NOT(I30269)
--	I30272 = NOT(g22797)
--	g23273 = NOT(I30272)
--	I30275 = NOT(g22156)
--	g23274 = NOT(I30275)
--	I30278 = NOT(g22691)
--	g23275 = NOT(I30278)
--	I30281 = NOT(g22635)
--	g23276 = NOT(I30281)
--	I30284 = NOT(g22662)
--	g23277 = NOT(I30284)
--	I30287 = NOT(g22692)
--	g23278 = NOT(I30287)
--	I30290 = NOT(g22663)
--	g23279 = NOT(I30290)
--	I30293 = NOT(g22693)
--	g23280 = NOT(I30293)
--	I30296 = NOT(g22723)
--	g23281 = NOT(I30296)
--	I30299 = NOT(g22694)
--	g23282 = NOT(I30299)
--	I30302 = NOT(g22724)
--	g23283 = NOT(I30302)
--	I30305 = NOT(g22746)
--	g23284 = NOT(I30305)
--	I30308 = NOT(g22725)
--	g23285 = NOT(I30308)
--	I30311 = NOT(g22747)
--	g23286 = NOT(I30311)
--	I30314 = NOT(g22772)
--	g23287 = NOT(I30314)
--	I30317 = NOT(g22748)
--	g23288 = NOT(I30317)
--	I30320 = NOT(g22773)
--	g23289 = NOT(I30320)
--	I30323 = NOT(g22799)
--	g23290 = NOT(I30323)
--	I30326 = NOT(g22774)
--	g23291 = NOT(I30326)
--	I30329 = NOT(g22800)
--	g23292 = NOT(I30329)
--	I30332 = NOT(g22836)
--	g23293 = NOT(I30332)
--	I30335 = NOT(g22801)
--	g23294 = NOT(I30335)
--	I30338 = NOT(g22837)
--	g23295 = NOT(I30338)
--	I30341 = NOT(g22871)
--	g23296 = NOT(I30341)
--	I30344 = NOT(g22838)
--	g23297 = NOT(I30344)
--	I30347 = NOT(g22872)
--	g23298 = NOT(I30347)
--	I30350 = NOT(g22901)
--	g23299 = NOT(I30350)
--	I30353 = NOT(g22873)
--	g23300 = NOT(I30353)
--	I30356 = NOT(g22902)
--	g23301 = NOT(I30356)
--	I30359 = NOT(g22934)
--	g23302 = NOT(I30359)
--	I30362 = NOT(g22636)
--	g23303 = NOT(I30362)
--	I30365 = NOT(g22664)
--	g23304 = NOT(I30365)
--	I30368 = NOT(g22695)
--	g23305 = NOT(I30368)
--	I30371 = NOT(g22749)
--	g23306 = NOT(I30371)
--	I30374 = NOT(g22775)
--	g23307 = NOT(I30374)
--	I30377 = NOT(g22802)
--	g23308 = NOT(I30377)
--	I30380 = NOT(g22776)
--	g23309 = NOT(I30380)
--	I30383 = NOT(g22803)
--	g23310 = NOT(I30383)
--	I30386 = NOT(g22839)
--	g23311 = NOT(I30386)
--	I30389 = NOT(g22225)
--	g23312 = NOT(I30389)
--	I30392 = NOT(g22226)
--	g23313 = NOT(I30392)
--	I30395 = NOT(g22253)
--	g23314 = NOT(I30395)
--	I30398 = NOT(g22840)
--	g23315 = NOT(I30398)
--	I30401 = NOT(g22444)
--	g23316 = NOT(I30401)
--	I30404 = NOT(g22948)
--	g23317 = NOT(I30404)
--	I30407 = NOT(g22970)
--	g23318 = NOT(I30407)
--	g23403 = NOT(g23052)
--	g23410 = NOT(g23071)
--	g23415 = NOT(g23084)
--	g23420 = NOT(g23089)
--	g23424 = NOT(g23100)
--	g23429 = NOT(g23107)
--	g23435 = NOT(g23120)
--	I30467 = NOT(g23000)
--	g23438 = NOT(I30467)
--	I30470 = NOT(g23117)
--	g23439 = NOT(I30470)
--	g23441 = NOT(g23129)
--	g23444 = NOT(g22945)
--	I30476 = NOT(g22876)
--	g23448 = NOT(I30476)
--	I30480 = NOT(g23014)
--	g23452 = NOT(I30480)
--	I30483 = NOT(g23126)
--	g23453 = NOT(I30483)
--	I30486 = NOT(g23022)
--	g23454 = NOT(I30486)
--	I30489 = NOT(g22911)
--	g23455 = NOT(I30489)
--	I30493 = NOT(g23030)
--	g23459 = NOT(I30493)
--	I30496 = NOT(g23137)
--	g23460 = NOT(I30496)
--	I30501 = NOT(g23039)
--	g23463 = NOT(I30501)
--	I30504 = NOT(g22936)
--	g23464 = NOT(I30504)
--	I30508 = NOT(g23047)
--	g23468 = NOT(I30508)
--	I30511 = NOT(g21970)
--	g23469 = NOT(I30511)
--	g23470 = NOT(g22188)
--	I30516 = NOT(g23058)
--	g23472 = NOT(I30516)
--	I30519 = NOT(g22942)
--	g23473 = NOT(I30519)
--	I30525 = NOT(g23067)
--	g23481 = NOT(I30525)
--	g23482 = NOT(g22197)
--	I30531 = NOT(g23076)
--	g23485 = NOT(I30531)
--	I30536 = NOT(g23081)
--	g23492 = NOT(I30536)
--	g23493 = NOT(g22203)
--	I30544 = NOT(g23092)
--	g23500 = NOT(I30544)
--	I30547 = NOT(g23093)
--	g23501 = NOT(I30547)
--	I30552 = NOT(g23097)
--	g23508 = NOT(I30552)
--	g23509 = NOT(g22209)
--	I30560 = NOT(g23110)
--	g23516 = NOT(I30560)
--	I30563 = NOT(g23111)
--	g23517 = NOT(I30563)
--	I30568 = NOT(g23114)
--	g23524 = NOT(I30568)
--	I30575 = NOT(g23123)
--	g23531 = NOT(I30575)
--	I30578 = NOT(g23124)
--	g23532 = NOT(I30578)
--	I30586 = NOT(g23132)
--	g23542 = NOT(I30586)
--	I30589 = NOT(g23133)
--	g23543 = NOT(I30589)
--	I30594 = NOT(g22025)
--	g23546 = NOT(I30594)
--	I30598 = NOT(g22027)
--	g23548 = NOT(I30598)
--	I30601 = NOT(g22028)
--	g23549 = NOT(I30601)
--	I30607 = NOT(g22029)
--	g23553 = NOT(I30607)
--	I30611 = NOT(g22030)
--	g23555 = NOT(I30611)
--	I30614 = NOT(g22031)
--	g23556 = NOT(I30614)
--	I30617 = NOT(g22032)
--	g23557 = NOT(I30617)
--	I30623 = NOT(g22033)
--	g23561 = NOT(I30623)
--	I30626 = NOT(g22034)
--	g23562 = NOT(I30626)
--	I30632 = NOT(g22035)
--	g23566 = NOT(I30632)
--	I30636 = NOT(g22037)
--	g23568 = NOT(I30636)
--	I30639 = NOT(g22038)
--	g23569 = NOT(I30639)
--	I30642 = NOT(g22039)
--	g23570 = NOT(I30642)
--	I30648 = NOT(g22040)
--	g23574 = NOT(I30648)
--	I30651 = NOT(g22041)
--	g23575 = NOT(I30651)
--	I30654 = NOT(g22042)
--	g23576 = NOT(I30654)
--	I30660 = NOT(g22043)
--	g23580 = NOT(I30660)
--	I30663 = NOT(g22044)
--	g23581 = NOT(I30663)
--	I30669 = NOT(g22045)
--	g23585 = NOT(I30669)
--	I30673 = NOT(g22047)
--	g23587 = NOT(I30673)
--	I30676 = NOT(g22048)
--	g23588 = NOT(I30676)
--	I30679 = NOT(g22049)
--	g23589 = NOT(I30679)
--	I30686 = NOT(g23136)
--	g23594 = NOT(I30686)
--	I30689 = NOT(g22054)
--	g23595 = NOT(I30689)
--	I30692 = NOT(g22055)
--	g23596 = NOT(I30692)
--	I30695 = NOT(g22056)
--	g23597 = NOT(I30695)
--	I30701 = NOT(g22057)
--	g23601 = NOT(I30701)
--	I30704 = NOT(g22058)
--	g23602 = NOT(I30704)
--	I30707 = NOT(g22059)
--	g23603 = NOT(I30707)
--	I30713 = NOT(g22060)
--	g23607 = NOT(I30713)
--	I30716 = NOT(g22061)
--	g23608 = NOT(I30716)
--	I30722 = NOT(g22063)
--	g23612 = NOT(I30722)
--	I30725 = NOT(g22064)
--	g23613 = NOT(I30725)
--	I30728 = NOT(g22065)
--	g23614 = NOT(I30728)
--	I30735 = NOT(g22066)
--	g23619 = NOT(I30735)
--	I30738 = NOT(g22067)
--	g23620 = NOT(I30738)
--	I30741 = NOT(g22068)
--	g23621 = NOT(I30741)
--	I30748 = NOT(g21969)
--	g23626 = NOT(I30748)
--	I30751 = NOT(g22073)
--	g23627 = NOT(I30751)
--	I30754 = NOT(g22074)
--	g23628 = NOT(I30754)
--	I30757 = NOT(g22075)
--	g23629 = NOT(I30757)
--	I30763 = NOT(g22076)
--	g23633 = NOT(I30763)
--	I30766 = NOT(g22077)
--	g23634 = NOT(I30766)
--	I30769 = NOT(g22078)
--	g23635 = NOT(I30769)
--	I30776 = NOT(g22079)
--	g23640 = NOT(I30776)
--	I30779 = NOT(g22080)
--	g23641 = NOT(I30779)
--	I30782 = NOT(g22081)
--	g23642 = NOT(I30782)
--	I30786 = NOT(g22454)
--	g23644 = NOT(I30786)
--	I30797 = NOT(g22087)
--	g23661 = NOT(I30797)
--	I30800 = NOT(g22088)
--	g23662 = NOT(I30800)
--	I30803 = NOT(g22089)
--	g23663 = NOT(I30803)
--	I30810 = NOT(g22090)
--	g23668 = NOT(I30810)
--	I30813 = NOT(g22091)
--	g23669 = NOT(I30813)
--	I30816 = NOT(g22092)
--	g23670 = NOT(I30816)
--	I30823 = NOT(g21972)
--	g23675 = NOT(I30823)
--	I30826 = NOT(g22097)
--	g23676 = NOT(I30826)
--	I30829 = NOT(g22098)
--	g23677 = NOT(I30829)
--	I30832 = NOT(g22099)
--	g23678 = NOT(I30832)
--	I30838 = NOT(g22100)
--	g23682 = NOT(I30838)
--	I30841 = NOT(g22101)
--	g23683 = NOT(I30841)
--	I30844 = NOT(g22102)
--	g23684 = NOT(I30844)
--	I30847 = NOT(g22103)
--	g23685 = NOT(I30847)
--	I30854 = NOT(g22104)
--	g23690 = NOT(I30854)
--	I30857 = NOT(g22105)
--	g23691 = NOT(I30857)
--	I30860 = NOT(g22106)
--	g23692 = NOT(I30860)
--	I30864 = NOT(g22493)
--	g23694 = NOT(I30864)
--	I30875 = NOT(g22112)
--	g23711 = NOT(I30875)
--	I30878 = NOT(g22113)
--	g23712 = NOT(I30878)
--	I30881 = NOT(g22114)
--	g23713 = NOT(I30881)
--	I30888 = NOT(g22115)
--	g23718 = NOT(I30888)
--	I30891 = NOT(g22116)
--	g23719 = NOT(I30891)
--	I30894 = NOT(g22117)
--	g23720 = NOT(I30894)
--	I30901 = NOT(g21974)
--	g23725 = NOT(I30901)
--	I30905 = NOT(g22122)
--	g23727 = NOT(I30905)
--	I30908 = NOT(g22123)
--	g23728 = NOT(I30908)
--	I30911 = NOT(g22124)
--	g23729 = NOT(I30911)
--	I30914 = NOT(g22125)
--	g23730 = NOT(I30914)
--	I30917 = NOT(g22806)
--	g23731 = NOT(I30917)
--	I30922 = NOT(g22126)
--	g23736 = NOT(I30922)
--	I30925 = NOT(g22127)
--	g23737 = NOT(I30925)
--	I30928 = NOT(g22128)
--	g23738 = NOT(I30928)
--	I30931 = NOT(g22129)
--	g23739 = NOT(I30931)
--	I30938 = NOT(g22130)
--	g23744 = NOT(I30938)
--	I30941 = NOT(g22131)
--	g23745 = NOT(I30941)
--	I30944 = NOT(g22132)
--	g23746 = NOT(I30944)
--	I30948 = NOT(g22536)
--	g23748 = NOT(I30948)
--	I30959 = NOT(g22138)
--	g23765 = NOT(I30959)
--	I30962 = NOT(g22139)
--	g23766 = NOT(I30962)
--	I30965 = NOT(g22140)
--	g23767 = NOT(I30965)
--	I30973 = NOT(g22141)
--	g23773 = NOT(I30973)
--	I30976 = NOT(g22142)
--	g23774 = NOT(I30976)
--	I30979 = NOT(g22143)
--	g23775 = NOT(I30979)
--	I30985 = NOT(g22992)
--	g23779 = NOT(I30985)
--	I30988 = NOT(g22145)
--	g23782 = NOT(I30988)
--	I30991 = NOT(g22146)
--	g23783 = NOT(I30991)
--	I30994 = NOT(g22147)
--	g23784 = NOT(I30994)
--	I30997 = NOT(g22148)
--	g23785 = NOT(I30997)
--	I31000 = NOT(g22847)
--	g23786 = NOT(I31000)
--	I31005 = NOT(g22149)
--	g23791 = NOT(I31005)
--	I31008 = NOT(g22150)
--	g23792 = NOT(I31008)
--	I31011 = NOT(g22151)
--	g23793 = NOT(I31011)
--	I31014 = NOT(g22152)
--	g23794 = NOT(I31014)
--	I31021 = NOT(g22153)
--	g23799 = NOT(I31021)
--	I31024 = NOT(g22154)
--	g23800 = NOT(I31024)
--	I31027 = NOT(g22155)
--	g23801 = NOT(I31027)
--	I31031 = NOT(g22576)
--	g23803 = NOT(I31031)
--	I31043 = NOT(g22161)
--	g23821 = NOT(I31043)
--	I31050 = NOT(g22162)
--	g23826 = NOT(I31050)
--	I31053 = NOT(g22163)
--	g23827 = NOT(I31053)
--	I31056 = NOT(g22164)
--	g23828 = NOT(I31056)
--	I31062 = NOT(g23003)
--	g23832 = NOT(I31062)
--	I31065 = NOT(g22166)
--	g23835 = NOT(I31065)
--	I31068 = NOT(g22167)
--	g23836 = NOT(I31068)
--	I31071 = NOT(g22168)
--	g23837 = NOT(I31071)
--	I31074 = NOT(g22169)
--	g23838 = NOT(I31074)
--	I31077 = NOT(g22882)
--	g23839 = NOT(I31077)
--	I31082 = NOT(g22170)
--	g23844 = NOT(I31082)
--	I31085 = NOT(g22171)
--	g23845 = NOT(I31085)
--	I31088 = NOT(g22172)
--	g23846 = NOT(I31088)
--	I31091 = NOT(g22173)
--	g23847 = NOT(I31091)
--	g23853 = NOT(g22300)
--	I31102 = NOT(g22177)
--	g23856 = NOT(I31102)
--	I31109 = NOT(g22178)
--	g23861 = NOT(I31109)
--	I31112 = NOT(g22179)
--	g23862 = NOT(I31112)
--	I31115 = NOT(g22180)
--	g23863 = NOT(I31115)
--	I31121 = NOT(g23017)
--	g23867 = NOT(I31121)
--	I31124 = NOT(g22182)
--	g23870 = NOT(I31124)
--	I31127 = NOT(g22183)
--	g23871 = NOT(I31127)
--	I31130 = NOT(g22184)
--	g23872 = NOT(I31130)
--	I31133 = NOT(g22185)
--	g23873 = NOT(I31133)
--	I31136 = NOT(g22917)
--	g23874 = NOT(I31136)
--	I31141 = NOT(g22777)
--	g23879 = NOT(I31141)
--	I31144 = NOT(g22935)
--	g23882 = NOT(I31144)
--	g23885 = NOT(g22062)
--	g23887 = NOT(g22328)
--	I31152 = NOT(g22191)
--	g23890 = NOT(I31152)
--	I31159 = NOT(g22192)
--	g23895 = NOT(I31159)
--	I31162 = NOT(g22193)
--	g23896 = NOT(I31162)
--	I31165 = NOT(g22194)
--	g23897 = NOT(I31165)
--	I31171 = NOT(g23033)
--	g23901 = NOT(I31171)
--	g23905 = NOT(g22046)
--	g23908 = NOT(g22353)
--	I31181 = NOT(g22200)
--	g23911 = NOT(I31181)
--	I31188 = NOT(g21989)
--	g23916 = NOT(I31188)
--	g23918 = NOT(g22036)
--	I31195 = NOT(g22578)
--	g23923 = NOT(I31195)
--	g23940 = NOT(g22376)
--	I31205 = NOT(g22002)
--	g23943 = NOT(I31205)
--	I31213 = NOT(g22615)
--	g23955 = NOT(I31213)
--	I31226 = NOT(g22651)
--	g23984 = NOT(I31226)
--	I31232 = NOT(g22026)
--	g24000 = NOT(I31232)
--	I31235 = NOT(g22218)
--	g24001 = NOT(I31235)
--	I31244 = NOT(g22687)
--	g24014 = NOT(I31244)
--	I31250 = NOT(g22953)
--	g24030 = NOT(I31250)
--	I31253 = NOT(g22231)
--	g24033 = NOT(I31253)
--	I31257 = NOT(g22234)
--	g24035 = NOT(I31257)
--	g24047 = NOT(g23023)
--	I31266 = NOT(g22242)
--	g24051 = NOT(I31266)
--	I31270 = NOT(g22247)
--	g24053 = NOT(I31270)
--	I31274 = NOT(g22249)
--	g24055 = NOT(I31274)
--	g24060 = NOT(g23040)
--	I31282 = NOT(g22263)
--	g24064 = NOT(I31282)
--	I31286 = NOT(g22267)
--	g24066 = NOT(I31286)
--	I31290 = NOT(g22269)
--	g24068 = NOT(I31290)
--	g24073 = NOT(g23059)
--	I31298 = NOT(g22280)
--	g24077 = NOT(I31298)
--	I31302 = NOT(g22284)
--	g24079 = NOT(I31302)
--	g24084 = NOT(g23077)
--	I31310 = NOT(g22299)
--	g24088 = NOT(I31310)
--	g24094 = NOT(g22339)
--	g24095 = NOT(g22362)
--	g24096 = NOT(g22405)
--	g24097 = NOT(g22382)
--	g24098 = NOT(g22409)
--	g24099 = NOT(g22412)
--	g24101 = NOT(g22415)
--	g24102 = NOT(g22418)
--	g24103 = NOT(g22397)
--	g24104 = NOT(g22422)
--	g24105 = NOT(g22425)
--	g24106 = NOT(g22428)
--	g24107 = NOT(g22431)
--	g24108 = NOT(g22434)
--	g24110 = NOT(g22437)
--	g24111 = NOT(g22440)
--	g24112 = NOT(g22445)
--	g24113 = NOT(g22448)
--	g24114 = NOT(g22451)
--	g24115 = NOT(g22381)
--	g24121 = NOT(g22455)
--	g24122 = NOT(g22458)
--	g24123 = NOT(g22461)
--	g24124 = NOT(g22464)
--	g24125 = NOT(g22467)
--	g24127 = NOT(g22470)
--	g24128 = NOT(g22473)
--	g24129 = NOT(g22477)
--	g24130 = NOT(g22480)
--	g24131 = NOT(g22484)
--	g24132 = NOT(g22487)
--	g24133 = NOT(g22490)
--	g24134 = NOT(g22396)
--	g24140 = NOT(g22494)
--	g24141 = NOT(g22497)
--	g24142 = NOT(g22500)
--	g24143 = NOT(g22503)
--	g24144 = NOT(g22506)
--	g24146 = NOT(g22509)
--	g24147 = NOT(g22512)
--	g24148 = NOT(g22520)
--	g24149 = NOT(g22523)
--	g24150 = NOT(g22527)
--	g24151 = NOT(g22530)
--	g24152 = NOT(g22533)
--	g24153 = NOT(g22399)
--	g24159 = NOT(g22537)
--	g24160 = NOT(g22540)
--	g24161 = NOT(g22543)
--	g24162 = NOT(g22552)
--	g24163 = NOT(g22560)
--	g24164 = NOT(g22563)
--	g24165 = NOT(g22567)
--	g24166 = NOT(g22570)
--	g24167 = NOT(g22573)
--	g24168 = NOT(g22400)
--	g24175 = NOT(g22592)
--	g24176 = NOT(g22600)
--	g24177 = NOT(g22603)
--	g24180 = NOT(g22629)
--	I31387 = NOT(g22811)
--	g24183 = NOT(I31387)
--	g24210 = NOT(g22696)
--	g24220 = NOT(g22750)
--	I31417 = NOT(g22578)
--	g24233 = NOT(I31417)
--	I31426 = NOT(g22615)
--	g24240 = NOT(I31426)
--	I31436 = NOT(g22651)
--	g24248 = NOT(I31436)
--	g24251 = NOT(g22903)
--	I31445 = NOT(g22687)
--	g24255 = NOT(I31445)
--	I31451 = NOT(g23682)
--	g24259 = NOT(I31451)
--	I31454 = NOT(g23727)
--	g24260 = NOT(I31454)
--	I31457 = NOT(g23773)
--	g24261 = NOT(I31457)
--	I31460 = NOT(g23728)
--	g24262 = NOT(I31460)
--	I31463 = NOT(g23774)
--	g24263 = NOT(I31463)
--	I31466 = NOT(g23821)
--	g24264 = NOT(I31466)
--	I31469 = NOT(g23546)
--	g24265 = NOT(I31469)
--	I31472 = NOT(g23548)
--	g24266 = NOT(I31472)
--	I31475 = NOT(g23555)
--	g24267 = NOT(I31475)
--	I31478 = NOT(g23549)
--	g24268 = NOT(I31478)
--	I31481 = NOT(g23556)
--	g24269 = NOT(I31481)
--	I31484 = NOT(g23568)
--	g24270 = NOT(I31484)
--	I31487 = NOT(g23557)
--	g24271 = NOT(I31487)
--	I31490 = NOT(g23569)
--	g24272 = NOT(I31490)
--	I31493 = NOT(g23587)
--	g24273 = NOT(I31493)
--	I31496 = NOT(g23570)
--	g24274 = NOT(I31496)
--	I31499 = NOT(g23588)
--	g24275 = NOT(I31499)
--	I31502 = NOT(g23612)
--	g24276 = NOT(I31502)
--	I31505 = NOT(g23589)
--	g24277 = NOT(I31505)
--	I31508 = NOT(g23613)
--	g24278 = NOT(I31508)
--	I31511 = NOT(g23640)
--	g24279 = NOT(I31511)
--	I31514 = NOT(g23614)
--	g24280 = NOT(I31514)
--	I31517 = NOT(g23641)
--	g24281 = NOT(I31517)
--	I31520 = NOT(g23683)
--	g24282 = NOT(I31520)
--	I31523 = NOT(g23642)
--	g24283 = NOT(I31523)
--	I31526 = NOT(g23684)
--	g24284 = NOT(I31526)
--	I31529 = NOT(g23729)
--	g24285 = NOT(I31529)
--	I31532 = NOT(g23685)
--	g24286 = NOT(I31532)
--	I31535 = NOT(g23730)
--	g24287 = NOT(I31535)
--	I31538 = NOT(g23775)
--	g24288 = NOT(I31538)
--	I31541 = NOT(g23500)
--	g24289 = NOT(I31541)
--	I31544 = NOT(g23438)
--	g24290 = NOT(I31544)
--	I31547 = NOT(g23454)
--	g24291 = NOT(I31547)
--	I31550 = NOT(g23481)
--	g24292 = NOT(I31550)
--	I31553 = NOT(g23501)
--	g24293 = NOT(I31553)
--	I31556 = NOT(g23439)
--	g24294 = NOT(I31556)
--	I31559 = NOT(g24233)
--	g24295 = NOT(I31559)
--	I31562 = NOT(g23594)
--	g24296 = NOT(I31562)
--	I31565 = NOT(g24001)
--	g24297 = NOT(I31565)
--	I31568 = NOT(g24033)
--	g24298 = NOT(I31568)
--	I31571 = NOT(g24051)
--	g24299 = NOT(I31571)
--	I31574 = NOT(g23736)
--	g24300 = NOT(I31574)
--	I31577 = NOT(g23782)
--	g24301 = NOT(I31577)
--	I31580 = NOT(g23826)
--	g24302 = NOT(I31580)
--	I31583 = NOT(g23783)
--	g24303 = NOT(I31583)
--	I31586 = NOT(g23827)
--	g24304 = NOT(I31586)
--	I31589 = NOT(g23856)
--	g24305 = NOT(I31589)
--	I31592 = NOT(g23553)
--	g24306 = NOT(I31592)
--	I31595 = NOT(g23561)
--	g24307 = NOT(I31595)
--	I31598 = NOT(g23574)
--	g24308 = NOT(I31598)
--	I31601 = NOT(g23562)
--	g24309 = NOT(I31601)
--	I31604 = NOT(g23575)
--	g24310 = NOT(I31604)
--	I31607 = NOT(g23595)
--	g24311 = NOT(I31607)
--	I31610 = NOT(g23576)
--	g24312 = NOT(I31610)
--	I31613 = NOT(g23596)
--	g24313 = NOT(I31613)
--	I31616 = NOT(g23619)
--	g24314 = NOT(I31616)
--	I31619 = NOT(g23597)
--	g24315 = NOT(I31619)
--	I31622 = NOT(g23620)
--	g24316 = NOT(I31622)
--	I31625 = NOT(g23661)
--	g24317 = NOT(I31625)
--	I31628 = NOT(g23621)
--	g24318 = NOT(I31628)
--	I31631 = NOT(g23662)
--	g24319 = NOT(I31631)
--	I31634 = NOT(g23690)
--	g24320 = NOT(I31634)
--	I31637 = NOT(g23663)
--	g24321 = NOT(I31637)
--	I31640 = NOT(g23691)
--	g24322 = NOT(I31640)
--	I31643 = NOT(g23737)
--	g24323 = NOT(I31643)
--	I31646 = NOT(g23692)
--	g24324 = NOT(I31646)
--	I31649 = NOT(g23738)
--	g24325 = NOT(I31649)
--	I31652 = NOT(g23784)
--	g24326 = NOT(I31652)
--	I31655 = NOT(g23739)
--	g24327 = NOT(I31655)
--	I31658 = NOT(g23785)
--	g24328 = NOT(I31658)
--	I31661 = NOT(g23828)
--	g24329 = NOT(I31661)
--	I31664 = NOT(g23516)
--	g24330 = NOT(I31664)
--	I31667 = NOT(g23452)
--	g24331 = NOT(I31667)
--	I31670 = NOT(g23463)
--	g24332 = NOT(I31670)
--	I31673 = NOT(g23492)
--	g24333 = NOT(I31673)
--	I31676 = NOT(g23517)
--	g24334 = NOT(I31676)
--	I31679 = NOT(g23453)
--	g24335 = NOT(I31679)
--	I31682 = NOT(g24240)
--	g24336 = NOT(I31682)
--	I31685 = NOT(g23626)
--	g24337 = NOT(I31685)
--	I31688 = NOT(g24035)
--	g24338 = NOT(I31688)
--	I31691 = NOT(g24053)
--	g24339 = NOT(I31691)
--	I31694 = NOT(g24064)
--	g24340 = NOT(I31694)
--	I31697 = NOT(g23791)
--	g24341 = NOT(I31697)
--	I31700 = NOT(g23835)
--	g24342 = NOT(I31700)
--	I31703 = NOT(g23861)
--	g24343 = NOT(I31703)
--	I31706 = NOT(g23836)
--	g24344 = NOT(I31706)
--	I31709 = NOT(g23862)
--	g24345 = NOT(I31709)
--	I31712 = NOT(g23890)
--	g24346 = NOT(I31712)
--	I31715 = NOT(g23566)
--	g24347 = NOT(I31715)
--	I31718 = NOT(g23580)
--	g24348 = NOT(I31718)
--	I31721 = NOT(g23601)
--	g24349 = NOT(I31721)
--	I31724 = NOT(g23581)
--	g24350 = NOT(I31724)
--	I31727 = NOT(g23602)
--	g24351 = NOT(I31727)
--	I31730 = NOT(g23627)
--	g24352 = NOT(I31730)
--	I31733 = NOT(g23603)
--	g24353 = NOT(I31733)
--	I31736 = NOT(g23628)
--	g24354 = NOT(I31736)
--	I31739 = NOT(g23668)
--	g24355 = NOT(I31739)
--	I31742 = NOT(g23629)
--	g24356 = NOT(I31742)
--	I31745 = NOT(g23669)
--	g24357 = NOT(I31745)
--	I31748 = NOT(g23711)
--	g24358 = NOT(I31748)
--	I31751 = NOT(g23670)
--	g24359 = NOT(I31751)
--	I31754 = NOT(g23712)
--	g24360 = NOT(I31754)
--	I31757 = NOT(g23744)
--	g24361 = NOT(I31757)
--	I31760 = NOT(g23713)
--	g24362 = NOT(I31760)
--	I31763 = NOT(g23745)
--	g24363 = NOT(I31763)
--	I31766 = NOT(g23792)
--	g24364 = NOT(I31766)
--	I31769 = NOT(g23746)
--	g24365 = NOT(I31769)
--	I31772 = NOT(g23793)
--	g24366 = NOT(I31772)
--	I31775 = NOT(g23837)
--	g24367 = NOT(I31775)
--	I31778 = NOT(g23794)
--	g24368 = NOT(I31778)
--	I31781 = NOT(g23838)
--	g24369 = NOT(I31781)
--	I31784 = NOT(g23863)
--	g24370 = NOT(I31784)
--	I31787 = NOT(g23531)
--	g24371 = NOT(I31787)
--	I31790 = NOT(g23459)
--	g24372 = NOT(I31790)
--	I31793 = NOT(g23472)
--	g24373 = NOT(I31793)
--	I31796 = NOT(g23508)
--	g24374 = NOT(I31796)
--	I31799 = NOT(g23532)
--	g24375 = NOT(I31799)
--	I31802 = NOT(g23460)
--	g24376 = NOT(I31802)
--	I31805 = NOT(g24248)
--	g24377 = NOT(I31805)
--	I31808 = NOT(g23675)
--	g24378 = NOT(I31808)
--	I31811 = NOT(g24055)
--	g24379 = NOT(I31811)
--	I31814 = NOT(g24066)
--	g24380 = NOT(I31814)
--	I31817 = NOT(g24077)
--	g24381 = NOT(I31817)
--	I31820 = NOT(g23844)
--	g24382 = NOT(I31820)
--	I31823 = NOT(g23870)
--	g24383 = NOT(I31823)
--	I31826 = NOT(g23895)
--	g24384 = NOT(I31826)
--	I31829 = NOT(g23871)
--	g24385 = NOT(I31829)
--	I31832 = NOT(g23896)
--	g24386 = NOT(I31832)
--	I31835 = NOT(g23911)
--	g24387 = NOT(I31835)
--	I31838 = NOT(g23585)
--	g24388 = NOT(I31838)
--	I31841 = NOT(g23607)
--	g24389 = NOT(I31841)
--	I31844 = NOT(g23633)
--	g24390 = NOT(I31844)
--	I31847 = NOT(g23608)
--	g24391 = NOT(I31847)
--	I31850 = NOT(g23634)
--	g24392 = NOT(I31850)
--	I31853 = NOT(g23676)
--	g24393 = NOT(I31853)
--	I31856 = NOT(g23635)
--	g24394 = NOT(I31856)
--	I31859 = NOT(g23677)
--	g24395 = NOT(I31859)
--	I31862 = NOT(g23718)
--	g24396 = NOT(I31862)
--	I31865 = NOT(g23678)
--	g24397 = NOT(I31865)
--	I31868 = NOT(g23719)
--	g24398 = NOT(I31868)
--	I31871 = NOT(g23765)
--	g24399 = NOT(I31871)
--	I31874 = NOT(g23720)
--	g24400 = NOT(I31874)
--	I31877 = NOT(g23766)
--	g24401 = NOT(I31877)
--	I31880 = NOT(g23799)
--	g24402 = NOT(I31880)
--	I31883 = NOT(g23767)
--	g24403 = NOT(I31883)
--	I31886 = NOT(g23800)
--	g24404 = NOT(I31886)
--	I31889 = NOT(g23845)
--	g24405 = NOT(I31889)
--	I31892 = NOT(g23801)
--	g24406 = NOT(I31892)
--	I31895 = NOT(g23846)
--	g24407 = NOT(I31895)
--	I31898 = NOT(g23872)
--	g24408 = NOT(I31898)
--	I31901 = NOT(g23847)
--	g24409 = NOT(I31901)
--	I31904 = NOT(g23873)
--	g24410 = NOT(I31904)
--	I31907 = NOT(g23897)
--	g24411 = NOT(I31907)
--	I31910 = NOT(g23542)
--	g24412 = NOT(I31910)
--	I31913 = NOT(g23468)
--	g24413 = NOT(I31913)
--	I31916 = NOT(g23485)
--	g24414 = NOT(I31916)
--	I31919 = NOT(g23524)
--	g24415 = NOT(I31919)
--	I31922 = NOT(g23543)
--	g24416 = NOT(I31922)
--	I31925 = NOT(g23469)
--	g24417 = NOT(I31925)
--	I31928 = NOT(g24255)
--	g24418 = NOT(I31928)
--	I31931 = NOT(g23725)
--	g24419 = NOT(I31931)
--	I31934 = NOT(g24068)
--	g24420 = NOT(I31934)
--	I31937 = NOT(g24079)
--	g24421 = NOT(I31937)
--	I31940 = NOT(g24088)
--	g24422 = NOT(I31940)
--	I31943 = NOT(g24000)
--	g24423 = NOT(I31943)
--	I31946 = NOT(g23916)
--	g24424 = NOT(I31946)
--	I31949 = NOT(g23943)
--	g24425 = NOT(I31949)
--	g24482 = NOT(g24183)
--	I32042 = NOT(g23399)
--	g24518 = NOT(I32042)
--	I32057 = NOT(g23406)
--	g24531 = NOT(I32057)
--	I32067 = NOT(g24174)
--	g24539 = NOT(I32067)
--	I32074 = NOT(g23413)
--	g24544 = NOT(I32074)
--	I32081 = NOT(g24178)
--	g24549 = NOT(I32081)
--	I32085 = NOT(g24179)
--	g24551 = NOT(I32085)
--	I32092 = NOT(g23418)
--	g24556 = NOT(I32092)
--	I32098 = NOT(g24181)
--	g24560 = NOT(I32098)
--	I32102 = NOT(g24182)
--	g24562 = NOT(I32102)
--	I32109 = NOT(g24206)
--	g24567 = NOT(I32109)
--	I32112 = NOT(g24207)
--	g24568 = NOT(I32112)
--	I32116 = NOT(g24208)
--	g24570 = NOT(I32116)
--	I32120 = NOT(g24209)
--	g24572 = NOT(I32120)
--	I32126 = NOT(g24212)
--	g24576 = NOT(I32126)
--	I32129 = NOT(g24213)
--	g24577 = NOT(I32129)
--	I32133 = NOT(g24214)
--	g24579 = NOT(I32133)
--	I32137 = NOT(g24215)
--	g24581 = NOT(I32137)
--	I32140 = NOT(g24216)
--	g24582 = NOT(I32140)
--	I32143 = NOT(g24218)
--	g24583 = NOT(I32143)
--	I32146 = NOT(g24219)
--	g24584 = NOT(I32146)
--	I32150 = NOT(g24222)
--	g24586 = NOT(I32150)
--	I32153 = NOT(g24223)
--	g24587 = NOT(I32153)
--	I32156 = NOT(g24225)
--	g24588 = NOT(I32156)
--	I32159 = NOT(g24226)
--	g24589 = NOT(I32159)
--	I32164 = NOT(g24228)
--	g24592 = NOT(I32164)
--	I32167 = NOT(g24230)
--	g24593 = NOT(I32167)
--	I32170 = NOT(g24231)
--	g24594 = NOT(I32170)
--	I32175 = NOT(g24235)
--	g24597 = NOT(I32175)
--	I32178 = NOT(g24237)
--	g24598 = NOT(I32178)
--	I32181 = NOT(g24238)
--	g24599 = NOT(I32181)
--	I32184 = NOT(g23497)
--	g24600 = NOT(I32184)
--	I32189 = NOT(g24243)
--	g24605 = NOT(I32189)
--	I32193 = NOT(g23513)
--	g24607 = NOT(I32193)
--	I32198 = NOT(g24250)
--	g24612 = NOT(I32198)
--	I32203 = NOT(g23528)
--	g24619 = NOT(I32203)
--	I32210 = NOT(g23539)
--	g24630 = NOT(I32210)
--	g24648 = NOT(g23470)
--	g24668 = NOT(g23482)
--	g24687 = NOT(g23493)
--	g24704 = NOT(g23509)
--	I32248 = NOT(g23919)
--	g24734 = NOT(I32248)
--	I32251 = NOT(g23919)
--	g24735 = NOT(I32251)
--	I32281 = NOT(g23950)
--	g24763 = NOT(I32281)
--	I32320 = NOT(g23979)
--	g24784 = NOT(I32320)
--	I32365 = NOT(g24009)
--	g24805 = NOT(I32365)
--	g24815 = NOT(g23448)
--	I32388 = NOT(g23385)
--	g24816 = NOT(I32388)
--	I32419 = NOT(g24043)
--	g24827 = NOT(I32419)
--	g24834 = NOT(g23455)
--	I32439 = NOT(g23392)
--	g24835 = NOT(I32439)
--	g24850 = NOT(g23464)
--	I32487 = NOT(g23400)
--	g24851 = NOT(I32487)
--	I32506 = NOT(g23324)
--	g24856 = NOT(I32506)
--	g24864 = NOT(g23473)
--	I32535 = NOT(g23407)
--	g24865 = NOT(I32535)
--	I32556 = NOT(g23329)
--	g24872 = NOT(I32556)
--	I32583 = NOT(g23330)
--	g24879 = NOT(I32583)
--	I32604 = NOT(g23339)
--	g24886 = NOT(I32604)
--	g24893 = NOT(g23486)
--	I32642 = NOT(g23348)
--	g24903 = NOT(I32642)
--	g24912 = NOT(g23495)
--	g24916 = NOT(g23502)
--	g24929 = NOT(g23511)
--	g24933 = NOT(g23518)
--	g24939 = NOT(g23660)
--	g24941 = NOT(g23526)
--	g24945 = NOT(g23533)
--	I32704 = NOT(g23357)
--	g24949 = NOT(I32704)
--	g24950 = NOT(g23710)
--	g24952 = NOT(g23537)
--	I32716 = NOT(g23358)
--	g24956 = NOT(I32716)
--	I32719 = NOT(g23359)
--	g24957 = NOT(I32719)
--	g24958 = NOT(g23478)
--	g24962 = NOT(g23764)
--	g24969 = NOT(g23489)
--	g24973 = NOT(g23819)
--	g24982 = NOT(g23505)
--	g24993 = NOT(g23521)
--	g25087 = NOT(g23731)
--	g25094 = NOT(g23779)
--	g25095 = NOT(g23786)
--	I32829 = NOT(g24059)
--	g25103 = NOT(I32829)
--	g25104 = NOT(g23832)
--	g25105 = NOT(g23839)
--	I32835 = NOT(g24072)
--	g25109 = NOT(I32835)
--	g25110 = NOT(g23867)
--	g25111 = NOT(g23874)
--	g25115 = NOT(g23879)
--	g25116 = NOT(g23882)
--	I32844 = NOT(g23644)
--	g25118 = NOT(I32844)
--	I32847 = NOT(g24083)
--	g25119 = NOT(I32847)
--	g25120 = NOT(g23901)
--	I32851 = NOT(g23694)
--	g25121 = NOT(I32851)
--	I32854 = NOT(g24092)
--	g25122 = NOT(I32854)
--	I32857 = NOT(g23748)
--	g25123 = NOT(I32857)
--	I32860 = NOT(g23803)
--	g25124 = NOT(I32860)
--	g25126 = NOT(g24030)
--	I32868 = NOT(g25118)
--	g25130 = NOT(I32868)
--	I32871 = NOT(g24518)
--	g25131 = NOT(I32871)
--	I32874 = NOT(g24539)
--	g25132 = NOT(I32874)
--	I32877 = NOT(g24567)
--	g25133 = NOT(I32877)
--	I32880 = NOT(g24581)
--	g25134 = NOT(I32880)
--	I32883 = NOT(g24592)
--	g25135 = NOT(I32883)
--	I32886 = NOT(g24549)
--	g25136 = NOT(I32886)
--	I32889 = NOT(g24568)
--	g25137 = NOT(I32889)
--	I32892 = NOT(g24582)
--	g25138 = NOT(I32892)
--	I32895 = NOT(g24816)
--	g25139 = NOT(I32895)
--	I32898 = NOT(g24856)
--	g25140 = NOT(I32898)
--	I32901 = NOT(g25121)
--	g25141 = NOT(I32901)
--	I32904 = NOT(g24531)
--	g25142 = NOT(I32904)
--	I32907 = NOT(g24551)
--	g25143 = NOT(I32907)
--	I32910 = NOT(g24576)
--	g25144 = NOT(I32910)
--	I32913 = NOT(g24586)
--	g25145 = NOT(I32913)
--	I32916 = NOT(g24597)
--	g25146 = NOT(I32916)
--	I32919 = NOT(g24560)
--	g25147 = NOT(I32919)
--	I32922 = NOT(g24577)
--	g25148 = NOT(I32922)
--	I32925 = NOT(g24587)
--	g25149 = NOT(I32925)
--	I32928 = NOT(g24835)
--	g25150 = NOT(I32928)
--	I32931 = NOT(g24872)
--	g25151 = NOT(I32931)
--	I32934 = NOT(g25123)
--	g25152 = NOT(I32934)
--	I32937 = NOT(g24544)
--	g25153 = NOT(I32937)
--	I32940 = NOT(g24562)
--	g25154 = NOT(I32940)
--	I32943 = NOT(g24583)
--	g25155 = NOT(I32943)
--	I32946 = NOT(g24593)
--	g25156 = NOT(I32946)
--	I32949 = NOT(g24605)
--	g25157 = NOT(I32949)
--	I32952 = NOT(g24570)
--	g25158 = NOT(I32952)
--	I32955 = NOT(g24584)
--	g25159 = NOT(I32955)
--	I32958 = NOT(g24594)
--	g25160 = NOT(I32958)
--	I32961 = NOT(g24851)
--	g25161 = NOT(I32961)
--	I32964 = NOT(g24886)
--	g25162 = NOT(I32964)
--	I32967 = NOT(g25124)
--	g25163 = NOT(I32967)
--	I32970 = NOT(g24556)
--	g25164 = NOT(I32970)
--	I32973 = NOT(g24572)
--	g25165 = NOT(I32973)
--	I32976 = NOT(g24588)
--	g25166 = NOT(I32976)
--	I32979 = NOT(g24598)
--	g25167 = NOT(I32979)
--	I32982 = NOT(g24612)
--	g25168 = NOT(I32982)
--	I32985 = NOT(g24579)
--	g25169 = NOT(I32985)
--	I32988 = NOT(g24589)
--	g25170 = NOT(I32988)
--	I32991 = NOT(g24599)
--	g25171 = NOT(I32991)
--	I32994 = NOT(g24865)
--	g25172 = NOT(I32994)
--	I32997 = NOT(g24903)
--	g25173 = NOT(I32997)
--	I33000 = NOT(g24949)
--	g25174 = NOT(I33000)
--	I33003 = NOT(g24956)
--	g25175 = NOT(I33003)
--	I33006 = NOT(g24957)
--	g25176 = NOT(I33006)
--	I33009 = NOT(g24879)
--	g25177 = NOT(I33009)
--	I33013 = NOT(g25119)
--	g25179 = NOT(I33013)
--	I33016 = NOT(g25122)
--	g25180 = NOT(I33016)
--	g25274 = NOT(g24912)
--	g25283 = NOT(g24929)
--	g25291 = NOT(g24941)
--	I33128 = NOT(g24975)
--	g25296 = NOT(I33128)
--	g25301 = NOT(g24952)
--	g25305 = NOT(g24880)
--	I33136 = NOT(g24986)
--	g25306 = NOT(I33136)
--	g25313 = NOT(g24868)
--	g25314 = NOT(g24897)
--	I33145 = NOT(g24997)
--	g25315 = NOT(I33145)
--	g25319 = NOT(g24857)
--	g25322 = NOT(g24883)
--	g25323 = NOT(g24920)
--	I33154 = NOT(g25005)
--	g25324 = NOT(I33154)
--	I33157 = NOT(g25027)
--	g25327 = NOT(I33157)
--	g25329 = NOT(g24844)
--	g25330 = NOT(g24873)
--	g25332 = NOT(g24900)
--	g25333 = NOT(g24937)
--	g25335 = NOT(g24832)
--	I33168 = NOT(g25042)
--	g25336 = NOT(I33168)
--	g25338 = NOT(g24860)
--	g25339 = NOT(g24887)
--	g25341 = NOT(g24923)
--	g25347 = NOT(g24817)
--	g25349 = NOT(g24848)
--	I33182 = NOT(g25056)
--	g25350 = NOT(I33182)
--	g25352 = NOT(g24875)
--	g25353 = NOT(g24904)
--	I33188 = NOT(g24814)
--	g25354 = NOT(I33188)
--	g25355 = NOT(g24797)
--	g25361 = NOT(g24837)
--	g25363 = NOT(g24862)
--	I33198 = NOT(g25067)
--	g25364 = NOT(I33198)
--	g25366 = NOT(g24889)
--	g25367 = NOT(g24676)
--	g25368 = NOT(g24778)
--	I33205 = NOT(g24833)
--	g25369 = NOT(I33205)
--	g25370 = NOT(g24820)
--	g25376 = NOT(g24852)
--	g25378 = NOT(g24877)
--	g25379 = NOT(g24893)
--	g25383 = NOT(g24766)
--	g25384 = NOT(g24695)
--	g25385 = NOT(g24801)
--	I33219 = NOT(g24849)
--	g25386 = NOT(I33219)
--	g25387 = NOT(g24839)
--	g25393 = NOT(g24866)
--	g25394 = NOT(g24753)
--	g25395 = NOT(g24916)
--	g25399 = NOT(g24787)
--	g25400 = NOT(g24712)
--	g25401 = NOT(g24823)
--	I33232 = NOT(g24863)
--	g25402 = NOT(I33232)
--	g25403 = NOT(g24854)
--	g25404 = NOT(g24771)
--	g25405 = NOT(g24933)
--	g25409 = NOT(g24808)
--	g25410 = NOT(g24723)
--	g25411 = NOT(g24842)
--	g25412 = NOT(g24791)
--	g25413 = NOT(g24945)
--	g25417 = NOT(g24830)
--	g25419 = NOT(g24812)
--	I33246 = NOT(g24890)
--	g25420 = NOT(I33246)
--	I33249 = NOT(g24890)
--	g25421 = NOT(I33249)
--	g25422 = NOT(g24958)
--	g25430 = NOT(g24616)
--	g25431 = NOT(g24969)
--	I33257 = NOT(g24909)
--	g25435 = NOT(I33257)
--	I33260 = NOT(g24909)
--	g25436 = NOT(I33260)
--	g25437 = NOT(g24627)
--	g25438 = NOT(g24982)
--	I33265 = NOT(g24925)
--	g25442 = NOT(I33265)
--	I33268 = NOT(g24925)
--	g25443 = NOT(I33268)
--	g25444 = NOT(g24641)
--	g25445 = NOT(g24993)
--	g25449 = NOT(g24660)
--	I33278 = NOT(g25088)
--	g25454 = NOT(I33278)
--	I33282 = NOT(g25096)
--	g25458 = NOT(I33282)
--	I33286 = NOT(g24426)
--	g25462 = NOT(I33286)
--	I33289 = NOT(g25106)
--	g25463 = NOT(I33289)
--	I33293 = NOT(g25008)
--	g25467 = NOT(I33293)
--	I33297 = NOT(g24430)
--	g25471 = NOT(I33297)
--	I33300 = NOT(g25112)
--	g25472 = NOT(I33300)
--	I33304 = NOT(g25004)
--	g25476 = NOT(I33304)
--	I33307 = NOT(g25011)
--	g25479 = NOT(I33307)
--	I33312 = NOT(g25014)
--	g25484 = NOT(I33312)
--	I33316 = NOT(g24434)
--	g25488 = NOT(I33316)
--	I33321 = NOT(g24442)
--	g25493 = NOT(I33321)
--	I33324 = NOT(g25009)
--	g25496 = NOT(I33324)
--	I33327 = NOT(g25017)
--	g25499 = NOT(I33327)
--	I33330 = NOT(g25019)
--	g25502 = NOT(I33330)
--	I33335 = NOT(g25010)
--	g25507 = NOT(I33335)
--	I33338 = NOT(g25021)
--	g25510 = NOT(I33338)
--	I33343 = NOT(g25024)
--	g25515 = NOT(I33343)
--	I33347 = NOT(g24438)
--	g25519 = NOT(I33347)
--	I33352 = NOT(g24443)
--	g25524 = NOT(I33352)
--	I33355 = NOT(g25012)
--	g25527 = NOT(I33355)
--	I33358 = NOT(g25028)
--	g25530 = NOT(I33358)
--	I33361 = NOT(g25013)
--	g25533 = NOT(I33361)
--	I33364 = NOT(g25029)
--	g25536 = NOT(I33364)
--	I33368 = NOT(g24444)
--	g25540 = NOT(I33368)
--	I33371 = NOT(g25015)
--	g25543 = NOT(I33371)
--	I33374 = NOT(g25031)
--	g25546 = NOT(I33374)
--	I33377 = NOT(g25033)
--	g25549 = NOT(I33377)
--	I33382 = NOT(g25016)
--	g25554 = NOT(I33382)
--	I33385 = NOT(g25035)
--	g25557 = NOT(I33385)
--	I33390 = NOT(g25038)
--	g25562 = NOT(I33390)
--	I33396 = NOT(g24447)
--	g25573 = NOT(I33396)
--	I33399 = NOT(g25018)
--	g25576 = NOT(I33399)
--	I33402 = NOT(g24448)
--	g25579 = NOT(I33402)
--	I33405 = NOT(g25020)
--	g25582 = NOT(I33405)
--	I33408 = NOT(g25040)
--	g25585 = NOT(I33408)
--	I33411 = NOT(g24491)
--	g25588 = NOT(I33411)
--	I33415 = NOT(g24449)
--	g25590 = NOT(I33415)
--	I33418 = NOT(g25022)
--	g25593 = NOT(I33418)
--	I33421 = NOT(g25043)
--	g25596 = NOT(I33421)
--	I33424 = NOT(g25023)
--	g25599 = NOT(I33424)
--	I33427 = NOT(g25044)
--	g25602 = NOT(I33427)
--	I33431 = NOT(g24450)
--	g25606 = NOT(I33431)
--	I33434 = NOT(g25025)
--	g25609 = NOT(I33434)
--	I33437 = NOT(g25046)
--	g25612 = NOT(I33437)
--	I33440 = NOT(g25048)
--	g25615 = NOT(I33440)
--	I33445 = NOT(g25026)
--	g25620 = NOT(I33445)
--	I33448 = NOT(g25050)
--	g25623 = NOT(I33448)
--	g25630 = NOT(g24478)
--	I33457 = NOT(g24451)
--	g25634 = NOT(I33457)
--	I33460 = NOT(g24452)
--	g25637 = NOT(I33460)
--	I33463 = NOT(g25030)
--	g25640 = NOT(I33463)
--	I33466 = NOT(g25053)
--	g25643 = NOT(I33466)
--	I33469 = NOT(g24498)
--	g25646 = NOT(I33469)
--	I33472 = NOT(g24499)
--	g25647 = NOT(I33472)
--	I33476 = NOT(g24453)
--	g25652 = NOT(I33476)
--	I33479 = NOT(g25032)
--	g25655 = NOT(I33479)
--	I33482 = NOT(g24454)
--	g25658 = NOT(I33482)
--	I33485 = NOT(g25034)
--	g25661 = NOT(I33485)
--	I33488 = NOT(g25054)
--	g25664 = NOT(I33488)
--	I33491 = NOT(g24501)
--	g25667 = NOT(I33491)
--	I33495 = NOT(g24455)
--	g25669 = NOT(I33495)
--	I33498 = NOT(g25036)
--	g25672 = NOT(I33498)
--	I33501 = NOT(g25057)
--	g25675 = NOT(I33501)
--	I33504 = NOT(g25037)
--	g25678 = NOT(I33504)
--	I33507 = NOT(g25058)
--	g25681 = NOT(I33507)
--	I33511 = NOT(g24456)
--	g25685 = NOT(I33511)
--	I33514 = NOT(g25039)
--	g25688 = NOT(I33514)
--	I33517 = NOT(g25060)
--	g25691 = NOT(I33517)
--	I33520 = NOT(g25062)
--	g25694 = NOT(I33520)
--	g25698 = NOT(g24600)
--	I33526 = NOT(g24457)
--	g25700 = NOT(I33526)
--	I33529 = NOT(g25041)
--	g25703 = NOT(I33529)
--	I33532 = NOT(g24507)
--	g25706 = NOT(I33532)
--	I33535 = NOT(g24508)
--	g25707 = NOT(I33535)
--	I33539 = NOT(g24458)
--	g25711 = NOT(I33539)
--	I33542 = NOT(g24459)
--	g25714 = NOT(I33542)
--	I33545 = NOT(g25045)
--	g25717 = NOT(I33545)
--	I33548 = NOT(g25064)
--	g25720 = NOT(I33548)
--	I33551 = NOT(g24510)
--	g25723 = NOT(I33551)
--	I33554 = NOT(g24511)
--	g25724 = NOT(I33554)
--	I33558 = NOT(g24460)
--	g25729 = NOT(I33558)
--	I33561 = NOT(g25047)
--	g25732 = NOT(I33561)
--	I33564 = NOT(g24461)
--	g25735 = NOT(I33564)
--	I33567 = NOT(g25049)
--	g25738 = NOT(I33567)
--	I33570 = NOT(g25065)
--	g25741 = NOT(I33570)
--	I33573 = NOT(g24513)
--	g25744 = NOT(I33573)
--	I33577 = NOT(g24462)
--	g25746 = NOT(I33577)
--	I33580 = NOT(g25051)
--	g25749 = NOT(I33580)
--	I33583 = NOT(g25068)
--	g25752 = NOT(I33583)
--	I33586 = NOT(g25052)
--	g25755 = NOT(I33586)
--	I33589 = NOT(g25069)
--	g25758 = NOT(I33589)
--	I33593 = NOT(g24445)
--	g25762 = NOT(I33593)
--	I33596 = NOT(g24446)
--	g25763 = NOT(I33596)
--	I33600 = NOT(g24463)
--	g25767 = NOT(I33600)
--	I33603 = NOT(g24519)
--	g25770 = NOT(I33603)
--	g25771 = NOT(g24607)
--	I33608 = NOT(g24464)
--	g25773 = NOT(I33608)
--	I33611 = NOT(g25055)
--	g25776 = NOT(I33611)
--	I33614 = NOT(g24521)
--	g25779 = NOT(I33614)
--	I33617 = NOT(g24522)
--	g25780 = NOT(I33617)
--	I33621 = NOT(g24465)
--	g25784 = NOT(I33621)
--	I33624 = NOT(g24466)
--	g25787 = NOT(I33624)
--	I33627 = NOT(g25059)
--	g25790 = NOT(I33627)
--	I33630 = NOT(g25071)
--	g25793 = NOT(I33630)
--	I33633 = NOT(g24524)
--	g25796 = NOT(I33633)
--	I33636 = NOT(g24525)
--	g25797 = NOT(I33636)
--	I33640 = NOT(g24467)
--	g25802 = NOT(I33640)
--	I33643 = NOT(g25061)
--	g25805 = NOT(I33643)
--	I33646 = NOT(g24468)
--	g25808 = NOT(I33646)
--	I33649 = NOT(g25063)
--	g25811 = NOT(I33649)
--	I33652 = NOT(g25072)
--	g25814 = NOT(I33652)
--	I33655 = NOT(g24527)
--	g25817 = NOT(I33655)
--	I33659 = NOT(g24469)
--	g25821 = NOT(I33659)
--	I33662 = NOT(g24532)
--	g25824 = NOT(I33662)
--	g25825 = NOT(g24619)
--	I33667 = NOT(g24470)
--	g25827 = NOT(I33667)
--	I33670 = NOT(g25066)
--	g25830 = NOT(I33670)
--	I33673 = NOT(g24534)
--	g25833 = NOT(I33673)
--	I33676 = NOT(g24535)
--	g25834 = NOT(I33676)
--	I33680 = NOT(g24471)
--	g25838 = NOT(I33680)
--	I33683 = NOT(g24472)
--	g25841 = NOT(I33683)
--	I33686 = NOT(g25070)
--	g25844 = NOT(I33686)
--	I33689 = NOT(g25074)
--	g25847 = NOT(I33689)
--	I33692 = NOT(g24537)
--	g25850 = NOT(I33692)
--	I33695 = NOT(g24538)
--	g25851 = NOT(I33695)
--	I33700 = NOT(g24474)
--	g25856 = NOT(I33700)
--	I33703 = NOT(g24545)
--	g25859 = NOT(I33703)
--	g25860 = NOT(g24630)
--	I33708 = NOT(g24475)
--	g25862 = NOT(I33708)
--	I33711 = NOT(g25073)
--	g25865 = NOT(I33711)
--	I33714 = NOT(g24547)
--	g25868 = NOT(I33714)
--	I33717 = NOT(g24548)
--	g25869 = NOT(I33717)
--	I33723 = NOT(g24477)
--	g25877 = NOT(I33723)
--	I33726 = NOT(g24557)
--	g25880 = NOT(I33726)
--	I33732 = NOT(g24473)
--	g25886 = NOT(I33732)
--	I33737 = NOT(g24476)
--	g25891 = NOT(I33737)
--	g25895 = NOT(g24939)
--	g25899 = NOT(g24928)
--	g25903 = NOT(g24950)
--	g25907 = NOT(g24940)
--	g25911 = NOT(g24962)
--	g25915 = NOT(g24951)
--	g25919 = NOT(g24973)
--	g25923 = NOT(g24963)
--	g25937 = NOT(g24763)
--	g25939 = NOT(g24784)
--	g25942 = NOT(g24805)
--	g25945 = NOT(g24827)
--	g25952 = NOT(g24735)
--	I33790 = NOT(g25103)
--	g25976 = NOT(I33790)
--	I33798 = NOT(g25109)
--	g25982 = NOT(I33798)
--	I33801 = NOT(g25327)
--	g25983 = NOT(I33801)
--	I33804 = NOT(g25976)
--	g25984 = NOT(I33804)
--	I33807 = NOT(g25588)
--	g25985 = NOT(I33807)
--	I33810 = NOT(g25646)
--	g25986 = NOT(I33810)
--	I33813 = NOT(g25706)
--	g25987 = NOT(I33813)
--	I33816 = NOT(g25647)
--	g25988 = NOT(I33816)
--	I33819 = NOT(g25707)
--	g25989 = NOT(I33819)
--	I33822 = NOT(g25770)
--	g25990 = NOT(I33822)
--	I33825 = NOT(g25462)
--	g25991 = NOT(I33825)
--	I33828 = NOT(g25336)
--	g25992 = NOT(I33828)
--	I33831 = NOT(g25982)
--	g25993 = NOT(I33831)
--	I33834 = NOT(g25667)
--	g25994 = NOT(I33834)
--	I33837 = NOT(g25723)
--	g25995 = NOT(I33837)
--	I33840 = NOT(g25779)
--	g25996 = NOT(I33840)
--	I33843 = NOT(g25724)
--	g25997 = NOT(I33843)
--	I33846 = NOT(g25780)
--	g25998 = NOT(I33846)
--	I33849 = NOT(g25824)
--	g25999 = NOT(I33849)
--	I33852 = NOT(g25471)
--	g26000 = NOT(I33852)
--	I33855 = NOT(g25350)
--	g26001 = NOT(I33855)
--	I33858 = NOT(g25179)
--	g26002 = NOT(I33858)
--	I33861 = NOT(g25744)
--	g26003 = NOT(I33861)
--	I33864 = NOT(g25796)
--	g26004 = NOT(I33864)
--	I33867 = NOT(g25833)
--	g26005 = NOT(I33867)
--	I33870 = NOT(g25797)
--	g26006 = NOT(I33870)
--	I33873 = NOT(g25834)
--	g26007 = NOT(I33873)
--	I33876 = NOT(g25859)
--	g26008 = NOT(I33876)
--	I33879 = NOT(g25488)
--	g26009 = NOT(I33879)
--	I33882 = NOT(g25364)
--	g26010 = NOT(I33882)
--	I33885 = NOT(g25180)
--	g26011 = NOT(I33885)
--	I33888 = NOT(g25817)
--	g26012 = NOT(I33888)
--	I33891 = NOT(g25850)
--	g26013 = NOT(I33891)
--	I33894 = NOT(g25868)
--	g26014 = NOT(I33894)
--	I33897 = NOT(g25851)
--	g26015 = NOT(I33897)
--	I33900 = NOT(g25869)
--	g26016 = NOT(I33900)
--	I33903 = NOT(g25880)
--	g26017 = NOT(I33903)
--	I33906 = NOT(g25519)
--	g26018 = NOT(I33906)
--	I33909 = NOT(g25886)
--	g26019 = NOT(I33909)
--	I33912 = NOT(g25891)
--	g26020 = NOT(I33912)
--	I33915 = NOT(g25762)
--	g26021 = NOT(I33915)
--	I33918 = NOT(g25763)
--	g26022 = NOT(I33918)
--	I33954 = NOT(g25343)
--	g26056 = NOT(I33954)
--	I33961 = NOT(g25357)
--	g26063 = NOT(I33961)
--	I33968 = NOT(g25372)
--	g26070 = NOT(I33968)
--	I33974 = NOT(g25389)
--	g26076 = NOT(I33974)
--	I33984 = NOT(g25932)
--	g26086 = NOT(I33984)
--	I33990 = NOT(g25870)
--	g26092 = NOT(I33990)
--	I33995 = NOT(g25935)
--	g26102 = NOT(I33995)
--	I33999 = NOT(g25490)
--	g26104 = NOT(I33999)
--	I34002 = NOT(g25490)
--	g26105 = NOT(I34002)
--	I34009 = NOT(g25882)
--	g26114 = NOT(I34009)
--	I34012 = NOT(g25938)
--	g26118 = NOT(I34012)
--	I34017 = NOT(g25887)
--	g26121 = NOT(I34017)
--	I34020 = NOT(g25940)
--	g26125 = NOT(I34020)
--	I34026 = NOT(g25892)
--	g26131 = NOT(I34026)
--	I34029 = NOT(g25520)
--	g26135 = NOT(I34029)
--	I34032 = NOT(g25520)
--	g26136 = NOT(I34032)
--	I34041 = NOT(g25566)
--	g26149 = NOT(I34041)
--	I34044 = NOT(g25566)
--	g26150 = NOT(I34044)
--	I34051 = NOT(g25204)
--	g26159 = NOT(I34051)
--	I34056 = NOT(g25206)
--	g26164 = NOT(I34056)
--	I34059 = NOT(g25207)
--	g26165 = NOT(I34059)
--	I34063 = NOT(g25209)
--	g26167 = NOT(I34063)
--	I34068 = NOT(g25211)
--	g26172 = NOT(I34068)
--	I34071 = NOT(g25212)
--	g26173 = NOT(I34071)
--	I34074 = NOT(g25213)
--	g26174 = NOT(I34074)
--	I34077 = NOT(g25954)
--	g26175 = NOT(I34077)
--	I34080 = NOT(g25539)
--	g26178 = NOT(I34080)
--	I34083 = NOT(g25214)
--	g26181 = NOT(I34083)
--	I34086 = NOT(g25215)
--	g26182 = NOT(I34086)
--	I34091 = NOT(g25217)
--	g26187 = NOT(I34091)
--	g26189 = NOT(g25952)
--	I34096 = NOT(g25218)
--	g26190 = NOT(I34096)
--	I34099 = NOT(g25219)
--	g26191 = NOT(I34099)
--	I34102 = NOT(g25220)
--	g26192 = NOT(I34102)
--	I34105 = NOT(g25221)
--	g26193 = NOT(I34105)
--	I34108 = NOT(g25222)
--	g26194 = NOT(I34108)
--	I34111 = NOT(g25223)
--	g26195 = NOT(I34111)
--	I34114 = NOT(g25958)
--	g26196 = NOT(I34114)
--	I34118 = NOT(g25605)
--	g26202 = NOT(I34118)
--	I34121 = NOT(g25224)
--	g26205 = NOT(I34121)
--	I34124 = NOT(g25225)
--	g26206 = NOT(I34124)
--	I34128 = NOT(g25227)
--	g26208 = NOT(I34128)
--	g26209 = NOT(g25296)
--	I34132 = NOT(g25228)
--	g26210 = NOT(I34132)
--	I34135 = NOT(g25229)
--	g26211 = NOT(I34135)
--	I34140 = NOT(g25230)
--	g26214 = NOT(I34140)
--	I34143 = NOT(g25231)
--	g26215 = NOT(I34143)
--	I34146 = NOT(g25232)
--	g26216 = NOT(I34146)
--	I34150 = NOT(g25233)
--	g26220 = NOT(I34150)
--	I34153 = NOT(g25234)
--	g26221 = NOT(I34153)
--	I34156 = NOT(g25235)
--	g26222 = NOT(I34156)
--	I34159 = NOT(g25964)
--	g26223 = NOT(I34159)
--	I34162 = NOT(g25684)
--	g26226 = NOT(I34162)
--	I34165 = NOT(g25236)
--	g26229 = NOT(I34165)
--	I34168 = NOT(g25237)
--	g26230 = NOT(I34168)
--	I34172 = NOT(g25239)
--	g26232 = NOT(I34172)
--	g26237 = NOT(g25306)
--	I34180 = NOT(g25240)
--	g26238 = NOT(I34180)
--	I34183 = NOT(g25241)
--	g26239 = NOT(I34183)
--	I34189 = NOT(g25242)
--	g26245 = NOT(I34189)
--	I34192 = NOT(g25243)
--	g26246 = NOT(I34192)
--	I34195 = NOT(g25244)
--	g26247 = NOT(I34195)
--	I34198 = NOT(g25245)
--	g26248 = NOT(I34198)
--	I34201 = NOT(g25246)
--	g26249 = NOT(I34201)
--	I34204 = NOT(g25247)
--	g26250 = NOT(I34204)
--	I34207 = NOT(g25969)
--	g26251 = NOT(I34207)
--	I34210 = NOT(g25761)
--	g26254 = NOT(I34210)
--	I34220 = NOT(g25248)
--	g26264 = NOT(I34220)
--	g26275 = NOT(g25315)
--	I34230 = NOT(g25249)
--	g26276 = NOT(I34230)
--	I34233 = NOT(g25250)
--	g26277 = NOT(I34233)
--	I34238 = NOT(g25251)
--	g26280 = NOT(I34238)
--	I34241 = NOT(g25252)
--	g26281 = NOT(I34241)
--	I34244 = NOT(g25253)
--	g26282 = NOT(I34244)
--	I34254 = NOT(g25185)
--	g26294 = NOT(I34254)
--	I34266 = NOT(g25255)
--	g26308 = NOT(I34266)
--	g26313 = NOT(g25324)
--	I34274 = NOT(g25256)
--	g26314 = NOT(I34274)
--	I34277 = NOT(g25257)
--	g26315 = NOT(I34277)
--	I34296 = NOT(g25189)
--	g26341 = NOT(I34296)
--	I34306 = NOT(g25259)
--	g26349 = NOT(I34306)
--	I34313 = NOT(g25265)
--	g26354 = NOT(I34313)
--	I34316 = NOT(g25191)
--	g26355 = NOT(I34316)
--	I34321 = NOT(g25928)
--	g26358 = NOT(I34321)
--	I34327 = NOT(g25260)
--	g26364 = NOT(I34327)
--	I34343 = NOT(g25194)
--	g26385 = NOT(I34343)
--	I34353 = NOT(g25927)
--	g26393 = NOT(I34353)
--	I34358 = NOT(g25262)
--	g26398 = NOT(I34358)
--	I34363 = NOT(g25930)
--	g26401 = NOT(I34363)
--	I34369 = NOT(g25263)
--	g26407 = NOT(I34369)
--	I34385 = NOT(g25197)
--	g26428 = NOT(I34385)
--	I34388 = NOT(g25200)
--	g26429 = NOT(I34388)
--	I34392 = NOT(g25266)
--	g26433 = NOT(I34392)
--	I34395 = NOT(g25929)
--	g26434 = NOT(I34395)
--	I34400 = NOT(g25267)
--	g26439 = NOT(I34400)
--	I34405 = NOT(g25933)
--	g26442 = NOT(I34405)
--	I34411 = NOT(g25268)
--	g26448 = NOT(I34411)
--	I34421 = NOT(g25203)
--	g26461 = NOT(I34421)
--	I34425 = NOT(g25270)
--	g26465 = NOT(I34425)
--	I34428 = NOT(g25931)
--	g26466 = NOT(I34428)
--	I34433 = NOT(g25271)
--	g26471 = NOT(I34433)
--	I34438 = NOT(g25936)
--	g26474 = NOT(I34438)
--	I34444 = NOT(g25272)
--	g26480 = NOT(I34444)
--	g26481 = NOT(g25764)
--	I34449 = NOT(g25205)
--	g26485 = NOT(I34449)
--	I34453 = NOT(g25279)
--	g26489 = NOT(I34453)
--	I34456 = NOT(g25934)
--	g26490 = NOT(I34456)
--	I34461 = NOT(g25280)
--	g26495 = NOT(I34461)
--	I34464 = NOT(g25199)
--	g26496 = NOT(I34464)
--	g26497 = NOT(g25818)
--	I34469 = NOT(g25210)
--	g26501 = NOT(I34469)
--	I34473 = NOT(g25288)
--	g26505 = NOT(I34473)
--	I34476 = NOT(g25201)
--	g26506 = NOT(I34476)
--	I34479 = NOT(g25202)
--	g26507 = NOT(I34479)
--	g26508 = NOT(g25312)
--	g26512 = NOT(g25853)
--	g26516 = NOT(g25320)
--	g26520 = NOT(g25874)
--	g26521 = NOT(g25331)
--	g26525 = NOT(g25340)
--	g26533 = NOT(g25454)
--	g26538 = NOT(g25458)
--	g26539 = NOT(g25463)
--	g26540 = NOT(g25467)
--	g26542 = NOT(g25472)
--	g26543 = NOT(g25476)
--	g26544 = NOT(g25479)
--	g26546 = NOT(g25484)
--	I34505 = NOT(g25450)
--	g26548 = NOT(I34505)
--	g26549 = NOT(g25421)
--	g26550 = NOT(g25493)
--	g26551 = NOT(g25496)
--	g26552 = NOT(g25499)
--	g26554 = NOT(g25502)
--	g26555 = NOT(g25507)
--	g26556 = NOT(g25510)
--	g26558 = NOT(g25515)
--	g26561 = NOT(g25524)
--	g26562 = NOT(g25527)
--	g26563 = NOT(g25530)
--	g26564 = NOT(g25533)
--	g26565 = NOT(g25536)
--	g26566 = NOT(g25540)
--	g26567 = NOT(g25543)
--	g26568 = NOT(g25546)
--	g26570 = NOT(g25549)
--	g26571 = NOT(g25554)
--	g26572 = NOT(g25557)
--	g26574 = NOT(g25562)
--	I34535 = NOT(g25451)
--	g26576 = NOT(I34535)
--	g26577 = NOT(g25436)
--	g26578 = NOT(g25573)
--	g26579 = NOT(g25576)
--	g26580 = NOT(g25579)
--	g26581 = NOT(g25582)
--	g26582 = NOT(g25585)
--	g26584 = NOT(g25590)
--	g26585 = NOT(g25593)
--	g26586 = NOT(g25596)
--	g26587 = NOT(g25599)
--	g26588 = NOT(g25602)
--	g26589 = NOT(g25606)
--	g26590 = NOT(g25609)
--	g26591 = NOT(g25612)
--	g26593 = NOT(g25615)
--	g26594 = NOT(g25620)
--	g26595 = NOT(g25623)
--	g26597 = NOT(g25443)
--	g26598 = NOT(g25634)
--	g26599 = NOT(g25637)
--	g26600 = NOT(g25640)
--	g26601 = NOT(g25643)
--	g26602 = NOT(g25652)
--	g26603 = NOT(g25655)
--	g26604 = NOT(g25658)
--	g26605 = NOT(g25661)
--	g26606 = NOT(g25664)
--	g26608 = NOT(g25669)
--	g26609 = NOT(g25672)
--	g26610 = NOT(g25675)
--	g26611 = NOT(g25678)
--	g26612 = NOT(g25681)
--	g26613 = NOT(g25685)
--	g26614 = NOT(g25688)
--	g26615 = NOT(g25691)
--	g26617 = NOT(g25694)
--	I34579 = NOT(g25452)
--	g26618 = NOT(I34579)
--	g26619 = NOT(g25700)
--	g26620 = NOT(g25703)
--	g26621 = NOT(g25711)
--	g26622 = NOT(g25714)
--	g26623 = NOT(g25717)
--	g26624 = NOT(g25720)
--	g26625 = NOT(g25729)
--	g26626 = NOT(g25732)
--	g26627 = NOT(g25735)
--	g26628 = NOT(g25738)
--	g26629 = NOT(g25741)
--	g26631 = NOT(g25746)
--	g26632 = NOT(g25749)
--	g26633 = NOT(g25752)
--	g26634 = NOT(g25755)
--	g26635 = NOT(g25758)
--	g26636 = NOT(g25767)
--	g26637 = NOT(g25773)
--	g26638 = NOT(g25776)
--	g26639 = NOT(g25784)
--	g26640 = NOT(g25787)
--	g26641 = NOT(g25790)
--	g26642 = NOT(g25793)
--	g26643 = NOT(g25802)
--	g26644 = NOT(g25805)
--	g26645 = NOT(g25808)
--	g26646 = NOT(g25811)
--	g26647 = NOT(g25814)
--	g26648 = NOT(g25821)
--	g26649 = NOT(g25827)
--	g26650 = NOT(g25830)
--	g26651 = NOT(g25838)
--	g26652 = NOT(g25841)
--	g26653 = NOT(g25844)
--	g26654 = NOT(g25847)
--	g26656 = NOT(g25856)
--	g26657 = NOT(g25862)
--	g26658 = NOT(g25865)
--	g26662 = NOT(g25877)
--	I34641 = NOT(g26086)
--	g26678 = NOT(I34641)
--	I34644 = NOT(g26159)
--	g26679 = NOT(I34644)
--	I34647 = NOT(g26164)
--	g26680 = NOT(I34647)
--	I34650 = NOT(g26172)
--	g26681 = NOT(I34650)
--	I34653 = NOT(g26165)
--	g26682 = NOT(I34653)
--	I34656 = NOT(g26173)
--	g26683 = NOT(I34656)
--	I34659 = NOT(g26190)
--	g26684 = NOT(I34659)
--	I34662 = NOT(g26174)
--	g26685 = NOT(I34662)
--	I34665 = NOT(g26191)
--	g26686 = NOT(I34665)
--	I34668 = NOT(g26210)
--	g26687 = NOT(I34668)
--	I34671 = NOT(g26192)
--	g26688 = NOT(I34671)
--	I34674 = NOT(g26211)
--	g26689 = NOT(I34674)
--	I34677 = NOT(g26232)
--	g26690 = NOT(I34677)
--	I34680 = NOT(g26294)
--	g26691 = NOT(I34680)
--	I34683 = NOT(g26364)
--	g26692 = NOT(I34683)
--	I34686 = NOT(g26398)
--	g26693 = NOT(I34686)
--	I34689 = NOT(g26433)
--	g26694 = NOT(I34689)
--	I34692 = NOT(g26102)
--	g26695 = NOT(I34692)
--	I34695 = NOT(g26167)
--	g26696 = NOT(I34695)
--	I34698 = NOT(g26181)
--	g26697 = NOT(I34698)
--	I34701 = NOT(g26193)
--	g26698 = NOT(I34701)
--	I34704 = NOT(g26182)
--	g26699 = NOT(I34704)
--	I34707 = NOT(g26194)
--	g26700 = NOT(I34707)
--	I34710 = NOT(g26214)
--	g26701 = NOT(I34710)
--	I34713 = NOT(g26195)
--	g26702 = NOT(I34713)
--	I34716 = NOT(g26215)
--	g26703 = NOT(I34716)
--	I34719 = NOT(g26238)
--	g26704 = NOT(I34719)
--	I34722 = NOT(g26216)
--	g26705 = NOT(I34722)
--	I34725 = NOT(g26239)
--	g26706 = NOT(I34725)
--	I34728 = NOT(g26264)
--	g26707 = NOT(I34728)
--	I34731 = NOT(g26341)
--	g26708 = NOT(I34731)
--	I34734 = NOT(g26407)
--	g26709 = NOT(I34734)
--	I34737 = NOT(g26439)
--	g26710 = NOT(I34737)
--	I34740 = NOT(g26465)
--	g26711 = NOT(I34740)
--	I34743 = NOT(g26118)
--	g26712 = NOT(I34743)
--	I34746 = NOT(g26187)
--	g26713 = NOT(I34746)
--	I34749 = NOT(g26205)
--	g26714 = NOT(I34749)
--	I34752 = NOT(g26220)
--	g26715 = NOT(I34752)
--	I34755 = NOT(g26206)
--	g26716 = NOT(I34755)
--	I34758 = NOT(g26221)
--	g26717 = NOT(I34758)
--	I34761 = NOT(g26245)
--	g26718 = NOT(I34761)
--	I34764 = NOT(g26222)
--	g26719 = NOT(I34764)
--	I34767 = NOT(g26246)
--	g26720 = NOT(I34767)
--	I34770 = NOT(g26276)
--	g26721 = NOT(I34770)
--	I34773 = NOT(g26247)
--	g26722 = NOT(I34773)
--	I34776 = NOT(g26277)
--	g26723 = NOT(I34776)
--	I34779 = NOT(g26308)
--	g26724 = NOT(I34779)
--	I34782 = NOT(g26385)
--	g26725 = NOT(I34782)
--	I34785 = NOT(g26448)
--	g26726 = NOT(I34785)
--	I34788 = NOT(g26471)
--	g26727 = NOT(I34788)
--	I34791 = NOT(g26489)
--	g26728 = NOT(I34791)
--	I34794 = NOT(g26125)
--	g26729 = NOT(I34794)
--	I34797 = NOT(g26208)
--	g26730 = NOT(I34797)
--	I34800 = NOT(g26229)
--	g26731 = NOT(I34800)
--	I34803 = NOT(g26248)
--	g26732 = NOT(I34803)
--	I34806 = NOT(g26230)
--	g26733 = NOT(I34806)
--	I34809 = NOT(g26249)
--	g26734 = NOT(I34809)
--	I34812 = NOT(g26280)
--	g26735 = NOT(I34812)
--	I34815 = NOT(g26250)
--	g26736 = NOT(I34815)
--	I34818 = NOT(g26281)
--	g26737 = NOT(I34818)
--	I34821 = NOT(g26314)
--	g26738 = NOT(I34821)
--	I34824 = NOT(g26282)
--	g26739 = NOT(I34824)
--	I34827 = NOT(g26315)
--	g26740 = NOT(I34827)
--	I34830 = NOT(g26349)
--	g26741 = NOT(I34830)
--	I34833 = NOT(g26428)
--	g26742 = NOT(I34833)
--	I34836 = NOT(g26480)
--	g26743 = NOT(I34836)
--	I34839 = NOT(g26495)
--	g26744 = NOT(I34839)
--	I34842 = NOT(g26505)
--	g26745 = NOT(I34842)
--	I34845 = NOT(g26496)
--	g26746 = NOT(I34845)
--	I34848 = NOT(g26506)
--	g26747 = NOT(I34848)
--	I34851 = NOT(g26354)
--	g26748 = NOT(I34851)
--	I34854 = NOT(g26507)
--	g26749 = NOT(I34854)
--	I34857 = NOT(g26355)
--	g26750 = NOT(I34857)
--	I34860 = NOT(g26548)
--	g26751 = NOT(I34860)
--	I34863 = NOT(g26576)
--	g26752 = NOT(I34863)
--	I34866 = NOT(g26618)
--	g26753 = NOT(I34866)
--	I34872 = NOT(g26217)
--	g26757 = NOT(I34872)
--	I34879 = NOT(g26240)
--	g26762 = NOT(I34879)
--	I34901 = NOT(g26295)
--	g26782 = NOT(I34901)
--	I34909 = NOT(g26265)
--	g26788 = NOT(I34909)
--	I34916 = NOT(g26240)
--	g26793 = NOT(I34916)
--	I34921 = NOT(g26217)
--	g26796 = NOT(I34921)
--	I34946 = NOT(g26534)
--	g26819 = NOT(I34946)
--	I34957 = NOT(g26541)
--	g26828 = NOT(I34957)
--	I34961 = NOT(g26545)
--	g26830 = NOT(I34961)
--	I34964 = NOT(g26547)
--	g26831 = NOT(I34964)
--	I34967 = NOT(g26553)
--	g26832 = NOT(I34967)
--	I34971 = NOT(g26557)
--	g26834 = NOT(I34971)
--	I34974 = NOT(g26168)
--	g26835 = NOT(I34974)
--	I34977 = NOT(g26559)
--	g26836 = NOT(I34977)
--	I34980 = NOT(g26458)
--	g26837 = NOT(I34980)
--	I34983 = NOT(g26569)
--	g26840 = NOT(I34983)
--	I34986 = NOT(g26160)
--	g26841 = NOT(I34986)
--	I34990 = NOT(g26573)
--	g26843 = NOT(I34990)
--	I34993 = NOT(g26575)
--	g26844 = NOT(I34993)
--	I34997 = NOT(g26482)
--	g26846 = NOT(I34997)
--	I35000 = NOT(g26336)
--	g26849 = NOT(I35000)
--	I35003 = NOT(g26592)
--	g26850 = NOT(I35003)
--	I35007 = NOT(g26596)
--	g26852 = NOT(I35007)
--	I35011 = NOT(g26304)
--	g26854 = NOT(I35011)
--	I35014 = NOT(g26498)
--	g26855 = NOT(I35014)
--	I35017 = NOT(g26616)
--	g26858 = NOT(I35017)
--	I35028 = NOT(g26513)
--	g26861 = NOT(I35028)
--	I35031 = NOT(g26529)
--	g26864 = NOT(I35031)
--	I35049 = NOT(g26530)
--	g26868 = NOT(I35049)
--	I35053 = NOT(g26655)
--	g26872 = NOT(I35053)
--	I35064 = NOT(g26531)
--	g26875 = NOT(I35064)
--	I35067 = NOT(g26659)
--	g26876 = NOT(I35067)
--	I35072 = NOT(g26661)
--	g26881 = NOT(I35072)
--	I35076 = NOT(g26532)
--	g26883 = NOT(I35076)
--	I35079 = NOT(g26664)
--	g26884 = NOT(I35079)
--	I35083 = NOT(g26665)
--	g26886 = NOT(I35083)
--	I35087 = NOT(g26667)
--	g26890 = NOT(I35087)
--	I35092 = NOT(g26669)
--	g26895 = NOT(I35092)
--	I35095 = NOT(g26670)
--	g26896 = NOT(I35095)
--	I35099 = NOT(g26672)
--	g26900 = NOT(I35099)
--	I35106 = NOT(g26675)
--	g26909 = NOT(I35106)
--	I35109 = NOT(g26676)
--	g26910 = NOT(I35109)
--	I35116 = NOT(g26025)
--	g26921 = NOT(I35116)
--	g26922 = NOT(g26283)
--	g26935 = NOT(g26327)
--	g26944 = NOT(g26374)
--	g26950 = NOT(g26417)
--	I35136 = NOT(g26660)
--	g26953 = NOT(I35136)
--	g26954 = NOT(g26549)
--	I35141 = NOT(g26666)
--	g26956 = NOT(I35141)
--	g26957 = NOT(g26577)
--	I35146 = NOT(g26671)
--	g26959 = NOT(I35146)
--	g26960 = NOT(g26597)
--	I35153 = NOT(g26677)
--	g26964 = NOT(I35153)
--	I35172 = NOT(g26272)
--	g26983 = NOT(I35172)
--	g26987 = NOT(g26056)
--	g27010 = NOT(g26063)
--	g27036 = NOT(g26070)
--	g27064 = NOT(g26076)
--	I35254 = NOT(g26048)
--	g27075 = NOT(I35254)
--	I35283 = NOT(g26031)
--	g27102 = NOT(I35283)
--	I35297 = NOT(g26199)
--	g27114 = NOT(I35297)
--	I35301 = NOT(g26037)
--	g27116 = NOT(I35301)
--	I35313 = NOT(g26534)
--	g27126 = NOT(I35313)
--	I35319 = NOT(g26183)
--	g27132 = NOT(I35319)
--	g27133 = NOT(g26105)
--	g27134 = NOT(g26175)
--	g27135 = NOT(g26178)
--	g27136 = NOT(g26196)
--	g27137 = NOT(g26202)
--	g27138 = NOT(g26223)
--	g27139 = NOT(g26226)
--	g27140 = NOT(g26136)
--	g27141 = NOT(g26251)
--	g27142 = NOT(g26254)
--	g27143 = NOT(g26150)
--	I35334 = NOT(g26106)
--	g27145 = NOT(I35334)
--	g27146 = NOT(g26358)
--	g27148 = NOT(g26393)
--	I35341 = NOT(g26120)
--	g27150 = NOT(I35341)
--	g27151 = NOT(g26401)
--	g27153 = NOT(g26429)
--	I35347 = NOT(g26265)
--	g27154 = NOT(I35347)
--	g27155 = NOT(g26434)
--	I35351 = NOT(g26272)
--	g27156 = NOT(I35351)
--	I35355 = NOT(g26130)
--	g27158 = NOT(I35355)
--	g27159 = NOT(g26442)
--	I35360 = NOT(g26295)
--	g27161 = NOT(I35360)
--	g27162 = NOT(g26461)
--	I35364 = NOT(g26304)
--	g27163 = NOT(I35364)
--	g27164 = NOT(g26466)
--	I35369 = NOT(g26144)
--	g27166 = NOT(I35369)
--	g27167 = NOT(g26474)
--	I35373 = NOT(g26189)
--	g27168 = NOT(I35373)
--	I35376 = NOT(g26336)
--	g27171 = NOT(I35376)
--	g27172 = NOT(g26485)
--	g27173 = NOT(g26490)
--	I35383 = NOT(g26160)
--	g27176 = NOT(I35383)
--	g27177 = NOT(g26501)
--	I35389 = NOT(g26168)
--	g27180 = NOT(I35389)
--	I35394 = NOT(g26183)
--	g27183 = NOT(I35394)
--	I35399 = NOT(g26199)
--	g27186 = NOT(I35399)
--	I35404 = NOT(g26864)
--	g27189 = NOT(I35404)
--	I35407 = NOT(g27145)
--	g27190 = NOT(I35407)
--	I35410 = NOT(g26872)
--	g27191 = NOT(I35410)
--	I35413 = NOT(g26876)
--	g27192 = NOT(I35413)
--	I35416 = NOT(g26884)
--	g27193 = NOT(I35416)
--	I35419 = NOT(g26828)
--	g27194 = NOT(I35419)
--	I35422 = NOT(g26830)
--	g27195 = NOT(I35422)
--	I35425 = NOT(g26832)
--	g27196 = NOT(I35425)
--	I35428 = NOT(g26953)
--	g27197 = NOT(I35428)
--	I35431 = NOT(g26868)
--	g27198 = NOT(I35431)
--	I35434 = NOT(g27150)
--	g27199 = NOT(I35434)
--	I35437 = NOT(g27183)
--	g27200 = NOT(I35437)
--	I35440 = NOT(g27186)
--	g27201 = NOT(I35440)
--	I35443 = NOT(g26757)
--	g27202 = NOT(I35443)
--	I35446 = NOT(g26762)
--	g27203 = NOT(I35446)
--	I35449 = NOT(g27154)
--	g27204 = NOT(I35449)
--	I35452 = NOT(g27161)
--	g27205 = NOT(I35452)
--	I35455 = NOT(g26881)
--	g27206 = NOT(I35455)
--	I35458 = NOT(g26886)
--	g27207 = NOT(I35458)
--	I35461 = NOT(g26895)
--	g27208 = NOT(I35461)
--	I35464 = NOT(g26831)
--	g27209 = NOT(I35464)
--	I35467 = NOT(g26834)
--	g27210 = NOT(I35467)
--	I35470 = NOT(g26840)
--	g27211 = NOT(I35470)
--	I35473 = NOT(g27156)
--	g27212 = NOT(I35473)
--	I35476 = NOT(g27163)
--	g27213 = NOT(I35476)
--	I35479 = NOT(g27171)
--	g27214 = NOT(I35479)
--	I35482 = NOT(g27176)
--	g27215 = NOT(I35482)
--	I35485 = NOT(g27180)
--	g27216 = NOT(I35485)
--	I35488 = NOT(g26819)
--	g27217 = NOT(I35488)
--	I35491 = NOT(g26956)
--	g27218 = NOT(I35491)
--	I35494 = NOT(g26875)
--	g27219 = NOT(I35494)
--	I35497 = NOT(g27158)
--	g27220 = NOT(I35497)
--	I35500 = NOT(g26890)
--	g27221 = NOT(I35500)
--	I35503 = NOT(g26896)
--	g27222 = NOT(I35503)
--	I35506 = NOT(g26909)
--	g27223 = NOT(I35506)
--	I35509 = NOT(g26836)
--	g27224 = NOT(I35509)
--	I35512 = NOT(g26843)
--	g27225 = NOT(I35512)
--	I35515 = NOT(g26850)
--	g27226 = NOT(I35515)
--	I35518 = NOT(g26959)
--	g27227 = NOT(I35518)
--	I35521 = NOT(g26883)
--	g27228 = NOT(I35521)
--	I35524 = NOT(g27166)
--	g27229 = NOT(I35524)
--	I35527 = NOT(g26900)
--	g27230 = NOT(I35527)
--	I35530 = NOT(g26910)
--	g27231 = NOT(I35530)
--	I35533 = NOT(g26921)
--	g27232 = NOT(I35533)
--	I35536 = NOT(g26844)
--	g27233 = NOT(I35536)
--	I35539 = NOT(g26852)
--	g27234 = NOT(I35539)
--	I35542 = NOT(g26858)
--	g27235 = NOT(I35542)
--	I35545 = NOT(g26964)
--	g27236 = NOT(I35545)
--	I35548 = NOT(g27116)
--	g27237 = NOT(I35548)
--	I35551 = NOT(g27075)
--	g27238 = NOT(I35551)
--	I35554 = NOT(g27102)
--	g27239 = NOT(I35554)
--	g27349 = NOT(g27126)
--	I35667 = NOT(g27120)
--	g27353 = NOT(I35667)
--	I35673 = NOT(g27123)
--	g27357 = NOT(I35673)
--	I35678 = NOT(g27129)
--	g27360 = NOT(I35678)
--	I35681 = NOT(g26869)
--	g27361 = NOT(I35681)
--	I35686 = NOT(g27131)
--	g27366 = NOT(I35686)
--	I35689 = NOT(g26878)
--	g27367 = NOT(I35689)
--	I35695 = NOT(g26887)
--	g27373 = NOT(I35695)
--	I35698 = NOT(g26897)
--	g27376 = NOT(I35698)
--	I35708 = NOT(g26974)
--	g27380 = NOT(I35708)
--	I35711 = NOT(g26974)
--	g27381 = NOT(I35711)
--	g27383 = NOT(g27133)
--	g27384 = NOT(g27140)
--	I35723 = NOT(g27168)
--	g27385 = NOT(I35723)
--	g27386 = NOT(g27143)
--	I35727 = NOT(g26902)
--	g27387 = NOT(I35727)
--	I35731 = NOT(g26892)
--	g27391 = NOT(I35731)
--	I35737 = NOT(g26915)
--	g27397 = NOT(I35737)
--	I35741 = NOT(g27118)
--	g27401 = NOT(I35741)
--	I35744 = NOT(g26906)
--	g27404 = NOT(I35744)
--	I35750 = NOT(g26928)
--	g27410 = NOT(I35750)
--	I35756 = NOT(g27117)
--	g27416 = NOT(I35756)
--	I35759 = NOT(g27121)
--	g27419 = NOT(I35759)
--	I35762 = NOT(g26918)
--	g27422 = NOT(I35762)
--	I35768 = NOT(g26941)
--	g27428 = NOT(I35768)
--	I35772 = NOT(g26772)
--	g27432 = NOT(I35772)
--	I35777 = NOT(g27119)
--	g27437 = NOT(I35777)
--	I35780 = NOT(g27124)
--	g27440 = NOT(I35780)
--	I35783 = NOT(g26931)
--	g27443 = NOT(I35783)
--	g27449 = NOT(g26837)
--	I35791 = NOT(g26779)
--	g27451 = NOT(I35791)
--	I35796 = NOT(g27122)
--	g27456 = NOT(I35796)
--	I35799 = NOT(g27130)
--	g27459 = NOT(I35799)
--	I35803 = NOT(g26803)
--	g27463 = NOT(I35803)
--	g27465 = NOT(g26846)
--	I35809 = NOT(g26785)
--	g27467 = NOT(I35809)
--	I35814 = NOT(g27125)
--	g27472 = NOT(I35814)
--	I35817 = NOT(g26922)
--	g27475 = NOT(I35817)
--	I35821 = NOT(g26804)
--	g27479 = NOT(I35821)
--	I35824 = NOT(g26805)
--	g27480 = NOT(I35824)
--	I35829 = NOT(g26806)
--	g27483 = NOT(I35829)
--	g27484 = NOT(g26855)
--	I35834 = NOT(g26792)
--	g27486 = NOT(I35834)
--	I35837 = NOT(g26911)
--	g27489 = NOT(I35837)
--	I35841 = NOT(g26807)
--	g27493 = NOT(I35841)
--	I35844 = NOT(g26808)
--	g27494 = NOT(I35844)
--	I35849 = NOT(g26776)
--	g27497 = NOT(I35849)
--	I35852 = NOT(g26935)
--	g27498 = NOT(I35852)
--	I35856 = NOT(g26809)
--	g27502 = NOT(I35856)
--	I35859 = NOT(g26810)
--	g27503 = NOT(I35859)
--	I35863 = NOT(g26811)
--	g27505 = NOT(I35863)
--	g27506 = NOT(g26861)
--	I35868 = NOT(g26812)
--	g27508 = NOT(I35868)
--	I35872 = NOT(g26925)
--	g27510 = NOT(I35872)
--	I35876 = NOT(g26813)
--	g27514 = NOT(I35876)
--	I35879 = NOT(g26814)
--	g27515 = NOT(I35879)
--	I35883 = NOT(g26781)
--	g27517 = NOT(I35883)
--	I35886 = NOT(g26944)
--	g27518 = NOT(I35886)
--	I35890 = NOT(g26815)
--	g27522 = NOT(I35890)
--	I35893 = NOT(g26816)
--	g27523 = NOT(I35893)
--	I35897 = NOT(g26817)
--	g27525 = NOT(I35897)
--	I35900 = NOT(g26786)
--	g27526 = NOT(I35900)
--	I35915 = NOT(g26818)
--	g27533 = NOT(I35915)
--	I35919 = NOT(g26938)
--	g27535 = NOT(I35919)
--	I35923 = NOT(g26820)
--	g27539 = NOT(I35923)
--	I35926 = NOT(g26821)
--	g27540 = NOT(I35926)
--	I35930 = NOT(g26789)
--	g27542 = NOT(I35930)
--	I35933 = NOT(g26950)
--	g27543 = NOT(I35933)
--	I35937 = NOT(g26822)
--	g27547 = NOT(I35937)
--	I35940 = NOT(g26823)
--	g27548 = NOT(I35940)
--	I35953 = NOT(g26824)
--	g27553 = NOT(I35953)
--	I35957 = NOT(g26947)
--	g27555 = NOT(I35957)
--	I35961 = NOT(g26825)
--	g27559 = NOT(I35961)
--	I35964 = NOT(g26826)
--	g27560 = NOT(I35964)
--	I35968 = NOT(g26795)
--	g27562 = NOT(I35968)
--	I35983 = NOT(g26827)
--	g27569 = NOT(I35983)
--	I36008 = NOT(g26798)
--	g27586 = NOT(I36008)
--	g27589 = NOT(g27168)
--	g27590 = NOT(g27144)
--	g27595 = NOT(g27149)
--	g27599 = NOT(g27147)
--	g27604 = NOT(g27157)
--	g27608 = NOT(g27152)
--	g27613 = NOT(g27165)
--	g27617 = NOT(g27160)
--	g27622 = NOT(g27174)
--	I36032 = NOT(g27113)
--	g27632 = NOT(I36032)
--	I36042 = NOT(g26960)
--	g27662 = NOT(I36042)
--	I36046 = NOT(g26957)
--	g27667 = NOT(I36046)
--	I36052 = NOT(g26954)
--	g27674 = NOT(I36052)
--	I36060 = NOT(g27353)
--	g27683 = NOT(I36060)
--	I36063 = NOT(g27463)
--	g27684 = NOT(I36063)
--	I36066 = NOT(g27479)
--	g27685 = NOT(I36066)
--	I36069 = NOT(g27493)
--	g27686 = NOT(I36069)
--	I36072 = NOT(g27480)
--	g27687 = NOT(I36072)
--	I36075 = NOT(g27494)
--	g27688 = NOT(I36075)
--	I36078 = NOT(g27508)
--	g27689 = NOT(I36078)
--	I36081 = NOT(g27497)
--	g27690 = NOT(I36081)
--	I36084 = NOT(g27357)
--	g27691 = NOT(I36084)
--	I36087 = NOT(g27483)
--	g27692 = NOT(I36087)
--	I36090 = NOT(g27502)
--	g27693 = NOT(I36090)
--	I36093 = NOT(g27514)
--	g27694 = NOT(I36093)
--	I36096 = NOT(g27503)
--	g27695 = NOT(I36096)
--	I36099 = NOT(g27515)
--	g27696 = NOT(I36099)
--	I36102 = NOT(g27533)
--	g27697 = NOT(I36102)
--	I36105 = NOT(g27517)
--	g27698 = NOT(I36105)
--	I36108 = NOT(g27360)
--	g27699 = NOT(I36108)
--	I36111 = NOT(g27505)
--	g27700 = NOT(I36111)
--	I36114 = NOT(g27522)
--	g27701 = NOT(I36114)
--	I36117 = NOT(g27539)
--	g27702 = NOT(I36117)
--	I36120 = NOT(g27523)
--	g27703 = NOT(I36120)
--	I36123 = NOT(g27540)
--	g27704 = NOT(I36123)
--	I36126 = NOT(g27553)
--	g27705 = NOT(I36126)
--	I36129 = NOT(g27542)
--	g27706 = NOT(I36129)
--	I36132 = NOT(g27366)
--	g27707 = NOT(I36132)
--	I36135 = NOT(g27525)
--	g27708 = NOT(I36135)
--	I36138 = NOT(g27547)
--	g27709 = NOT(I36138)
--	I36141 = NOT(g27559)
--	g27710 = NOT(I36141)
--	I36144 = NOT(g27548)
--	g27711 = NOT(I36144)
--	I36147 = NOT(g27560)
--	g27712 = NOT(I36147)
--	I36150 = NOT(g27569)
--	g27713 = NOT(I36150)
--	I36153 = NOT(g27562)
--	g27714 = NOT(I36153)
--	I36156 = NOT(g27586)
--	g27715 = NOT(I36156)
--	I36159 = NOT(g27526)
--	g27716 = NOT(I36159)
--	I36162 = NOT(g27385)
--	g27717 = NOT(I36162)
--	g27748 = NOT(g27632)
--	I36213 = NOT(g27571)
--	g27776 = NOT(I36213)
--	I36217 = NOT(g27580)
--	g27780 = NOT(I36217)
--	I36221 = NOT(g27662)
--	g27784 = NOT(I36221)
--	I36224 = NOT(g27589)
--	g27785 = NOT(I36224)
--	I36227 = NOT(g27594)
--	g27786 = NOT(I36227)
--	I36230 = NOT(g27583)
--	g27787 = NOT(I36230)
--	I36234 = NOT(g27667)
--	g27791 = NOT(I36234)
--	I36237 = NOT(g27662)
--	g27792 = NOT(I36237)
--	I36240 = NOT(g27603)
--	g27793 = NOT(I36240)
--	I36243 = NOT(g27587)
--	g27794 = NOT(I36243)
--	I36246 = NOT(g27674)
--	g27797 = NOT(I36246)
--	I36250 = NOT(g27612)
--	g27799 = NOT(I36250)
--	I36253 = NOT(g27674)
--	g27800 = NOT(I36253)
--	I36264 = NOT(g27621)
--	g27805 = NOT(I36264)
--	I36267 = NOT(g27395)
--	g27806 = NOT(I36267)
--	I36280 = NOT(g27390)
--	g27817 = NOT(I36280)
--	I36283 = NOT(g27408)
--	g27820 = NOT(I36283)
--	I36296 = NOT(g27626)
--	g27831 = NOT(I36296)
--	I36307 = NOT(g27400)
--	g27839 = NOT(I36307)
--	I36311 = NOT(g27426)
--	g27843 = NOT(I36311)
--	I36321 = NOT(g27627)
--	g27847 = NOT(I36321)
--	I36327 = NOT(g27413)
--	g27858 = NOT(I36327)
--	I36330 = NOT(g27447)
--	g27861 = NOT(I36330)
--	I36337 = NOT(g27628)
--	g27872 = NOT(I36337)
--	I36341 = NOT(g27431)
--	g27879 = NOT(I36341)
--	I36347 = NOT(g27630)
--	g27889 = NOT(I36347)
--	I36354 = NOT(g27662)
--	g27903 = NOT(I36354)
--	I36358 = NOT(g27672)
--	g27905 = NOT(I36358)
--	I36362 = NOT(g27667)
--	g27907 = NOT(I36362)
--	I36367 = NOT(g27678)
--	g27910 = NOT(I36367)
--	I36371 = NOT(g27674)
--	g27912 = NOT(I36371)
--	I36379 = NOT(g27682)
--	g27918 = NOT(I36379)
--	I36382 = NOT(g27563)
--	g27919 = NOT(I36382)
--	I36390 = NOT(g27243)
--	g27927 = NOT(I36390)
--	I36393 = NOT(g27572)
--	g27928 = NOT(I36393)
--	I36397 = NOT(g27574)
--	g27932 = NOT(I36397)
--	I36404 = NOT(g27450)
--	g27939 = NOT(I36404)
--	I36407 = NOT(g27581)
--	g27942 = NOT(I36407)
--	I36411 = NOT(g27582)
--	g27946 = NOT(I36411)
--	I36417 = NOT(g27462)
--	g27952 = NOT(I36417)
--	I36420 = NOT(g27253)
--	g27955 = NOT(I36420)
--	I36423 = NOT(g27466)
--	g27956 = NOT(I36423)
--	I36426 = NOT(g27584)
--	g27959 = NOT(I36426)
--	I36432 = NOT(g27585)
--	g27965 = NOT(I36432)
--	g27969 = NOT(g27361)
--	I36438 = NOT(g27255)
--	g27971 = NOT(I36438)
--	I36441 = NOT(g27256)
--	g27972 = NOT(I36441)
--	I36444 = NOT(g27482)
--	g27973 = NOT(I36444)
--	I36447 = NOT(g27257)
--	g27976 = NOT(I36447)
--	I36450 = NOT(g27485)
--	g27977 = NOT(I36450)
--	I36454 = NOT(g27588)
--	g27981 = NOT(I36454)
--	I36459 = NOT(g27258)
--	g27986 = NOT(I36459)
--	I36462 = NOT(g27259)
--	g27987 = NOT(I36462)
--	I36465 = NOT(g27260)
--	g27988 = NOT(I36465)
--	I36468 = NOT(g27261)
--	g27989 = NOT(I36468)
--	g27990 = NOT(g27367)
--	I36473 = NOT(g27262)
--	g27992 = NOT(I36473)
--	I36476 = NOT(g27263)
--	g27993 = NOT(I36476)
--	I36479 = NOT(g27504)
--	g27994 = NOT(I36479)
--	I36483 = NOT(g27264)
--	g27998 = NOT(I36483)
--	I36486 = NOT(g27507)
--	g27999 = NOT(I36486)
--	I36490 = NOT(g27265)
--	g28003 = NOT(I36490)
--	I36493 = NOT(g27266)
--	g28004 = NOT(I36493)
--	I36496 = NOT(g27267)
--	g28005 = NOT(I36496)
--	I36499 = NOT(g27268)
--	g28006 = NOT(I36499)
--	I36502 = NOT(g27269)
--	g28007 = NOT(I36502)
--	I36507 = NOT(g27270)
--	g28010 = NOT(I36507)
--	I36510 = NOT(g27271)
--	g28011 = NOT(I36510)
--	I36513 = NOT(g27272)
--	g28012 = NOT(I36513)
--	I36516 = NOT(g27273)
--	g28013 = NOT(I36516)
--	g28014 = NOT(g27373)
--	I36521 = NOT(g27274)
--	g28016 = NOT(I36521)
--	I36524 = NOT(g27275)
--	g28017 = NOT(I36524)
--	I36527 = NOT(g27524)
--	g28018 = NOT(I36527)
--	I36530 = NOT(g27276)
--	g28021 = NOT(I36530)
--	I36533 = NOT(g27277)
--	g28022 = NOT(I36533)
--	I36536 = NOT(g27278)
--	g28023 = NOT(I36536)
--	I36539 = NOT(g27279)
--	g28024 = NOT(I36539)
--	I36542 = NOT(g27280)
--	g28025 = NOT(I36542)
--	I36545 = NOT(g27281)
--	g28026 = NOT(I36545)
--	I36551 = NOT(g27282)
--	g28030 = NOT(I36551)
--	I36554 = NOT(g27283)
--	g28031 = NOT(I36554)
--	I36557 = NOT(g27284)
--	g28032 = NOT(I36557)
--	I36560 = NOT(g27285)
--	g28033 = NOT(I36560)
--	I36563 = NOT(g27286)
--	g28034 = NOT(I36563)
--	I36568 = NOT(g27287)
--	g28037 = NOT(I36568)
--	I36571 = NOT(g27288)
--	g28038 = NOT(I36571)
--	I36574 = NOT(g27289)
--	g28039 = NOT(I36574)
--	I36577 = NOT(g27290)
--	g28040 = NOT(I36577)
--	g28041 = NOT(g27376)
--	I36582 = NOT(g27291)
--	g28043 = NOT(I36582)
--	I36585 = NOT(g27292)
--	g28044 = NOT(I36585)
--	I36588 = NOT(g27293)
--	g28045 = NOT(I36588)
--	I36598 = NOT(g27294)
--	g28047 = NOT(I36598)
--	I36601 = NOT(g27295)
--	g28048 = NOT(I36601)
--	I36604 = NOT(g27296)
--	g28049 = NOT(I36604)
--	I36609 = NOT(g27297)
--	g28052 = NOT(I36609)
--	I36612 = NOT(g27298)
--	g28053 = NOT(I36612)
--	I36615 = NOT(g27299)
--	g28054 = NOT(I36615)
--	I36618 = NOT(g27300)
--	g28055 = NOT(I36618)
--	I36621 = NOT(g27301)
--	g28056 = NOT(I36621)
--	I36627 = NOT(g27302)
--	g28060 = NOT(I36627)
--	I36630 = NOT(g27303)
--	g28061 = NOT(I36630)
--	I36633 = NOT(g27304)
--	g28062 = NOT(I36633)
--	I36636 = NOT(g27305)
--	g28063 = NOT(I36636)
--	I36639 = NOT(g27306)
--	g28064 = NOT(I36639)
--	I36644 = NOT(g27307)
--	g28067 = NOT(I36644)
--	I36647 = NOT(g27308)
--	g28068 = NOT(I36647)
--	I36650 = NOT(g27309)
--	g28069 = NOT(I36650)
--	I36653 = NOT(g27310)
--	g28070 = NOT(I36653)
--	I36656 = NOT(g27311)
--	g28071 = NOT(I36656)
--	I36659 = NOT(g27312)
--	g28072 = NOT(I36659)
--	I36663 = NOT(g27313)
--	g28074 = NOT(I36663)
--	I36673 = NOT(g27314)
--	g28076 = NOT(I36673)
--	I36676 = NOT(g27315)
--	g28077 = NOT(I36676)
--	I36679 = NOT(g27316)
--	g28078 = NOT(I36679)
--	I36684 = NOT(g27317)
--	g28081 = NOT(I36684)
--	I36687 = NOT(g27318)
--	g28082 = NOT(I36687)
--	I36690 = NOT(g27319)
--	g28083 = NOT(I36690)
--	I36693 = NOT(g27320)
--	g28084 = NOT(I36693)
--	I36696 = NOT(g27321)
--	g28085 = NOT(I36696)
--	I36702 = NOT(g27322)
--	g28089 = NOT(I36702)
--	I36705 = NOT(g27323)
--	g28090 = NOT(I36705)
--	I36708 = NOT(g27324)
--	g28091 = NOT(I36708)
--	I36711 = NOT(g27325)
--	g28092 = NOT(I36711)
--	I36714 = NOT(g27326)
--	g28093 = NOT(I36714)
--	I36718 = NOT(g27327)
--	g28095 = NOT(I36718)
--	I36721 = NOT(g27328)
--	g28096 = NOT(I36721)
--	I36724 = NOT(g27329)
--	g28097 = NOT(I36724)
--	I36728 = NOT(g27330)
--	g28099 = NOT(I36728)
--	I36738 = NOT(g27331)
--	g28101 = NOT(I36738)
--	I36741 = NOT(g27332)
--	g28102 = NOT(I36741)
--	I36744 = NOT(g27333)
--	g28103 = NOT(I36744)
--	I36749 = NOT(g27334)
--	g28106 = NOT(I36749)
--	I36752 = NOT(g27335)
--	g28107 = NOT(I36752)
--	I36755 = NOT(g27336)
--	g28108 = NOT(I36755)
--	I36758 = NOT(g27337)
--	g28109 = NOT(I36758)
--	I36761 = NOT(g27338)
--	g28110 = NOT(I36761)
--	I36766 = NOT(g27339)
--	g28113 = NOT(I36766)
--	I36769 = NOT(g27340)
--	g28114 = NOT(I36769)
--	I36772 = NOT(g27341)
--	g28115 = NOT(I36772)
--	I36776 = NOT(g27342)
--	g28117 = NOT(I36776)
--	I36786 = NOT(g27343)
--	g28119 = NOT(I36786)
--	I36789 = NOT(g27344)
--	g28120 = NOT(I36789)
--	I36792 = NOT(g27345)
--	g28121 = NOT(I36792)
--	I36797 = NOT(g27346)
--	g28124 = NOT(I36797)
--	I36800 = NOT(g27347)
--	g28125 = NOT(I36800)
--	I36803 = NOT(g27348)
--	g28126 = NOT(I36803)
--	g28128 = NOT(g27528)
--	I36808 = NOT(g27354)
--	g28132 = NOT(I36808)
--	g28133 = NOT(g27550)
--	g28137 = NOT(g27566)
--	g28141 = NOT(g27576)
--	g28149 = NOT(g27667)
--	g28150 = NOT(g27387)
--	g28151 = NOT(g27381)
--	g28152 = NOT(g27391)
--	g28153 = NOT(g27397)
--	g28154 = NOT(g27401)
--	g28155 = NOT(g27404)
--	g28156 = NOT(g27410)
--	g28158 = NOT(g27416)
--	g28159 = NOT(g27419)
--	g28160 = NOT(g27422)
--	g28161 = NOT(g27428)
--	g28162 = NOT(g27432)
--	g28163 = NOT(g27437)
--	g28164 = NOT(g27440)
--	g28165 = NOT(g27443)
--	g28166 = NOT(g27451)
--	g28167 = NOT(g27456)
--	g28168 = NOT(g27459)
--	g28169 = NOT(g27467)
--	g28170 = NOT(g27472)
--	g28172 = NOT(g27475)
--	g28173 = NOT(g27486)
--	g28174 = NOT(g27489)
--	g28175 = NOT(g27498)
--	g28177 = NOT(g27510)
--	g28178 = NOT(g27518)
--	I36848 = NOT(g27383)
--	g28179 = NOT(I36848)
--	g28186 = NOT(g27535)
--	g28187 = NOT(g27543)
--	g28190 = NOT(g27555)
--	I36860 = NOT(g27386)
--	g28194 = NOT(I36860)
--	I36864 = NOT(g27384)
--	g28200 = NOT(I36864)
--	I36867 = NOT(g27786)
--	g28206 = NOT(I36867)
--	I36870 = NOT(g27955)
--	g28207 = NOT(I36870)
--	I36873 = NOT(g27971)
--	g28208 = NOT(I36873)
--	I36876 = NOT(g27986)
--	g28209 = NOT(I36876)
--	I36879 = NOT(g27972)
--	g28210 = NOT(I36879)
--	I36882 = NOT(g27987)
--	g28211 = NOT(I36882)
--	I36885 = NOT(g28003)
--	g28212 = NOT(I36885)
--	I36888 = NOT(g27988)
--	g28213 = NOT(I36888)
--	I36891 = NOT(g28004)
--	g28214 = NOT(I36891)
--	I36894 = NOT(g28022)
--	g28215 = NOT(I36894)
--	I36897 = NOT(g28005)
--	g28216 = NOT(I36897)
--	I36900 = NOT(g28023)
--	g28217 = NOT(I36900)
--	I36903 = NOT(g28045)
--	g28218 = NOT(I36903)
--	I36906 = NOT(g27989)
--	g28219 = NOT(I36906)
--	I36909 = NOT(g28006)
--	g28220 = NOT(I36909)
--	I36912 = NOT(g28024)
--	g28221 = NOT(I36912)
--	I36915 = NOT(g28007)
--	g28222 = NOT(I36915)
--	I36918 = NOT(g28025)
--	g28223 = NOT(I36918)
--	I36921 = NOT(g28047)
--	g28224 = NOT(I36921)
--	I36924 = NOT(g28026)
--	g28225 = NOT(I36924)
--	I36927 = NOT(g28048)
--	g28226 = NOT(I36927)
--	I36930 = NOT(g28071)
--	g28227 = NOT(I36930)
--	I36933 = NOT(g28049)
--	g28228 = NOT(I36933)
--	I36936 = NOT(g28072)
--	g28229 = NOT(I36936)
--	I36939 = NOT(g28095)
--	g28230 = NOT(I36939)
--	I36942 = NOT(g27905)
--	g28231 = NOT(I36942)
--	I36945 = NOT(g27793)
--	g28232 = NOT(I36945)
--	I36948 = NOT(g27976)
--	g28233 = NOT(I36948)
--	I36951 = NOT(g27992)
--	g28234 = NOT(I36951)
--	I36954 = NOT(g28010)
--	g28235 = NOT(I36954)
--	I36957 = NOT(g27993)
--	g28236 = NOT(I36957)
--	I36960 = NOT(g28011)
--	g28237 = NOT(I36960)
--	I36963 = NOT(g28030)
--	g28238 = NOT(I36963)
--	I36966 = NOT(g28012)
--	g28239 = NOT(I36966)
--	I36969 = NOT(g28031)
--	g28240 = NOT(I36969)
--	I36972 = NOT(g28052)
--	g28241 = NOT(I36972)
--	I36975 = NOT(g28032)
--	g28242 = NOT(I36975)
--	I36978 = NOT(g28053)
--	g28243 = NOT(I36978)
--	I36981 = NOT(g28074)
--	g28244 = NOT(I36981)
--	I36984 = NOT(g28013)
--	g28245 = NOT(I36984)
--	I36987 = NOT(g28033)
--	g28246 = NOT(I36987)
--	I36990 = NOT(g28054)
--	g28247 = NOT(I36990)
--	I36993 = NOT(g28034)
--	g28248 = NOT(I36993)
--	I36996 = NOT(g28055)
--	g28249 = NOT(I36996)
--	I36999 = NOT(g28076)
--	g28250 = NOT(I36999)
--	I37002 = NOT(g28056)
--	g28251 = NOT(I37002)
--	I37005 = NOT(g28077)
--	g28252 = NOT(I37005)
--	I37008 = NOT(g28096)
--	g28253 = NOT(I37008)
--	I37011 = NOT(g28078)
--	g28254 = NOT(I37011)
--	I37014 = NOT(g28097)
--	g28255 = NOT(I37014)
--	I37017 = NOT(g28113)
--	g28256 = NOT(I37017)
--	I37020 = NOT(g27910)
--	g28257 = NOT(I37020)
--	I37023 = NOT(g27799)
--	g28258 = NOT(I37023)
--	I37026 = NOT(g27998)
--	g28259 = NOT(I37026)
--	I37029 = NOT(g28016)
--	g28260 = NOT(I37029)
--	I37032 = NOT(g28037)
--	g28261 = NOT(I37032)
--	I37035 = NOT(g28017)
--	g28262 = NOT(I37035)
--	I37038 = NOT(g28038)
--	g28263 = NOT(I37038)
--	I37041 = NOT(g28060)
--	g28264 = NOT(I37041)
--	I37044 = NOT(g28039)
--	g28265 = NOT(I37044)
--	I37047 = NOT(g28061)
--	g28266 = NOT(I37047)
--	I37050 = NOT(g28081)
--	g28267 = NOT(I37050)
--	I37053 = NOT(g28062)
--	g28268 = NOT(I37053)
--	I37056 = NOT(g28082)
--	g28269 = NOT(I37056)
--	I37059 = NOT(g28099)
--	g28270 = NOT(I37059)
--	I37062 = NOT(g28040)
--	g28271 = NOT(I37062)
--	I37065 = NOT(g28063)
--	g28272 = NOT(I37065)
--	I37068 = NOT(g28083)
--	g28273 = NOT(I37068)
--	I37071 = NOT(g28064)
--	g28274 = NOT(I37071)
--	I37074 = NOT(g28084)
--	g28275 = NOT(I37074)
--	I37077 = NOT(g28101)
--	g28276 = NOT(I37077)
--	I37080 = NOT(g28085)
--	g28277 = NOT(I37080)
--	I37083 = NOT(g28102)
--	g28278 = NOT(I37083)
--	I37086 = NOT(g28114)
--	g28279 = NOT(I37086)
--	I37089 = NOT(g28103)
--	g28280 = NOT(I37089)
--	I37092 = NOT(g28115)
--	g28281 = NOT(I37092)
--	I37095 = NOT(g28124)
--	g28282 = NOT(I37095)
--	I37098 = NOT(g27918)
--	g28283 = NOT(I37098)
--	I37101 = NOT(g27805)
--	g28284 = NOT(I37101)
--	I37104 = NOT(g28021)
--	g28285 = NOT(I37104)
--	I37107 = NOT(g28043)
--	g28286 = NOT(I37107)
--	I37110 = NOT(g28067)
--	g28287 = NOT(I37110)
--	I37113 = NOT(g28044)
--	g28288 = NOT(I37113)
--	I37116 = NOT(g28068)
--	g28289 = NOT(I37116)
--	I37119 = NOT(g28089)
--	g28290 = NOT(I37119)
--	I37122 = NOT(g28069)
--	g28291 = NOT(I37122)
--	I37125 = NOT(g28090)
--	g28292 = NOT(I37125)
--	I37128 = NOT(g28106)
--	g28293 = NOT(I37128)
--	I37131 = NOT(g28091)
--	g28294 = NOT(I37131)
--	I37134 = NOT(g28107)
--	g28295 = NOT(I37134)
--	I37137 = NOT(g28117)
--	g28296 = NOT(I37137)
--	I37140 = NOT(g28070)
--	g28297 = NOT(I37140)
--	I37143 = NOT(g28092)
--	g28298 = NOT(I37143)
--	I37146 = NOT(g28108)
--	g28299 = NOT(I37146)
--	I37149 = NOT(g28093)
--	g28300 = NOT(I37149)
--	I37152 = NOT(g28109)
--	g28301 = NOT(I37152)
--	I37155 = NOT(g28119)
--	g28302 = NOT(I37155)
--	I37158 = NOT(g28110)
--	g28303 = NOT(I37158)
--	I37161 = NOT(g28120)
--	g28304 = NOT(I37161)
--	I37164 = NOT(g28125)
--	g28305 = NOT(I37164)
--	I37167 = NOT(g28121)
--	g28306 = NOT(I37167)
--	I37170 = NOT(g28126)
--	g28307 = NOT(I37170)
--	I37173 = NOT(g28132)
--	g28308 = NOT(I37173)
--	I37176 = NOT(g27927)
--	g28309 = NOT(I37176)
--	I37179 = NOT(g27784)
--	g28310 = NOT(I37179)
--	I37182 = NOT(g27791)
--	g28311 = NOT(I37182)
--	I37185 = NOT(g27797)
--	g28312 = NOT(I37185)
--	I37188 = NOT(g27785)
--	g28313 = NOT(I37188)
--	I37191 = NOT(g27792)
--	g28314 = NOT(I37191)
--	I37194 = NOT(g27800)
--	g28315 = NOT(I37194)
--	I37197 = NOT(g27903)
--	g28316 = NOT(I37197)
--	I37200 = NOT(g27907)
--	g28317 = NOT(I37200)
--	I37203 = NOT(g27912)
--	g28318 = NOT(I37203)
--	I37228 = NOT(g28194)
--	g28341 = NOT(I37228)
--	I37232 = NOT(g28200)
--	g28343 = NOT(I37232)
--	I37238 = NOT(g28179)
--	g28347 = NOT(I37238)
--	I37252 = NOT(g28200)
--	g28359 = NOT(I37252)
--	I37260 = NOT(g28179)
--	g28365 = NOT(I37260)
--	I37266 = NOT(g28200)
--	g28369 = NOT(I37266)
--	I37269 = NOT(g28145)
--	g28370 = NOT(I37269)
--	I37273 = NOT(g28179)
--	g28372 = NOT(I37273)
--	I37277 = NOT(g28146)
--	g28374 = NOT(I37277)
--	I37280 = NOT(g28179)
--	g28375 = NOT(I37280)
--	I37284 = NOT(g28147)
--	g28377 = NOT(I37284)
--	I37291 = NOT(g28148)
--	g28382 = NOT(I37291)
--	I37319 = NOT(g28149)
--	g28390 = NOT(I37319)
--	I37330 = NOT(g28194)
--	g28393 = NOT(I37330)
--	I37334 = NOT(g28194)
--	g28395 = NOT(I37334)
--	g28419 = NOT(g28151)
--	I37379 = NOT(g28199)
--	g28432 = NOT(I37379)
--	I37386 = NOT(g28194)
--	g28437 = NOT(I37386)
--	I37394 = NOT(g27718)
--	g28443 = NOT(I37394)
--	I37400 = NOT(g28200)
--	g28447 = NOT(I37400)
--	I37410 = NOT(g27722)
--	g28455 = NOT(I37410)
--	I37415 = NOT(g28179)
--	g28458 = NOT(I37415)
--	I37426 = NOT(g27724)
--	g28467 = NOT(I37426)
--	g28483 = NOT(g27776)
--	g28491 = NOT(g27780)
--	g28496 = NOT(g27787)
--	I37459 = NOT(g27759)
--	g28498 = NOT(I37459)
--	g28500 = NOT(g27794)
--	I37467 = NOT(g27760)
--	g28524 = NOT(I37467)
--	I37471 = NOT(g27761)
--	g28526 = NOT(I37471)
--	I37474 = NOT(g27762)
--	g28527 = NOT(I37474)
--	I37481 = NOT(g27763)
--	g28552 = NOT(I37481)
--	I37484 = NOT(g27764)
--	g28553 = NOT(I37484)
--	g28554 = NOT(g27806)
--	I37488 = NOT(g27765)
--	g28555 = NOT(I37488)
--	I37494 = NOT(g27766)
--	g28579 = NOT(I37494)
--	I37497 = NOT(g27767)
--	g28580 = NOT(I37497)
--	g28581 = NOT(g27817)
--	g28582 = NOT(g27820)
--	I37502 = NOT(g27768)
--	g28583 = NOT(I37502)
--	I37508 = NOT(g27769)
--	g28607 = NOT(I37508)
--	g28608 = NOT(g27831)
--	g28609 = NOT(g27839)
--	g28610 = NOT(g27843)
--	I37514 = NOT(g27771)
--	g28611 = NOT(I37514)
--	g28612 = NOT(g28046)
--	g28616 = NOT(g27847)
--	g28617 = NOT(g27858)
--	g28618 = NOT(g27861)
--	g28619 = NOT(g28075)
--	g28623 = NOT(g27872)
--	g28624 = NOT(g27879)
--	g28625 = NOT(g28100)
--	g28629 = NOT(g27889)
--	g28630 = NOT(g28118)
--	g28638 = NOT(g28200)
--	g28639 = NOT(g27919)
--	g28640 = NOT(g27928)
--	g28641 = NOT(g27932)
--	g28642 = NOT(g27939)
--	g28643 = NOT(g27942)
--	g28644 = NOT(g27946)
--	g28645 = NOT(g27952)
--	g28646 = NOT(g27956)
--	g28647 = NOT(g27959)
--	g28648 = NOT(g27965)
--	g28649 = NOT(g27973)
--	g28650 = NOT(g27977)
--	g28651 = NOT(g27981)
--	g28652 = NOT(g27994)
--	g28653 = NOT(g27999)
--	g28655 = NOT(g28018)
--	I37566 = NOT(g28370)
--	g28673 = NOT(I37566)
--	I37569 = NOT(g28498)
--	g28674 = NOT(I37569)
--	I37572 = NOT(g28524)
--	g28675 = NOT(I37572)
--	I37575 = NOT(g28527)
--	g28676 = NOT(I37575)
--	I37578 = NOT(g28432)
--	g28677 = NOT(I37578)
--	I37581 = NOT(g28374)
--	g28678 = NOT(I37581)
--	I37584 = NOT(g28526)
--	g28679 = NOT(I37584)
--	I37587 = NOT(g28552)
--	g28680 = NOT(I37587)
--	I37590 = NOT(g28555)
--	g28681 = NOT(I37590)
--	I37593 = NOT(g28443)
--	g28682 = NOT(I37593)
--	I37596 = NOT(g28377)
--	g28683 = NOT(I37596)
--	I37599 = NOT(g28553)
--	g28684 = NOT(I37599)
--	I37602 = NOT(g28579)
--	g28685 = NOT(I37602)
--	I37605 = NOT(g28583)
--	g28686 = NOT(I37605)
--	I37608 = NOT(g28455)
--	g28687 = NOT(I37608)
--	I37611 = NOT(g28382)
--	g28688 = NOT(I37611)
--	I37614 = NOT(g28580)
--	g28689 = NOT(I37614)
--	I37617 = NOT(g28607)
--	g28690 = NOT(I37617)
--	I37620 = NOT(g28611)
--	g28691 = NOT(I37620)
--	I37623 = NOT(g28467)
--	g28692 = NOT(I37623)
--	I37626 = NOT(g28393)
--	g28693 = NOT(I37626)
--	I37629 = NOT(g28369)
--	g28694 = NOT(I37629)
--	I37632 = NOT(g28372)
--	g28695 = NOT(I37632)
--	I37635 = NOT(g28390)
--	g28696 = NOT(I37635)
--	I37638 = NOT(g28395)
--	g28697 = NOT(I37638)
--	I37641 = NOT(g28375)
--	g28698 = NOT(I37641)
--	I37644 = NOT(g28341)
--	g28699 = NOT(I37644)
--	I37647 = NOT(g28343)
--	g28700 = NOT(I37647)
--	I37650 = NOT(g28347)
--	g28701 = NOT(I37650)
--	I37653 = NOT(g28359)
--	g28702 = NOT(I37653)
--	I37656 = NOT(g28365)
--	g28703 = NOT(I37656)
--	I37659 = NOT(g28437)
--	g28704 = NOT(I37659)
--	I37662 = NOT(g28447)
--	g28705 = NOT(I37662)
--	I37665 = NOT(g28458)
--	g28706 = NOT(I37665)
--	g28720 = NOT(g28495)
--	g28721 = NOT(g28490)
--	g28723 = NOT(g28528)
--	g28725 = NOT(g28499)
--	g28727 = NOT(g28489)
--	g28730 = NOT(g28470)
--	g28734 = NOT(g28525)
--	g28740 = NOT(g28488)
--	I37702 = NOT(g28512)
--	g28741 = NOT(I37702)
--	I37712 = NOT(g28512)
--	g28751 = NOT(I37712)
--	I37716 = NOT(g28540)
--	g28755 = NOT(I37716)
--	I37725 = NOT(g28540)
--	g28764 = NOT(I37725)
--	I37729 = NOT(g28567)
--	g28768 = NOT(I37729)
--	I37736 = NOT(g28567)
--	g28775 = NOT(I37736)
--	I37740 = NOT(g28595)
--	g28779 = NOT(I37740)
--	I37746 = NOT(g28595)
--	g28785 = NOT(I37746)
--	I37752 = NOT(g28512)
--	g28791 = NOT(I37752)
--	I37757 = NOT(g28512)
--	g28796 = NOT(I37757)
--	I37760 = NOT(g28540)
--	g28799 = NOT(I37760)
--	I37765 = NOT(g28512)
--	g28804 = NOT(I37765)
--	I37768 = NOT(g28540)
--	g28807 = NOT(I37768)
--	I37771 = NOT(g28567)
--	g28810 = NOT(I37771)
--	I37775 = NOT(g28540)
--	g28814 = NOT(I37775)
--	I37778 = NOT(g28567)
--	g28817 = NOT(I37778)
--	I37781 = NOT(g28595)
--	g28820 = NOT(I37781)
--	I37784 = NOT(g28567)
--	g28823 = NOT(I37784)
--	I37787 = NOT(g28595)
--	g28826 = NOT(I37787)
--	I37790 = NOT(g28595)
--	g28829 = NOT(I37790)
--	I37793 = NOT(g28638)
--	g28832 = NOT(I37793)
--	I37796 = NOT(g28634)
--	g28833 = NOT(I37796)
--	I37800 = NOT(g28635)
--	g28835 = NOT(I37800)
--	I37804 = NOT(g28636)
--	g28837 = NOT(I37804)
--	I37808 = NOT(g28637)
--	g28839 = NOT(I37808)
--	g28855 = NOT(g28409)
--	g28859 = NOT(g28413)
--	g28863 = NOT(g28417)
--	g28867 = NOT(g28418)
--	I37842 = NOT(g28501)
--	g28871 = NOT(I37842)
--	I37846 = NOT(g28501)
--	g28877 = NOT(I37846)
--	I37851 = NOT(g28668)
--	g28882 = NOT(I37851)
--	I37854 = NOT(g28529)
--	g28883 = NOT(I37854)
--	I37858 = NOT(g28501)
--	g28889 = NOT(I37858)
--	I37863 = NOT(g28529)
--	g28894 = NOT(I37863)
--	I37868 = NOT(g28321)
--	g28899 = NOT(I37868)
--	I37871 = NOT(g28556)
--	g28900 = NOT(I37871)
--	I37875 = NOT(g28501)
--	g28906 = NOT(I37875)
--	I37880 = NOT(g28529)
--	g28911 = NOT(I37880)
--	I37885 = NOT(g28556)
--	g28916 = NOT(I37885)
--	I37891 = NOT(g28325)
--	g28924 = NOT(I37891)
--	I37894 = NOT(g28584)
--	g28925 = NOT(I37894)
--	I37897 = NOT(g28501)
--	g28928 = NOT(I37897)
--	I37901 = NOT(g28529)
--	g28932 = NOT(I37901)
--	I37906 = NOT(g28556)
--	g28937 = NOT(I37906)
--	I37912 = NOT(g28584)
--	g28945 = NOT(I37912)
--	I37917 = NOT(g28328)
--	g28950 = NOT(I37917)
--	I37920 = NOT(g28501)
--	g28951 = NOT(I37920)
--	I37924 = NOT(g28529)
--	g28955 = NOT(I37924)
--	I37928 = NOT(g28556)
--	g28959 = NOT(I37928)
--	I37934 = NOT(g28584)
--	g28967 = NOT(I37934)
--	I37939 = NOT(g28501)
--	g28972 = NOT(I37939)
--	I37942 = NOT(g28501)
--	g28975 = NOT(I37942)
--	I37946 = NOT(g28529)
--	g28979 = NOT(I37946)
--	I37950 = NOT(g28556)
--	g28983 = NOT(I37950)
--	I37956 = NOT(g28584)
--	g28993 = NOT(I37956)
--	I37961 = NOT(g28501)
--	g28998 = NOT(I37961)
--	I37965 = NOT(g28529)
--	g29002 = NOT(I37965)
--	I37968 = NOT(g28529)
--	g29005 = NOT(I37968)
--	I37973 = NOT(g28556)
--	g29010 = NOT(I37973)
--	I37978 = NOT(g28584)
--	g29019 = NOT(I37978)
--	I37982 = NOT(g28501)
--	g29023 = NOT(I37982)
--	I37986 = NOT(g28529)
--	g29027 = NOT(I37986)
--	I37991 = NOT(g28556)
--	g29032 = NOT(I37991)
--	I37994 = NOT(g28556)
--	g29035 = NOT(I37994)
--	I37999 = NOT(g28584)
--	g29042 = NOT(I37999)
--	I38003 = NOT(g28529)
--	g29046 = NOT(I38003)
--	I38007 = NOT(g28556)
--	g29050 = NOT(I38007)
--	I38011 = NOT(g28584)
--	g29054 = NOT(I38011)
--	I38014 = NOT(g28584)
--	g29057 = NOT(I38014)
--	I38018 = NOT(g28342)
--	g29061 = NOT(I38018)
--	I38024 = NOT(g28556)
--	g29065 = NOT(I38024)
--	I38028 = NOT(g28584)
--	g29069 = NOT(I38028)
--	I38032 = NOT(g28344)
--	g29073 = NOT(I38032)
--	I38035 = NOT(g28345)
--	g29074 = NOT(I38035)
--	I38038 = NOT(g28346)
--	g29075 = NOT(I38038)
--	I38042 = NOT(g28584)
--	g29077 = NOT(I38042)
--	I38046 = NOT(g28348)
--	g29081 = NOT(I38046)
--	I38049 = NOT(g28349)
--	g29082 = NOT(I38049)
--	I38053 = NOT(g28350)
--	g29084 = NOT(I38053)
--	I38056 = NOT(g28351)
--	g29085 = NOT(I38056)
--	I38059 = NOT(g28352)
--	g29086 = NOT(I38059)
--	I38064 = NOT(g28353)
--	g29089 = NOT(I38064)
--	I38068 = NOT(g28354)
--	g29091 = NOT(I38068)
--	I38071 = NOT(g28355)
--	g29092 = NOT(I38071)
--	I38074 = NOT(g28356)
--	g29093 = NOT(I38074)
--	I38077 = NOT(g28357)
--	g29094 = NOT(I38077)
--	I38080 = NOT(g28358)
--	g29095 = NOT(I38080)
--	I38085 = NOT(g28360)
--	g29098 = NOT(I38085)
--	I38088 = NOT(g28361)
--	g29099 = NOT(I38088)
--	I38091 = NOT(g28362)
--	g29100 = NOT(I38091)
--	I38094 = NOT(g28363)
--	g29101 = NOT(I38094)
--	I38097 = NOT(g28364)
--	g29102 = NOT(I38097)
--	I38101 = NOT(g28366)
--	g29104 = NOT(I38101)
--	I38104 = NOT(g28367)
--	g29105 = NOT(I38104)
--	I38107 = NOT(g28368)
--	g29106 = NOT(I38107)
--	I38111 = NOT(g28371)
--	g29108 = NOT(I38111)
--	I38119 = NOT(g28420)
--	g29117 = NOT(I38119)
--	I38122 = NOT(g28421)
--	g29118 = NOT(I38122)
--	I38125 = NOT(g28425)
--	g29119 = NOT(I38125)
--	I38128 = NOT(g28419)
--	g29120 = NOT(I38128)
--	I38136 = NOT(g28833)
--	g29131 = NOT(I38136)
--	I38139 = NOT(g29061)
--	g29132 = NOT(I38139)
--	I38142 = NOT(g29073)
--	g29133 = NOT(I38142)
--	I38145 = NOT(g29081)
--	g29134 = NOT(I38145)
--	I38148 = NOT(g29074)
--	g29135 = NOT(I38148)
--	I38151 = NOT(g29082)
--	g29136 = NOT(I38151)
--	I38154 = NOT(g29089)
--	g29137 = NOT(I38154)
--	I38157 = NOT(g28882)
--	g29138 = NOT(I38157)
--	I38160 = NOT(g28835)
--	g29139 = NOT(I38160)
--	I38163 = NOT(g29075)
--	g29140 = NOT(I38163)
--	I38166 = NOT(g29084)
--	g29141 = NOT(I38166)
--	I38169 = NOT(g29091)
--	g29142 = NOT(I38169)
--	I38172 = NOT(g29085)
--	g29143 = NOT(I38172)
--	I38175 = NOT(g29092)
--	g29144 = NOT(I38175)
--	I38178 = NOT(g29098)
--	g29145 = NOT(I38178)
--	I38181 = NOT(g28899)
--	g29146 = NOT(I38181)
--	I38184 = NOT(g28837)
--	g29147 = NOT(I38184)
--	I38187 = NOT(g29086)
--	g29148 = NOT(I38187)
--	I38190 = NOT(g29093)
--	g29149 = NOT(I38190)
--	I38193 = NOT(g29099)
--	g29150 = NOT(I38193)
--	I38196 = NOT(g29094)
--	g29151 = NOT(I38196)
--	I38199 = NOT(g29100)
--	g29152 = NOT(I38199)
--	I38202 = NOT(g29104)
--	g29153 = NOT(I38202)
--	I38205 = NOT(g28924)
--	g29154 = NOT(I38205)
--	I38208 = NOT(g28839)
--	g29155 = NOT(I38208)
--	I38211 = NOT(g29095)
--	g29156 = NOT(I38211)
--	I38214 = NOT(g29101)
--	g29157 = NOT(I38214)
--	I38217 = NOT(g29105)
--	g29158 = NOT(I38217)
--	I38220 = NOT(g29102)
--	g29159 = NOT(I38220)
--	I38223 = NOT(g29106)
--	g29160 = NOT(I38223)
--	I38226 = NOT(g29108)
--	g29161 = NOT(I38226)
--	I38229 = NOT(g28950)
--	g29162 = NOT(I38229)
--	I38232 = NOT(g29117)
--	g29163 = NOT(I38232)
--	I38235 = NOT(g29118)
--	g29164 = NOT(I38235)
--	I38238 = NOT(g29119)
--	g29165 = NOT(I38238)
--	I38241 = NOT(g28832)
--	g29166 = NOT(I38241)
--	I38245 = NOT(g28920)
--	g29168 = NOT(I38245)
--	I38250 = NOT(g28941)
--	g29171 = NOT(I38250)
--	I38258 = NOT(g28963)
--	g29177 = NOT(I38258)
--	I38272 = NOT(g29013)
--	g29189 = NOT(I38272)
--	I38275 = NOT(g28987)
--	g29190 = NOT(I38275)
--	I38278 = NOT(g28963)
--	g29191 = NOT(I38278)
--	g29192 = NOT(g28954)
--	I38282 = NOT(g28941)
--	g29193 = NOT(I38282)
--	I38321 = NOT(g29113)
--	g29230 = NOT(I38321)
--	I38330 = NOT(g29120)
--	g29237 = NOT(I38330)
--	I38339 = NOT(g29120)
--	g29244 = NOT(I38339)
--	I38342 = NOT(g28886)
--	g29245 = NOT(I38342)
--	I38345 = NOT(g29109)
--	g29246 = NOT(I38345)
--	I38348 = NOT(g28874)
--	g29247 = NOT(I38348)
--	I38352 = NOT(g29110)
--	g29249 = NOT(I38352)
--	I38355 = NOT(g29039)
--	g29250 = NOT(I38355)
--	I38360 = NOT(g29111)
--	g29253 = NOT(I38360)
--	I38363 = NOT(g29016)
--	g29254 = NOT(I38363)
--	I38369 = NOT(g29112)
--	g29258 = NOT(I38369)
--	g29266 = NOT(g28741)
--	I38386 = NOT(g28734)
--	g29267 = NOT(I38386)
--	g29268 = NOT(g28751)
--	g29269 = NOT(g28755)
--	I38391 = NOT(g28730)
--	g29270 = NOT(I38391)
--	g29271 = NOT(g28764)
--	g29272 = NOT(g28768)
--	I38396 = NOT(g28727)
--	g29273 = NOT(I38396)
--	g29274 = NOT(g28775)
--	g29275 = NOT(g28779)
--	I38401 = NOT(g28725)
--	g29276 = NOT(I38401)
--	g29277 = NOT(g28785)
--	I38405 = NOT(g28723)
--	g29278 = NOT(I38405)
--	I38408 = NOT(g28721)
--	g29279 = NOT(I38408)
--	g29280 = NOT(g28791)
--	I38412 = NOT(g28720)
--	g29281 = NOT(I38412)
--	g29282 = NOT(g28796)
--	g29283 = NOT(g28799)
--	g29285 = NOT(g28804)
--	g29286 = NOT(g28807)
--	g29287 = NOT(g28810)
--	I38421 = NOT(g28740)
--	g29288 = NOT(I38421)
--	g29290 = NOT(g28814)
--	g29291 = NOT(g28817)
--	g29292 = NOT(g28820)
--	I38428 = NOT(g28732)
--	g29293 = NOT(I38428)
--	g29295 = NOT(g28823)
--	g29296 = NOT(g28826)
--	I38434 = NOT(g28735)
--	g29297 = NOT(I38434)
--	I38437 = NOT(g28736)
--	g29298 = NOT(I38437)
--	I38440 = NOT(g28738)
--	g29299 = NOT(I38440)
--	g29301 = NOT(g28829)
--	I38447 = NOT(g28744)
--	g29304 = NOT(I38447)
--	I38450 = NOT(g28745)
--	g29305 = NOT(I38450)
--	I38453 = NOT(g28746)
--	g29306 = NOT(I38453)
--	I38456 = NOT(g28747)
--	g29307 = NOT(I38456)
--	I38459 = NOT(g28749)
--	g29308 = NOT(I38459)
--	I38462 = NOT(g29120)
--	g29309 = NOT(I38462)
--	I38466 = NOT(g28754)
--	g29311 = NOT(I38466)
--	I38471 = NOT(g28758)
--	g29314 = NOT(I38471)
--	I38474 = NOT(g28759)
--	g29315 = NOT(I38474)
--	I38477 = NOT(g28760)
--	g29316 = NOT(I38477)
--	I38480 = NOT(g28761)
--	g29317 = NOT(I38480)
--	I38483 = NOT(g28990)
--	g29318 = NOT(I38483)
--	I38486 = NOT(g28763)
--	g29319 = NOT(I38486)
--	I38491 = NOT(g28767)
--	g29322 = NOT(I38491)
--	I38496 = NOT(g28771)
--	g29325 = NOT(I38496)
--	I38499 = NOT(g28772)
--	g29326 = NOT(I38499)
--	I38502 = NOT(g28773)
--	g29327 = NOT(I38502)
--	I38505 = NOT(g28774)
--	g29328 = NOT(I38505)
--	I38510 = NOT(g28778)
--	g29331 = NOT(I38510)
--	I38515 = NOT(g28782)
--	g29334 = NOT(I38515)
--	I38518 = NOT(g28783)
--	g29335 = NOT(I38518)
--	I38524 = NOT(g28788)
--	g29339 = NOT(I38524)
--	I38536 = NOT(g28920)
--	g29349 = NOT(I38536)
--	I38539 = NOT(g29113)
--	g29350 = NOT(I38539)
--	g29356 = NOT(g29120)
--	g29358 = NOT(g29120)
--	I38548 = NOT(g28903)
--	g29359 = NOT(I38548)
--	g29360 = NOT(g28871)
--	g29361 = NOT(g28877)
--	g29362 = NOT(g28883)
--	g29363 = NOT(g28889)
--	g29364 = NOT(g28894)
--	g29365 = NOT(g28900)
--	g29366 = NOT(g28906)
--	g29367 = NOT(g28911)
--	g29368 = NOT(g28916)
--	g29369 = NOT(g28925)
--	g29370 = NOT(g28928)
--	g29371 = NOT(g28932)
--	g29372 = NOT(g28937)
--	g29373 = NOT(g28945)
--	g29374 = NOT(g28951)
--	g29375 = NOT(g28955)
--	g29376 = NOT(g28959)
--	g29377 = NOT(g28967)
--	g29378 = NOT(g28972)
--	g29379 = NOT(g28975)
--	g29380 = NOT(g28979)
--	g29381 = NOT(g28983)
--	g29382 = NOT(g28993)
--	g29383 = NOT(g28998)
--	g29384 = NOT(g29002)
--	g29385 = NOT(g29005)
--	g29386 = NOT(g29010)
--	g29387 = NOT(g29019)
--	g29388 = NOT(g29023)
--	g29389 = NOT(g29027)
--	g29390 = NOT(g29032)
--	g29391 = NOT(g29035)
--	g29392 = NOT(g29042)
--	g29393 = NOT(g29046)
--	g29394 = NOT(g29050)
--	g29395 = NOT(g29054)
--	g29396 = NOT(g29057)
--	g29397 = NOT(g29065)
--	g29398 = NOT(g29069)
--	I38591 = NOT(g28987)
--	g29400 = NOT(I38591)
--	I38594 = NOT(g28990)
--	g29401 = NOT(I38594)
--	g29402 = NOT(g29077)
--	I38599 = NOT(g29013)
--	g29404 = NOT(I38599)
--	I38602 = NOT(g29016)
--	g29405 = NOT(I38602)
--	I38606 = NOT(g29039)
--	g29407 = NOT(I38606)
--	I38609 = NOT(g28874)
--	g29408 = NOT(I38609)
--	I38613 = NOT(g28886)
--	g29410 = NOT(I38613)
--	I38617 = NOT(g28903)
--	g29412 = NOT(I38617)
--	I38620 = NOT(g29246)
--	g29413 = NOT(I38620)
--	I38623 = NOT(g29293)
--	g29414 = NOT(I38623)
--	I38626 = NOT(g29297)
--	g29415 = NOT(I38626)
--	I38629 = NOT(g29304)
--	g29416 = NOT(I38629)
--	I38632 = NOT(g29298)
--	g29417 = NOT(I38632)
--	I38635 = NOT(g29305)
--	g29418 = NOT(I38635)
--	I38638 = NOT(g29311)
--	g29419 = NOT(I38638)
--	I38641 = NOT(g29249)
--	g29420 = NOT(I38641)
--	I38644 = NOT(g29299)
--	g29421 = NOT(I38644)
--	I38647 = NOT(g29306)
--	g29422 = NOT(I38647)
--	I38650 = NOT(g29314)
--	g29423 = NOT(I38650)
--	I38653 = NOT(g29307)
--	g29424 = NOT(I38653)
--	I38656 = NOT(g29315)
--	g29425 = NOT(I38656)
--	I38659 = NOT(g29322)
--	g29426 = NOT(I38659)
--	I38662 = NOT(g29253)
--	g29427 = NOT(I38662)
--	I38665 = NOT(g29412)
--	g29428 = NOT(I38665)
--	I38668 = NOT(g29168)
--	g29429 = NOT(I38668)
--	I38671 = NOT(g29171)
--	g29430 = NOT(I38671)
--	I38674 = NOT(g29177)
--	g29431 = NOT(I38674)
--	I38677 = NOT(g29400)
--	g29432 = NOT(I38677)
--	I38680 = NOT(g29404)
--	g29433 = NOT(I38680)
--	I38683 = NOT(g29308)
--	g29434 = NOT(I38683)
--	I38686 = NOT(g29316)
--	g29435 = NOT(I38686)
--	I38689 = NOT(g29325)
--	g29436 = NOT(I38689)
--	I38692 = NOT(g29317)
--	g29437 = NOT(I38692)
--	I38695 = NOT(g29326)
--	g29438 = NOT(I38695)
--	I38698 = NOT(g29331)
--	g29439 = NOT(I38698)
--	I38701 = NOT(g29401)
--	g29440 = NOT(I38701)
--	I38704 = NOT(g29405)
--	g29441 = NOT(I38704)
--	I38707 = NOT(g29407)
--	g29442 = NOT(I38707)
--	I38710 = NOT(g29408)
--	g29443 = NOT(I38710)
--	I38713 = NOT(g29410)
--	g29444 = NOT(I38713)
--	I38716 = NOT(g29230)
--	g29445 = NOT(I38716)
--	I38719 = NOT(g29258)
--	g29446 = NOT(I38719)
--	I38722 = NOT(g29319)
--	g29447 = NOT(I38722)
--	I38725 = NOT(g29327)
--	g29448 = NOT(I38725)
--	I38728 = NOT(g29334)
--	g29449 = NOT(I38728)
--	I38731 = NOT(g29328)
--	g29450 = NOT(I38731)
--	I38734 = NOT(g29335)
--	g29451 = NOT(I38734)
--	I38737 = NOT(g29339)
--	g29452 = NOT(I38737)
--	I38740 = NOT(g29288)
--	g29453 = NOT(I38740)
--	I38743 = NOT(g29267)
--	g29454 = NOT(I38743)
--	I38746 = NOT(g29270)
--	g29455 = NOT(I38746)
--	I38749 = NOT(g29273)
--	g29456 = NOT(I38749)
--	I38752 = NOT(g29276)
--	g29457 = NOT(I38752)
--	I38755 = NOT(g29278)
--	g29458 = NOT(I38755)
--	I38758 = NOT(g29279)
--	g29459 = NOT(I38758)
--	I38761 = NOT(g29281)
--	g29460 = NOT(I38761)
--	I38764 = NOT(g29237)
--	g29461 = NOT(I38764)
--	I38767 = NOT(g29244)
--	g29462 = NOT(I38767)
--	I38770 = NOT(g29309)
--	g29463 = NOT(I38770)
--	g29491 = NOT(g29350)
--	I38801 = NOT(g29358)
--	g29495 = NOT(I38801)
--	I38804 = NOT(g29353)
--	g29496 = NOT(I38804)
--	I38807 = NOT(g29356)
--	g29497 = NOT(I38807)
--	I38817 = NOT(g29354)
--	g29499 = NOT(I38817)
--	I38827 = NOT(g29355)
--	g29501 = NOT(I38827)
--	I38838 = NOT(g29357)
--	g29504 = NOT(I38838)
--	I38848 = NOT(g29167)
--	g29506 = NOT(I38848)
--	I38851 = NOT(g29169)
--	g29507 = NOT(I38851)
--	I38854 = NOT(g29170)
--	g29508 = NOT(I38854)
--	I38857 = NOT(g29172)
--	g29509 = NOT(I38857)
--	I38860 = NOT(g29173)
--	g29510 = NOT(I38860)
--	I38863 = NOT(g29178)
--	g29511 = NOT(I38863)
--	I38866 = NOT(g29179)
--	g29512 = NOT(I38866)
--	I38869 = NOT(g29181)
--	g29513 = NOT(I38869)
--	I38872 = NOT(g29182)
--	g29514 = NOT(I38872)
--	I38875 = NOT(g29184)
--	g29515 = NOT(I38875)
--	I38878 = NOT(g29185)
--	g29516 = NOT(I38878)
--	I38881 = NOT(g29187)
--	g29517 = NOT(I38881)
--	I38885 = NOT(g29192)
--	g29519 = NOT(I38885)
--	I38898 = NOT(g29194)
--	g29530 = NOT(I38898)
--	I38905 = NOT(g29197)
--	g29535 = NOT(I38905)
--	I38909 = NOT(g29198)
--	g29537 = NOT(I38909)
--	I38916 = NOT(g29201)
--	g29542 = NOT(I38916)
--	I38920 = NOT(g29204)
--	g29544 = NOT(I38920)
--	I38924 = NOT(g29205)
--	g29546 = NOT(I38924)
--	I38931 = NOT(g29209)
--	g29551 = NOT(I38931)
--	I38936 = NOT(g29212)
--	g29554 = NOT(I38936)
--	I38940 = NOT(g29213)
--	g29556 = NOT(I38940)
--	I38947 = NOT(g29218)
--	g29561 = NOT(I38947)
--	I38951 = NOT(g29221)
--	g29563 = NOT(I38951)
--	I38958 = NOT(g29226)
--	g29568 = NOT(I38958)
--	I38975 = NOT(g29348)
--	g29583 = NOT(I38975)
--	I38999 = NOT(g29496)
--	g29627 = NOT(I38999)
--	I39002 = NOT(g29506)
--	g29628 = NOT(I39002)
--	I39005 = NOT(g29507)
--	g29629 = NOT(I39005)
--	I39008 = NOT(g29509)
--	g29630 = NOT(I39008)
--	I39011 = NOT(g29530)
--	g29631 = NOT(I39011)
--	I39014 = NOT(g29535)
--	g29632 = NOT(I39014)
--	I39017 = NOT(g29542)
--	g29633 = NOT(I39017)
--	I39020 = NOT(g29499)
--	g29634 = NOT(I39020)
--	I39023 = NOT(g29508)
--	g29635 = NOT(I39023)
--	I39026 = NOT(g29510)
--	g29636 = NOT(I39026)
--	I39029 = NOT(g29512)
--	g29637 = NOT(I39029)
--	I39032 = NOT(g29537)
--	g29638 = NOT(I39032)
--	I39035 = NOT(g29544)
--	g29639 = NOT(I39035)
--	I39038 = NOT(g29551)
--	g29640 = NOT(I39038)
--	I39041 = NOT(g29501)
--	g29641 = NOT(I39041)
--	I39044 = NOT(g29511)
--	g29642 = NOT(I39044)
--	I39047 = NOT(g29513)
--	g29643 = NOT(I39047)
--	I39050 = NOT(g29515)
--	g29644 = NOT(I39050)
--	I39053 = NOT(g29546)
--	g29645 = NOT(I39053)
--	I39056 = NOT(g29554)
--	g29646 = NOT(I39056)
--	I39059 = NOT(g29561)
--	g29647 = NOT(I39059)
--	I39062 = NOT(g29504)
--	g29648 = NOT(I39062)
--	I39065 = NOT(g29514)
--	g29649 = NOT(I39065)
--	I39068 = NOT(g29516)
--	g29650 = NOT(I39068)
--	I39071 = NOT(g29517)
--	g29651 = NOT(I39071)
--	I39074 = NOT(g29556)
--	g29652 = NOT(I39074)
--	I39077 = NOT(g29563)
--	g29653 = NOT(I39077)
--	I39080 = NOT(g29568)
--	g29654 = NOT(I39080)
--	I39083 = NOT(g29519)
--	g29655 = NOT(I39083)
--	I39086 = NOT(g29497)
--	g29656 = NOT(I39086)
--	I39089 = NOT(g29495)
--	g29657 = NOT(I39089)
--	g29658 = NOT(g29574)
--	g29659 = NOT(g29571)
--	g29660 = NOT(g29578)
--	g29661 = NOT(g29576)
--	g29662 = NOT(g29570)
--	g29664 = NOT(g29552)
--	g29666 = NOT(g29577)
--	g29668 = NOT(g29569)
--	g29673 = NOT(g29583)
--	I39121 = NOT(g29579)
--	g29689 = NOT(I39121)
--	I39124 = NOT(g29606)
--	g29690 = NOT(I39124)
--	I39127 = NOT(g29608)
--	g29691 = NOT(I39127)
--	I39130 = NOT(g29580)
--	g29692 = NOT(I39130)
--	I39133 = NOT(g29609)
--	g29693 = NOT(I39133)
--	I39136 = NOT(g29611)
--	g29694 = NOT(I39136)
--	I39139 = NOT(g29612)
--	g29695 = NOT(I39139)
--	I39142 = NOT(g29581)
--	g29696 = NOT(I39142)
--	I39145 = NOT(g29613)
--	g29697 = NOT(I39145)
--	I39148 = NOT(g29616)
--	g29698 = NOT(I39148)
--	I39151 = NOT(g29617)
--	g29699 = NOT(I39151)
--	I39154 = NOT(g29582)
--	g29700 = NOT(I39154)
--	I39157 = NOT(g29618)
--	g29701 = NOT(I39157)
--	I39160 = NOT(g29620)
--	g29702 = NOT(I39160)
--	I39164 = NOT(g29621)
--	g29704 = NOT(I39164)
--	I39168 = NOT(g29623)
--	g29708 = NOT(I39168)
--	g29716 = NOT(g29498)
--	g29724 = NOT(g29500)
--	g29726 = NOT(g29503)
--	g29739 = NOT(g29505)
--	I39234 = NOT(g29689)
--	g29794 = NOT(I39234)
--	I39237 = NOT(g29690)
--	g29795 = NOT(I39237)
--	I39240 = NOT(g29691)
--	g29796 = NOT(I39240)
--	I39243 = NOT(g29694)
--	g29797 = NOT(I39243)
--	I39246 = NOT(g29692)
--	g29798 = NOT(I39246)
--	I39249 = NOT(g29693)
--	g29799 = NOT(I39249)
--	I39252 = NOT(g29695)
--	g29800 = NOT(I39252)
--	I39255 = NOT(g29698)
--	g29801 = NOT(I39255)
--	I39258 = NOT(g29696)
--	g29802 = NOT(I39258)
--	I39261 = NOT(g29697)
--	g29803 = NOT(I39261)
--	I39264 = NOT(g29699)
--	g29804 = NOT(I39264)
--	I39267 = NOT(g29702)
--	g29805 = NOT(I39267)
--	I39270 = NOT(g29700)
--	g29806 = NOT(I39270)
--	I39273 = NOT(g29701)
--	g29807 = NOT(I39273)
--	I39276 = NOT(g29704)
--	g29808 = NOT(I39276)
--	I39279 = NOT(g29708)
--	g29809 = NOT(I39279)
--	g29823 = NOT(g29663)
--	g29829 = NOT(g29665)
--	g29835 = NOT(g29667)
--	g29840 = NOT(g29669)
--	g29844 = NOT(g29670)
--	g29848 = NOT(g29761)
--	g29849 = NOT(g29671)
--	g29853 = NOT(g29672)
--	g29857 = NOT(g29676)
--	g29861 = NOT(g29677)
--	g29865 = NOT(g29678)
--	g29869 = NOT(g29679)
--	g29873 = NOT(g29680)
--	g29877 = NOT(g29681)
--	g29881 = NOT(g29682)
--	g29885 = NOT(g29683)
--	g29889 = NOT(g29684)
--	g29893 = NOT(g29685)
--	g29897 = NOT(g29686)
--	g29901 = NOT(g29687)
--	g29905 = NOT(g29688)
--	I39398 = NOT(g29664)
--	g29932 = NOT(I39398)
--	I39401 = NOT(g29662)
--	g29933 = NOT(I39401)
--	I39404 = NOT(g29661)
--	g29934 = NOT(I39404)
--	I39407 = NOT(g29660)
--	g29935 = NOT(I39407)
--	I39411 = NOT(g29659)
--	g29937 = NOT(I39411)
--	I39414 = NOT(g29658)
--	g29938 = NOT(I39414)
--	I39418 = NOT(g29668)
--	g29940 = NOT(I39418)
--	I39423 = NOT(g29666)
--	g29943 = NOT(I39423)
--	I39454 = NOT(g29940)
--	g29972 = NOT(I39454)
--	I39457 = NOT(g29943)
--	g29973 = NOT(I39457)
--	I39460 = NOT(g29932)
--	g29974 = NOT(I39460)
--	I39463 = NOT(g29933)
--	g29975 = NOT(I39463)
--	I39466 = NOT(g29934)
--	g29976 = NOT(I39466)
--	I39469 = NOT(g29935)
--	g29977 = NOT(I39469)
--	I39472 = NOT(g29937)
--	g29978 = NOT(I39472)
--	I39475 = NOT(g29938)
--	g29979 = NOT(I39475)
--	g30036 = NOT(g29912)
--	g30040 = NOT(g29914)
--	g30044 = NOT(g29916)
--	g30048 = NOT(g29920)
--	I39550 = NOT(g29848)
--	g30052 = NOT(I39550)
--	I39573 = NOT(g29936)
--	g30076 = NOT(I39573)
--	I39577 = NOT(g29939)
--	g30078 = NOT(I39577)
--	I39585 = NOT(g29941)
--	g30084 = NOT(I39585)
--	I39622 = NOT(g30052)
--	g30119 = NOT(I39622)
--	I39625 = NOT(g30076)
--	g30120 = NOT(I39625)
--	I39628 = NOT(g30078)
--	g30121 = NOT(I39628)
--	I39631 = NOT(g30084)
--	g30122 = NOT(I39631)
--	I39635 = NOT(g30055)
--	g30124 = NOT(I39635)
--	I39638 = NOT(g30056)
--	g30125 = NOT(I39638)
--	I39641 = NOT(g30057)
--	g30126 = NOT(I39641)
--	I39647 = NOT(g30058)
--	g30130 = NOT(I39647)
--	g30134 = NOT(g30010)
--	g30139 = NOT(g30011)
--	g30143 = NOT(g30012)
--	g30147 = NOT(g30013)
--	g30151 = NOT(g30014)
--	g30155 = NOT(g30015)
--	g30159 = NOT(g30016)
--	g30163 = NOT(g30017)
--	g30167 = NOT(g30018)
--	g30171 = NOT(g30019)
--	g30175 = NOT(g30020)
--	g30179 = NOT(g30021)
--	g30183 = NOT(g30022)
--	g30187 = NOT(g30023)
--	g30191 = NOT(g30024)
--	g30195 = NOT(g30025)
--	g30199 = NOT(g30026)
--	g30203 = NOT(g30027)
--	g30207 = NOT(g30028)
--	g30211 = NOT(g30029)
--	I39674 = NOT(g30072)
--	g30215 = NOT(I39674)
--	g30229 = NOT(g30030)
--	g30233 = NOT(g30031)
--	g30237 = NOT(g30032)
--	g30241 = NOT(g30033)
--	I39761 = NOT(g30072)
--	g30306 = NOT(I39761)
--	I39764 = NOT(g30060)
--	g30307 = NOT(I39764)
--	I39767 = NOT(g30061)
--	g30308 = NOT(I39767)
--	I39770 = NOT(g30063)
--	g30309 = NOT(I39770)
--	I39773 = NOT(g30064)
--	g30310 = NOT(I39773)
--	I39776 = NOT(g30066)
--	g30311 = NOT(I39776)
--	I39779 = NOT(g30053)
--	g30312 = NOT(I39779)
--	I39782 = NOT(g30054)
--	g30313 = NOT(I39782)
--	I39785 = NOT(g30124)
--	g30314 = NOT(I39785)
--	I39788 = NOT(g30125)
--	g30315 = NOT(I39788)
--	I39791 = NOT(g30126)
--	g30316 = NOT(I39791)
--	I39794 = NOT(g30130)
--	g30317 = NOT(I39794)
--	I39797 = NOT(g30307)
--	g30318 = NOT(I39797)
--	I39800 = NOT(g30309)
--	g30319 = NOT(I39800)
--	I39803 = NOT(g30308)
--	g30320 = NOT(I39803)
--	I39806 = NOT(g30310)
--	g30321 = NOT(I39806)
--	I39809 = NOT(g30311)
--	g30322 = NOT(I39809)
--	I39812 = NOT(g30312)
--	g30323 = NOT(I39812)
--	I39815 = NOT(g30313)
--	g30324 = NOT(I39815)
--	I39818 = NOT(g30215)
--	g30325 = NOT(I39818)
--	I39821 = NOT(g30267)
--	g30326 = NOT(I39821)
--	I39825 = NOT(g30268)
--	g30328 = NOT(I39825)
--	I39828 = NOT(g30269)
--	g30329 = NOT(I39828)
--	I39832 = NOT(g30270)
--	g30331 = NOT(I39832)
--	I39835 = NOT(g30271)
--	g30332 = NOT(I39835)
--	I39840 = NOT(g30272)
--	g30335 = NOT(I39840)
--	I39843 = NOT(g30273)
--	g30336 = NOT(I39843)
--	I39848 = NOT(g30274)
--	g30339 = NOT(I39848)
--	I39853 = NOT(g30275)
--	g30342 = NOT(I39853)
--	I39856 = NOT(g30276)
--	g30343 = NOT(I39856)
--	I39859 = NOT(g30277)
--	g30344 = NOT(I39859)
--	I39863 = NOT(g30278)
--	g30346 = NOT(I39863)
--	I39866 = NOT(g30279)
--	g30347 = NOT(I39866)
--	I39870 = NOT(g30280)
--	g30349 = NOT(I39870)
--	I39873 = NOT(g30281)
--	g30350 = NOT(I39873)
--	I39878 = NOT(g30282)
--	g30353 = NOT(I39878)
--	I39881 = NOT(g30283)
--	g30354 = NOT(I39881)
--	I39886 = NOT(g30284)
--	g30357 = NOT(I39886)
--	I39889 = NOT(g30285)
--	g30358 = NOT(I39889)
--	I39892 = NOT(g30286)
--	g30359 = NOT(I39892)
--	I39895 = NOT(g30287)
--	g30360 = NOT(I39895)
--	I39899 = NOT(g30288)
--	g30362 = NOT(I39899)
--	I39902 = NOT(g30289)
--	g30363 = NOT(I39902)
--	I39906 = NOT(g30290)
--	g30365 = NOT(I39906)
--	I39909 = NOT(g30291)
--	g30366 = NOT(I39909)
--	I39913 = NOT(g30292)
--	g30368 = NOT(I39913)
--	I39916 = NOT(g30293)
--	g30369 = NOT(I39916)
--	I39919 = NOT(g30294)
--	g30370 = NOT(I39919)
--	I39922 = NOT(g30295)
--	g30371 = NOT(I39922)
--	I39926 = NOT(g30296)
--	g30373 = NOT(I39926)
--	I39930 = NOT(g30297)
--	g30375 = NOT(I39930)
--	I39933 = NOT(g30298)
--	g30376 = NOT(I39933)
--	I39936 = NOT(g30299)
--	g30377 = NOT(I39936)
--	I39939 = NOT(g30300)
--	g30378 = NOT(I39939)
--	I39942 = NOT(g30301)
--	g30379 = NOT(I39942)
--	I39945 = NOT(g30302)
--	g30380 = NOT(I39945)
--	I39948 = NOT(g30303)
--	g30381 = NOT(I39948)
--	I39951 = NOT(g30304)
--	g30382 = NOT(I39951)
--	g30383 = NOT(g30306)
--	I39976 = NOT(g30245)
--	g30408 = NOT(I39976)
--	I39982 = NOT(g30305)
--	g30412 = NOT(I39982)
--	I39985 = NOT(g30246)
--	g30435 = NOT(I39985)
--	I39991 = NOT(g30247)
--	g30439 = NOT(I39991)
--	I39997 = NOT(g30248)
--	g30443 = NOT(I39997)
--	I40002 = NOT(g30249)
--	g30446 = NOT(I40002)
--	I40008 = NOT(g30250)
--	g30450 = NOT(I40008)
--	I40016 = NOT(g30251)
--	g30456 = NOT(I40016)
--	I40021 = NOT(g30252)
--	g30459 = NOT(I40021)
--	I40027 = NOT(g30253)
--	g30463 = NOT(I40027)
--	I40032 = NOT(g30254)
--	g30466 = NOT(I40032)
--	I40039 = NOT(g30255)
--	g30471 = NOT(I40039)
--	I40044 = NOT(g30256)
--	g30474 = NOT(I40044)
--	I40051 = NOT(g30257)
--	g30479 = NOT(I40051)
--	I40054 = NOT(g30258)
--	g30480 = NOT(I40054)
--	I40059 = NOT(g30259)
--	g30483 = NOT(I40059)
--	I40066 = NOT(g30260)
--	g30488 = NOT(I40066)
--	I40071 = NOT(g30261)
--	g30491 = NOT(I40071)
--	I40075 = NOT(g30262)
--	g30493 = NOT(I40075)
--	I40078 = NOT(g30263)
--	g30494 = NOT(I40078)
--	I40083 = NOT(g30264)
--	g30497 = NOT(I40083)
--	I40086 = NOT(g30265)
--	g30498 = NOT(I40086)
--	I40091 = NOT(g30266)
--	g30501 = NOT(I40091)
--	I40098 = NOT(g30491)
--	g30506 = NOT(I40098)
--	I40101 = NOT(g30326)
--	g30507 = NOT(I40101)
--	I40104 = NOT(g30342)
--	g30508 = NOT(I40104)
--	I40107 = NOT(g30343)
--	g30509 = NOT(I40107)
--	I40110 = NOT(g30357)
--	g30510 = NOT(I40110)
--	I40113 = NOT(g30368)
--	g30511 = NOT(I40113)
--	I40116 = NOT(g30408)
--	g30512 = NOT(I40116)
--	I40119 = NOT(g30435)
--	g30513 = NOT(I40119)
--	I40122 = NOT(g30443)
--	g30514 = NOT(I40122)
--	I40125 = NOT(g30466)
--	g30515 = NOT(I40125)
--	I40128 = NOT(g30479)
--	g30516 = NOT(I40128)
--	I40131 = NOT(g30493)
--	g30517 = NOT(I40131)
--	I40134 = NOT(g30480)
--	g30518 = NOT(I40134)
--	I40137 = NOT(g30494)
--	g30519 = NOT(I40137)
--	I40140 = NOT(g30328)
--	g30520 = NOT(I40140)
--	I40143 = NOT(g30329)
--	g30521 = NOT(I40143)
--	I40146 = NOT(g30344)
--	g30522 = NOT(I40146)
--	I40149 = NOT(g30358)
--	g30523 = NOT(I40149)
--	I40152 = NOT(g30359)
--	g30524 = NOT(I40152)
--	I40155 = NOT(g30369)
--	g30525 = NOT(I40155)
--	I40158 = NOT(g30376)
--	g30526 = NOT(I40158)
--	I40161 = NOT(g30439)
--	g30527 = NOT(I40161)
--	I40164 = NOT(g30446)
--	g30528 = NOT(I40164)
--	I40167 = NOT(g30456)
--	g30529 = NOT(I40167)
--	I40170 = NOT(g30483)
--	g30530 = NOT(I40170)
--	I40173 = NOT(g30497)
--	g30531 = NOT(I40173)
--	I40176 = NOT(g30331)
--	g30532 = NOT(I40176)
--	I40179 = NOT(g30498)
--	g30533 = NOT(I40179)
--	I40182 = NOT(g30332)
--	g30534 = NOT(I40182)
--	I40185 = NOT(g30346)
--	g30535 = NOT(I40185)
--	I40188 = NOT(g30347)
--	g30536 = NOT(I40188)
--	I40191 = NOT(g30360)
--	g30537 = NOT(I40191)
--	I40194 = NOT(g30370)
--	g30538 = NOT(I40194)
--	I40197 = NOT(g30371)
--	g30539 = NOT(I40197)
--	I40200 = NOT(g30377)
--	g30540 = NOT(I40200)
--	I40203 = NOT(g30380)
--	g30541 = NOT(I40203)
--	I40206 = NOT(g30450)
--	g30542 = NOT(I40206)
--	I40209 = NOT(g30459)
--	g30543 = NOT(I40209)
--	I40212 = NOT(g30471)
--	g30544 = NOT(I40212)
--	I40215 = NOT(g30501)
--	g30545 = NOT(I40215)
--	I40218 = NOT(g30335)
--	g30546 = NOT(I40218)
--	I40221 = NOT(g30349)
--	g30547 = NOT(I40221)
--	I40224 = NOT(g30336)
--	g30548 = NOT(I40224)
--	I40227 = NOT(g30350)
--	g30549 = NOT(I40227)
--	I40230 = NOT(g30362)
--	g30550 = NOT(I40230)
--	I40233 = NOT(g30363)
--	g30551 = NOT(I40233)
--	I40236 = NOT(g30373)
--	g30552 = NOT(I40236)
--	I40239 = NOT(g30378)
--	g30553 = NOT(I40239)
--	I40242 = NOT(g30379)
--	g30554 = NOT(I40242)
--	I40245 = NOT(g30381)
--	g30555 = NOT(I40245)
--	I40248 = NOT(g30382)
--	g30556 = NOT(I40248)
--	I40251 = NOT(g30463)
--	g30557 = NOT(I40251)
--	I40254 = NOT(g30474)
--	g30558 = NOT(I40254)
--	I40257 = NOT(g30488)
--	g30559 = NOT(I40257)
--	I40260 = NOT(g30339)
--	g30560 = NOT(I40260)
--	I40263 = NOT(g30353)
--	g30561 = NOT(I40263)
--	I40266 = NOT(g30365)
--	g30562 = NOT(I40266)
--	I40269 = NOT(g30354)
--	g30563 = NOT(I40269)
--	I40272 = NOT(g30366)
--	g30564 = NOT(I40272)
--	I40275 = NOT(g30375)
--	g30565 = NOT(I40275)
--	g30567 = NOT(g30403)
--	g30568 = NOT(g30402)
--	g30569 = NOT(g30406)
--	g30570 = NOT(g30404)
--	g30571 = NOT(g30401)
--	g30572 = NOT(g30399)
--	g30573 = NOT(g30405)
--	g30574 = NOT(g30400)
--	g30575 = NOT(g30412)
--	I40288 = NOT(g30455)
--	g30578 = NOT(I40288)
--	I40291 = NOT(g30468)
--	g30579 = NOT(I40291)
--	I40294 = NOT(g30470)
--	g30580 = NOT(I40294)
--	I40297 = NOT(g30482)
--	g30581 = NOT(I40297)
--	I40300 = NOT(g30485)
--	g30582 = NOT(I40300)
--	I40303 = NOT(g30487)
--	g30583 = NOT(I40303)
--	I40307 = NOT(g30500)
--	g30585 = NOT(I40307)
--	I40310 = NOT(g30503)
--	g30586 = NOT(I40310)
--	I40313 = NOT(g30505)
--	g30587 = NOT(I40313)
--	I40317 = NOT(g30338)
--	g30591 = NOT(I40317)
--	I40320 = NOT(g30341)
--	g30592 = NOT(I40320)
--	I40326 = NOT(g30356)
--	g30600 = NOT(I40326)
--	I40420 = NOT(g30578)
--	g30710 = NOT(I40420)
--	I40423 = NOT(g30579)
--	g30711 = NOT(I40423)
--	I40426 = NOT(g30581)
--	g30712 = NOT(I40426)
--	I40429 = NOT(g30580)
--	g30713 = NOT(I40429)
--	I40432 = NOT(g30582)
--	g30714 = NOT(I40432)
--	I40435 = NOT(g30585)
--	g30715 = NOT(I40435)
--	I40438 = NOT(g30583)
--	g30716 = NOT(I40438)
--	I40441 = NOT(g30586)
--	g30717 = NOT(I40441)
--	I40444 = NOT(g30591)
--	g30718 = NOT(I40444)
--	I40447 = NOT(g30587)
--	g30719 = NOT(I40447)
--	I40450 = NOT(g30592)
--	g30720 = NOT(I40450)
--	I40453 = NOT(g30600)
--	g30721 = NOT(I40453)
--	I40456 = NOT(g30668)
--	g30722 = NOT(I40456)
--	I40459 = NOT(g30669)
--	g30723 = NOT(I40459)
--	I40462 = NOT(g30670)
--	g30724 = NOT(I40462)
--	I40465 = NOT(g30671)
--	g30725 = NOT(I40465)
--	I40468 = NOT(g30672)
--	g30726 = NOT(I40468)
--	I40471 = NOT(g30673)
--	g30727 = NOT(I40471)
--	I40475 = NOT(g30674)
--	g30729 = NOT(I40475)
--	I40478 = NOT(g30675)
--	g30730 = NOT(I40478)
--	I40481 = NOT(g30676)
--	g30731 = NOT(I40481)
--	I40484 = NOT(g30677)
--	g30732 = NOT(I40484)
--	I40487 = NOT(g30678)
--	g30733 = NOT(I40487)
--	I40490 = NOT(g30679)
--	g30734 = NOT(I40490)
--	I40495 = NOT(g30680)
--	g30737 = NOT(I40495)
--	I40498 = NOT(g30681)
--	g30738 = NOT(I40498)
--	I40501 = NOT(g30682)
--	g30739 = NOT(I40501)
--	I40504 = NOT(g30683)
--	g30740 = NOT(I40504)
--	I40507 = NOT(g30684)
--	g30741 = NOT(I40507)
--	I40510 = NOT(g30686)
--	g30742 = NOT(I40510)
--	I40515 = NOT(g30687)
--	g30745 = NOT(I40515)
--	I40518 = NOT(g30688)
--	g30746 = NOT(I40518)
--	I40521 = NOT(g30689)
--	g30747 = NOT(I40521)
--	I40524 = NOT(g30690)
--	g30748 = NOT(I40524)
--	I40527 = NOT(g30691)
--	g30749 = NOT(I40527)
--	I40531 = NOT(g30692)
--	g30751 = NOT(I40531)
--	I40534 = NOT(g30693)
--	g30752 = NOT(I40534)
--	I40537 = NOT(g30694)
--	g30753 = NOT(I40537)
--	I40542 = NOT(g30695)
--	g30756 = NOT(I40542)
--	g30765 = NOT(g30685)
--	I40555 = NOT(g30699)
--	g30767 = NOT(I40555)
--	I40565 = NOT(g30700)
--	g30769 = NOT(I40565)
--	I40568 = NOT(g30701)
--	g30770 = NOT(I40568)
--	I40578 = NOT(g30702)
--	g30772 = NOT(I40578)
--	I40581 = NOT(g30703)
--	g30773 = NOT(I40581)
--	I40584 = NOT(g30704)
--	g30774 = NOT(I40584)
--	I40594 = NOT(g30705)
--	g30776 = NOT(I40594)
--	I40597 = NOT(g30706)
--	g30777 = NOT(I40597)
--	I40600 = NOT(g30707)
--	g30778 = NOT(I40600)
--	I40611 = NOT(g30708)
--	g30781 = NOT(I40611)
--	I40614 = NOT(g30709)
--	g30782 = NOT(I40614)
--	I40618 = NOT(g30566)
--	g30784 = NOT(I40618)
--	I40634 = NOT(g30571)
--	g30792 = NOT(I40634)
--	I40637 = NOT(g30570)
--	g30793 = NOT(I40637)
--	I40640 = NOT(g30569)
--	g30794 = NOT(I40640)
--	I40643 = NOT(g30568)
--	g30795 = NOT(I40643)
--	I40647 = NOT(g30567)
--	g30797 = NOT(I40647)
--	I40651 = NOT(g30574)
--	g30799 = NOT(I40651)
--	I40654 = NOT(g30573)
--	g30800 = NOT(I40654)
--	I40658 = NOT(g30572)
--	g30802 = NOT(I40658)
--	I40661 = NOT(g30635)
--	g30803 = NOT(I40661)
--	I40664 = NOT(g30636)
--	g30804 = NOT(I40664)
--	I40667 = NOT(g30637)
--	g30805 = NOT(I40667)
--	I40670 = NOT(g30638)
--	g30806 = NOT(I40670)
--	I40673 = NOT(g30639)
--	g30807 = NOT(I40673)
--	I40676 = NOT(g30640)
--	g30808 = NOT(I40676)
--	I40679 = NOT(g30641)
--	g30809 = NOT(I40679)
--	I40682 = NOT(g30642)
--	g30810 = NOT(I40682)
--	I40685 = NOT(g30643)
--	g30811 = NOT(I40685)
--	I40688 = NOT(g30644)
--	g30812 = NOT(I40688)
--	I40691 = NOT(g30645)
--	g30813 = NOT(I40691)
--	I40694 = NOT(g30646)
--	g30814 = NOT(I40694)
--	I40697 = NOT(g30647)
--	g30815 = NOT(I40697)
--	I40700 = NOT(g30648)
--	g30816 = NOT(I40700)
--	I40703 = NOT(g30649)
--	g30817 = NOT(I40703)
--	I40706 = NOT(g30650)
--	g30818 = NOT(I40706)
--	I40709 = NOT(g30651)
--	g30819 = NOT(I40709)
--	I40712 = NOT(g30652)
--	g30820 = NOT(I40712)
--	I40715 = NOT(g30653)
--	g30821 = NOT(I40715)
--	I40718 = NOT(g30654)
--	g30822 = NOT(I40718)
--	I40721 = NOT(g30655)
--	g30823 = NOT(I40721)
--	I40724 = NOT(g30656)
--	g30824 = NOT(I40724)
--	I40727 = NOT(g30657)
--	g30825 = NOT(I40727)
--	I40730 = NOT(g30658)
--	g30826 = NOT(I40730)
--	I40733 = NOT(g30659)
--	g30827 = NOT(I40733)
--	I40736 = NOT(g30660)
--	g30828 = NOT(I40736)
--	I40739 = NOT(g30661)
--	g30829 = NOT(I40739)
--	I40742 = NOT(g30662)
--	g30830 = NOT(I40742)
--	I40745 = NOT(g30663)
--	g30831 = NOT(I40745)
--	I40748 = NOT(g30664)
--	g30832 = NOT(I40748)
--	I40751 = NOT(g30665)
--	g30833 = NOT(I40751)
--	I40754 = NOT(g30666)
--	g30834 = NOT(I40754)
--	I40757 = NOT(g30667)
--	g30835 = NOT(I40757)
--	I40760 = NOT(g30722)
--	g30836 = NOT(I40760)
--	I40763 = NOT(g30729)
--	g30837 = NOT(I40763)
--	I40766 = NOT(g30737)
--	g30838 = NOT(I40766)
--	I40769 = NOT(g30803)
--	g30839 = NOT(I40769)
--	I40772 = NOT(g30804)
--	g30840 = NOT(I40772)
--	I40775 = NOT(g30807)
--	g30841 = NOT(I40775)
--	I40778 = NOT(g30805)
--	g30842 = NOT(I40778)
--	I40781 = NOT(g30808)
--	g30843 = NOT(I40781)
--	I40784 = NOT(g30813)
--	g30844 = NOT(I40784)
--	I40787 = NOT(g30809)
--	g30845 = NOT(I40787)
--	I40790 = NOT(g30814)
--	g30846 = NOT(I40790)
--	I40793 = NOT(g30821)
--	g30847 = NOT(I40793)
--	I40796 = NOT(g30829)
--	g30848 = NOT(I40796)
--	I40799 = NOT(g30723)
--	g30849 = NOT(I40799)
--	I40802 = NOT(g30730)
--	g30850 = NOT(I40802)
--	I40805 = NOT(g30767)
--	g30851 = NOT(I40805)
--	I40808 = NOT(g30769)
--	g30852 = NOT(I40808)
--	I40811 = NOT(g30772)
--	g30853 = NOT(I40811)
--	I40814 = NOT(g30731)
--	g30854 = NOT(I40814)
--	I40817 = NOT(g30738)
--	g30855 = NOT(I40817)
--	I40820 = NOT(g30745)
--	g30856 = NOT(I40820)
--	I40823 = NOT(g30806)
--	g30857 = NOT(I40823)
--	I40826 = NOT(g30810)
--	g30858 = NOT(I40826)
--	I40829 = NOT(g30815)
--	g30859 = NOT(I40829)
--	I40832 = NOT(g30811)
--	g30860 = NOT(I40832)
--	I40835 = NOT(g30816)
--	g30861 = NOT(I40835)
--	I40838 = NOT(g30822)
--	g30862 = NOT(I40838)
--	I40841 = NOT(g30817)
--	g30863 = NOT(I40841)
--	I40844 = NOT(g30823)
--	g30864 = NOT(I40844)
--	I40847 = NOT(g30830)
--	g30865 = NOT(I40847)
--	I40850 = NOT(g30724)
--	g30866 = NOT(I40850)
--	I40853 = NOT(g30732)
--	g30867 = NOT(I40853)
--	I40856 = NOT(g30739)
--	g30868 = NOT(I40856)
--	I40859 = NOT(g30770)
--	g30869 = NOT(I40859)
--	I40862 = NOT(g30773)
--	g30870 = NOT(I40862)
--	I40865 = NOT(g30776)
--	g30871 = NOT(I40865)
--	I40868 = NOT(g30740)
--	g30872 = NOT(I40868)
--	I40871 = NOT(g30746)
--	g30873 = NOT(I40871)
--	I40874 = NOT(g30751)
--	g30874 = NOT(I40874)
--	I40877 = NOT(g30812)
--	g30875 = NOT(I40877)
--	I40880 = NOT(g30818)
--	g30876 = NOT(I40880)
--	I40883 = NOT(g30824)
--	g30877 = NOT(I40883)
--	I40886 = NOT(g30819)
--	g30878 = NOT(I40886)
--	I40889 = NOT(g30825)
--	g30879 = NOT(I40889)
--	I40892 = NOT(g30831)
--	g30880 = NOT(I40892)
--	I40895 = NOT(g30826)
--	g30881 = NOT(I40895)
--	I40898 = NOT(g30832)
--	g30882 = NOT(I40898)
--	I40901 = NOT(g30725)
--	g30883 = NOT(I40901)
--	I40904 = NOT(g30733)
--	g30884 = NOT(I40904)
--	I40907 = NOT(g30741)
--	g30885 = NOT(I40907)
--	I40910 = NOT(g30747)
--	g30886 = NOT(I40910)
--	I40913 = NOT(g30774)
--	g30887 = NOT(I40913)
--	I40916 = NOT(g30777)
--	g30888 = NOT(I40916)
--	I40919 = NOT(g30781)
--	g30889 = NOT(I40919)
--	I40922 = NOT(g30748)
--	g30890 = NOT(I40922)
--	I40925 = NOT(g30752)
--	g30891 = NOT(I40925)
--	I40928 = NOT(g30756)
--	g30892 = NOT(I40928)
--	I40931 = NOT(g30820)
--	g30893 = NOT(I40931)
--	I40934 = NOT(g30827)
--	g30894 = NOT(I40934)
--	I40937 = NOT(g30833)
--	g30895 = NOT(I40937)
--	I40940 = NOT(g30828)
--	g30896 = NOT(I40940)
--	I40943 = NOT(g30834)
--	g30897 = NOT(I40943)
--	I40946 = NOT(g30726)
--	g30898 = NOT(I40946)
--	I40949 = NOT(g30835)
--	g30899 = NOT(I40949)
--	I40952 = NOT(g30727)
--	g30900 = NOT(I40952)
--	I40955 = NOT(g30734)
--	g30901 = NOT(I40955)
--	I40958 = NOT(g30742)
--	g30902 = NOT(I40958)
--	I40961 = NOT(g30749)
--	g30903 = NOT(I40961)
--	I40964 = NOT(g30753)
--	g30904 = NOT(I40964)
--	I40967 = NOT(g30778)
--	g30905 = NOT(I40967)
--	I40970 = NOT(g30782)
--	g30906 = NOT(I40970)
--	I40973 = NOT(g30784)
--	g30907 = NOT(I40973)
--	I40976 = NOT(g30799)
--	g30908 = NOT(I40976)
--	I40979 = NOT(g30800)
--	g30909 = NOT(I40979)
--	I40982 = NOT(g30802)
--	g30910 = NOT(I40982)
--	I40985 = NOT(g30792)
--	g30911 = NOT(I40985)
--	I40988 = NOT(g30793)
--	g30912 = NOT(I40988)
--	I40991 = NOT(g30794)
--	g30913 = NOT(I40991)
--	I40994 = NOT(g30795)
--	g30914 = NOT(I40994)
--	I40997 = NOT(g30797)
--	g30915 = NOT(I40997)
--	I41024 = NOT(g30765)
--	g30928 = NOT(I41024)
--	I41035 = NOT(g30796)
--	g30937 = NOT(I41035)
--	I41038 = NOT(g30798)
--	g30938 = NOT(I41038)
--	I41041 = NOT(g30801)
--	g30939 = NOT(I41041)
--	I41044 = NOT(g30928)
--	g30940 = NOT(I41044)
--	I41047 = NOT(g30937)
--	g30941 = NOT(I41047)
--	I41050 = NOT(g30938)
--	g30942 = NOT(I41050)
--	I41053 = NOT(g30939)
--	g30943 = NOT(I41053)
--	g30962 = NOT(g30958)
--	g30963 = NOT(g30957)
--	g30964 = NOT(g30961)
--	g30965 = NOT(g30959)
--	g30966 = NOT(g30956)
--	g30967 = NOT(g30954)
--	g30968 = NOT(g30960)
--	g30969 = NOT(g30955)
--	g30971 = NOT(g30970)
--	I41090 = NOT(g30965)
--	g30972 = NOT(I41090)
--	I41093 = NOT(g30964)
--	g30973 = NOT(I41093)
--	I41096 = NOT(g30963)
--	g30974 = NOT(I41096)
--	I41099 = NOT(g30962)
--	g30975 = NOT(I41099)
--	I41102 = NOT(g30969)
--	g30976 = NOT(I41102)
--	I41105 = NOT(g30968)
--	g30977 = NOT(I41105)
--	I41108 = NOT(g30967)
--	g30978 = NOT(I41108)
--	I41111 = NOT(g30966)
--	g30979 = NOT(I41111)
--	I41114 = NOT(g30976)
--	g30980 = NOT(I41114)
--	I41117 = NOT(g30977)
--	g30981 = NOT(I41117)
--	I41120 = NOT(g30978)
--	g30982 = NOT(I41120)
--	I41123 = NOT(g30979)
--	g30983 = NOT(I41123)
--	I41126 = NOT(g30972)
--	g30984 = NOT(I41126)
--	I41129 = NOT(g30973)
--	g30985 = NOT(I41129)
--	I41132 = NOT(g30974)
--	g30986 = NOT(I41132)
--	I41135 = NOT(g30975)
--	g30987 = NOT(I41135)
--	I41138 = NOT(g30971)
--	g30988 = NOT(I41138)
--	I41141 = NOT(g30988)
--	g30989 = NOT(I41141)
--	
--	g5630 = AND(g325, g349)
--	g5649 = AND(g331, g351)
--	g5650 = AND(g325, g364)
--	g5658 = AND(g1012, g1036)
--	g5676 = AND(g337, g353)
--	g5677 = AND(g331, g366)
--	g5678 = AND(g325, g379)
--	g5687 = AND(g1018, g1038)
--	g5688 = AND(g1012, g1051)
--	g5696 = AND(g1706, g1730)
--	g5709 = AND(g337, g368)
--	g5710 = AND(g331, g381)
--	g5711 = AND(g325, g394)
--	g5728 = AND(g1024, g1040)
--	g5729 = AND(g1018, g1053)
--	g5730 = AND(g1012, g1066)
--	g5739 = AND(g1712, g1732)
--	g5740 = AND(g1706, g1745)
--	g5748 = AND(g2400, g2424)
--	g5757 = AND(g337, g383)
--	g5758 = AND(g331, g396)
--	g5767 = AND(g1024, g1055)
--	g5768 = AND(g1018, g1068)
--	g5769 = AND(g1012, g1081)
--	g5786 = AND(g1718, g1734)
--	g5787 = AND(g1712, g1747)
--	g5788 = AND(g1706, g1760)
--	g5797 = AND(g2406, g2426)
--	g5798 = AND(g2400, g2439)
--	g5807 = AND(g337, g324)
--	g5816 = AND(g1024, g1070)
--	g5817 = AND(g1018, g1083)
--	g5826 = AND(g1718, g1749)
--	g5827 = AND(g1712, g1762)
--	g5828 = AND(g1706, g1775)
--	g5845 = AND(g2412, g2428)
--	g5846 = AND(g2406, g2441)
--	g5847 = AND(g2400, g2454)
--	g5863 = AND(g1024, g1011)
--	g5872 = AND(g1718, g1764)
--	g5873 = AND(g1712, g1777)
--	g5882 = AND(g2412, g2443)
--	g5883 = AND(g2406, g2456)
--	g5884 = AND(g2400, g2469)
--	g5910 = AND(g1718, g1705)
--	g5919 = AND(g2412, g2458)
--	g5920 = AND(g2406, g2471)
--	g5949 = AND(g2412, g2399)
--	g8327 = AND(g3254, g219)
--	g8328 = AND(g6314, g225)
--	g8329 = AND(g6232, g231)
--	g8339 = AND(g6519, g903)
--	g8340 = AND(g6369, g909)
--	g8350 = AND(g6574, g1594)
--	g8385 = AND(g3254, g228)
--	g8386 = AND(g6314, g234)
--	g8387 = AND(g6232, g240)
--	g8394 = AND(g3410, g906)
--	g8395 = AND(g6519, g912)
--	g8396 = AND(g6369, g918)
--	g8406 = AND(g6783, g1597)
--	g8407 = AND(g6574, g1603)
--	g8417 = AND(g6838, g2288)
--	g8431 = AND(g3254, g237)
--	g8432 = AND(g6314, g243)
--	g8433 = AND(g6232, g249)
--	g8437 = AND(g3410, g915)
--	g8438 = AND(g6519, g921)
--	g8439 = AND(g6369, g927)
--	g8446 = AND(g3566, g1600)
--	g8447 = AND(g6783, g1606)
--	g8448 = AND(g6574, g1612)
--	g8458 = AND(g7085, g2291)
--	g8459 = AND(g6838, g2297)
--	g8463 = AND(g3254, g246)
--	g8464 = AND(g6314, g252)
--	g8465 = AND(g6232, g258)
--	g8466 = AND(g3410, g924)
--	g8467 = AND(g6519, g930)
--	g8468 = AND(g6369, g936)
--	g8472 = AND(g3566, g1609)
--	g8473 = AND(g6783, g1615)
--	g8474 = AND(g6574, g1621)
--	g8481 = AND(g3722, g2294)
--	g8482 = AND(g7085, g2300)
--	g8483 = AND(g6838, g2306)
--	g8484 = AND(g6232, g186)
--	g8485 = AND(g3254, g255)
--	g8486 = AND(g6314, g261)
--	g8487 = AND(g6232, g267)
--	g8488 = AND(g3410, g933)
--	g8489 = AND(g6519, g939)
--	g8490 = AND(g6369, g945)
--	g8491 = AND(g3566, g1618)
--	g8492 = AND(g6783, g1624)
--	g8493 = AND(g6574, g1630)
--	g8497 = AND(g3722, g2303)
--	g8498 = AND(g7085, g2309)
--	g8499 = AND(g6838, g2315)
--	g8500 = AND(g6314, g189)
--	g8501 = AND(g6232, g195)
--	g8502 = AND(g3254, g264)
--	g8503 = AND(g6314, g270)
--	g8504 = AND(g6369, g873)
--	g8505 = AND(g3410, g942)
--	g8506 = AND(g6519, g948)
--	g8507 = AND(g6369, g954)
--	g8508 = AND(g3566, g1627)
--	g8509 = AND(g6783, g1633)
--	g8510 = AND(g6574, g1639)
--	g8511 = AND(g3722, g2312)
--	g8512 = AND(g7085, g2318)
--	g8513 = AND(g6838, g2324)
--	g8515 = AND(g3254, g192)
--	g8516 = AND(g6314, g198)
--	g8517 = AND(g6232, g204)
--	g8518 = AND(g3254, g273)
--	g8519 = AND(g6519, g876)
--	g8520 = AND(g6369, g882)
--	g8521 = AND(g3410, g951)
--	g8522 = AND(g6519, g957)
--	g8523 = AND(g6574, g1567)
--	g8524 = AND(g3566, g1636)
--	g8525 = AND(g6783, g1642)
--	g8526 = AND(g6574, g1648)
--	g8527 = AND(g3722, g2321)
--	g8528 = AND(g7085, g2327)
--	g8529 = AND(g6838, g2333)
--	g8531 = AND(g3254, g201)
--	g8532 = AND(g6314, g207)
--	g8534 = AND(g3410, g879)
--	g8535 = AND(g6519, g885)
--	g8536 = AND(g6369, g891)
--	g8537 = AND(g3410, g960)
--	g8538 = AND(g6783, g1570)
--	g8539 = AND(g6574, g1576)
--	g8540 = AND(g3566, g1645)
--	g8541 = AND(g6783, g1651)
--	g8542 = AND(g6838, g2261)
--	g8543 = AND(g3722, g2330)
--	g8544 = AND(g7085, g2336)
--	g8545 = AND(g6838, g2342)
--	g8546 = AND(g3254, g210)
--	g8548 = AND(g3410, g888)
--	g8549 = AND(g6519, g894)
--	g8551 = AND(g3566, g1573)
--	g8552 = AND(g6783, g1579)
--	g8553 = AND(g6574, g1585)
--	g8554 = AND(g3566, g1654)
--	g8555 = AND(g7085, g2264)
--	g8556 = AND(g6838, g2270)
--	g8557 = AND(g3722, g2339)
--	g8558 = AND(g7085, g2345)
--	g8559 = AND(g3410, g897)
--	g8561 = AND(g3566, g1582)
--	g8562 = AND(g6783, g1588)
--	g8564 = AND(g3722, g2267)
--	g8565 = AND(g7085, g2273)
--	g8566 = AND(g6838, g2279)
--	g8567 = AND(g3722, g2348)
--	g8570 = AND(g3566, g1591)
--	g8572 = AND(g3722, g2276)
--	g8573 = AND(g7085, g2282)
--	g8576 = AND(g3722, g2285)
--	g8601 = AND(g6643, g7153)
--	g8612 = AND(g3338, g6908)
--	g8613 = AND(g6945, g7349)
--	g8621 = AND(g6486, g6672)
--	g8625 = AND(g3494, g7158)
--	g8626 = AND(g7195, g7479)
--	g8631 = AND(g6751, g6974)
--	g8635 = AND(g3650, g7354)
--	g8636 = AND(g7391, g7535)
--	g8650 = AND(g7053, g7224)
--	g8654 = AND(g3806, g7484)
--	g8666 = AND(g7303, g7420)
--	g8676 = AND(g6643, g7838)
--	g8687 = AND(g3338, g7827)
--	g8688 = AND(g6945, g7858)
--	g8703 = AND(g6486, g7819)
--	g8704 = AND(g6643, g7996)
--	g8705 = AND(g3494, g7842)
--	g8706 = AND(g7195, g7888)
--	g8717 = AND(g3338, g7953)
--	g8722 = AND(g6751, g7830)
--	g8723 = AND(g6945, g8071)
--	g8724 = AND(g3650, g7862)
--	g8725 = AND(g7391, g7912)
--	g8751 = AND(g6486, g7906)
--	g8755 = AND(g3494, g8004)
--	g8760 = AND(g7053, g7845)
--	g8761 = AND(g7195, g8156)
--	g8762 = AND(g3806, g7892)
--	g8774 = AND(g6751, g7958)
--	g8778 = AND(g3650, g8079)
--	g8783 = AND(g7303, g7865)
--	g8784 = AND(g7391, g8242)
--	g8797 = AND(g7053, g8009)
--	g8801 = AND(g3806, g8164)
--	g8816 = AND(g7303, g8084)
--	g8841 = AND(g6486, g490)
--	g8842 = AND(g6512, g5508)
--	g8861 = AND(g6643, g493)
--	g8868 = AND(g6751, g1177)
--	g8869 = AND(g6776, g5552)
--	g8892 = AND(g3338, g496)
--	g8899 = AND(g6945, g1180)
--	g8906 = AND(g7053, g1871)
--	g8907 = AND(g7078, g5598)
--	g8932 = AND(g3494, g1183)
--	g8939 = AND(g7195, g1874)
--	g8946 = AND(g7303, g2565)
--	g8947 = AND(g7328, g5615)
--	g8972 = AND(g3650, g1877)
--	g8979 = AND(g7391, g2568)
--	g9004 = AND(g3806, g2571)
--	g9009 = AND(g6486, g565)
--	g9026 = AND(g5438, g7610)
--	g9033 = AND(g6643, g567)
--	g9034 = AND(g6751, g1251)
--	g9047 = AND(g6448, g7616)
--	g9048 = AND(g3338, g489)
--	g9049 = AND(g5473, g7619)
--	g9056 = AND(g6945, g1253)
--	g9057 = AND(g7053, g1945)
--	g9061 = AND(g3306, g7623)
--	g9062 = AND(g5438, g7626)
--	g9063 = AND(g5438, g7629)
--	g9064 = AND(g6713, g7632)
--	g9065 = AND(g3494, g1176)
--	g9066 = AND(g5512, g7635)
--	g9073 = AND(g7195, g1947)
--	g9074 = AND(g7303, g2639)
--	g9075 = AND(g6448, g7643)
--	g9076 = AND(g5438, g7646)
--	g9077 = AND(g6448, g7649)
--	g9078 = AND(g3462, g7652)
--	g9079 = AND(g5473, g7655)
--	g9080 = AND(g5473, g7658)
--	g9081 = AND(g7015, g7661)
--	g9082 = AND(g3650, g1870)
--	g9083 = AND(g5556, g7664)
--	g9090 = AND(g7391, g2641)
--	g9091 = AND(g3306, g7670)
--	g9092 = AND(g6448, g7673)
--	g9093 = AND(g3306, g7676)
--	g9094 = AND(g6713, g7679)
--	g9095 = AND(g5473, g7682)
--	g9096 = AND(g6713, g7685)
--	g9097 = AND(g3618, g7688)
--	g9098 = AND(g5512, g7691)
--	g9099 = AND(g5512, g7694)
--	g9100 = AND(g7265, g7697)
--	g9101 = AND(g3806, g2564)
--	g9102 = AND(g3306, g7703)
--	g9103 = AND(g3462, g7706)
--	g9104 = AND(g6713, g7709)
--	g9105 = AND(g3462, g7712)
--	g9106 = AND(g7015, g7715)
--	g9107 = AND(g5512, g7718)
--	g9108 = AND(g7015, g7721)
--	g9109 = AND(g3774, g7724)
--	g9110 = AND(g5556, g7727)
--	g9111 = AND(g5556, g7730)
--	g9112 = AND(g3462, g7733)
--	g9113 = AND(g3618, g7736)
--	g9114 = AND(g7015, g7739)
--	g9115 = AND(g3618, g7742)
--	g9116 = AND(g7265, g7745)
--	g9117 = AND(g5556, g7748)
--	g9118 = AND(g7265, g7751)
--	g9119 = AND(g5438, g7754)
--	g9120 = AND(g3618, g7757)
--	g9121 = AND(g3774, g7760)
--	g9122 = AND(g7265, g7763)
--	g9123 = AND(g3774, g7766)
--	g9124 = AND(g6448, g7769)
--	g9125 = AND(g5473, g7776)
--	g9126 = AND(g3774, g7779)
--	g9127 = AND(g3306, g7782)
--	g9131 = AND(g6713, g7785)
--	g9132 = AND(g5512, g7792)
--	g9133 = AND(g3462, g7796)
--	g9137 = AND(g7015, g7799)
--	g9138 = AND(g5556, g7806)
--	g9139 = AND(g3618, g7809)
--	g9143 = AND(g7265, g7812)
--	g9145 = AND(g3774, g7823)
--	g9241 = AND(g6232, g7950)
--	g9301 = AND(g6314, g7990)
--	g9302 = AND(g6232, g7993)
--	g9319 = AND(g6369, g8001)
--	g9364 = AND(g3254, g8053)
--	g9365 = AND(g6314, g8056)
--	g9366 = AND(g6232, g8059)
--	g9367 = AND(g6232, g8062)
--	g9382 = AND(g6519, g8065)
--	g9383 = AND(g6369, g8068)
--	g9400 = AND(g6574, g8076)
--	g9438 = AND(g3254, g8123)
--	g9439 = AND(g6314, g8126)
--	g9440 = AND(g6232, g8129)
--	g9441 = AND(g6314, g8132)
--	g9442 = AND(g6232, g8135)
--	g9461 = AND(g3410, g8138)
--	g9462 = AND(g6519, g8141)
--	g9463 = AND(g6369, g8144)
--	g9464 = AND(g6369, g8147)
--	g9479 = AND(g6783, g8150)
--	g9480 = AND(g6574, g8153)
--	g9497 = AND(g6838, g8161)
--	g9518 = AND(g3254, g8191)
--	g9519 = AND(g6314, g8194)
--	g9520 = AND(g6232, g8197)
--	g9521 = AND(g3254, g8200)
--	g9522 = AND(g6314, g8203)
--	g9523 = AND(g6232, g8206)
--	g9534 = AND(g7772, g6135, g538)
--	g9580 = AND(g3410, g8209)
--	g9581 = AND(g6519, g8212)
--	g9582 = AND(g6369, g8215)
--	g9583 = AND(g6519, g8218)
--	g9584 = AND(g6369, g8221)
--	g9603 = AND(g3566, g8224)
--	g9604 = AND(g6783, g8227)
--	g9605 = AND(g6574, g8230)
--	g9606 = AND(g6574, g8233)
--	g9621 = AND(g7085, g8236)
--	g9622 = AND(g6838, g8239)
--	g9630 = AND(g3254, g3922)
--	g9631 = AND(g6314, g3925)
--	g9632 = AND(g6232, g3928)
--	g9633 = AND(g3254, g3931)
--	g9634 = AND(g6314, g3934)
--	g9635 = AND(g6232, g3937)
--	I16735 = AND(g5856, g4338, g4339, g5141)
--	I16736 = AND(g5713, g5958, g4735, g4736)
--	g9636 = AND(I16735, I16736)
--	g9639 = AND(g5438, g408)
--	g9647 = AND(g6678, g3942)
--	g9648 = AND(g6678, g3945)
--	g9660 = AND(g3410, g3948)
--	g9661 = AND(g6519, g3951)
--	g9662 = AND(g6369, g3954)
--	g9663 = AND(g3410, g3957)
--	g9664 = AND(g6519, g3960)
--	g9665 = AND(g6369, g3963)
--	g9676 = AND(g7788, g6145, g1224)
--	g9722 = AND(g3566, g3966)
--	g9723 = AND(g6783, g3969)
--	g9724 = AND(g6574, g3972)
--	g9725 = AND(g6783, g3975)
--	g9726 = AND(g6574, g3978)
--	g9745 = AND(g3722, g3981)
--	g9746 = AND(g7085, g3984)
--	g9747 = AND(g6838, g3987)
--	g9748 = AND(g6838, g3990)
--	g9759 = AND(g3254, g4000)
--	g9760 = AND(g6314, g4003)
--	g9761 = AND(g6232, g4006)
--	g9762 = AND(g3254, g4009)
--	g9763 = AND(g6314, g4012)
--	g9764 = AND(g6448, g411)
--	g9765 = AND(g5438, g417)
--	g9766 = AND(g5438, g4017)
--	g9773 = AND(g6912, g4020)
--	g9774 = AND(g6678, g4023)
--	g9775 = AND(g6912, g4026)
--	g9776 = AND(g3410, g4029)
--	g9777 = AND(g6519, g4032)
--	g9778 = AND(g6369, g4035)
--	g9779 = AND(g3410, g4038)
--	g9780 = AND(g6519, g4041)
--	g9781 = AND(g6369, g4044)
--	I16826 = AND(g5903, g4507, g4508, g5234)
--	I16827 = AND(g5771, g5987, g4911, g4912)
--	g9782 = AND(I16826, I16827)
--	g9785 = AND(g5473, g1095)
--	g9793 = AND(g6980, g4049)
--	g9794 = AND(g6980, g4052)
--	g9806 = AND(g3566, g4055)
--	g9807 = AND(g6783, g4058)
--	g9808 = AND(g6574, g4061)
--	g9809 = AND(g3566, g4064)
--	g9810 = AND(g6783, g4067)
--	g9811 = AND(g6574, g4070)
--	g9822 = AND(g7802, g6166, g1918)
--	g9868 = AND(g3722, g4073)
--	g9869 = AND(g7085, g4076)
--	g9870 = AND(g6838, g4079)
--	g9871 = AND(g7085, g4082)
--	g9872 = AND(g6838, g4085)
--	g9887 = AND(g6232, g4095)
--	g9888 = AND(g3254, g4098)
--	g9889 = AND(g6314, g4101)
--	g9890 = AND(g6232, g4104)
--	g9891 = AND(g3254, g4107)
--	g9892 = AND(g3306, g414)
--	g9893 = AND(g6448, g420)
--	g9894 = AND(g6448, g4112)
--	g9901 = AND(g3366, g4115)
--	g9902 = AND(g6912, g4118)
--	g9903 = AND(g6678, g4121)
--	g9904 = AND(g3366, g4124)
--	g9905 = AND(g3410, g4127)
--	g9906 = AND(g6519, g4130)
--	g9907 = AND(g6369, g4133)
--	g9908 = AND(g3410, g4136)
--	g9909 = AND(g6519, g4139)
--	g9910 = AND(g6713, g1098)
--	g9911 = AND(g5473, g1104)
--	g9912 = AND(g5473, g4144)
--	g9919 = AND(g7162, g4147)
--	g9920 = AND(g6980, g4150)
--	g9921 = AND(g7162, g4153)
--	g9922 = AND(g3566, g4156)
--	g9923 = AND(g6783, g4159)
--	g9924 = AND(g6574, g4162)
--	g9925 = AND(g3566, g4165)
--	g9926 = AND(g6783, g4168)
--	g9927 = AND(g6574, g4171)
--	I16930 = AND(g5942, g4683, g4684, g5297)
--	I16931 = AND(g5830, g6024, g5070, g5071)
--	g9928 = AND(I16930, I16931)
--	g9931 = AND(g5512, g1789)
--	g9939 = AND(g7230, g4176)
--	g9940 = AND(g7230, g4179)
--	g9952 = AND(g3722, g4182)
--	g9953 = AND(g7085, g4185)
--	g9954 = AND(g6838, g4188)
--	g9955 = AND(g3722, g4191)
--	g9956 = AND(g7085, g4194)
--	g9957 = AND(g6838, g4197)
--	g9968 = AND(g7815, g6193, g2612)
--	g10007 = AND(g6314, g4205)
--	g10008 = AND(g6232, g4208)
--	g10009 = AND(g3254, g4211)
--	g10010 = AND(g6314, g4214)
--	g10011 = AND(g5438, g4217)
--	g10012 = AND(g3306, g423)
--	g10013 = AND(g3306, g4221)
--	g10014 = AND(g5438, g429)
--	g10024 = AND(g3398, g6912)
--	g10035 = AND(g3366, g4225)
--	g10036 = AND(g6912, g4228)
--	g10037 = AND(g6678, g4231)
--	g10041 = AND(g6369, g4234)
--	g10042 = AND(g3410, g4237)
--	g10043 = AND(g6519, g4240)
--	g10044 = AND(g6369, g4243)
--	g10045 = AND(g3410, g4246)
--	g10046 = AND(g3462, g1101)
--	g10047 = AND(g6713, g1107)
--	g10048 = AND(g6713, g4251)
--	g10055 = AND(g3522, g4254)
--	g10056 = AND(g7162, g4257)
--	g10057 = AND(g6980, g4260)
--	g10058 = AND(g3522, g4263)
--	g10059 = AND(g3566, g4266)
--	g10060 = AND(g6783, g4269)
--	g10061 = AND(g6574, g4272)
--	g10062 = AND(g3566, g4275)
--	g10063 = AND(g6783, g4278)
--	g10064 = AND(g7015, g1792)
--	g10065 = AND(g5512, g1798)
--	g10066 = AND(g5512, g4283)
--	g10073 = AND(g7358, g4286)
--	g10074 = AND(g7230, g4289)
--	g10075 = AND(g7358, g4292)
--	g10076 = AND(g3722, g4295)
--	g10077 = AND(g7085, g4298)
--	g10078 = AND(g6838, g4301)
--	g10079 = AND(g3722, g4304)
--	g10080 = AND(g7085, g4307)
--	g10081 = AND(g6838, g4310)
--	I17042 = AND(g5976, g4860, g4861, g5334)
--	I17043 = AND(g5886, g6040, g5199, g5200)
--	g10082 = AND(I17042, I17043)
--	g10085 = AND(g5556, g2483)
--	g10093 = AND(g7426, g4315)
--	g10094 = AND(g7426, g4318)
--	g10101 = AND(g3254, g4329)
--	g10102 = AND(g6314, g4332)
--	g10103 = AND(g3254, g4335)
--	g10104 = AND(g6448, g4340)
--	g10105 = AND(g5438, g4343)
--	g10106 = AND(g6448, g432)
--	g10107 = AND(g5438, g438)
--	g10108 = AND(g6486, g569)
--	g10112 = AND(g3366, g4348)
--	g10113 = AND(g6912, g4351)
--	g10114 = AND(g6678, g4354)
--	g10115 = AND(g6678, g4357)
--	g10116 = AND(g6519, g4360)
--	g10117 = AND(g6369, g4363)
--	g10118 = AND(g3410, g4366)
--	g10119 = AND(g6519, g4369)
--	g10120 = AND(g5473, g4372)
--	g10121 = AND(g3462, g1110)
--	g10122 = AND(g3462, g4376)
--	g10123 = AND(g5473, g1116)
--	g10133 = AND(g3554, g7162)
--	g10144 = AND(g3522, g4380)
--	g10145 = AND(g7162, g4383)
--	g10146 = AND(g6980, g4386)
--	g10150 = AND(g6574, g4389)
--	g10151 = AND(g3566, g4392)
--	g10152 = AND(g6783, g4395)
--	g10153 = AND(g6574, g4398)
--	g10154 = AND(g3566, g4401)
--	g10155 = AND(g3618, g1795)
--	g10156 = AND(g7015, g1801)
--	g10157 = AND(g7015, g4406)
--	g10164 = AND(g3678, g4409)
--	g10165 = AND(g7358, g4412)
--	g10166 = AND(g7230, g4415)
--	g10167 = AND(g3678, g4418)
--	g10168 = AND(g3722, g4421)
--	g10169 = AND(g7085, g4424)
--	g10170 = AND(g6838, g4427)
--	g10171 = AND(g3722, g4430)
--	g10172 = AND(g7085, g4433)
--	g10173 = AND(g7265, g2486)
--	g10174 = AND(g5556, g2492)
--	g10175 = AND(g5556, g4438)
--	g10182 = AND(g7488, g4441)
--	g10183 = AND(g7426, g4444)
--	g10184 = AND(g7488, g4447)
--	I17156 = AND(g6898, g2998, g6901, g3002)
--	g10186 = AND(g3013, g7466, g3024, I17156)
--	g10192 = AND(g3254, g4453)
--	g10193 = AND(g3306, g4465)
--	g10194 = AND(g6448, g4468)
--	g10195 = AND(g5438, g4471)
--	g10196 = AND(g3306, g435)
--	g10197 = AND(g6448, g441)
--	g10198 = AND(g6643, g571)
--	g10199 = AND(g6486, g4476)
--	g10200 = AND(g6486, g587)
--	g10201 = AND(g3366, g4480)
--	g10202 = AND(g6912, g4483)
--	g10203 = AND(g6678, g4486)
--	g10204 = AND(g6912, g4489)
--	g10205 = AND(g6678, g4492)
--	g10206 = AND(g3410, g4498)
--	g10207 = AND(g6519, g4501)
--	g10208 = AND(g3410, g4504)
--	g10209 = AND(g6713, g4509)
--	g10210 = AND(g5473, g4512)
--	g10211 = AND(g6713, g1119)
--	g10212 = AND(g5473, g1125)
--	g10213 = AND(g6751, g1255)
--	g10217 = AND(g3522, g4517)
--	g10218 = AND(g7162, g4520)
--	g10219 = AND(g6980, g4523)
--	g10220 = AND(g6980, g4526)
--	g10221 = AND(g6783, g4529)
--	g10222 = AND(g6574, g4532)
--	g10223 = AND(g3566, g4535)
--	g10224 = AND(g6783, g4538)
--	g10225 = AND(g5512, g4541)
--	g10226 = AND(g3618, g1804)
--	g10227 = AND(g3618, g4545)
--	g10228 = AND(g5512, g1810)
--	g10238 = AND(g3710, g7358)
--	g10249 = AND(g3678, g4549)
--	g10250 = AND(g7358, g4552)
--	g10251 = AND(g7230, g4555)
--	g10255 = AND(g6838, g4558)
--	g10256 = AND(g3722, g4561)
--	g10257 = AND(g7085, g4564)
--	g10258 = AND(g6838, g4567)
--	g10259 = AND(g3722, g4570)
--	g10260 = AND(g3774, g2489)
--	g10261 = AND(g7265, g2495)
--	g10262 = AND(g7265, g4575)
--	g10269 = AND(g3834, g4578)
--	g10270 = AND(g7488, g4581)
--	g10271 = AND(g7426, g4584)
--	g10272 = AND(g3834, g4587)
--	g10279 = AND(g3306, g4592)
--	g10280 = AND(g6448, g4595)
--	g10281 = AND(g5438, g4598)
--	g10282 = AND(g3306, g444)
--	g10283 = AND(g3338, g573)
--	g10284 = AND(g6643, g4603)
--	g10285 = AND(g6486, g4606)
--	g10286 = AND(g6643, g590)
--	g10287 = AND(g6486, g596)
--	g10288 = AND(g3366, g4611)
--	g10289 = AND(g6912, g4614)
--	g10290 = AND(g6678, g4617)
--	g10291 = AND(g3366, g4620)
--	g10292 = AND(g6912, g4623)
--	g10293 = AND(g6678, g4626)
--	g10294 = AND(g3410, g4629)
--	g10295 = AND(g3462, g4641)
--	g10296 = AND(g6713, g4644)
--	g10297 = AND(g5473, g4647)
--	g10298 = AND(g3462, g1122)
--	g10299 = AND(g6713, g1128)
--	g10300 = AND(g6945, g1257)
--	g10301 = AND(g6751, g4652)
--	g10302 = AND(g6751, g1273)
--	g10303 = AND(g3522, g4656)
--	g10304 = AND(g7162, g4659)
--	g10305 = AND(g6980, g4662)
--	g10306 = AND(g7162, g4665)
--	g10307 = AND(g6980, g4668)
--	g10308 = AND(g3566, g4674)
--	g10309 = AND(g6783, g4677)
--	g10310 = AND(g3566, g4680)
--	g10311 = AND(g7015, g4685)
--	g10312 = AND(g5512, g4688)
--	g10313 = AND(g7015, g1813)
--	g10314 = AND(g5512, g1819)
--	g10315 = AND(g7053, g1949)
--	g10319 = AND(g3678, g4693)
--	g10320 = AND(g7358, g4696)
--	g10321 = AND(g7230, g4699)
--	g10322 = AND(g7230, g4702)
--	g10323 = AND(g7085, g4705)
--	g10324 = AND(g6838, g4708)
--	g10325 = AND(g3722, g4711)
--	g10326 = AND(g7085, g4714)
--	g10327 = AND(g5556, g4717)
--	g10328 = AND(g3774, g2498)
--	g10329 = AND(g3774, g4721)
--	g10330 = AND(g5556, g2504)
--	g10340 = AND(g3866, g7488)
--	g10351 = AND(g3834, g4725)
--	g10352 = AND(g7488, g4728)
--	g10353 = AND(g7426, g4731)
--	g10360 = AND(g3306, g4737)
--	g10361 = AND(g6448, g4740)
--	g10362 = AND(g3338, g4743)
--	g10363 = AND(g6643, g4746)
--	g10364 = AND(g6486, g4749)
--	g10365 = AND(g3338, g593)
--	g10366 = AND(g6643, g599)
--	g10367 = AND(g3366, g4754)
--	g10368 = AND(g6912, g4757)
--	g10369 = AND(g6678, g4760)
--	g10370 = AND(g3366, g4763)
--	g10371 = AND(g6912, g4766)
--	g10372 = AND(g3462, g4769)
--	g10373 = AND(g6713, g4772)
--	g10374 = AND(g5473, g4775)
--	g10375 = AND(g3462, g1131)
--	g10376 = AND(g3494, g1259)
--	g10377 = AND(g6945, g4780)
--	g10378 = AND(g6751, g4783)
--	g10379 = AND(g6945, g1276)
--	g10380 = AND(g6751, g1282)
--	g10381 = AND(g3522, g4788)
--	g10382 = AND(g7162, g4791)
--	g10383 = AND(g6980, g4794)
--	g10384 = AND(g3522, g4797)
--	g10385 = AND(g7162, g4800)
--	g10386 = AND(g6980, g4803)
--	g10387 = AND(g3566, g4806)
--	g10388 = AND(g3618, g4818)
--	g10389 = AND(g7015, g4821)
--	g10390 = AND(g5512, g4824)
--	g10391 = AND(g3618, g1816)
--	g10392 = AND(g7015, g1822)
--	g10393 = AND(g7195, g1951)
--	g10394 = AND(g7053, g4829)
--	g10395 = AND(g7053, g1967)
--	g10396 = AND(g3678, g4833)
--	g10397 = AND(g7358, g4836)
--	g10398 = AND(g7230, g4839)
--	g10399 = AND(g7358, g4842)
--	g10400 = AND(g7230, g4845)
--	g10401 = AND(g3722, g4851)
--	g10402 = AND(g7085, g4854)
--	g10403 = AND(g3722, g4857)
--	g10404 = AND(g7265, g4862)
--	g10405 = AND(g5556, g4865)
--	g10406 = AND(g7265, g2507)
--	g10407 = AND(g5556, g2513)
--	g10408 = AND(g7303, g2643)
--	g10412 = AND(g3834, g4870)
--	g10413 = AND(g7488, g4873)
--	g10414 = AND(g7426, g4876)
--	g10415 = AND(g7426, g4879)
--	g10422 = AND(g3306, g4882)
--	g10423 = AND(g5438, g4885)
--	g10430 = AND(g3338, g4888)
--	g10431 = AND(g6643, g4891)
--	g10432 = AND(g6486, g4894)
--	g10433 = AND(g3338, g602)
--	g10434 = AND(g6486, g605)
--	g10435 = AND(g3366, g4899)
--	g10436 = AND(g6912, g4902)
--	g10437 = AND(g6678, g4905)
--	g10438 = AND(g3366, g4908)
--	g10439 = AND(g3462, g4913)
--	g10440 = AND(g6713, g4916)
--	g10441 = AND(g3494, g4919)
--	g10442 = AND(g6945, g4922)
--	g10443 = AND(g6751, g4925)
--	g10444 = AND(g3494, g1279)
--	g10445 = AND(g6945, g1285)
--	g10446 = AND(g3522, g4930)
--	g10447 = AND(g7162, g4933)
--	g10448 = AND(g6980, g4936)
--	g10449 = AND(g3522, g4939)
--	g10450 = AND(g7162, g4942)
--	g10451 = AND(g3618, g4945)
--	g10452 = AND(g7015, g4948)
--	g10453 = AND(g5512, g4951)
--	g10454 = AND(g3618, g1825)
--	g10455 = AND(g3650, g1953)
--	g10456 = AND(g7195, g4956)
--	g10457 = AND(g7053, g4959)
--	g10458 = AND(g7195, g1970)
--	g10459 = AND(g7053, g1976)
--	g10460 = AND(g3678, g4964)
--	g10461 = AND(g7358, g4967)
--	g10462 = AND(g7230, g4970)
--	g10463 = AND(g3678, g4973)
--	g10464 = AND(g7358, g4976)
--	g10465 = AND(g7230, g4979)
--	g10466 = AND(g3722, g4982)
--	g10467 = AND(g3774, g4994)
--	g10468 = AND(g7265, g4997)
--	g10469 = AND(g5556, g5000)
--	g10470 = AND(g3774, g2510)
--	g10471 = AND(g7265, g2516)
--	g10472 = AND(g7391, g2645)
--	g10473 = AND(g7303, g5005)
--	g10474 = AND(g7303, g2661)
--	g10475 = AND(g3834, g5009)
--	g10476 = AND(g7488, g5012)
--	g10477 = AND(g7426, g5015)
--	g10478 = AND(g7488, g5018)
--	g10479 = AND(g7426, g5021)
--	I17429 = AND(g6901, g7338, g7146)
--	g10480 = AND(g7466, g7342, I17429)
--	g10485 = AND(g6448, g5024)
--	g10492 = AND(g3338, g5027)
--	g10493 = AND(g6643, g5030)
--	g10494 = AND(g6643, g608)
--	g10495 = AND(g6486, g614)
--	g10496 = AND(g3366, g5035)
--	g10497 = AND(g6912, g5038)
--	g10498 = AND(g3462, g5041)
--	g10499 = AND(g5473, g5044)
--	g10506 = AND(g3494, g5047)
--	g10507 = AND(g6945, g5050)
--	g10508 = AND(g6751, g5053)
--	g10509 = AND(g3494, g1288)
--	g10510 = AND(g6751, g1291)
--	g10511 = AND(g3522, g5058)
--	g10512 = AND(g7162, g5061)
--	g10513 = AND(g6980, g5064)
--	g10514 = AND(g3522, g5067)
--	g10515 = AND(g3618, g5072)
--	g10516 = AND(g7015, g5075)
--	g10517 = AND(g3650, g5078)
--	g10518 = AND(g7195, g5081)
--	g10519 = AND(g7053, g5084)
--	g10520 = AND(g3650, g1973)
--	g10521 = AND(g7195, g1979)
--	g10522 = AND(g3678, g5089)
--	g10523 = AND(g7358, g5092)
--	g10524 = AND(g7230, g5095)
--	g10525 = AND(g3678, g5098)
--	g10526 = AND(g7358, g5101)
--	g10527 = AND(g3774, g5104)
--	g10528 = AND(g7265, g5107)
--	g10529 = AND(g5556, g5110)
--	g10530 = AND(g3774, g2519)
--	g10531 = AND(g3806, g2647)
--	g10532 = AND(g7391, g5115)
--	g10533 = AND(g7303, g5118)
--	g10534 = AND(g7391, g2664)
--	g10535 = AND(g7303, g2670)
--	g10536 = AND(g3834, g5123)
--	g10537 = AND(g7488, g5126)
--	g10538 = AND(g7426, g5129)
--	g10539 = AND(g3834, g5132)
--	g10540 = AND(g7488, g5135)
--	g10541 = AND(g7426, g5138)
--	g10548 = AND(g3306, g5142)
--	g10555 = AND(g3338, g5145)
--	g10556 = AND(g3338, g611)
--	g10557 = AND(g6643, g617)
--	g10558 = AND(g3366, g5150)
--	g10559 = AND(g6713, g5153)
--	g10566 = AND(g3494, g5156)
--	g10567 = AND(g6945, g5159)
--	g10568 = AND(g6945, g1294)
--	g10569 = AND(g6751, g1300)
--	g10570 = AND(g3522, g5164)
--	g10571 = AND(g7162, g5167)
--	g10572 = AND(g3618, g5170)
--	g10573 = AND(g5512, g5173)
--	g10580 = AND(g3650, g5176)
--	g10581 = AND(g7195, g5179)
--	g10582 = AND(g7053, g5182)
--	g10583 = AND(g3650, g1982)
--	g10584 = AND(g7053, g1985)
--	g10585 = AND(g3678, g5187)
--	g10586 = AND(g7358, g5190)
--	g10587 = AND(g7230, g5193)
--	g10588 = AND(g3678, g5196)
--	g10589 = AND(g3774, g5201)
--	g10590 = AND(g7265, g5204)
--	g10591 = AND(g3806, g5207)
--	g10592 = AND(g7391, g5210)
--	g10593 = AND(g7303, g5213)
--	g10594 = AND(g3806, g2667)
--	g10595 = AND(g7391, g2673)
--	g10596 = AND(g3834, g5218)
--	g10597 = AND(g7488, g5221)
--	g10598 = AND(g7426, g5224)
--	g10599 = AND(g3834, g5227)
--	g10600 = AND(g7488, g5230)
--	g10604 = AND(g3338, g620)
--	g10605 = AND(g3462, g5235)
--	g10612 = AND(g3494, g5238)
--	g10613 = AND(g3494, g1297)
--	g10614 = AND(g6945, g1303)
--	g10615 = AND(g3522, g5243)
--	g10616 = AND(g7015, g5246)
--	g10623 = AND(g3650, g5249)
--	g10624 = AND(g7195, g5252)
--	g10625 = AND(g7195, g1988)
--	g10626 = AND(g7053, g1994)
--	g10627 = AND(g3678, g5257)
--	g10628 = AND(g7358, g5260)
--	g10629 = AND(g3774, g5263)
--	g10630 = AND(g5556, g5266)
--	g10637 = AND(g3806, g5269)
--	g10638 = AND(g7391, g5272)
--	g10639 = AND(g7303, g5275)
--	g10640 = AND(g3806, g2676)
--	g10641 = AND(g7303, g2679)
--	g10642 = AND(g3834, g5280)
--	g10643 = AND(g7488, g5283)
--	g10644 = AND(g7426, g5286)
--	g10645 = AND(g3834, g5289)
--	g10650 = AND(g6678, g5293)
--	g10651 = AND(g3494, g1306)
--	g10652 = AND(g3618, g5298)
--	g10659 = AND(g3650, g5301)
--	g10660 = AND(g3650, g1991)
--	g10661 = AND(g7195, g1997)
--	g10662 = AND(g3678, g5306)
--	g10663 = AND(g7265, g5309)
--	g10670 = AND(g3806, g5312)
--	g10671 = AND(g7391, g5315)
--	g10672 = AND(g7391, g2682)
--	g10673 = AND(g7303, g2688)
--	g10674 = AND(g3834, g5320)
--	g10675 = AND(g7488, g5323)
--	g10678 = AND(g6912, g5327)
--	g10680 = AND(g6980, g5330)
--	g10681 = AND(g3650, g2000)
--	g10682 = AND(g3774, g5335)
--	g10689 = AND(g3806, g5338)
--	g10690 = AND(g3806, g2685)
--	g10691 = AND(g7391, g2691)
--	g10692 = AND(g3834, g5343)
--	g10693 = AND(g7462, g7522, g2924, g7545)
--	g10704 = AND(g3366, g5352)
--	g10707 = AND(g7162, g5355)
--	g10709 = AND(g7230, g5358)
--	g10710 = AND(g3806, g2694)
--	I17599 = AND(g7566, g7583, g7587)
--	g10711 = AND(g7595, g7600, I17599)
--	g10724 = AND(g3522, g5369)
--	g10727 = AND(g7358, g5372)
--	g10729 = AND(g7426, g5375)
--	g10745 = AND(g3678, g5382)
--	g10748 = AND(g7488, g5385)
--	g10764 = AND(g3834, g5391)
--	g11347 = AND(g6232, g213)
--	g11420 = AND(g6314, g216)
--	g11421 = AND(g6232, g222)
--	g11431 = AND(g6369, g900)
--	g11607 = AND(g5871, g8360)
--	g11612 = AND(g5881, g8378)
--	g11637 = AND(g5918, g8427)
--	g11771 = AND(g554, g8622)
--	g11788 = AND(g1240, g8632)
--	g11805 = AND(g6173, g8643)
--	g11814 = AND(g1934, g8651)
--	g11816 = AND(g7869, g8655)
--	g11838 = AND(g6205, g8659)
--	g11847 = AND(g2628, g8667)
--	g11851 = AND(g7849, g8670)
--	g11880 = AND(g6294, g8678)
--	g11885 = AND(g7834, g8684)
--	g11922 = AND(g6431, g8690)
--	g11926 = AND(g8169, g8696)
--	g11966 = AND(g8090, g8708)
--	g11967 = AND(g7967, g8711)
--	g12012 = AND(g8015, g8745)
--	g12069 = AND(g7964, g8763)
--	g12070 = AND(g8018, g8766)
--	g12128 = AND(g7916, g8785)
--	g12129 = AND(g7872, g8788)
--	g12186 = AND(g8093, g8805)
--	g12273 = AND(g8172, g8829)
--	g12274 = AND(g7900, g8832)
--	g12307 = AND(g7919, g8853)
--	g12330 = AND(g8246, g8879)
--	g12331 = AND(g7927, g8882)
--	g12353 = AND(g7852, g8915)
--	g12376 = AND(g7974, g8949)
--	g12419 = AND(g8028, g9006)
--	g12429 = AND(g8101, g9044)
--	g12477 = AND(g7822, g9128)
--	g12494 = AND(g7833, g9134)
--	g12514 = AND(g7848, g9140)
--	g12531 = AND(g7868, g9146)
--	g12650 = AND(g6149, g9290)
--	I19937 = AND(g9507, g9427, g9356, g9293)
--	I19938 = AND(g9232, g9187, g9161, g9150)
--	g12876 = AND(I19937, I19938)
--	g12908 = AND(g7899, g10004)
--	I19971 = AND(g9649, g9569, g9453, g9374)
--	I19972 = AND(g9310, g9248, g9203, g9174)
--	g12916 = AND(I19971, I19972)
--	g12938 = AND(g8179, g10096)
--	I19996 = AND(g9795, g9711, g9595, g9471)
--	I19997 = AND(g9391, g9326, g9264, g9216)
--	g12945 = AND(I19996, I19997)
--	g12966 = AND(g7926, g10189)
--	I20021 = AND(g9941, g9857, g9737, g9613)
--	I20022 = AND(g9488, g9407, g9342, g9277)
--	g12974 = AND(I20021, I20022)
--	g12989 = AND(g8254, g10273)
--	g12990 = AND(g8180, g10276)
--	g13000 = AND(g7973, g10357)
--	g13004 = AND(g10186, g8317)
--	g13009 = AND(g3995, g10416)
--	g13010 = AND(g8255, g10419)
--	g13023 = AND(g8027, g10482)
--	g13031 = AND(g7879, g10542)
--	g13032 = AND(g3996, g10545)
--	g13042 = AND(g8100, g10601)
--	I20100 = AND(g10186, g3018, g3028)
--	g13055 = AND(g7471, g7570, I20100)
--	g13056 = AND(g4092, g10646)
--	I20131 = AND(g8313, g7542, g2888, g7566)
--	I20132 = AND(g2892, g2903, g7595, g2908)
--	g13082 = AND(I20131, I20132)
--	g13110 = AND(g10693, g2883, g7562, g10711)
--	g13247 = AND(g298, g11032)
--	g13266 = AND(g5628, g11088)
--	g13270 = AND(g985, g11102)
--	g13289 = AND(g5647, g11141)
--	g13291 = AND(g5656, g11154)
--	g13295 = AND(g1679, g11170)
--	g13316 = AND(g5675, g11210)
--	g13320 = AND(g5685, g11225)
--	g13322 = AND(g5694, g11240)
--	g13326 = AND(g2373, g11256)
--	g13335 = AND(g5708, g11278)
--	g13340 = AND(g5727, g11294)
--	g13343 = AND(g5737, g11309)
--	g13345 = AND(g5746, g11324)
--	g13355 = AND(g5756, g11355)
--	g13360 = AND(g5766, g11373)
--	g13365 = AND(g5785, g11389)
--	g13368 = AND(g5795, g11404)
--	g13385 = AND(g5815, g11441)
--	g13390 = AND(g5825, g11459)
--	g13395 = AND(g5844, g11475)
--	g13477 = AND(g6016, g12191)
--	g13479 = AND(g6017, g12196)
--	g13480 = AND(g6018, g12197)
--	g13481 = AND(g5864, g11603)
--	g13483 = AND(g6020, g12209)
--	g13484 = AND(g6021, g12210)
--	g13485 = AND(g6022, g12211)
--	g13486 = AND(g6023, g12212)
--	g13487 = AND(g5874, g11608)
--	g13488 = AND(g6025, g12218)
--	g13489 = AND(g6026, g12219)
--	g13490 = AND(g6027, g12220)
--	g13491 = AND(g6028, g12221)
--	g13492 = AND(g2371, g12222)
--	g13493 = AND(g5887, g11613)
--	g13496 = AND(g6032, g12246)
--	g13498 = AND(g6033, g12251)
--	g13499 = AND(g6034, g12252)
--	g13500 = AND(g5911, g11633)
--	g13502 = AND(g6036, g12264)
--	g13503 = AND(g6037, g12265)
--	g13504 = AND(g6038, g12266)
--	g13505 = AND(g6039, g12267)
--	g13506 = AND(g5921, g11638)
--	g13513 = AND(g6043, g12289)
--	g13515 = AND(g6044, g12294)
--	g13516 = AND(g6045, g12295)
--	g13517 = AND(g5950, g11656)
--	g13527 = AND(g6047, g12325)
--	g13609 = AND(g6141, g12456)
--	g13619 = AND(g6162, g12466)
--	g13623 = AND(g5428, g12472)
--	g13625 = AND(g6173, g12476)
--	g13631 = AND(g6189, g12481)
--	g13634 = AND(g12776, g8617)
--	g13636 = AND(g6205, g12493)
--	g13642 = AND(g6221, g12498)
--	g13643 = AND(g5431, g12502)
--	g13645 = AND(g6281, g12504)
--	g13646 = AND(g7772, g12505)
--	g13648 = AND(g6294, g12513)
--	g13654 = AND(g8093, g11791)
--	g13655 = AND(g7540, g12518)
--	g13656 = AND(g12776, g8640)
--	g13671 = AND(g6418, g12521)
--	g13672 = AND(g7788, g12522)
--	g13674 = AND(g6431, g12530)
--	g13675 = AND(g7561, g12532)
--	g13676 = AND(g5434, g12533)
--	g13701 = AND(g6623, g12536)
--	g13702 = AND(g7802, g12537)
--	g13703 = AND(g8018, g11848)
--	g13704 = AND(g7581, g12542)
--	g13705 = AND(g12776, g8673)
--	g13738 = AND(g6887, g12545)
--	g13739 = AND(g7815, g12546)
--	g13740 = AND(g6636, g12547)
--	g13755 = AND(g7347, g12551)
--	g13787 = AND(g7967, g11923)
--	g13788 = AND(g6897, g12553)
--	g13789 = AND(g7140, g12554)
--	g13790 = AND(g7475, g12558)
--	g13796 = AND(g7477, g12559)
--	g13815 = AND(g7139, g12560)
--	g13816 = AND(g7530, g12596)
--	g13818 = AND(g7531, g12597)
--	g13824 = AND(g7533, g12598)
--	g13833 = AND(g7919, g12009)
--	g13834 = AND(g7336, g12599)
--	g13835 = AND(g7461, g12600)
--	g13837 = AND(g7556, g12642)
--	g13839 = AND(g7557, g12643)
--	g13845 = AND(g7559, g12644)
--	g13846 = AND(g7460, g12645)
--	g13847 = AND(g7521, g12646)
--	g13851 = AND(g7579, g12688)
--	g13853 = AND(g7580, g12689)
--	g13854 = AND(g5349, g12690)
--	g13855 = AND(g7541, g12691)
--	g13860 = AND(g7593, g12742)
--	g13862 = AND(g5366, g12743)
--	g13865 = AND(g548, g12748)
--	g13870 = AND(g7582, g12768)
--	g13871 = AND(g7898, g12775)
--	g13878 = AND(g7610, g12782)
--	g13880 = AND(g1234, g12790)
--	g13884 = AND(g7594, g12807)
--	g13892 = AND(g7616, g12815)
--	g13900 = AND(g7619, g12821)
--	g13902 = AND(g1928, g12829)
--	g13904 = AND(g7337, g12843)
--	g13905 = AND(g7925, g12847)
--	g13913 = AND(g7623, g12850)
--	g13914 = AND(g7626, g12851)
--	g13933 = AND(g7632, g12853)
--	g13941 = AND(g7635, g12859)
--	g13943 = AND(g2622, g12867)
--	g13944 = AND(g7141, g12874)
--	g13952 = AND(g7643, g12881)
--	g13953 = AND(g7646, g12882)
--	g13969 = AND(g7652, g12891)
--	g13970 = AND(g7655, g12892)
--	g13989 = AND(g7661, g12894)
--	g13997 = AND(g7664, g12900)
--	g13998 = AND(g7972, g12907)
--	g14006 = AND(g7670, g12914)
--	g14007 = AND(g7673, g12915)
--	g14022 = AND(g7679, g12921)
--	g14023 = AND(g7682, g12922)
--	g14039 = AND(g7688, g12931)
--	g14040 = AND(g7691, g12932)
--	g14059 = AND(g7697, g12934)
--	g14067 = AND(g7703, g12940)
--	g14097 = AND(g7706, g12943)
--	g14098 = AND(g7709, g12944)
--	g14113 = AND(g7715, g12950)
--	g14114 = AND(g7718, g12951)
--	g14130 = AND(g7724, g12960)
--	g14131 = AND(g7727, g12961)
--	g14143 = AND(g8026, g12965)
--	g14182 = AND(g7733, g12969)
--	g14212 = AND(g7736, g12972)
--	g14213 = AND(g7739, g12973)
--	g14228 = AND(g7745, g12979)
--	g14229 = AND(g7748, g12980)
--	g14297 = AND(g7757, g12993)
--	g14327 = AND(g7760, g12996)
--	g14328 = AND(g7763, g12997)
--	g14336 = AND(g8099, g12998)
--	g14419 = AND(g7779, g13003)
--	g14690 = AND(g7841, g13101)
--	g14724 = AND(g7861, g13117)
--	g14752 = AND(g7891, g13130)
--	g14767 = AND(g13245, g10765)
--	g14773 = AND(g7915, g13141)
--	g14884 = AND(g8169, g12548)
--	g14894 = AND(g3940, g13148)
--	g14956 = AND(g11059, g13151)
--	g14957 = AND(g4015, g13152)
--	g14958 = AND(g4016, g13153)
--	g14975 = AND(g4047, g13154)
--	g15020 = AND(g8090, g12561)
--	g15030 = AND(g4110, g13158)
--	g15031 = AND(g4111, g13159)
--	g15046 = AND(g4142, g13161)
--	g15047 = AND(g4143, g13162)
--	g15064 = AND(g4174, g13163)
--	g15093 = AND(g7869, g12601)
--	g15094 = AND(g7872, g12604)
--	g15104 = AND(g4220, g13167)
--	g15105 = AND(g4224, g13168)
--	g15126 = AND(g4249, g13169)
--	g15127 = AND(g4250, g13170)
--	g15142 = AND(g4281, g13172)
--	g15143 = AND(g4282, g13173)
--	g15160 = AND(g4313, g13174)
--	g15171 = AND(g8015, g12647)
--	g15172 = AND(g4346, g13176)
--	g15173 = AND(g4347, g13177)
--	g15178 = AND(g640, g12651)
--	g15196 = AND(g4375, g13178)
--	g15197 = AND(g4379, g13179)
--	g15218 = AND(g4404, g13180)
--	g15219 = AND(g4405, g13181)
--	g15234 = AND(g4436, g13183)
--	g15235 = AND(g4437, g13184)
--	g15243 = AND(g7849, g12692)
--	g15244 = AND(g7852, g12695)
--	g15245 = AND(g4474, g13185)
--	g15246 = AND(g4475, g13186)
--	g15247 = AND(g4479, g13187)
--	g15257 = AND(g4357, g12702)
--	g15258 = AND(g4515, g13188)
--	g15259 = AND(g4516, g13189)
--	g15264 = AND(g1326, g12705)
--	g15282 = AND(g4544, g13190)
--	g15283 = AND(g4548, g13191)
--	g15304 = AND(g4573, g13192)
--	g15305 = AND(g4574, g13193)
--	g15320 = AND(g7964, g12744)
--	g15321 = AND(g4601, g13195)
--	g15324 = AND(g4609, g13196)
--	g15325 = AND(g4610, g13197)
--	g15335 = AND(g4489, g12749)
--	g15336 = AND(g4492, g12752)
--	g15337 = AND(g4650, g13198)
--	g15338 = AND(g4651, g13199)
--	g15339 = AND(g4655, g13200)
--	g15349 = AND(g4526, g12759)
--	g15350 = AND(g4691, g13201)
--	g15351 = AND(g4692, g13202)
--	g15356 = AND(g2020, g12762)
--	g15374 = AND(g4720, g13203)
--	g15375 = AND(g4724, g13204)
--	g15388 = AND(g7834, g12769)
--	g15389 = AND(g8246, g12772)
--	g15391 = AND(g4752, g13205)
--	g15392 = AND(g4753, g13206)
--	g15402 = AND(g4620, g12783)
--	g15403 = AND(g4623, g12786)
--	g15407 = AND(g4778, g13207)
--	g15410 = AND(g4786, g13208)
--	g15411 = AND(g4787, g13209)
--	g15421 = AND(g4665, g12791)
--	g15422 = AND(g4668, g12794)
--	g15423 = AND(g4827, g13210)
--	g15424 = AND(g4828, g13211)
--	g15425 = AND(g4832, g13212)
--	g15435 = AND(g4702, g12801)
--	g15436 = AND(g4868, g13213)
--	g15437 = AND(g4869, g13214)
--	g15442 = AND(g2714, g12804)
--	g15452 = AND(g7916, g12808)
--	g15453 = AND(g6898, g12811)
--	g15459 = AND(g4897, g13218)
--	g15460 = AND(g4898, g13219)
--	g15470 = AND(g4763, g12816)
--	g15475 = AND(g4928, g13220)
--	g15476 = AND(g4929, g13221)
--	g15486 = AND(g4797, g12822)
--	g15487 = AND(g4800, g12825)
--	g15491 = AND(g4954, g13222)
--	g15494 = AND(g4962, g13223)
--	g15495 = AND(g4963, g13224)
--	g15505 = AND(g4842, g12830)
--	g15506 = AND(g4845, g12833)
--	g15507 = AND(g5003, g13225)
--	g15508 = AND(g5004, g13226)
--	g15509 = AND(g5008, g13227)
--	g15519 = AND(g4879, g12840)
--	g15520 = AND(g8172, g12844)
--	g15526 = AND(g5033, g13232)
--	g15527 = AND(g5034, g13233)
--	g15545 = AND(g5056, g13237)
--	g15546 = AND(g5057, g13238)
--	g15556 = AND(g4939, g12854)
--	g15561 = AND(g5087, g13239)
--	g15562 = AND(g5088, g13240)
--	g15572 = AND(g4973, g12860)
--	g15573 = AND(g4976, g12863)
--	g15577 = AND(g5113, g13241)
--	g15580 = AND(g5121, g13242)
--	g15581 = AND(g5122, g13243)
--	g15591 = AND(g5018, g12868)
--	g15592 = AND(g5021, g12871)
--	g15593 = AND(g7897, g13244)
--	g15594 = AND(g5148, g13249)
--	g15595 = AND(g5149, g13250)
--	g15604 = AND(g5162, g13255)
--	g15605 = AND(g5163, g13256)
--	g15623 = AND(g5185, g13260)
--	g15624 = AND(g5186, g13261)
--	g15634 = AND(g5098, g12895)
--	g15639 = AND(g5216, g13262)
--	g15640 = AND(g5217, g13263)
--	g15650 = AND(g5132, g12901)
--	g15651 = AND(g5135, g12904)
--	g15658 = AND(g8177, g13264)
--	g15666 = AND(g5233, g13268)
--	g15670 = AND(g5241, g13272)
--	g15671 = AND(g5242, g13273)
--	g15680 = AND(g5255, g13278)
--	g15681 = AND(g5256, g13279)
--	g15699 = AND(g5278, g13283)
--	g15700 = AND(g5279, g13284)
--	g15710 = AND(g5227, g12935)
--	g15717 = AND(g7924, g13285)
--	g15725 = AND(g5296, g13293)
--	g15729 = AND(g5304, g13297)
--	g15730 = AND(g5305, g13298)
--	g15739 = AND(g5318, g13303)
--	g15740 = AND(g5319, g13304)
--	g15753 = AND(g7542, g12962)
--	g15754 = AND(g7837, g13308)
--	g15755 = AND(g8178, g13309)
--	g15765 = AND(g5333, g13324)
--	g15769 = AND(g5341, g13328)
--	g15770 = AND(g5342, g13329)
--	I22028 = AND(g13004, g3018, g7549)
--	g15780 = AND(g7471, g3032, I22028)
--	g15781 = AND(g7971, g13330)
--	g15793 = AND(g5361, g13347)
--	g15801 = AND(g7856, g13351)
--	g15802 = AND(g8253, g13352)
--	g15817 = AND(g8025, g13373)
--	g15828 = AND(g7877, g13398)
--	g15829 = AND(g7857, g13400)
--	g15840 = AND(g8098, g11620)
--	g15852 = AND(g7878, g11642)
--	I22136 = AND(g13082, g2912, g7522)
--	g15902 = AND(g7607, g2920, I22136)
--	g15998 = AND(g5469, g11732)
--	g16003 = AND(g12013, g10826)
--	g16004 = AND(g5587, g11734)
--	g16008 = AND(g5504, g11735)
--	g16009 = AND(g12071, g10843)
--	g16010 = AND(g7639, g11736)
--	g16015 = AND(g12013, g10859)
--	g16016 = AND(g5601, g11740)
--	g16017 = AND(g12130, g10862)
--	g16018 = AND(g6149, g11741)
--	g16019 = AND(g5507, g11742)
--	g16028 = AND(g5543, g11745)
--	g16029 = AND(g12071, g10877)
--	g16030 = AND(g7667, g11746)
--	g16031 = AND(g6227, g11747)
--	g16032 = AND(g12187, g10883)
--	g16033 = AND(g5546, g11748)
--	g16045 = AND(g12013, g10892)
--	g16046 = AND(g5618, g11761)
--	g16047 = AND(g12130, g10895)
--	g16048 = AND(g6170, g11762)
--	g16049 = AND(g6638, g11763)
--	g16050 = AND(g5590, g11764)
--	g16051 = AND(g12235, g10901)
--	g16052 = AND(g5591, g11765)
--	g16053 = AND(g297, g11770)
--	g16066 = AND(g12071, g10912)
--	g16067 = AND(g7700, g11774)
--	g16068 = AND(g6310, g11775)
--	g16069 = AND(g5346, g11776)
--	g16070 = AND(g12187, g10921)
--	g16071 = AND(g5604, g11777)
--	g16072 = AND(g12275, g10924)
--	g16073 = AND(g5605, g11778)
--	g16074 = AND(g5646, g11782)
--	g16081 = AND(g3304, g11783)
--	g16089 = AND(g984, g11787)
--	g16100 = AND(g12130, g10937)
--	g16101 = AND(g6197, g11794)
--	g16102 = AND(g6905, g11795)
--	g16103 = AND(g5621, g11796)
--	g16104 = AND(g12235, g10946)
--	g16105 = AND(g5622, g11797)
--	g16106 = AND(g12308, g10949)
--	g16107 = AND(g5666, g11801)
--	g16108 = AND(g5667, g11802)
--	g16109 = AND(g8277, g11803)
--	g16110 = AND(g516, g11804)
--	g16111 = AND(g5551, g13215)
--	g16112 = AND(g5684, g11808)
--	g16119 = AND(g3460, g11809)
--	g16127 = AND(g1678, g11813)
--	g16133 = AND(g6444, g11817)
--	g16134 = AND(g5363, g11818)
--	g16135 = AND(g12187, g10980)
--	g16136 = AND(g5640, g11819)
--	g16137 = AND(g12275, g10983)
--	g16138 = AND(g5641, g11820)
--	g16139 = AND(g5704, g11824)
--	g16140 = AND(g5705, g11825)
--	g16141 = AND(g5706, g11826)
--	g16152 = AND(g517, g11829)
--	g16153 = AND(g5592, g13229)
--	g16158 = AND(g5718, g11834)
--	g16159 = AND(g5719, g11835)
--	g16160 = AND(g8286, g11836)
--	g16161 = AND(g1202, g11837)
--	g16162 = AND(g5597, g13234)
--	g16163 = AND(g5736, g11841)
--	g16170 = AND(g3616, g11842)
--	g16178 = AND(g2372, g11846)
--	g16182 = AND(g7149, g11852)
--	g16183 = AND(g12235, g11014)
--	g16184 = AND(g5663, g11853)
--	g16185 = AND(g12308, g11017)
--	g16186 = AND(g5753, g11856)
--	g16187 = AND(g5754, g11857)
--	g16188 = AND(g5755, g11858)
--	g16197 = AND(g518, g11862)
--	g16198 = AND(g5762, g11866)
--	g16199 = AND(g5763, g11867)
--	g16200 = AND(g5764, g11868)
--	g16211 = AND(g1203, g11871)
--	g16212 = AND(g5609, g13252)
--	g16217 = AND(g5776, g11876)
--	g16218 = AND(g5777, g11877)
--	g16219 = AND(g8295, g11878)
--	g16220 = AND(g1896, g11879)
--	g16221 = AND(g5614, g13257)
--	g16222 = AND(g5794, g11883)
--	g16229 = AND(g3772, g11884)
--	g16237 = AND(g5379, g11886)
--	g16238 = AND(g12275, g11066)
--	g16239 = AND(g5700, g11887)
--	g16240 = AND(g5804, g11891)
--	g16241 = AND(g5805, g11892)
--	g16242 = AND(g5806, g11893)
--	g16250 = AND(g519, g11895)
--	g16251 = AND(g5812, g11898)
--	g16252 = AND(g5813, g11899)
--	g16253 = AND(g5814, g11900)
--	g16262 = AND(g1204, g11904)
--	g16263 = AND(g5821, g11908)
--	g16264 = AND(g5822, g11909)
--	g16265 = AND(g5823, g11910)
--	g16276 = AND(g1897, g11913)
--	g16277 = AND(g5634, g13275)
--	g16282 = AND(g5835, g11918)
--	g16283 = AND(g5836, g11919)
--	g16284 = AND(g8304, g11920)
--	g16285 = AND(g2590, g11921)
--	g16286 = AND(g5639, g13280)
--	g16288 = AND(g12308, g11129)
--	g16289 = AND(g5853, g11929)
--	g16290 = AND(g5854, g11930)
--	g16291 = AND(g5855, g11931)
--	g16292 = AND(g294, g11932)
--	g16298 = AND(g520, g11936)
--	g16299 = AND(g5860, g11941)
--	g16300 = AND(g5861, g11942)
--	g16301 = AND(g5862, g11943)
--	g16309 = AND(g1205, g11945)
--	g16310 = AND(g5868, g11948)
--	g16311 = AND(g5869, g11949)
--	g16312 = AND(g5870, g11950)
--	g16321 = AND(g1898, g11954)
--	g16322 = AND(g5877, g11958)
--	g16323 = AND(g5878, g11959)
--	g16324 = AND(g5879, g11960)
--	g16335 = AND(g2591, g11963)
--	g16336 = AND(g5662, g13300)
--	g16342 = AND(g5894, g11968)
--	g16343 = AND(g5895, g11969)
--	g16344 = AND(g5896, g11970)
--	g16345 = AND(g5897, g11971)
--	g16346 = AND(g295, g11972)
--	g16347 = AND(g5900, g11982)
--	g16348 = AND(g5901, g11983)
--	g16349 = AND(g5902, g11984)
--	g16350 = AND(g981, g11985)
--	g16356 = AND(g1206, g11989)
--	g16357 = AND(g5907, g11994)
--	g16358 = AND(g5908, g11995)
--	g16359 = AND(g5909, g11996)
--	g16367 = AND(g1899, g11998)
--	g16368 = AND(g5915, g12001)
--	g16369 = AND(g5916, g12002)
--	g16370 = AND(g5917, g12003)
--	g16379 = AND(g2592, g12007)
--	g16380 = AND(g5925, g12020)
--	g16381 = AND(g5926, g12021)
--	g16382 = AND(g5927, g12022)
--	g16383 = AND(g5928, g12023)
--	g16384 = AND(g296, g12024)
--	g16385 = AND(g5714, g13336)
--	g16386 = AND(g5933, g12037)
--	g16387 = AND(g5934, g12038)
--	g16388 = AND(g5935, g12039)
--	g16389 = AND(g5936, g12040)
--	g16390 = AND(g982, g12041)
--	g16391 = AND(g5939, g12051)
--	g16392 = AND(g5940, g12052)
--	g16393 = AND(g5941, g12053)
--	g16394 = AND(g1675, g12054)
--	g16400 = AND(g1900, g12058)
--	g16401 = AND(g5946, g12063)
--	g16402 = AND(g5947, g12064)
--	g16403 = AND(g5948, g12065)
--	g16411 = AND(g2593, g12067)
--	g16413 = AND(g5954, g12075)
--	g16414 = AND(g5955, g12076)
--	g16415 = AND(g5956, g12077)
--	g16416 = AND(g5957, g12078)
--	g16417 = AND(g5759, g13356)
--	g16418 = AND(g5959, g12084)
--	g16419 = AND(g5960, g12085)
--	g16420 = AND(g5961, g12086)
--	g16421 = AND(g5962, g12087)
--	g16422 = AND(g983, g12088)
--	g16423 = AND(g5772, g13361)
--	g16424 = AND(g5967, g12101)
--	g16425 = AND(g5968, g12102)
--	g16426 = AND(g5969, g12103)
--	g16427 = AND(g5970, g12104)
--	g16428 = AND(g1676, g12105)
--	g16429 = AND(g5973, g12115)
--	g16430 = AND(g5974, g12116)
--	g16431 = AND(g5975, g12117)
--	g16432 = AND(g2369, g12118)
--	g16438 = AND(g2594, g12122)
--	g16443 = AND(g5980, g12134)
--	g16444 = AND(g5981, g12135)
--	g16445 = AND(g5808, g13381)
--	g16447 = AND(g5983, g12147)
--	g16448 = AND(g5984, g12148)
--	g16449 = AND(g5985, g12149)
--	g16450 = AND(g5986, g12150)
--	g16451 = AND(g5818, g13386)
--	g16452 = AND(g5988, g12156)
--	g16453 = AND(g5989, g12157)
--	g16454 = AND(g5990, g12158)
--	g16455 = AND(g5991, g12159)
--	g16456 = AND(g1677, g12160)
--	g16457 = AND(g5831, g13391)
--	g16458 = AND(g5996, g12173)
--	g16459 = AND(g5997, g12174)
--	g16460 = AND(g5998, g12175)
--	g16461 = AND(g5999, g12176)
--	g16462 = AND(g2370, g12177)
--	g16505 = AND(g14776, g14797, g16142, g16243)
--	g16513 = AND(g15065, g13724, g13764, g13797)
--	g16527 = AND(g14811, g14849, g16201, g16302)
--	g16535 = AND(g15161, g13774, g13805, g13825)
--	g16558 = AND(g14863, g14922, g16266, g16360)
--	g16590 = AND(g14936, g15003, g16325, g16404)
--	g16607 = AND(g15022, g15096)
--	g16625 = AND(g15118, g15188)
--	g16639 = AND(g15210, g15274)
--	g16650 = AND(g15296, g15366)
--	g16850 = AND(g6226, g14764)
--	g16855 = AND(g15722, g8646)
--	g16856 = AND(g6443, g14794)
--	g16859 = AND(g15762, g8662)
--	g16864 = AND(g15790, g8681)
--	g16865 = AND(g6896, g14881)
--	g16879 = AND(g15813, g8693)
--	g16894 = AND(g7156, g14959)
--	g16907 = AND(g7335, g15017)
--	g16908 = AND(g7838, g15032)
--	g16909 = AND(g6908, g15033)
--	g16923 = AND(g7352, g15048)
--	g16938 = AND(g7858, g15128)
--	g16939 = AND(g7158, g15129)
--	g16953 = AND(g7482, g15144)
--	g16964 = AND(g7520, g15170)
--	g16966 = AND(g7529, g15174)
--	g16967 = AND(g7827, g15175)
--	g16968 = AND(g6672, g15176)
--	g16969 = AND(g7888, g15220)
--	g16970 = AND(g7354, g15221)
--	g16984 = AND(g7538, g15236)
--	g16987 = AND(g7555, g15260)
--	g16988 = AND(g7842, g15261)
--	g16989 = AND(g6974, g15262)
--	g16990 = AND(g7912, g15306)
--	g16991 = AND(g7484, g15307)
--	g16993 = AND(g7576, g15322)
--	g16994 = AND(g7819, g15323)
--	g16997 = AND(g7578, g15352)
--	g16998 = AND(g7862, g15353)
--	g16999 = AND(g7224, g15354)
--	g17001 = AND(g3254, g10694, g14144)
--	g17015 = AND(g7996, g15390)
--	g17017 = AND(g7590, g15408)
--	g17018 = AND(g7830, g15409)
--	g17021 = AND(g7592, g15438)
--	g17022 = AND(g7892, g15439)
--	g17023 = AND(g7420, g15440)
--	g17028 = AND(g7604, g15458)
--	g17031 = AND(g3410, g10714, g14259)
--	g17045 = AND(g8071, g15474)
--	g17047 = AND(g7605, g15492)
--	g17048 = AND(g7845, g15493)
--	g17055 = AND(g7153, g15524)
--	g17056 = AND(g7953, g15525)
--	g17062 = AND(g7613, g15544)
--	g17065 = AND(g3566, g10735, g14381)
--	g17079 = AND(g8156, g15560)
--	g17081 = AND(g7614, g15578)
--	g17082 = AND(g7865, g15579)
--	g17084 = AND(g7629, g13954)
--	g17090 = AND(g7349, g15602)
--	g17091 = AND(g8004, g15603)
--	g17097 = AND(g7622, g15622)
--	g17100 = AND(g3722, g10754, g14493)
--	g17114 = AND(g8242, g15638)
--	g17116 = AND(g7649, g14008)
--	g17117 = AND(g7906, g15665)
--	g17122 = AND(g7658, g14024)
--	g17128 = AND(g7479, g15678)
--	g17129 = AND(g8079, g15679)
--	g17135 = AND(g7638, g15698)
--	g17138 = AND(g7676, g14068)
--	g17143 = AND(g7685, g14099)
--	g17144 = AND(g7958, g15724)
--	g17149 = AND(g7694, g14115)
--	g17155 = AND(g7535, g15737)
--	g17156 = AND(g8164, g15738)
--	g17161 = AND(g7712, g14183)
--	g17166 = AND(g7721, g14214)
--	g17167 = AND(g8009, g15764)
--	g17172 = AND(g7730, g14230)
--	g17176 = AND(g7742, g14298)
--	g17181 = AND(g7751, g14329)
--	g17182 = AND(g8084, g15792)
--	g17193 = AND(g7766, g14420)
--	g17268 = AND(g8024, g15991)
--	g17301 = AND(g8097, g15994)
--	g17339 = AND(g8176, g15997)
--	g17352 = AND(g3942, g14960)
--	g17353 = AND(g3945, g14963)
--	g17381 = AND(g8250, g16001)
--	g17382 = AND(g8252, g16002)
--	g17393 = AND(g3941, g16005)
--	g17395 = AND(g6177, g15034)
--	g17396 = AND(g4020, g15037)
--	g17397 = AND(g4023, g15040)
--	g17398 = AND(g4026, g15043)
--	g17408 = AND(g4049, g15049)
--	g17409 = AND(g4052, g15052)
--	g17428 = AND(g3994, g16007)
--	g17446 = AND(g6284, g16011)
--	g17447 = AND(g4115, g15106)
--	g17448 = AND(g4118, g15109)
--	g17449 = AND(g4121, g15112)
--	g17450 = AND(g4124, g15115)
--	g17460 = AND(g4048, g16012)
--	g17461 = AND(g6209, g15130)
--	g17462 = AND(g4147, g15133)
--	g17463 = AND(g4150, g15136)
--	g17464 = AND(g4153, g15139)
--	g17474 = AND(g4176, g15145)
--	g17475 = AND(g4179, g15148)
--	g17485 = AND(g4089, g16013)
--	g17486 = AND(g4091, g16014)
--	g17506 = AND(g6675, g16023)
--	g17508 = AND(g4225, g15179)
--	g17509 = AND(g4228, g15182)
--	g17510 = AND(g4231, g15185)
--	g17526 = AND(g6421, g16025)
--	g17527 = AND(g4254, g15198)
--	g17528 = AND(g4257, g15201)
--	g17529 = AND(g4260, g15204)
--	g17530 = AND(g4263, g15207)
--	g17540 = AND(g4175, g16026)
--	g17541 = AND(g6298, g15222)
--	g17542 = AND(g4286, g15225)
--	g17543 = AND(g4289, g15228)
--	g17544 = AND(g4292, g15231)
--	g17554 = AND(g4315, g15237)
--	g17555 = AND(g4318, g15240)
--	g17556 = AND(g4201, g16027)
--	g17576 = AND(g4348, g15248)
--	g17577 = AND(g4351, g15251)
--	g17578 = AND(g4354, g15254)
--	g17597 = AND(g6977, g16039)
--	g17598 = AND(g4380, g15265)
--	g17599 = AND(g4383, g15268)
--	g17600 = AND(g4386, g15271)
--	g17616 = AND(g6626, g16041)
--	g17617 = AND(g4409, g15284)
--	g17618 = AND(g4412, g15287)
--	g17619 = AND(g4415, g15290)
--	g17620 = AND(g4418, g15293)
--	g17630 = AND(g4314, g16042)
--	g17631 = AND(g6435, g15308)
--	g17632 = AND(g4441, g15311)
--	g17633 = AND(g4444, g15314)
--	g17634 = AND(g4447, g15317)
--	g17635 = AND(g4322, g16043)
--	g17636 = AND(g4324, g16044)
--	g17652 = AND(g4480, g15326)
--	g17653 = AND(g4483, g15329)
--	g17654 = AND(g4486, g15332)
--	g17673 = AND(g4517, g15340)
--	g17674 = AND(g4520, g15343)
--	g17675 = AND(g4523, g15346)
--	g17694 = AND(g7227, g16061)
--	g17695 = AND(g4549, g15357)
--	g17696 = AND(g4552, g15360)
--	g17697 = AND(g4555, g15363)
--	g17713 = AND(g6890, g16063)
--	g17714 = AND(g4578, g15376)
--	g17715 = AND(g4581, g15379)
--	g17716 = AND(g4584, g15382)
--	g17717 = AND(g4587, g15385)
--	g17718 = AND(g4451, g16064)
--	g17719 = AND(g2993, g16065)
--	g17734 = AND(g4611, g15393)
--	g17735 = AND(g4614, g15396)
--	g17736 = AND(g4617, g15399)
--	g17737 = AND(g4626, g15404)
--	g17752 = AND(g4656, g15412)
--	g17753 = AND(g4659, g15415)
--	g17754 = AND(g4662, g15418)
--	g17773 = AND(g4693, g15426)
--	g17774 = AND(g4696, g15429)
--	g17775 = AND(g4699, g15432)
--	g17794 = AND(g7423, g16097)
--	g17795 = AND(g4725, g15443)
--	g17796 = AND(g4728, g15446)
--	g17797 = AND(g4731, g15449)
--	g17798 = AND(g4591, g16099)
--	g17812 = AND(g4754, g15461)
--	g17813 = AND(g4757, g15464)
--	g17814 = AND(g4760, g15467)
--	g17824 = AND(g4766, g15471)
--	g17835 = AND(g4788, g15477)
--	g17836 = AND(g4791, g15480)
--	g17837 = AND(g4794, g15483)
--	g17838 = AND(g4803, g15488)
--	g17853 = AND(g4833, g15496)
--	g17854 = AND(g4836, g15499)
--	g17855 = AND(g4839, g15502)
--	g17874 = AND(g4870, g15510)
--	g17875 = AND(g4873, g15513)
--	g17876 = AND(g4876, g15516)
--	g17877 = AND(g2998, g15521)
--	g17900 = AND(g4899, g15528)
--	g17901 = AND(g4902, g15531)
--	g17902 = AND(g4905, g15534)
--	g17912 = AND(g4908, g15537)
--	g17924 = AND(g4930, g15547)
--	g17925 = AND(g4933, g15550)
--	g17926 = AND(g4936, g15553)
--	g17936 = AND(g4942, g15557)
--	g17947 = AND(g4964, g15563)
--	g17948 = AND(g4967, g15566)
--	g17949 = AND(g4970, g15569)
--	g17950 = AND(g4979, g15574)
--	g17965 = AND(g5009, g15582)
--	g17966 = AND(g5012, g15585)
--	g17967 = AND(g5015, g15588)
--	g17989 = AND(g5035, g15596)
--	g17990 = AND(g5038, g15599)
--	g18011 = AND(g5058, g15606)
--	g18012 = AND(g5061, g15609)
--	g18013 = AND(g5064, g15612)
--	g18023 = AND(g5067, g15615)
--	g18035 = AND(g5089, g15625)
--	g18036 = AND(g5092, g15628)
--	g18037 = AND(g5095, g15631)
--	g18047 = AND(g5101, g15635)
--	g18058 = AND(g5123, g15641)
--	g18059 = AND(g5126, g15644)
--	g18060 = AND(g5129, g15647)
--	g18061 = AND(g5138, g15652)
--	g18062 = AND(g7462, g15655)
--	g18088 = AND(g5150, g15667)
--	g18106 = AND(g5164, g15672)
--	g18107 = AND(g5167, g15675)
--	g18128 = AND(g5187, g15682)
--	g18129 = AND(g5190, g15685)
--	g18130 = AND(g5193, g15688)
--	g18140 = AND(g5196, g15691)
--	g18152 = AND(g5218, g15701)
--	g18153 = AND(g5221, g15704)
--	g18154 = AND(g5224, g15707)
--	g18164 = AND(g5230, g15711)
--	g18165 = AND(g2883, g16287)
--	g18169 = AND(g7527, g15714)
--	g18204 = AND(g5243, g15726)
--	g18222 = AND(g5257, g15731)
--	g18223 = AND(g5260, g15734)
--	g18244 = AND(g5280, g15741)
--	g18245 = AND(g5283, g15744)
--	g18246 = AND(g5286, g15747)
--	g18256 = AND(g5289, g15750)
--	g18311 = AND(g5306, g15766)
--	g18329 = AND(g5320, g15771)
--	g18330 = AND(g5323, g15774)
--	g18333 = AND(g2888, g15777)
--	g18404 = AND(g5343, g15794)
--	I24619 = AND(g14776, g14837, g16142)
--	g18547 = AND(g13677, g13750, I24619)
--	I24689 = AND(g14811, g14910, g16201)
--	g18597 = AND(g13714, g13791, I24689)
--	I24738 = AND(g14863, g14991, g16266)
--	g18629 = AND(g13764, g13819, I24738)
--	I24758 = AND(g14936, g15080, g16325)
--	g18638 = AND(g13805, g13840, I24758)
--	g18645 = AND(g14776, g14895, g16142, g13750)
--	g18647 = AND(g14895, g16142, g16243)
--	g18648 = AND(g14811, g14976, g16201, g13791)
--	g18649 = AND(g14776, g14837, g13657, g16189)
--	g18650 = AND(g14976, g16201, g16302)
--	g18651 = AND(g14863, g15065, g16266, g13819)
--	g18652 = AND(g14797, g13657, g13677, g16243)
--	g18653 = AND(g14811, g14910, g13687, g16254)
--	g18654 = AND(g15065, g16266, g16360)
--	g18655 = AND(g14936, g15161, g16325, g13840)
--	g18665 = AND(g14776, g14837, g16189, g13706)
--	g18666 = AND(g14849, g13687, g13714, g16302)
--	g18667 = AND(g14863, g14991, g13724, g16313)
--	g18668 = AND(g15161, g16325, g16404)
--	g18688 = AND(g14811, g14910, g16254, g13756)
--	g18689 = AND(g14922, g13724, g13764, g16360)
--	g18690 = AND(g14936, g15080, g13774, g16371)
--	g18717 = AND(g14863, g14991, g16313, g13797)
--	g18718 = AND(g15003, g13774, g13805, g16404)
--	g18753 = AND(g14936, g15080, g16371, g13825)
--	g18982 = AND(g13519, g16154)
--	g18990 = AND(g13530, g16213)
--	g18994 = AND(g14895, g13657, g13677, g13706)
--	g18997 = AND(g13541, g16278)
--	g19007 = AND(g14976, g13687, g13714, g13756)
--	g19010 = AND(g13552, g16337)
--	g19063 = AND(g18679, g14910, g13687, g16254)
--	g19079 = AND(g14797, g18692, g16142, g16189)
--	g19080 = AND(g18708, g14991, g13724, g16313)
--	g19087 = AND(g17215, g16540)
--	g19088 = AND(g18656, g14797, g16189, g13706)
--	g19089 = AND(g14849, g18728, g16201, g16254)
--	g19090 = AND(g18744, g15080, g13774, g16371)
--	g19092 = AND(g14776, g18670, g18692, g16293)
--	g19093 = AND(g17218, g16572)
--	g19094 = AND(g18679, g14849, g16254, g13756)
--	g19095 = AND(g14922, g18765, g16266, g16313)
--	I25280 = AND(g18656, g18670, g18720)
--	g19097 = AND(g13657, g16243, I25280)
--	g19099 = AND(g14811, g18699, g18728, g16351)
--	g19100 = AND(g17220, g16596)
--	g19101 = AND(g18708, g14922, g16313, g13797)
--	g19102 = AND(g15003, g18796, g16325, g16371)
--	I25291 = AND(g18679, g18699, g18758)
--	g19104 = AND(g13687, g16302, I25291)
--	g19106 = AND(g14863, g18735, g18765, g16395)
--	g19107 = AND(g17223, g16616)
--	g19108 = AND(g18744, g15003, g16371, g13825)
--	I25300 = AND(g18708, g18735, g18789)
--	g19109 = AND(g13724, g16360, I25300)
--	g19111 = AND(g14936, g18772, g18796, g16433)
--	g19112 = AND(g14657, g16633)
--	I25311 = AND(g18744, g18772, g18815)
--	g19116 = AND(g13774, g16404, I25311)
--	g19117 = AND(g14691, g16644)
--	g19124 = AND(g14725, g16656)
--	g19131 = AND(g14753, g16673)
--	g19142 = AND(g17159, g16719)
--	g19143 = AND(g17174, g16761)
--	g19146 = AND(g17191, g16788)
--	g19148 = AND(g17202, g16817)
--	g19150 = AND(g17189, g8602)
--	g19155 = AND(g17200, g8614)
--	g19161 = AND(g17207, g8627)
--	g19166 = AND(g17212, g8637)
--	g19228 = AND(g16662, g12125)
--	g19236 = AND(g16935, g8802)
--	g19241 = AND(g16867, g14158, g14071)
--	g19248 = AND(g16662, g8817)
--	g19252 = AND(g18725, g9527)
--	g19254 = AND(g16895, g14273, g14186)
--	g19260 = AND(g16749, g3124)
--	g19267 = AND(g16924, g14395, g14301)
--	g19282 = AND(g16954, g14507, g14423)
--	g19284 = AND(g18063, g3111)
--	g19285 = AND(g16749, g7642)
--	g19289 = AND(g17029, g8580)
--	g19303 = AND(g16867, g16543, g14071)
--	g19307 = AND(g17063, g8587)
--	g19316 = AND(g18063, g3110)
--	g19317 = AND(g16749, g3126)
--	g19320 = AND(g16867, g16515, g14158)
--	g19324 = AND(g16895, g16575, g14186)
--	g19328 = AND(g17098, g8594)
--	g19347 = AND(g16895, g16546, g14273)
--	g19351 = AND(g16924, g16599, g14301)
--	g19355 = AND(g17136, g8605)
--	g19356 = AND(g18063, g3112)
--	g19381 = AND(g16924, g16578, g14395)
--	g19385 = AND(g16954, g16619, g14423)
--	g19413 = AND(g16954, g16602, g14507)
--	g19449 = AND(g16884, g14797, g14776)
--	g19476 = AND(g16913, g14849, g14811)
--	g19499 = AND(g16943, g14922, g14863)
--	g19520 = AND(g16974, g15003, g14936)
--	g19531 = AND(g16884, g16722, g14776)
--	g19540 = AND(g16884, g16697, g14797)
--	g19541 = AND(g16913, g16764, g14811)
--	g19544 = AND(g16913, g16728, g14849)
--	g19545 = AND(g16943, g16791, g14863)
--	g19547 = AND(g16943, g16770, g14922)
--	g19548 = AND(g16974, g16820, g14936)
--	g19549 = AND(g7950, g17230)
--	g19551 = AND(g16974, g16797, g15003)
--	g19552 = AND(g16829, g6048)
--	g19553 = AND(g7990, g17237)
--	g19554 = AND(g7993, g17240)
--	g19555 = AND(g8001, g17243)
--	g19557 = AND(g8053, g17249)
--	g19558 = AND(g8056, g17252)
--	g19559 = AND(g8059, g17255)
--	g19560 = AND(g8065, g17259)
--	g19561 = AND(g8068, g17262)
--	g19562 = AND(g8076, g17265)
--	g19564 = AND(g8123, g17272)
--	g19565 = AND(g8126, g17275)
--	g19566 = AND(g8129, g17278)
--	g19567 = AND(g8138, g17282)
--	g19568 = AND(g8141, g17285)
--	g19569 = AND(g8144, g17288)
--	g19570 = AND(g8150, g17291)
--	g19571 = AND(g8153, g17294)
--	g19572 = AND(g8161, g17297)
--	g19574 = AND(g8191, g17304)
--	g19575 = AND(g8194, g17307)
--	g19576 = AND(g8197, g17310)
--	g19584 = AND(g640, g18756)
--	g19585 = AND(g692, g18757)
--	g19586 = AND(g8209, g17315)
--	g19587 = AND(g8212, g17318)
--	g19588 = AND(g8215, g17321)
--	g19589 = AND(g8224, g17324)
--	g19590 = AND(g8227, g17327)
--	g19591 = AND(g8230, g17330)
--	g19592 = AND(g8236, g17333)
--	g19593 = AND(g8239, g17336)
--	g19594 = AND(g16935, g12555)
--	g19597 = AND(g3922, g17342)
--	g19598 = AND(g3925, g17345)
--	g19599 = AND(g3928, g17348)
--	g19600 = AND(g633, g18783)
--	g19601 = AND(g640, g18784)
--	g19602 = AND(g633, g18785)
--	g19603 = AND(g692, g18786)
--	g19604 = AND(g3948, g17354)
--	g19605 = AND(g3951, g17357)
--	g19606 = AND(g3954, g17360)
--	g19614 = AND(g1326, g18787)
--	g19615 = AND(g1378, g18788)
--	g19616 = AND(g3966, g17363)
--	g19617 = AND(g3969, g17366)
--	g19618 = AND(g3972, g17369)
--	g19619 = AND(g3981, g17372)
--	g19620 = AND(g3984, g17375)
--	g19621 = AND(g3987, g17378)
--	g19623 = AND(g4000, g17384)
--	g19624 = AND(g4003, g17387)
--	g19625 = AND(g4006, g17390)
--	g19626 = AND(g640, g18805)
--	g19627 = AND(g633, g18806)
--	g19628 = AND(g653, g18807)
--	g19629 = AND(g692, g18808)
--	g19630 = AND(g4029, g17399)
--	g19631 = AND(g4032, g17402)
--	g19632 = AND(g4035, g17405)
--	g19633 = AND(g1319, g18809)
--	g19634 = AND(g1326, g18810)
--	g19635 = AND(g1319, g18811)
--	g19636 = AND(g1378, g18812)
--	g19637 = AND(g4055, g17410)
--	g19638 = AND(g4058, g17413)
--	g19639 = AND(g4061, g17416)
--	g19647 = AND(g2020, g18813)
--	g19648 = AND(g2072, g18814)
--	g19649 = AND(g4073, g17419)
--	g19650 = AND(g4076, g17422)
--	g19651 = AND(g4079, g17425)
--	g19653 = AND(g4095, g17430)
--	g19654 = AND(g4098, g17433)
--	g19655 = AND(g4101, g17436)
--	g19656 = AND(g4104, g17439)
--	g19660 = AND(g633, g18822)
--	g19661 = AND(g653, g18823)
--	g19662 = AND(g646, g18824)
--	g19663 = AND(g4127, g17451)
--	g19664 = AND(g4130, g17454)
--	g19665 = AND(g4133, g17457)
--	g19666 = AND(g1326, g18825)
--	g19667 = AND(g1319, g18826)
--	g19668 = AND(g1339, g18827)
--	g19669 = AND(g1378, g18828)
--	g19670 = AND(g4156, g17465)
--	g19671 = AND(g4159, g17468)
--	g19672 = AND(g4162, g17471)
--	g19673 = AND(g2013, g18829)
--	g19674 = AND(g2020, g18830)
--	g19675 = AND(g2013, g18831)
--	g19676 = AND(g2072, g18832)
--	g19677 = AND(g4182, g17476)
--	g19678 = AND(g4185, g17479)
--	g19679 = AND(g4188, g17482)
--	g19687 = AND(g2714, g18833)
--	g19688 = AND(g2766, g18834)
--	g19691 = AND(g16841, g10865)
--	g19692 = AND(g4205, g17487)
--	g19693 = AND(g4208, g17490)
--	g19694 = AND(g4211, g17493)
--	g19695 = AND(g4214, g17496)
--	g19697 = AND(g653, g18838)
--	g19698 = AND(g646, g18839)
--	g19699 = AND(g660, g18840)
--	g19700 = AND(g17815, g16024)
--	g19701 = AND(g4234, g17511)
--	g19702 = AND(g4237, g17514)
--	g19703 = AND(g4240, g17517)
--	g19704 = AND(g4243, g17520)
--	g19708 = AND(g1319, g18841)
--	g19709 = AND(g1339, g18842)
--	g19710 = AND(g1332, g18843)
--	g19711 = AND(g4266, g17531)
--	g19712 = AND(g4269, g17534)
--	g19713 = AND(g4272, g17537)
--	g19714 = AND(g2020, g18844)
--	g19715 = AND(g2013, g18845)
--	g19716 = AND(g2033, g18846)
--	g19717 = AND(g2072, g18847)
--	g19718 = AND(g4295, g17545)
--	g19719 = AND(g4298, g17548)
--	g19720 = AND(g4301, g17551)
--	g19721 = AND(g2707, g18848)
--	g19722 = AND(g2714, g18849)
--	g19723 = AND(g2707, g18850)
--	g19724 = AND(g2766, g18851)
--	g19726 = AND(g16847, g6131)
--	g19727 = AND(g4329, g17557)
--	g19728 = AND(g4332, g17560)
--	g19729 = AND(g4335, g17563)
--	g19730 = AND(g653, g17573)
--	g19731 = AND(g646, g18853)
--	g19732 = AND(g660, g18854)
--	g19733 = AND(g672, g18855)
--	g19734 = AND(g17815, g16034)
--	g19735 = AND(g17903, g16035)
--	g19736 = AND(g4360, g17579)
--	g19737 = AND(g4363, g17582)
--	g19738 = AND(g4366, g17585)
--	g19739 = AND(g4369, g17588)
--	g19741 = AND(g1339, g18856)
--	g19742 = AND(g1332, g18857)
--	g19743 = AND(g1346, g18858)
--	g19744 = AND(g17927, g16040)
--	g19745 = AND(g4389, g17601)
--	g19746 = AND(g4392, g17604)
--	g19747 = AND(g4395, g17607)
--	g19748 = AND(g4398, g17610)
--	g19752 = AND(g2013, g18859)
--	g19753 = AND(g2033, g18860)
--	g19754 = AND(g2026, g18861)
--	g19755 = AND(g4421, g17621)
--	g19756 = AND(g4424, g17624)
--	g19757 = AND(g4427, g17627)
--	g19758 = AND(g2714, g18862)
--	g19759 = AND(g2707, g18863)
--	g19760 = AND(g2727, g18864)
--	g19761 = AND(g2766, g18865)
--	g19764 = AND(g4453, g17637)
--	g19765 = AND(g660, g18870)
--	g19766 = AND(g672, g18871)
--	g19767 = AND(g666, g18872)
--	g19768 = AND(g17815, g16054)
--	g19769 = AND(g17903, g16055)
--	g19770 = AND(g4498, g17655)
--	g19771 = AND(g4501, g17658)
--	g19772 = AND(g4504, g17661)
--	g19773 = AND(g1339, g17670)
--	g19774 = AND(g1332, g18874)
--	g19775 = AND(g1346, g18875)
--	g19776 = AND(g1358, g18876)
--	g19777 = AND(g17927, g16056)
--	g19778 = AND(g18014, g16057)
--	g19779 = AND(g4529, g17676)
--	g19780 = AND(g4532, g17679)
--	g19781 = AND(g4535, g17682)
--	g19782 = AND(g4538, g17685)
--	g19784 = AND(g2033, g18877)
--	g19785 = AND(g2026, g18878)
--	g19786 = AND(g2040, g18879)
--	g19787 = AND(g18038, g16062)
--	g19788 = AND(g4558, g17698)
--	g19789 = AND(g4561, g17701)
--	g19790 = AND(g4564, g17704)
--	g19791 = AND(g4567, g17707)
--	g19795 = AND(g2707, g18880)
--	g19796 = AND(g2727, g18881)
--	g19797 = AND(g2720, g18882)
--	I26240 = AND(g18174, g18341, g17974)
--	g19799 = AND(g17640, g18074, I26240)
--	g19802 = AND(g672, g18891)
--	g19803 = AND(g666, g18892)
--	g19804 = AND(g679, g18893)
--	g19805 = AND(g17903, g16088)
--	g19806 = AND(g4629, g17738)
--	g19807 = AND(g1346, g18896)
--	g19808 = AND(g1358, g18897)
--	g19809 = AND(g1352, g18898)
--	g19810 = AND(g17927, g16090)
--	g19811 = AND(g18014, g16091)
--	g19812 = AND(g4674, g17755)
--	g19813 = AND(g4677, g17758)
--	g19814 = AND(g4680, g17761)
--	g19815 = AND(g2033, g17770)
--	g19816 = AND(g2026, g18900)
--	g19817 = AND(g2040, g18901)
--	g19818 = AND(g2052, g18902)
--	g19819 = AND(g18038, g16092)
--	g19820 = AND(g18131, g16093)
--	g19821 = AND(g4705, g17776)
--	g19822 = AND(g4708, g17779)
--	g19823 = AND(g4711, g17782)
--	g19824 = AND(g4714, g17785)
--	g19826 = AND(g2727, g18903)
--	g19827 = AND(g2720, g18904)
--	g19828 = AND(g2734, g18905)
--	g19829 = AND(g18155, g16098)
--	g19836 = AND(g7143, g18908)
--	g19837 = AND(g6901, g17799)
--	g19839 = AND(g666, g18909)
--	g19840 = AND(g679, g18910)
--	g19841 = AND(g686, g18911)
--	I26282 = AND(g18188, g18089, g17991)
--	g19842 = AND(g14525, g13922, I26282)
--	I26285 = AND(g18281, g18436, g18091)
--	g19843 = AND(g17741, g18190, I26285)
--	g19846 = AND(g1358, g18914)
--	g19847 = AND(g1352, g18915)
--	g19848 = AND(g1365, g18916)
--	g19849 = AND(g18014, g16126)
--	g19850 = AND(g4806, g17839)
--	g19851 = AND(g2040, g18919)
--	g19852 = AND(g2052, g18920)
--	g19853 = AND(g2046, g18921)
--	g19854 = AND(g18038, g16128)
--	g19855 = AND(g18131, g16129)
--	g19856 = AND(g4851, g17856)
--	g19857 = AND(g4854, g17859)
--	g19858 = AND(g4857, g17862)
--	g19859 = AND(g2727, g17871)
--	g19860 = AND(g2720, g18923)
--	g19861 = AND(g2734, g18924)
--	g19862 = AND(g2746, g18925)
--	g19863 = AND(g18155, g16130)
--	g19864 = AND(g18247, g16131)
--	g19868 = AND(g16498, g16867, g19001)
--	g19869 = AND(g679, g18926)
--	g19870 = AND(g686, g18927)
--	I26311 = AND(g18353, g13958, g14011)
--	g19871 = AND(g14086, g18275, I26311)
--	g19872 = AND(g1352, g18928)
--	g19873 = AND(g1365, g18929)
--	g19874 = AND(g1372, g18930)
--	I26317 = AND(g18295, g18205, g18108)
--	g19875 = AND(g14580, g13978, I26317)
--	I26320 = AND(g18374, g18509, g18207)
--	g19876 = AND(g17842, g18297, I26320)
--	g19879 = AND(g2052, g18933)
--	g19880 = AND(g2046, g18934)
--	g19881 = AND(g2059, g18935)
--	g19882 = AND(g18131, g16177)
--	g19883 = AND(g4982, g17951)
--	g19884 = AND(g2734, g18938)
--	g19885 = AND(g2746, g18939)
--	g19886 = AND(g2740, g18940)
--	g19887 = AND(g18155, g16179)
--	g19888 = AND(g18247, g16180)
--	g19889 = AND(g2912, g18943)
--	g19895 = AND(g686, g18945)
--	g19899 = AND(g16520, g16895, g16507)
--	g19900 = AND(g1365, g18946)
--	g19901 = AND(g1372, g18947)
--	I26348 = AND(g18448, g14028, g14102)
--	g19902 = AND(g14201, g18368, I26348)
--	g19903 = AND(g2046, g18948)
--	g19904 = AND(g2059, g18949)
--	g19905 = AND(g2066, g18950)
--	I26354 = AND(g18388, g18312, g18224)
--	g19906 = AND(g14614, g14048, I26354)
--	I26357 = AND(g18469, g18573, g18314)
--	g19907 = AND(g17954, g18390, I26357)
--	g19910 = AND(g2746, g18953)
--	g19911 = AND(g2740, g18954)
--	g19912 = AND(g2753, g18955)
--	g19913 = AND(g18247, g16236)
--	g19914 = AND(g3018, g18958)
--	g19920 = AND(g1372, g18961)
--	g19924 = AND(g16551, g16924, g16529)
--	g19925 = AND(g2059, g18962)
--	g19926 = AND(g2066, g18963)
--	I26377 = AND(g18521, g14119, g14217)
--	g19927 = AND(g14316, g18463, I26377)
--	g19928 = AND(g2740, g18964)
--	g19929 = AND(g2753, g18965)
--	g19930 = AND(g2760, g18966)
--	I26383 = AND(g18483, g18405, g18331)
--	g19931 = AND(g14637, g14139, I26383)
--	g19932 = AND(g2917, g18166)
--	g19935 = AND(g2066, g18972)
--	g19939 = AND(g16583, g16954, g16560)
--	g19940 = AND(g2753, g18973)
--	g19941 = AND(g2760, g18974)
--	I26396 = AND(g18585, g14234, g14332)
--	g19942 = AND(g14438, g18536, I26396)
--	g19943 = AND(g7562, g18976)
--	g19944 = AND(g3028, g18258)
--	g19949 = AND(g5293, g18278)
--	g19952 = AND(g2760, g18987)
--	g19953 = AND(g7566, g18334)
--	I26416 = AND(g18553, g18491, g18431)
--	g19970 = AND(g18354, g18276, I26416)
--	g19971 = AND(g5327, g18355)
--	g19976 = AND(g5330, g18371)
--	I26432 = AND(g18277, g18189, g18090)
--	g19982 = AND(g17992, g17913, I26432)
--	g19983 = AND(g5352, g18432)
--	I26440 = AND(g18603, g18555, g18504)
--	g20000 = AND(g18449, g18369, I26440)
--	g20001 = AND(g5355, g18450)
--	g20006 = AND(g5358, g18466)
--	g20011 = AND(g18063, g3113)
--	g20012 = AND(g16804, g3135)
--	g20013 = AND(g17720, g12848)
--	g20014 = AND(g7615, g16749)
--	I26464 = AND(g18370, g18296, g18206)
--	g20020 = AND(g18109, g18024, I26464)
--	g20021 = AND(g5369, g18505)
--	I26472 = AND(g18635, g18605, g18568)
--	g20038 = AND(g18522, g18464, I26472)
--	g20039 = AND(g5372, g18523)
--	g20044 = AND(g5375, g18539)
--	g20048 = AND(g16749, g3127)
--	g20049 = AND(g17878, g3155)
--	g20050 = AND(g18070, g3161)
--	g20051 = AND(g18063, g3114)
--	g20052 = AND(g16804, g3134)
--	g20053 = AND(g17720, g12875)
--	I26500 = AND(g18465, g18389, g18313)
--	g20062 = AND(g18225, g18141, I26500)
--	g20063 = AND(g5382, g18569)
--	I26508 = AND(g18644, g18637, g18618)
--	g20080 = AND(g18586, g18537, I26508)
--	g20081 = AND(g5385, g18587)
--	g20084 = AND(g17969, g3158)
--	g20085 = AND(g18170, g3164)
--	g20086 = AND(g18337, g3170)
--	g20087 = AND(g16749, g7574)
--	g20088 = AND(g16836, g3147)
--	g20089 = AND(g17969, g9160)
--	g20090 = AND(g18063, g3120)
--	g20091 = AND(g16804, g3136)
--	g20092 = AND(g16749, g7603)
--	I26525 = AND(g18656, g18670, g18692)
--	g20093 = AND(g13657, g13677, g13750, I26525)
--	I26528 = AND(g18656, g14837, g13657)
--	g20094 = AND(g13677, g13706, I26528)
--	I26541 = AND(g18538, g18484, g18406)
--	g20103 = AND(g18332, g18257, I26541)
--	g20104 = AND(g5391, g18619)
--	g20106 = AND(g18261, g3167)
--	g20107 = AND(g18415, g3173)
--	g20108 = AND(g18543, g3179)
--	g20109 = AND(g17878, g9504)
--	g20110 = AND(g18070, g9286)
--	g20111 = AND(g18261, g9884)
--	g20112 = AND(g16749, g3132)
--	g20113 = AND(g16836, g3142)
--	g20114 = AND(g17969, g9755)
--	g20115 = AND(g16804, g3139)
--	I26558 = AND(g14776, g18670, g18720)
--	g20116 = AND(g16142, g13677, g13706, I26558)
--	I26561 = AND(g14776, g18720, g13657)
--	g20117 = AND(g16189, g13706, I26561)
--	I26564 = AND(g18679, g18699, g18728)
--	g20118 = AND(g13687, g13714, g13791, I26564)
--	I26567 = AND(g18679, g14910, g13687)
--	g20119 = AND(g13714, g13756, I26567)
--	g20131 = AND(g18486, g3176)
--	g20132 = AND(g18593, g3182)
--	g20133 = AND(g18170, g9505)
--	g20134 = AND(g18337, g9506)
--	g20135 = AND(g18486, g9885)
--	g20136 = AND(g17878, g9423)
--	g20137 = AND(g18070, g9226)
--	g20138 = AND(g18261, g9756)
--	g20139 = AND(g16836, g3151)
--	g20144 = AND(g16679, g16884, g16665)
--	g20145 = AND(g14776, g18670, g16142, g16189)
--	I26590 = AND(g14811, g18699, g18758)
--	g20146 = AND(g16201, g13714, g13756, I26590)
--	I26593 = AND(g14811, g18758, g13687)
--	g20147 = AND(g16254, g13756, I26593)
--	I26596 = AND(g18708, g18735, g18765)
--	g20148 = AND(g13724, g13764, g13819, I26596)
--	I26599 = AND(g18708, g14991, g13724)
--	g20149 = AND(g13764, g13797, I26599)
--	g20156 = AND(g16809, g3185)
--	g20157 = AND(g18415, g9287)
--	g20158 = AND(g18543, g9886)
--	g20159 = AND(g16809, g9288)
--	g20160 = AND(g18170, g9424)
--	g20161 = AND(g18337, g9426)
--	g20162 = AND(g18486, g9757)
--	I26615 = AND(g14797, g18692, g13657)
--	g20177 = AND(g13677, g13750, I26615)
--	g20182 = AND(g16705, g16913, g16686)
--	g20183 = AND(g14811, g18699, g16201, g16254)
--	I26621 = AND(g14863, g18735, g18789)
--	g20184 = AND(g16266, g13764, g13797, I26621)
--	I26624 = AND(g14863, g18789, g13724)
--	g20185 = AND(g16313, g13797, I26624)
--	I26627 = AND(g18744, g18772, g18796)
--	g20186 = AND(g13774, g13805, g13840, I26627)
--	I26630 = AND(g18744, g15080, g13774)
--	g20187 = AND(g13805, g13825, I26630)
--	g20188 = AND(g18593, g9425)
--	g20189 = AND(g16825, g9289)
--	g20190 = AND(g18415, g9227)
--	g20191 = AND(g18543, g9758)
--	g20192 = AND(g16809, g9228)
--	I26639 = AND(g18656, g18670, g16142)
--	g20197 = AND(g13677, g13706, I26639)
--	I26645 = AND(g14849, g18728, g13687)
--	g20211 = AND(g13714, g13791, I26645)
--	g20216 = AND(g16736, g16943, g16712)
--	g20217 = AND(g14863, g18735, g16266, g16313)
--	I26651 = AND(g14936, g18772, g18815)
--	g20218 = AND(g16325, g13805, g13825, I26651)
--	I26654 = AND(g14936, g18815, g13774)
--	g20219 = AND(g16371, g13825, I26654)
--	g20220 = AND(g18593, g9355)
--	g20221 = AND(g16825, g10099)
--	g20222 = AND(g18656, g18720, g13657, g16293)
--	I26661 = AND(g18679, g18699, g16201)
--	g20227 = AND(g13714, g13756, I26661)
--	I26667 = AND(g14922, g18765, g13724)
--	g20241 = AND(g13764, g13819, I26667)
--	g20246 = AND(g16778, g16974, g16743)
--	g20247 = AND(g14936, g18772, g16325, g16371)
--	g20248 = AND(g18656, g14837, g16293)
--	g20249 = AND(g18679, g18758, g13687, g16351)
--	I26676 = AND(g18708, g18735, g16266)
--	g20254 = AND(g13764, g13797, I26676)
--	I26682 = AND(g15003, g18796, g13774)
--	g20268 = AND(g13805, g13840, I26682)
--	g20270 = AND(g14797, g18692, g13657, g16243)
--	g20271 = AND(g18679, g14910, g16351)
--	g20272 = AND(g18708, g18789, g13724, g16395)
--	I26690 = AND(g18744, g18772, g16325)
--	g20277 = AND(g13805, g13825, I26690)
--	I26695 = AND(g18670, g18692, g16142)
--	g20280 = AND(g13677, g16243, I26695)
--	g20282 = AND(g14849, g18728, g13687, g16302)
--	g20283 = AND(g18708, g14991, g16395)
--	g20284 = AND(g18744, g18815, g13774, g16433)
--	g20285 = AND(g16846, g8103)
--	I26708 = AND(g18699, g18728, g16201)
--	g20291 = AND(g13714, g16302, I26708)
--	g20293 = AND(g14922, g18765, g13724, g16360)
--	g20294 = AND(g18744, g15080, g16433)
--	I26726 = AND(g18735, g18765, g16266)
--	g20307 = AND(g13764, g16360, I26726)
--	g20309 = AND(g15003, g18796, g13774, g16404)
--	I26745 = AND(g18772, g18796, g16325)
--	g20326 = AND(g13805, g16404, I26745)
--	g20460 = AND(g17351, g13644)
--	g20472 = AND(g17314, g13669)
--	g20480 = AND(g17313, g11827)
--	g20486 = AND(g17281, g11859)
--	g20492 = AND(g17258, g11894)
--	g20499 = AND(g17648, g11933)
--	g20502 = AND(g17566, g11973)
--	g20503 = AND(g17507, g13817)
--	g20506 = AND(g17499, g12025)
--	g20512 = AND(g17445, g13836)
--	g20525 = AND(g17394, g13849)
--	g20538 = AND(g18656, g14837, g13657, g16189)
--	g20640 = AND(g4809, g19064)
--	g20647 = AND(g5888, g19075)
--	g20665 = AND(g4985, g19081)
--	g20809 = AND(g5712, g19113)
--	g20826 = AND(g5770, g19118)
--	g20836 = AND(g5829, g19125)
--	g20840 = AND(g5885, g19132)
--	g21049 = AND(g20016, g14079, g14165)
--	g21067 = AND(g20193, g12030)
--	g21068 = AND(g20058, g14194, g14280)
--	g21077 = AND(g20223, g12094)
--	g21078 = AND(g20099, g14309, g14402)
--	g21085 = AND(g19484, g14158, g19001)
--	g21086 = AND(g20193, g12142)
--	g21091 = AND(g20250, g12166)
--	g21092 = AND(g20124, g14431, g14514)
--	g21097 = AND(g19505, g14273, g16507)
--	g21098 = AND(g20223, g12204)
--	g21103 = AND(g20273, g12228)
--	g21107 = AND(g19444, g17893, g14079)
--	g21111 = AND(g19524, g14395, g16529)
--	g21112 = AND(g20250, g12259)
--	g21121 = AND(g20054, g14244)
--	g21122 = AND(g20140, g12279)
--	g21123 = AND(g19970, g19982)
--	g21124 = AND(g19471, g18004, g14194)
--	g21128 = AND(g19534, g14507, g16560)
--	g21129 = AND(g20273, g12302)
--	I27695 = AND(g19318, g19300, g19286)
--	g21136 = AND(g19271, g19261, I27695)
--	g21137 = AND(g5750, g19272)
--	g21138 = AND(g19484, g14347)
--	g21140 = AND(g20095, g14366)
--	g21141 = AND(g20178, g12315)
--	g21142 = AND(g20000, g20020)
--	g21143 = AND(g19494, g18121, g14309)
--	I27711 = AND(g19262, g19414, g19386)
--	g21152 = AND(g19357, g19334, I27711)
--	g21153 = AND(g20054, g16543, g16501)
--	g21154 = AND(g20193, g12333)
--	g21155 = AND(g20140, g12336)
--	I27717 = AND(g19345, g19321, g19304)
--	g21156 = AND(g19290, g19276, I27717)
--	g21157 = AND(g5809, g19291)
--	g21158 = AND(g19505, g14459)
--	g21160 = AND(g20120, g14478)
--	g21161 = AND(g20212, g12343)
--	g21162 = AND(g20038, g20062)
--	g21163 = AND(g19515, g18237, g14431)
--	I27733 = AND(g19277, g19451, g19416)
--	g21172 = AND(g19389, g19368, I27733)
--	g21173 = AND(g20095, g16575, g16523)
--	g21174 = AND(g20223, g12363)
--	g21175 = AND(g20178, g12366)
--	I27739 = AND(g19379, g19348, g19325)
--	g21176 = AND(g19308, g19295, I27739)
--	g21177 = AND(g5865, g19309)
--	g21178 = AND(g19524, g14546)
--	g21180 = AND(g20150, g14565)
--	g21181 = AND(g20242, g12373)
--	g21182 = AND(g20080, g20103)
--	g21188 = AND(g20140, g12379)
--	I27755 = AND(g19296, g19478, g19453)
--	g21192 = AND(g19419, g19400, I27755)
--	g21193 = AND(g20120, g16599, g16554)
--	g21194 = AND(g20250, g12382)
--	g21195 = AND(g20212, g12385)
--	I27761 = AND(g19411, g19382, g19352)
--	g21196 = AND(g19329, g19313, I27761)
--	g21197 = AND(g5912, g19330)
--	g21198 = AND(g19534, g14601)
--	g21203 = AND(g20178, g12409)
--	I27772 = AND(g19314, g19501, g19480)
--	g21207 = AND(g19456, g19430, I27772)
--	g21208 = AND(g20150, g16619, g16586)
--	g21209 = AND(g20273, g12412)
--	g21210 = AND(g20242, g12415)
--	g21218 = AND(g20212, g12421)
--	g21226 = AND(g20242, g12426)
--	g21229 = AND(g19578, g14797, g16665)
--	g21234 = AND(g19608, g14849, g16686)
--	g21243 = AND(g19641, g14922, g16712)
--	g21245 = AND(g20299, g14837)
--	g21251 = AND(g19681, g15003, g16743)
--	g21252 = AND(g19578, g14895)
--	g21254 = AND(g20318, g14910)
--	g21259 = AND(g20299, g16722, g16682)
--	g21260 = AND(g19608, g14976)
--	g21262 = AND(g20337, g14991)
--	g21267 = AND(g20318, g16764, g16708)
--	g21268 = AND(g19641, g15065)
--	g21270 = AND(g20357, g15080)
--	g21276 = AND(g20337, g16791, g16739)
--	g21277 = AND(g19681, g15161)
--	g21283 = AND(g20357, g16820, g16781)
--	g21284 = AND(g9356, g20269)
--	g21290 = AND(g9356, g20278)
--	g21291 = AND(g9293, g20279)
--	g21292 = AND(g9453, g20281)
--	g21298 = AND(g9356, g20286)
--	g21299 = AND(g9293, g20287)
--	g21300 = AND(g9232, g20288)
--	g21301 = AND(g9453, g20289)
--	g21302 = AND(g9374, g20290)
--	g21303 = AND(g9595, g20292)
--	g21304 = AND(g9293, g20296)
--	g21305 = AND(g9232, g20297)
--	g21306 = AND(g9187, g20298)
--	g21307 = AND(g9453, g20302)
--	g21308 = AND(g9374, g20303)
--	g21309 = AND(g9310, g20304)
--	g21310 = AND(g9595, g20305)
--	g21311 = AND(g9471, g20306)
--	g21312 = AND(g9737, g20308)
--	g21313 = AND(g9232, g20311)
--	g21314 = AND(g9187, g20312)
--	g21315 = AND(g9161, g20313)
--	g21319 = AND(g9374, g20315)
--	g21320 = AND(g9310, g20316)
--	g21321 = AND(g9248, g20317)
--	g21322 = AND(g9595, g20321)
--	g21323 = AND(g9471, g20322)
--	g21324 = AND(g9391, g20323)
--	g21325 = AND(g9737, g20324)
--	g21326 = AND(g9613, g20325)
--	g21328 = AND(g9187, g20327)
--	g21329 = AND(g9161, g20328)
--	g21330 = AND(g9150, g20329)
--	g21334 = AND(g9310, g20330)
--	g21335 = AND(g9248, g20331)
--	g21336 = AND(g9203, g20332)
--	g21337 = AND(g9471, g20334)
--	g21338 = AND(g9391, g20335)
--	g21339 = AND(g9326, g20336)
--	g21340 = AND(g9737, g20340)
--	g21341 = AND(g9613, g20341)
--	g21342 = AND(g9488, g20342)
--	g21343 = AND(g9161, g20344)
--	g21344 = AND(g9150, g20345)
--	g21345 = AND(g15096, g20346)
--	g21349 = AND(g9248, g20347)
--	g21350 = AND(g9203, g20348)
--	g21351 = AND(g9174, g20349)
--	g21352 = AND(g9391, g20350)
--	g21353 = AND(g9326, g20351)
--	g21354 = AND(g9264, g20352)
--	g21355 = AND(g9613, g20354)
--	g21356 = AND(g9488, g20355)
--	g21357 = AND(g9407, g20356)
--	g21360 = AND(g9507, g20361)
--	g21361 = AND(g9150, g20362)
--	g21362 = AND(g15096, g20363)
--	g21363 = AND(g15022, g20364)
--	g21367 = AND(g9203, g20366)
--	g21368 = AND(g9174, g20367)
--	g21369 = AND(g15188, g20368)
--	g21370 = AND(g9326, g20369)
--	g21371 = AND(g9264, g20370)
--	g21372 = AND(g9216, g20371)
--	g21373 = AND(g9488, g20372)
--	g21374 = AND(g9407, g20373)
--	g21375 = AND(g9342, g20374)
--	g21378 = AND(g9507, g20378)
--	g21379 = AND(g9427, g20379)
--	g21380 = AND(g15096, g20380)
--	g21381 = AND(g15022, g20381)
--	g21388 = AND(g6201, g19657)
--	g21389 = AND(g9649, g20384)
--	g21390 = AND(g9174, g20385)
--	g21391 = AND(g15188, g20386)
--	g21392 = AND(g15118, g20387)
--	g21393 = AND(g9264, g20389)
--	g21394 = AND(g9216, g20390)
--	g21395 = AND(g15274, g20391)
--	g21396 = AND(g9407, g20392)
--	g21397 = AND(g9342, g20393)
--	g21398 = AND(g9277, g20394)
--	g21401 = AND(g9507, g20397)
--	g21402 = AND(g9427, g20398)
--	g21403 = AND(g15022, g20399)
--	g21410 = AND(g6363, g20402)
--	g21411 = AND(g9649, g20403)
--	g21412 = AND(g9569, g20404)
--	g21413 = AND(g15188, g20405)
--	g21414 = AND(g15118, g20406)
--	g21418 = AND(g6290, g19705)
--	g21419 = AND(g9795, g20409)
--	g21420 = AND(g9216, g20410)
--	g21421 = AND(g15274, g20411)
--	g21422 = AND(g15210, g20412)
--	g21423 = AND(g9342, g20414)
--	g21424 = AND(g9277, g20415)
--	g21425 = AND(g15366, g20416)
--	g21428 = AND(g9427, g20420)
--	g21438 = AND(g9649, g20422)
--	g21439 = AND(g9569, g20423)
--	g21440 = AND(g15118, g20424)
--	g21444 = AND(g6568, g20427)
--	g21445 = AND(g9795, g20428)
--	g21446 = AND(g9711, g20429)
--	g21447 = AND(g15274, g20430)
--	g21448 = AND(g15210, g20431)
--	g21452 = AND(g6427, g19749)
--	g21453 = AND(g9941, g20434)
--	g21454 = AND(g9277, g20435)
--	g21455 = AND(g15366, g20436)
--	g21456 = AND(g15296, g20437)
--	g21476 = AND(g9569, g20442)
--	g21480 = AND(g9795, g20444)
--	g21481 = AND(g9711, g20445)
--	g21482 = AND(g15210, g20446)
--	g21486 = AND(g6832, g20449)
--	g21487 = AND(g9941, g20450)
--	g21488 = AND(g9857, g20451)
--	g21489 = AND(g15366, g20452)
--	g21490 = AND(g15296, g20453)
--	g21494 = AND(g6632, g19792)
--	g21497 = AND(g3006, g20456)
--	g21517 = AND(g9711, g20461)
--	g21521 = AND(g9941, g20463)
--	g21522 = AND(g9857, g20464)
--	g21523 = AND(g15296, g20465)
--	g21527 = AND(g7134, g20468)
--	I28068 = AND(g17802, g18265, g17882)
--	g21533 = AND(g17724, g18179, g19799, I28068)
--	g21553 = AND(g9857, g20476)
--	I28096 = AND(g13907, g14238, g13946)
--	g21564 = AND(g13886, g14153, g19799, I28096)
--	I28103 = AND(g17914, g18358, g17993)
--	g21569 = AND(g17825, g18286, g19843, I28103)
--	g21589 = AND(g3002, g19890)
--	g21593 = AND(g16498, g19484, g14071)
--	I28126 = AND(g13963, g14360, g14016)
--	g21597 = AND(g13927, g14268, g19843, I28126)
--	I28133 = AND(g18025, g18453, g18110)
--	g21602 = AND(g17937, g18379, g19876, I28133)
--	g21610 = AND(g7522, g20490)
--	g21611 = AND(g7471, g19915)
--	g21622 = AND(g16520, g19505, g14186)
--	I28155 = AND(g14033, g14472, g14107)
--	g21626 = AND(g13983, g14390, g19876, I28155)
--	I28162 = AND(g18142, g18526, g18226)
--	g21631 = AND(g18048, g18474, g19907, I28162)
--	g21635 = AND(g7549, g20496)
--	g21639 = AND(g3398, g20500)
--	g21650 = AND(g16551, g19524, g14301)
--	I28181 = AND(g14124, g14559, g14222)
--	g21654 = AND(g14053, g14502, g19907, I28181)
--	g21658 = AND(g2896, g20501)
--	g21666 = AND(g3398, g20504)
--	g21670 = AND(g3554, g20505)
--	g21681 = AND(g16583, g19534, g14423)
--	g21687 = AND(g3398, g20516)
--	g21695 = AND(g3554, g20517)
--	g21699 = AND(g3710, g20518)
--	g21707 = AND(g2892, g19978)
--	g21723 = AND(g3554, g20534)
--	g21731 = AND(g3710, g20535)
--	g21735 = AND(g3866, g20536)
--	g21749 = AND(g3710, g20553)
--	g21757 = AND(g3866, g20554)
--	g21758 = AND(g7607, g20045)
--	g21773 = AND(g3866, g19078)
--	g21805 = AND(g16679, g19578, g14776)
--	g21812 = AND(g16705, g19608, g14811)
--	g21818 = AND(g16736, g19641, g14863)
--	g21822 = AND(g16778, g19681, g14936)
--	g21891 = AND(g19302, g11749)
--	g21892 = AND(g19288, g13011)
--	g21899 = AND(g19323, g11749)
--	g21900 = AND(g19306, g13011)
--	g21906 = AND(g5715, g20513)
--	g21911 = AND(g19350, g11749)
--	g21912 = AND(g19327, g13011)
--	g21913 = AND(g4456, g20519)
--	g21920 = AND(g5773, g20531)
--	g21925 = AND(g19384, g11749)
--	g21926 = AND(g19354, g13011)
--	g21931 = AND(g4632, g20539)
--	g21938 = AND(g5832, g20550)
--	g21990 = AND(g291, g21187)
--	g22004 = AND(g978, g21202)
--	g22015 = AND(g1672, g21217)
--	g22020 = AND(g2366, g21225)
--	I28582 = AND(g19141, g21133, g21116)
--	g22036 = AND(g21104, g21095, g21084, I28582)
--	I28594 = AND(g21167, g21147, g21134)
--	g22046 = AND(g21117, g21105, g21096, I28594)
--	I28609 = AND(g21183, g21168, g21148)
--	g22062 = AND(g21135, g21118, g21106, I28609)
--	g22187 = AND(g21564, g20986)
--	g22196 = AND(g21597, g21012)
--	g22201 = AND(g21271, g16881)
--	g22202 = AND(g21626, g21036)
--	g22206 = AND(g21895, g11976)
--	g22207 = AND(g21278, g16910)
--	g22208 = AND(g21654, g21057)
--	g22211 = AND(g21661, g12027)
--	g22214 = AND(g21907, g12045)
--	g22215 = AND(g21285, g16940)
--	g22220 = AND(g21690, g12091)
--	g22223 = AND(g21921, g12109)
--	g22224 = AND(g21293, g16971)
--	g22228 = AND(g21716, g12136)
--	g22229 = AND(g21661, g12139)
--	g22235 = AND(g21726, g12163)
--	g22238 = AND(g21939, g12181)
--	g22244 = AND(g21742, g12198)
--	g22245 = AND(g21690, g12201)
--	g22250 = AND(g21752, g12225)
--	g22254 = AND(g21716, g12239)
--	g22255 = AND(g21661, g12242)
--	g22264 = AND(g21766, g12253)
--	g22265 = AND(g21726, g12256)
--	g22270 = AND(g92, g21529)
--	g22272 = AND(g21742, g12282)
--	g22273 = AND(g21690, g12285)
--	g22281 = AND(g21782, g12296)
--	g22282 = AND(g21752, g12299)
--	g22285 = AND(g21716, g12312)
--	g22289 = AND(g780, g21565)
--	g22291 = AND(g21766, g12318)
--	g22292 = AND(g21726, g12321)
--	g22305 = AND(g21742, g12340)
--	g22309 = AND(g1466, g21598)
--	g22311 = AND(g21782, g12346)
--	g22312 = AND(g21752, g12349)
--	g22333 = AND(g21766, g12370)
--	g22337 = AND(g2160, g21627)
--	g22340 = AND(g88, g21184)
--	g22358 = AND(g21782, g12389)
--	g22363 = AND(g776, g21199)
--	g22383 = AND(g1462, g21214)
--	g22398 = AND(g2156, g21222)
--	g22483 = AND(g646, g21861)
--	g22515 = AND(g13873, g21382)
--	g22516 = AND(g20885, g17442)
--	g22517 = AND(g21895, g12608)
--	g22526 = AND(g1332, g21867)
--	g22546 = AND(g13886, g21404)
--	g22555 = AND(g13895, g21415)
--	g22556 = AND(g20904, g17523)
--	g22557 = AND(g21907, g12654)
--	g22566 = AND(g2026, g21872)
--	g22577 = AND(g13907, g21429)
--	g22581 = AND(g21895, g12699)
--	g22587 = AND(g13927, g21441)
--	g22595 = AND(g13936, g21449)
--	g22596 = AND(g20928, g17613)
--	g22597 = AND(g21921, g12708)
--	g22606 = AND(g2720, g21876)
--	g22607 = AND(g13946, g21458)
--	g22610 = AND(g660, g21473)
--	g22614 = AND(g13963, g21477)
--	g22618 = AND(g21907, g12756)
--	g22624 = AND(g13983, g21483)
--	g22632 = AND(g13992, g21491)
--	g22633 = AND(g20956, g17710)
--	g22634 = AND(g21939, g12765)
--	g22637 = AND(g20841, g10927)
--	g22638 = AND(g14001, g21498)
--	g22643 = AND(g14016, g21505)
--	g22646 = AND(g1346, g21514)
--	g22650 = AND(g14033, g21518)
--	g22654 = AND(g21921, g12798)
--	g22660 = AND(g14053, g21524)
--	g22665 = AND(g20920, g6153)
--	g22666 = AND(g21825, g20014)
--	g22667 = AND(g14062, g21530)
--	g22674 = AND(g14092, g21537)
--	g22679 = AND(g14107, g21541)
--	g22682 = AND(g2040, g21550)
--	g22686 = AND(g14124, g21554)
--	g22690 = AND(g21939, g12837)
--	g22699 = AND(g7338, g21883)
--	g22700 = AND(g7146, g21558)
--	g22701 = AND(g18174, g21561)
--	g22707 = AND(g14177, g21566)
--	g22714 = AND(g14207, g21573)
--	g22719 = AND(g14222, g21577)
--	g22722 = AND(g2734, g21586)
--	g22726 = AND(g3036, g21886)
--	g22727 = AND(g14238, g21590)
--	g22732 = AND(g18281, g21594)
--	g22738 = AND(g14292, g21599)
--	g22745 = AND(g14322, g21606)
--	g22754 = AND(g14342, g21612)
--	g22759 = AND(g14360, g21619)
--	g22764 = AND(g18374, g21623)
--	g22770 = AND(g14414, g21628)
--	g22788 = AND(g14454, g21640)
--	g22793 = AND(g14472, g21647)
--	g22798 = AND(g18469, g21651)
--	g22804 = AND(g2920, g21655)
--	g22830 = AND(g14541, g21671)
--	g22835 = AND(g14559, g21678)
--	g22841 = AND(g7583, g21902)
--	g22842 = AND(g3032, g21682)
--	g22869 = AND(g14596, g21700)
--	g22874 = AND(g7587, g21708)
--	g22906 = AND(g2924, g21927)
--	g22984 = AND(g16840, g21400)
--	g23104 = AND(g20842, g15859)
--	g23106 = AND(g5857, g21050)
--	g23118 = AND(g20850, g15890)
--	g23119 = AND(g5904, g21069)
--	g23127 = AND(g20858, g15923)
--	g23128 = AND(g5943, g21079)
--	g23138 = AND(g20866, g15952)
--	g23139 = AND(g5977, g21093)
--	g23409 = AND(g21533, g22408)
--	g23414 = AND(g21569, g22421)
--	g23419 = AND(g22755, g19577)
--	g23423 = AND(g21602, g22443)
--	g23428 = AND(g22789, g19607)
--	g23432 = AND(g21631, g22476)
--	g23434 = AND(g22831, g19640)
--	g23440 = AND(g22870, g19680)
--	g23451 = AND(g18552, g22547)
--	g23458 = AND(g18602, g22588)
--	g23462 = AND(g17988, g22609)
--	g23467 = AND(g18634, g22625)
--	g23471 = AND(g18105, g22645)
--	g23476 = AND(g18643, g22661)
--	g23483 = AND(g22945, g8847)
--	g23484 = AND(g18221, g22681)
--	g23494 = AND(g18328, g22721)
--	g23496 = AND(g5802, g22300)
--	g23510 = AND(g5890, g22753)
--	g23512 = AND(g5858, g22328)
--	g23525 = AND(g5929, g22787)
--	g23527 = AND(g5905, g22353)
--	g23536 = AND(g5963, g22829)
--	g23538 = AND(g5944, g22376)
--	g23544 = AND(g5992, g22868)
--	g23547 = AND(g8062, g22405)
--	g23550 = AND(g8132, g22409)
--	g23551 = AND(g8135, g22412)
--	g23552 = AND(g6136, g22415)
--	g23554 = AND(g8147, g22418)
--	g23558 = AND(g8200, g22422)
--	g23559 = AND(g8203, g22425)
--	g23560 = AND(g8206, g22428)
--	g23563 = AND(g8218, g22431)
--	g23564 = AND(g8221, g22434)
--	g23565 = AND(g6146, g22437)
--	g23567 = AND(g8233, g22440)
--	g23571 = AND(g3931, g22445)
--	g23572 = AND(g3934, g22448)
--	g23573 = AND(g3937, g22451)
--	g23577 = AND(g3957, g22455)
--	g23578 = AND(g3960, g22458)
--	g23579 = AND(g3963, g22461)
--	g23582 = AND(g3975, g22464)
--	g23583 = AND(g3978, g22467)
--	g23584 = AND(g6167, g22470)
--	g23586 = AND(g3990, g22473)
--	g23590 = AND(g4009, g22477)
--	g23591 = AND(g4012, g22480)
--	g23592 = AND(g17640, g22986)
--	g23593 = AND(g22845, g20365)
--	g23598 = AND(g4038, g22484)
--	g23599 = AND(g4041, g22487)
--	g23600 = AND(g4044, g22490)
--	g23604 = AND(g4064, g22494)
--	g23605 = AND(g4067, g22497)
--	g23606 = AND(g4070, g22500)
--	g23609 = AND(g4082, g22503)
--	g23610 = AND(g4085, g22506)
--	g23611 = AND(g6194, g22509)
--	g23615 = AND(g4107, g22512)
--	g23616 = AND(g17724, g22988)
--	g23617 = AND(g22810, g20382)
--	g23618 = AND(g22608, g20383)
--	g23622 = AND(g4136, g22520)
--	g23623 = AND(g4139, g22523)
--	g23624 = AND(g17741, g22989)
--	g23625 = AND(g22880, g20388)
--	g23630 = AND(g4165, g22527)
--	g23631 = AND(g4168, g22530)
--	g23632 = AND(g4171, g22533)
--	g23636 = AND(g4191, g22537)
--	g23637 = AND(g4194, g22540)
--	g23638 = AND(g4197, g22543)
--	g23639 = AND(g21825, g22805)
--	g23643 = AND(g17802, g22991)
--	g23659 = AND(g22784, g17500)
--	g23664 = AND(g4246, g22552)
--	g23665 = AND(g17825, g22995)
--	g23666 = AND(g22851, g20407)
--	g23667 = AND(g22644, g20408)
--	g23671 = AND(g4275, g22560)
--	g23672 = AND(g4278, g22563)
--	g23673 = AND(g17842, g22996)
--	g23674 = AND(g22915, g20413)
--	g23679 = AND(g4304, g22567)
--	g23680 = AND(g4307, g22570)
--	g23681 = AND(g4310, g22573)
--	g23686 = AND(g17882, g22998)
--	g23687 = AND(g22668, g17570)
--	g23689 = AND(g6513, g23001)
--	g23693 = AND(g17914, g23002)
--	g23709 = AND(g22826, g17591)
--	g23714 = AND(g4401, g22592)
--	g23715 = AND(g17937, g23006)
--	g23716 = AND(g22886, g20432)
--	g23717 = AND(g22680, g20433)
--	g23721 = AND(g4430, g22600)
--	g23722 = AND(g4433, g22603)
--	g23723 = AND(g17954, g23007)
--	g23724 = AND(g22940, g20438)
--	g23726 = AND(g21825, g22843)
--	g23734 = AND(g17974, g23008)
--	g23735 = AND(g22949, g9450)
--	g23740 = AND(g17993, g23012)
--	g23741 = AND(g22708, g17667)
--	g23743 = AND(g6777, g23015)
--	g23747 = AND(g18025, g23016)
--	g23763 = AND(g22865, g17688)
--	g23768 = AND(g4570, g22629)
--	g23769 = AND(g18048, g23020)
--	g23770 = AND(g22921, g20454)
--	g23771 = AND(g22720, g20455)
--	g23772 = AND(g21825, g22875)
--	g23776 = AND(g18074, g23021)
--	g23777 = AND(g22949, g9528)
--	g23778 = AND(g22954, g9531)
--	g23789 = AND(g18091, g23024)
--	g23790 = AND(g22958, g9592)
--	g23795 = AND(g18110, g23028)
--	g23796 = AND(g22739, g17767)
--	g23798 = AND(g7079, g23031)
--	g23802 = AND(g18142, g23032)
--	g23818 = AND(g22900, g17788)
--	g23820 = AND(g3013, g23036)
--	g23822 = AND(g14148, g23037)
--	g23824 = AND(g22949, g9641)
--	g23825 = AND(g22954, g9644)
--	g23829 = AND(g18190, g23038)
--	g23830 = AND(g22958, g9670)
--	g23831 = AND(g22962, g9673)
--	g23842 = AND(g18207, g23041)
--	g23843 = AND(g22966, g9734)
--	g23848 = AND(g18226, g23045)
--	g23849 = AND(g22771, g17868)
--	g23851 = AND(g7329, g23048)
--	g23852 = AND(g19179, g22696)
--	g23854 = AND(g18265, g23049)
--	g23855 = AND(g22954, g9767)
--	g23857 = AND(g14263, g23056)
--	g23859 = AND(g22958, g9787)
--	g23860 = AND(g22962, g9790)
--	g23864 = AND(g18297, g23057)
--	g23865 = AND(g22966, g9816)
--	g23866 = AND(g22971, g9819)
--	g23877 = AND(g18314, g23060)
--	g23878 = AND(g22975, g9880)
--	g23886 = AND(g18341, g23064)
--	g23888 = AND(g18358, g23069)
--	g23889 = AND(g22962, g9913)
--	g23891 = AND(g14385, g23074)
--	g23893 = AND(g22966, g9933)
--	g23894 = AND(g22971, g9936)
--	g23898 = AND(g18390, g23075)
--	g23899 = AND(g22975, g9962)
--	g23900 = AND(g22980, g9965)
--	g23904 = AND(g3010, g22750)
--	g23907 = AND(g18436, g23079)
--	g23909 = AND(g18453, g23082)
--	g23910 = AND(g22971, g10067)
--	g23912 = AND(g14497, g23087)
--	g23914 = AND(g22975, g10087)
--	g23915 = AND(g22980, g10090)
--	g23917 = AND(g7545, g23088)
--	g23939 = AND(g18509, g23095)
--	g23941 = AND(g18526, g23098)
--	g23942 = AND(g22980, g10176)
--	g23944 = AND(g7570, g23103)
--	g23971 = AND(g18573, g23112)
--	g23972 = AND(g2903, g23115)
--	g24029 = AND(g2900, g22903)
--	g24211 = AND(g22014, g10969)
--	g24217 = AND(g22825, g10999)
--	g24221 = AND(g22979, g11042)
--	g24224 = AND(g22219, g11045)
--	g24229 = AND(g22232, g11105)
--	g24236 = AND(g22243, g11157)
--	g24241 = AND(g22259, g11228)
--	g24246 = AND(g21982, g11291)
--	g24247 = AND(g22551, g11297)
--	g24253 = AND(g21995, g11370)
--	g24256 = AND(g22003, g11438)
--	g24427 = AND(g17086, g24134, g13626)
--	g24429 = AND(g24115, g13614)
--	g24431 = AND(g17124, g24153, g13637)
--	g24432 = AND(g14642, g15904, g24115)
--	g24433 = AND(g24134, g13626)
--	g24435 = AND(g17151, g24168, g13649)
--	g24436 = AND(g14669, g15933, g24134)
--	g24437 = AND(g24153, g13637)
--	g24439 = AND(g14703, g15962, g24153)
--	g24440 = AND(g24168, g13649)
--	g24441 = AND(g14737, g15981, g24168)
--	g24478 = AND(g23545, g21119, g21227)
--	g24529 = AND(g19933, g17896, g23403)
--	g24540 = AND(g18548, g23089, g23403)
--	g24541 = AND(g23420, g17896, g23052)
--	g24542 = AND(g19950, g18007, g23410)
--	g24550 = AND(g18548, g23420, g19948)
--	g24552 = AND(g18598, g23107, g23410)
--	g24553 = AND(g23429, g18007, g23071)
--	g24554 = AND(g19977, g18124, g23415)
--	g24559 = AND(g79, g23448)
--	g24561 = AND(g18598, g23429, g19975)
--	g24563 = AND(g18630, g23120, g23415)
--	g24564 = AND(g23435, g18124, g23084)
--	g24565 = AND(g20007, g18240, g23424)
--	g24569 = AND(g767, g23455)
--	g24571 = AND(g18630, g23435, g20005)
--	g24573 = AND(g18639, g23129, g23424)
--	g24574 = AND(g23441, g18240, g23100)
--	g24578 = AND(g1453, g23464)
--	g24580 = AND(g18639, g23441, g20043)
--	g24585 = AND(g2147, g23473)
--	g24590 = AND(g23486, g23478)
--	g24591 = AND(g83, g23853)
--	g24595 = AND(g23502, g23489)
--	g24596 = AND(g771, g23887)
--	g24603 = AND(g23518, g23505)
--	g24604 = AND(g1457, g23908)
--	g24610 = AND(g23533, g23521)
--	g24611 = AND(g2151, g23940)
--	g24644 = AND(g17203, g24115)
--	g24664 = AND(g17208, g24134)
--	g24676 = AND(g13568, g24115)
--	g24683 = AND(g17214, g24153)
--	g24695 = AND(g13576, g24134)
--	g24700 = AND(g17217, g24168)
--	g24712 = AND(g13585, g24153)
--	g24723 = AND(g13605, g24168)
--	g24745 = AND(g15454, g24096)
--	g24746 = AND(g15454, g24098)
--	g24747 = AND(g9427, g24099)
--	g24748 = AND(g672, g24101)
--	g24749 = AND(g15540, g24102)
--	g24750 = AND(g15454, g24104)
--	g24751 = AND(g9427, g24105)
--	g24752 = AND(g9507, g24106)
--	g24754 = AND(g15540, g24107)
--	g24755 = AND(g9569, g24108)
--	g24757 = AND(g1358, g24110)
--	g24758 = AND(g15618, g24111)
--	g24759 = AND(g21825, g23885)
--	g24760 = AND(g9427, g24112)
--	g24761 = AND(g9507, g24113)
--	g24762 = AND(g12876, g24114)
--	g24767 = AND(g15540, g24121)
--	g24768 = AND(g9569, g24122)
--	g24769 = AND(g9649, g24123)
--	g24772 = AND(g15618, g24124)
--	g24773 = AND(g9711, g24125)
--	g24774 = AND(g2052, g24127)
--	g24775 = AND(g15694, g24128)
--	g24776 = AND(g9507, g24129)
--	g24777 = AND(g12876, g24130)
--	g24779 = AND(g9569, g24131)
--	g24780 = AND(g9649, g24132)
--	g24781 = AND(g12916, g24133)
--	g24788 = AND(g15618, g24140)
--	g24789 = AND(g9711, g24141)
--	g24790 = AND(g9795, g24142)
--	g24792 = AND(g15694, g24143)
--	g24793 = AND(g9857, g24144)
--	g24794 = AND(g2746, g24146)
--	g24795 = AND(g12017, g24232)
--	g24796 = AND(g12876, g24147)
--	g24798 = AND(g9649, g24148)
--	g24799 = AND(g12916, g24149)
--	g24802 = AND(g9711, g24150)
--	g24803 = AND(g9795, g24151)
--	g24804 = AND(g12945, g24152)
--	g24809 = AND(g15694, g24159)
--	g24810 = AND(g9857, g24160)
--	g24811 = AND(g9941, g24161)
--	g24813 = AND(g21825, g23905)
--	g24818 = AND(g12916, g24162)
--	g24821 = AND(g9795, g24163)
--	g24822 = AND(g12945, g24164)
--	g24824 = AND(g9857, g24165)
--	g24825 = AND(g9941, g24166)
--	g24826 = AND(g12974, g24167)
--	g24831 = AND(g24100, g20401)
--	g24838 = AND(g12945, g24175)
--	g24840 = AND(g9941, g24176)
--	g24841 = AND(g12974, g24177)
--	g24843 = AND(g21825, g23918)
--	g24846 = AND(g24109, g20426)
--	g24853 = AND(g12974, g24180)
--	g24855 = AND(g18174, g23731)
--	g24858 = AND(g24047, g18873)
--	g24861 = AND(g24126, g20448)
--	g24867 = AND(g666, g23779)
--	g24869 = AND(g24047, g18894)
--	g24870 = AND(g18281, g23786)
--	g24874 = AND(g24060, g18899)
--	g24876 = AND(g24145, g20467)
--	g24878 = AND(g19830, g24210)
--	g24881 = AND(g24047, g18912)
--	g24882 = AND(g1352, g23832)
--	g24884 = AND(g24060, g18917)
--	g24885 = AND(g18374, g23839)
--	g24888 = AND(g24073, g18922)
--	g24898 = AND(g24060, g18931)
--	g24899 = AND(g2046, g23867)
--	g24901 = AND(g24073, g18936)
--	g24902 = AND(g18469, g23874)
--	g24905 = AND(g24084, g18941)
--	g24906 = AND(g18886, g23879)
--	g24907 = AND(g7466, g24220)
--	g24908 = AND(g7342, g23882)
--	g24921 = AND(g24073, g18951)
--	g24922 = AND(g2740, g23901)
--	g24924 = AND(g24084, g18956)
--	g24938 = AND(g24084, g18967)
--	g24964 = AND(g7595, g24251)
--	g24974 = AND(g7600, g24030)
--	g25086 = AND(g23444, g10880)
--	g25102 = AND(g23444, g10915)
--	g25117 = AND(g23444, g10974)
--	g25128 = AND(g17051, g24115, g13614)
--	g25178 = AND(g24623, g20634)
--	g25181 = AND(g24636, g20673)
--	g25182 = AND(g24681, g20676)
--	g25184 = AND(g24694, g20735)
--	g25187 = AND(g24633, g16608)
--	g25188 = AND(g24652, g20763)
--	g25192 = AND(g24711, g20790)
--	g25193 = AND(g24653, g16626)
--	g25196 = AND(g24672, g16640)
--	g25198 = AND(g24691, g16651)
--	g25269 = AND(g24648, g8700)
--	g25277 = AND(g24648, g8714)
--	g25278 = AND(g24668, g8719)
--	g25281 = AND(g5606, g24815)
--	g25282 = AND(g24648, g8748)
--	g25286 = AND(g24668, g8752)
--	g25287 = AND(g24687, g8757)
--	g25289 = AND(g5631, g24834)
--	g25290 = AND(g24668, g8771)
--	g25294 = AND(g24687, g8775)
--	g25295 = AND(g24704, g8780)
--	g25299 = AND(g5659, g24850)
--	g25300 = AND(g24687, g8794)
--	g25304 = AND(g24704, g8798)
--	g25309 = AND(g5697, g24864)
--	g25310 = AND(g24704, g8813)
--	g25318 = AND(g24682, g19358, g19335)
--	g25321 = AND(g25075, g9669)
--	g25328 = AND(g24644, g17892)
--	g25334 = AND(g24644, g17984)
--	g25337 = AND(g24664, g18003)
--	g25342 = AND(g5851, g24600)
--	g25346 = AND(g24644, g18084)
--	g25348 = AND(g24664, g18101)
--	g25351 = AND(g24683, g18120)
--	g25356 = AND(g5898, g24607)
--	g25360 = AND(g24664, g18200)
--	g25362 = AND(g24683, g18217)
--	g25365 = AND(g24700, g18236)
--	g25371 = AND(g5937, g24619)
--	g25375 = AND(g24683, g18307)
--	g25377 = AND(g24700, g18324)
--	g25388 = AND(g5971, g24630)
--	g25392 = AND(g24700, g18400)
--	g25453 = AND(g6142, g24763)
--	g25457 = AND(g6163, g24784)
--	g25461 = AND(g6190, g24805)
--	g25466 = AND(g6222, g24827)
--	g25470 = AND(g24479, g20400)
--	g25475 = AND(g14148, g25087)
--	g25482 = AND(g24480, g17567)
--	g25483 = AND(g24481, g20421)
--	g25487 = AND(g24485, g20425)
--	g25505 = AND(g6707, g25094)
--	g25506 = AND(g14263, g25095)
--	g25513 = AND(g24487, g17664)
--	g25514 = AND(g24488, g20443)
--	g25518 = AND(g24489, g20447)
--	g25552 = AND(g7009, g25104)
--	g25553 = AND(g14385, g25105)
--	g25560 = AND(g24494, g17764)
--	g25561 = AND(g24495, g20462)
--	g25565 = AND(g24496, g20466)
--	g25618 = AND(g7259, g25110)
--	g25619 = AND(g14497, g25111)
--	g25626 = AND(g24504, g17865)
--	g25627 = AND(g24505, g20477)
--	g25628 = AND(g21008, g25115)
--	g25629 = AND(g3024, g25116)
--	g25697 = AND(g7455, g25120)
--	g25881 = AND(g2908, g25126)
--	g25951 = AND(g24800, g13670)
--	g25953 = AND(g24783, g13699)
--	g25957 = AND(g24782, g11869)
--	g25961 = AND(g24770, g11901)
--	g25963 = AND(g24756, g11944)
--	g25968 = AND(g24871, g11986)
--	g25972 = AND(g24859, g12042)
--	g25973 = AND(g24847, g13838)
--	g25975 = AND(g24606, g21917)
--	g25977 = AND(g24845, g12089)
--	g25978 = AND(g24836, g13850)
--	g25980 = AND(g24663, g21928)
--	g25981 = AND(g24819, g13858)
--	g26023 = AND(g25422, g24912)
--	g26024 = AND(g25301, g21102)
--	g26026 = AND(g25431, g24929)
--	g26027 = AND(g25418, g22271)
--	g26028 = AND(g25438, g24941)
--	g26029 = AND(g25445, g24952)
--	g26030 = AND(g25429, g22304)
--	g26032 = AND(g25379, g19415)
--	g26033 = AND(g25395, g19452)
--	g26034 = AND(g25405, g19479)
--	g26035 = AND(g25523, g19483)
--	g26036 = AND(g25413, g19502)
--	g26038 = AND(g25589, g19504)
--	g26039 = AND(g25668, g19523)
--	g26040 = AND(g25745, g19533)
--	g26051 = AND(g70, g25296)
--	g26052 = AND(g25941, g21087)
--	g26053 = AND(g758, g25306)
--	g26054 = AND(g25944, g21099)
--	g26060 = AND(g25943, g21108)
--	g26061 = AND(g1444, g25315)
--	g26062 = AND(g25947, g21113)
--	g26067 = AND(g25946, g21125)
--	g26068 = AND(g2138, g25324)
--	g26069 = AND(g25949, g21130)
--	g26074 = AND(g25948, g21144)
--	g26075 = AND(g74, g25698)
--	g26080 = AND(g25950, g21164)
--	g26082 = AND(g762, g25771)
--	g26085 = AND(g1448, g25825)
--	g26091 = AND(g2142, g25860)
--	g26157 = AND(g21825, g25630)
--	g26158 = AND(g679, g25937)
--	g26163 = AND(g1365, g25939)
--	g26166 = AND(g686, g25454)
--	g26171 = AND(g2059, g25942)
--	g26186 = AND(g1372, g25458)
--	g26188 = AND(g2753, g25945)
--	g26207 = AND(g2066, g25463)
--	g26212 = AND(g4217, g25467)
--	g26213 = AND(g25895, g9306)
--	g26231 = AND(g2760, g25472)
--	g26233 = AND(g4340, g25476)
--	g26234 = AND(g4343, g25479)
--	g26235 = AND(g25895, g9368)
--	g26236 = AND(g25899, g9371)
--	g26243 = AND(g4372, g25484)
--	g26244 = AND(g25903, g9387)
--	g26257 = AND(g4465, g25493)
--	g26258 = AND(g4468, g25496)
--	g26259 = AND(g4471, g25499)
--	g26260 = AND(g25254, g17649)
--	g26261 = AND(g25895, g9443)
--	g26262 = AND(g25899, g9446)
--	g26263 = AND(g4476, g25502)
--	g26268 = AND(g4509, g25507)
--	g26269 = AND(g4512, g25510)
--	g26270 = AND(g25903, g9465)
--	g26271 = AND(g25907, g9468)
--	g26278 = AND(g4541, g25515)
--	g26279 = AND(g25911, g9484)
--	g26288 = AND(g4592, g25524)
--	g26289 = AND(g4595, g25527)
--	g26290 = AND(g4598, g25530)
--	g26291 = AND(g25899, g9524)
--	g26292 = AND(g4603, g25533)
--	g26293 = AND(g4606, g25536)
--	g26298 = AND(g4641, g25540)
--	g26299 = AND(g4644, g25543)
--	g26300 = AND(g4647, g25546)
--	g26301 = AND(g25258, g17749)
--	g26302 = AND(g25903, g9585)
--	g26303 = AND(g25907, g9588)
--	g26307 = AND(g4652, g25549)
--	g26309 = AND(g4685, g25554)
--	g26310 = AND(g4688, g25557)
--	g26311 = AND(g25911, g9607)
--	g26312 = AND(g25915, g9610)
--	g26316 = AND(g4717, g25562)
--	g26317 = AND(g25919, g9626)
--	g26318 = AND(g4737, g25573)
--	g26319 = AND(g4740, g25576)
--	g26324 = AND(g4743, g25579)
--	g26325 = AND(g4746, g25582)
--	g26326 = AND(g4749, g25585)
--	g26332 = AND(g4769, g25590)
--	g26333 = AND(g4772, g25593)
--	g26334 = AND(g4775, g25596)
--	g26335 = AND(g25907, g9666)
--	g26339 = AND(g4780, g25599)
--	g26340 = AND(g4783, g25602)
--	g26342 = AND(g4818, g25606)
--	g26343 = AND(g4821, g25609)
--	g26344 = AND(g4824, g25612)
--	g26345 = AND(g25261, g17850)
--	g26346 = AND(g25911, g9727)
--	g26347 = AND(g25915, g9730)
--	g26348 = AND(g4829, g25615)
--	g26350 = AND(g4862, g25620)
--	g26351 = AND(g4865, g25623)
--	g26352 = AND(g25919, g9749)
--	g26353 = AND(g25923, g9752)
--	g26357 = AND(g4882, g25634)
--	g26361 = AND(g4888, g25637)
--	g26362 = AND(g4891, g25640)
--	g26363 = AND(g4894, g25643)
--	g26365 = AND(g4913, g25652)
--	g26366 = AND(g4916, g25655)
--	g26371 = AND(g4919, g25658)
--	g26372 = AND(g4922, g25661)
--	g26373 = AND(g4925, g25664)
--	g26379 = AND(g4945, g25669)
--	g26380 = AND(g4948, g25672)
--	g26381 = AND(g4951, g25675)
--	g26382 = AND(g25915, g9812)
--	g26383 = AND(g4956, g25678)
--	g26384 = AND(g4959, g25681)
--	g26386 = AND(g4994, g25685)
--	g26387 = AND(g4997, g25688)
--	g26388 = AND(g5000, g25691)
--	g26389 = AND(g25264, g17962)
--	g26390 = AND(g25919, g9873)
--	g26391 = AND(g25923, g9876)
--	g26392 = AND(g5005, g25694)
--	g26396 = AND(g5027, g25700)
--	g26397 = AND(g5030, g25703)
--	g26400 = AND(g5041, g25711)
--	g26404 = AND(g5047, g25714)
--	g26405 = AND(g5050, g25717)
--	g26406 = AND(g5053, g25720)
--	g26408 = AND(g5072, g25729)
--	g26409 = AND(g5075, g25732)
--	g26414 = AND(g5078, g25735)
--	g26415 = AND(g5081, g25738)
--	g26416 = AND(g5084, g25741)
--	g26422 = AND(g5104, g25746)
--	g26423 = AND(g5107, g25749)
--	g26424 = AND(g5110, g25752)
--	g26425 = AND(g25923, g9958)
--	g26426 = AND(g5115, g25755)
--	g26427 = AND(g5118, g25758)
--	g26432 = AND(g5145, g25767)
--	g26437 = AND(g5156, g25773)
--	g26438 = AND(g5159, g25776)
--	g26441 = AND(g5170, g25784)
--	g26445 = AND(g5176, g25787)
--	g26446 = AND(g5179, g25790)
--	g26447 = AND(g5182, g25793)
--	g26449 = AND(g5201, g25802)
--	g26450 = AND(g5204, g25805)
--	g26455 = AND(g5207, g25808)
--	g26456 = AND(g5210, g25811)
--	g26457 = AND(g5213, g25814)
--	g26464 = AND(g5238, g25821)
--	g26469 = AND(g5249, g25827)
--	g26470 = AND(g5252, g25830)
--	g26473 = AND(g5263, g25838)
--	g26477 = AND(g5269, g25841)
--	g26478 = AND(g5272, g25844)
--	g26479 = AND(g5275, g25847)
--	g26488 = AND(g5301, g25856)
--	g26493 = AND(g5312, g25862)
--	g26494 = AND(g5315, g25865)
--	g26504 = AND(g5338, g25877)
--	g26663 = AND(g25274, g21066)
--	g26668 = AND(g25283, g21076)
--	g26673 = AND(g12431, g25318)
--	g26674 = AND(g25291, g21090)
--	g26754 = AND(g14657, g26508)
--	g26755 = AND(g26083, g22239)
--	g26756 = AND(g26113, g22240)
--	g26758 = AND(g16614, g26521, g13637)
--	g26759 = AND(g26356, g19251)
--	g26760 = AND(g26137, g22256)
--	g26761 = AND(g26154, g22257)
--	g26763 = AND(g14691, g26516)
--	g26764 = AND(g16632, g26525, g13649)
--	g26765 = AND(g26399, g19265)
--	g26766 = AND(g14725, g26521)
--	g26767 = AND(g26087, g22287)
--	g26768 = AND(g26440, g19280)
--	g26769 = AND(g14753, g26525)
--	g26770 = AND(g26059, g19287)
--	g26771 = AND(g24912, g26508, g13614)
--	g26773 = AND(g26145, g22303)
--	g26774 = AND(g26472, g19299)
--	g26775 = AND(g26099, g22318)
--	g26777 = AND(g26066, g19305)
--	g26778 = AND(g24929, g26516, g13626)
--	g26780 = AND(g26119, g16622)
--	g26783 = AND(g26073, g19326)
--	g26784 = AND(g24941, g26521, g13637)
--	g26787 = AND(g26129, g16636)
--	g26790 = AND(g26079, g19353)
--	g26791 = AND(g24952, g26525, g13649)
--	g26794 = AND(g26143, g16647)
--	g26797 = AND(g26148, g16659)
--	g26829 = AND(g5623, g26209)
--	g26833 = AND(g5651, g26237)
--	g26842 = AND(g5689, g26275)
--	g26845 = AND(g5664, g26056)
--	g26851 = AND(g5741, g26313)
--	g26853 = AND(g5716, g26063)
--	g26860 = AND(g5774, g26070)
--	g26866 = AND(g5833, g26076)
--	g26955 = AND(g6157, g26533)
--	g26958 = AND(g6184, g26538)
--	g26961 = AND(g13907, g26175)
--	g26962 = AND(g6180, g26178)
--	g26963 = AND(g6216, g26539)
--	g26965 = AND(g23320, g26540)
--	g26966 = AND(g13963, g26196)
--	g26967 = AND(g6212, g26202)
--	g26968 = AND(g6305, g26542)
--	g26969 = AND(g23320, g26543)
--	g26970 = AND(g21976, g26544)
--	g26971 = AND(g23325, g26546)
--	g26972 = AND(g14033, g26223)
--	g26973 = AND(g6301, g26226)
--	g26977 = AND(g23320, g26550)
--	g26978 = AND(g21976, g26551)
--	g26979 = AND(g23331, g26552)
--	g26980 = AND(g23360, g26554)
--	g26981 = AND(g23325, g26555)
--	g26982 = AND(g21983, g26556)
--	g26984 = AND(g23335, g26558)
--	g26985 = AND(g14124, g26251)
--	g26986 = AND(g6438, g26254)
--	g26993 = AND(g21976, g26561)
--	g26994 = AND(g23331, g26562)
--	g26995 = AND(g21991, g26563)
--	g26996 = AND(g23360, g26564)
--	g26997 = AND(g22050, g26565)
--	g26998 = AND(g23325, g26566)
--	g26999 = AND(g21983, g26567)
--	g27000 = AND(g23340, g26568)
--	g27001 = AND(g23364, g26570)
--	g27002 = AND(g23335, g26571)
--	g27003 = AND(g21996, g26572)
--	g27004 = AND(g23344, g26574)
--	g27005 = AND(g23331, g26578)
--	g27006 = AND(g21991, g26579)
--	g27007 = AND(g23360, g26580)
--	g27008 = AND(g22050, g26581)
--	g27009 = AND(g23368, g26582)
--	g27016 = AND(g21983, g26584)
--	g27017 = AND(g23340, g26585)
--	g27018 = AND(g22005, g26586)
--	g27019 = AND(g23364, g26587)
--	g27020 = AND(g22069, g26588)
--	g27021 = AND(g23335, g26589)
--	g27022 = AND(g21996, g26590)
--	g27023 = AND(g23349, g26591)
--	g27024 = AND(g23372, g26593)
--	g27025 = AND(g23344, g26594)
--	g27026 = AND(g22009, g26595)
--	g27027 = AND(g21991, g26598)
--	g27028 = AND(g22050, g26599)
--	g27029 = AND(g23368, g26600)
--	g27030 = AND(g22083, g26601)
--	g27031 = AND(g23340, g26602)
--	g27032 = AND(g22005, g26603)
--	g27033 = AND(g23364, g26604)
--	g27034 = AND(g22069, g26605)
--	g27035 = AND(g23377, g26606)
--	g27042 = AND(g21996, g26608)
--	g27043 = AND(g23349, g26609)
--	g27044 = AND(g22016, g26610)
--	g27045 = AND(g23372, g26611)
--	g27046 = AND(g22093, g26612)
--	g27047 = AND(g23344, g26613)
--	g27048 = AND(g22009, g26614)
--	g27049 = AND(g23353, g26615)
--	g27050 = AND(g23381, g26617)
--	g27052 = AND(g4885, g26358)
--	g27053 = AND(g23368, g26619)
--	g27054 = AND(g22083, g26620)
--	g27055 = AND(g22005, g26621)
--	g27056 = AND(g22069, g26622)
--	g27057 = AND(g23377, g26623)
--	g27058 = AND(g22108, g26624)
--	g27059 = AND(g23349, g26625)
--	g27060 = AND(g22016, g26626)
--	g27061 = AND(g23372, g26627)
--	g27062 = AND(g22093, g26628)
--	g27063 = AND(g23388, g26629)
--	g27070 = AND(g22009, g26631)
--	g27071 = AND(g23353, g26632)
--	g27072 = AND(g22021, g26633)
--	g27073 = AND(g23381, g26634)
--	g27074 = AND(g22118, g26635)
--	g27076 = AND(g5024, g26393)
--	g27077 = AND(g22083, g26636)
--	g27079 = AND(g5044, g26401)
--	g27080 = AND(g23377, g26637)
--	g27081 = AND(g22108, g26638)
--	g27082 = AND(g22016, g26639)
--	g27083 = AND(g22093, g26640)
--	g27084 = AND(g23388, g26641)
--	g27085 = AND(g22134, g26642)
--	g27086 = AND(g23353, g26643)
--	g27087 = AND(g22021, g26644)
--	g27088 = AND(g23381, g26645)
--	g27089 = AND(g22118, g26646)
--	g27090 = AND(g23395, g26647)
--	g27091 = AND(g5142, g26429)
--	g27092 = AND(g5153, g26434)
--	g27093 = AND(g22108, g26648)
--	g27095 = AND(g5173, g26442)
--	g27096 = AND(g23388, g26649)
--	g27097 = AND(g22134, g26650)
--	g27098 = AND(g22021, g26651)
--	g27099 = AND(g22118, g26652)
--	g27100 = AND(g23395, g26653)
--	g27101 = AND(g22157, g26654)
--	g27103 = AND(g5235, g26461)
--	g27104 = AND(g5246, g26466)
--	g27105 = AND(g22134, g26656)
--	g27107 = AND(g5266, g26474)
--	g27108 = AND(g23395, g26657)
--	g27109 = AND(g22157, g26658)
--	g27110 = AND(g5298, g26485)
--	g27111 = AND(g5309, g26490)
--	g27112 = AND(g22157, g26662)
--	g27115 = AND(g5335, g26501)
--	g27178 = AND(g26110, g22213)
--	g27181 = AND(g16570, g26508, g13614)
--	g27182 = AND(g26151, g22217)
--	g27185 = AND(g26126, g22230)
--	g27187 = AND(g16594, g26516, g13626)
--	g27240 = AND(g26905, g22241)
--	g27241 = AND(g10730, g26934)
--	g27242 = AND(g26793, g8357)
--	g27244 = AND(g26914, g22258)
--	g27245 = AND(g26877, g22286)
--	g27246 = AND(g26988, g16676)
--	g27247 = AND(g27011, g16702)
--	g27248 = AND(g27037, g16733)
--	g27249 = AND(g27065, g16775)
--	g27355 = AND(g61, g26837)
--	g27356 = AND(g65, g26987)
--	g27358 = AND(g749, g26846)
--	g27359 = AND(g753, g27010)
--	g27364 = AND(g1435, g26855)
--	g27365 = AND(g1439, g27036)
--	g27370 = AND(g27126, g8874)
--	g27371 = AND(g2129, g26861)
--	g27372 = AND(g2133, g27064)
--	g27394 = AND(g17802, g27134)
--	g27396 = AND(g692, g27135)
--	g27407 = AND(g17914, g27136)
--	g27409 = AND(g1378, g27137)
--	g27425 = AND(g18025, g27138)
--	g27427 = AND(g2072, g27139)
--	g27446 = AND(g18142, g27141)
--	g27448 = AND(g2766, g27142)
--	g27495 = AND(g23945, g27146)
--	g27509 = AND(g23945, g27148)
--	g27516 = AND(g23974, g27151)
--	g27530 = AND(g23945, g27153)
--	g27534 = AND(g23974, g27155)
--	g27541 = AND(g24004, g27159)
--	g27552 = AND(g23974, g27162)
--	g27554 = AND(g24004, g27164)
--	g27561 = AND(g24038, g27167)
--	g27568 = AND(g24004, g27172)
--	g27570 = AND(g24038, g27173)
--	g27578 = AND(g24038, g27177)
--	g27656 = AND(g26796, g11004)
--	g27657 = AND(g27114, g11051)
--	g27659 = AND(g27132, g11114)
--	g27660 = AND(g26835, g11117)
--	g27661 = AND(g26841, g11173)
--	g27666 = AND(g26849, g11243)
--	g27671 = AND(g26885, g22212)
--	g27673 = AND(g26854, g11312)
--	g27679 = AND(g26782, g11386)
--	g27680 = AND(g26983, g11392)
--	g27681 = AND(g26788, g11456)
--	g27719 = AND(g27496, g20649)
--	g27720 = AND(g27481, g20652)
--	g27721 = AND(g27579, g20655)
--	g27723 = AND(g27464, g20679)
--	g27725 = AND(g27532, g20704)
--	g27726 = AND(g27531, g20732)
--	g27727 = AND(g27414, g19301)
--	g27728 = AND(g27564, g20766)
--	g27729 = AND(g27435, g19322)
--	g27730 = AND(g27454, g19349)
--	g27731 = AND(g27470, g19383)
--	g27732 = AND(g27492, g16758)
--	g27733 = AND(g27513, g16785)
--	g27734 = AND(g27538, g16814)
--	g27737 = AND(g27558, g16832)
--	g27770 = AND(g5642, g27449)
--	g27772 = AND(g5680, g27465)
--	g27773 = AND(g5732, g27484)
--	g27774 = AND(g5702, g27361)
--	g27775 = AND(g5790, g27506)
--	g27779 = AND(g5760, g27367)
--	g27783 = AND(g5819, g27373)
--	g27790 = AND(g5875, g27376)
--	g27904 = AND(g13873, g27387)
--	g27908 = AND(g13886, g27391)
--	g27909 = AND(g13895, g27397)
--	g27913 = AND(g4017, g27401)
--	g27914 = AND(g13927, g27404)
--	g27915 = AND(g13936, g27410)
--	g27922 = AND(g4112, g27416)
--	g27923 = AND(g4144, g27419)
--	g27924 = AND(g13983, g27422)
--	g27926 = AND(g13992, g27428)
--	g27931 = AND(g4221, g27432)
--	g27935 = AND(g4251, g27437)
--	g27936 = AND(g4283, g27440)
--	g27938 = AND(g14053, g27443)
--	g27945 = AND(g4376, g27451)
--	g27949 = AND(g4406, g27456)
--	g27951 = AND(g4438, g27459)
--	g27963 = AND(g4545, g27467)
--	g27968 = AND(g4575, g27472)
--	g27970 = AND(g14238, g27475)
--	g27984 = AND(g4721, g27486)
--	g27985 = AND(g14342, g27489)
--	g27991 = AND(g14360, g27498)
--	g28008 = AND(g27590, g9770)
--	g28009 = AND(g14454, g27510)
--	g28015 = AND(g14472, g27518)
--	g28027 = AND(g27590, g9895)
--	g28028 = AND(g27595, g9898)
--	g28035 = AND(g27599, g9916)
--	g28036 = AND(g14541, g27535)
--	g28042 = AND(g14559, g27543)
--	g28050 = AND(g27590, g10018)
--	g28051 = AND(g27595, g10021)
--	g28057 = AND(g27599, g10049)
--	g28058 = AND(g27604, g10052)
--	g28065 = AND(g27608, g10070)
--	g28066 = AND(g14596, g27555)
--	g28073 = AND(g27595, g10109)
--	g28079 = AND(g27599, g10127)
--	g28080 = AND(g27604, g10130)
--	g28086 = AND(g27608, g10158)
--	g28087 = AND(g27613, g10161)
--	g28094 = AND(g27617, g10179)
--	g28098 = AND(g27604, g10214)
--	g28104 = AND(g27608, g10232)
--	g28105 = AND(g27613, g10235)
--	g28111 = AND(g27617, g10263)
--	g28112 = AND(g27622, g10266)
--	g28116 = AND(g27613, g10316)
--	g28122 = AND(g27617, g10334)
--	g28123 = AND(g27622, g10337)
--	g28127 = AND(g27622, g10409)
--	g28171 = AND(g27349, g10898)
--	g28176 = AND(g27349, g10940)
--	g28188 = AND(g27349, g11008)
--	g28193 = AND(g27573, g21914)
--	g28319 = AND(g27855, g22246)
--	g28320 = AND(g27854, g20637)
--	g28322 = AND(g27937, g13868)
--	g28323 = AND(g8580, g27838)
--	g28324 = AND(g27810, g20659)
--	g28326 = AND(g27865, g22274)
--	g28327 = AND(g27900, g22275)
--	g28329 = AND(g27823, g20708)
--	g28330 = AND(g27864, g20711)
--	g28331 = AND(g27802, g22307)
--	g28332 = AND(g27883, g22331)
--	g28333 = AND(g27882, g20772)
--	g28334 = AND(g27842, g20793)
--	g28335 = AND(g27814, g22343)
--	g28336 = AND(g27896, g20810)
--	g28337 = AND(g28002, g19448)
--	g28338 = AND(g28029, g19475)
--	g28339 = AND(g28059, g19498)
--	g28340 = AND(g28088, g19519)
--	g28373 = AND(g56, g27969)
--	g28376 = AND(g744, g27990)
--	g28378 = AND(g52, g27776)
--	g28379 = AND(g27868, g19390, g19369)
--	g28380 = AND(g1430, g28014)
--	g28381 = AND(g28157, g9815)
--	g28383 = AND(g740, g27780)
--	g28385 = AND(g2124, g28041)
--	g28387 = AND(g1426, g27787)
--	g28389 = AND(g2120, g27794)
--	g28396 = AND(g7754, g27806)
--	g28398 = AND(g7769, g27817)
--	g28399 = AND(g7776, g27820)
--	g28401 = AND(g7782, g27831)
--	g28402 = AND(g7785, g27839)
--	g28404 = AND(g7792, g27843)
--	g28405 = AND(g7796, g27847)
--	g28407 = AND(g7799, g27858)
--	g28408 = AND(g7806, g27861)
--	g28411 = AND(g7809, g27872)
--	g28412 = AND(g7812, g27879)
--	g28416 = AND(g7823, g27889)
--	g28422 = AND(g17640, g28150)
--	g28423 = AND(g17724, g28152)
--	g28424 = AND(g17741, g28153)
--	g28426 = AND(g28128, g9170)
--	g28427 = AND(g26092, g28154)
--	g28428 = AND(g17825, g28155)
--	g28429 = AND(g17842, g28156)
--	g28430 = AND(g28128, g9196)
--	g28431 = AND(g26092, g28158)
--	g28433 = AND(g28133, g9212)
--	g28434 = AND(g26114, g28159)
--	g28435 = AND(g17937, g28160)
--	g28436 = AND(g17954, g28161)
--	g28438 = AND(g17882, g27919)
--	g28439 = AND(g28128, g9242)
--	g28440 = AND(g26092, g28162)
--	g28441 = AND(g28133, g9257)
--	g28442 = AND(g26114, g28163)
--	g28444 = AND(g28137, g9273)
--	g28445 = AND(g26121, g28164)
--	g28446 = AND(g18048, g28165)
--	g28448 = AND(g17974, g27928)
--	g28450 = AND(g17993, g27932)
--	g28451 = AND(g28133, g9320)
--	g28452 = AND(g26114, g28166)
--	g28453 = AND(g28137, g9335)
--	g28454 = AND(g26121, g28167)
--	g28456 = AND(g28141, g9351)
--	g28457 = AND(g26131, g28168)
--	g28459 = AND(g18074, g27939)
--	g28460 = AND(g18091, g27942)
--	g28462 = AND(g18110, g27946)
--	g28463 = AND(g28137, g9401)
--	g28464 = AND(g26121, g28169)
--	g28465 = AND(g28141, g9416)
--	g28466 = AND(g26131, g28170)
--	g28468 = AND(g18265, g28172)
--	g28469 = AND(g18179, g27952)
--	g28471 = AND(g18190, g27956)
--	g28472 = AND(g18207, g27959)
--	g28474 = AND(g18226, g27965)
--	g28475 = AND(g28141, g9498)
--	g28476 = AND(g26131, g28173)
--	g28477 = AND(g18341, g28174)
--	g28478 = AND(g18358, g28175)
--	g28479 = AND(g18286, g27973)
--	g28480 = AND(g18297, g27977)
--	g28481 = AND(g18314, g27981)
--	g28484 = AND(g18436, g28177)
--	g28485 = AND(g18453, g28178)
--	g28486 = AND(g18379, g27994)
--	g28487 = AND(g18390, g27999)
--	g28492 = AND(g18509, g28186)
--	g28493 = AND(g18526, g28187)
--	g28494 = AND(g18474, g28018)
--	g28497 = AND(g18573, g28190)
--	g28657 = AND(g27925, g13700)
--	g28659 = AND(g27917, g13736)
--	g28660 = AND(g27916, g11911)
--	g28662 = AND(g27911, g11951)
--	g28663 = AND(g27906, g11997)
--	g28664 = AND(g27997, g12055)
--	g28665 = AND(g27827, g22222)
--	g28666 = AND(g27980, g12106)
--	g28667 = AND(g27964, g13852)
--	g28669 = AND(g27897, g22233)
--	g28670 = AND(g27798, g21935)
--	g28671 = AND(g27962, g12161)
--	g28672 = AND(g27950, g13859)
--	g28707 = AND(g12436, g28379)
--	g28708 = AND(g28392, g22260)
--	g28709 = AND(g28400, g22261)
--	g28710 = AND(g28403, g22262)
--	g28711 = AND(g10749, g28415)
--	g28712 = AND(g28406, g22276)
--	g28713 = AND(g28410, g22290)
--	g28714 = AND(g28394, g22306)
--	g28715 = AND(g28414, g22332)
--	g28716 = AND(g28449, g19319)
--	g28717 = AND(g28461, g19346)
--	g28718 = AND(g28473, g19380)
--	g28719 = AND(g28482, g19412)
--	g28722 = AND(g28523, g16694)
--	g28724 = AND(g28551, g16725)
--	g28726 = AND(g28578, g16767)
--	g28729 = AND(g28606, g16794)
--	g28834 = AND(g5751, g28483)
--	g28836 = AND(g5810, g28491)
--	g28838 = AND(g5866, g28496)
--	g28840 = AND(g5913, g28500)
--	g28841 = AND(g27834, g28554)
--	g28843 = AND(g27834, g28581)
--	g28844 = AND(g27850, g28582)
--	g28846 = AND(g27834, g28608)
--	g28847 = AND(g27850, g28609)
--	g28848 = AND(g27875, g28610)
--	g28849 = AND(g27850, g28616)
--	g28850 = AND(g27875, g28617)
--	g28851 = AND(g27892, g28618)
--	g28852 = AND(g27875, g28623)
--	g28853 = AND(g27892, g28624)
--	g28854 = AND(g27892, g28629)
--	g28880 = AND(g13946, g28639)
--	g28881 = AND(g28612, g9199)
--	g28892 = AND(g14001, g28640)
--	g28893 = AND(g28612, g9245)
--	g28897 = AND(g14016, g28641)
--	g28898 = AND(g28619, g9260)
--	g28909 = AND(g14062, g28642)
--	g28910 = AND(g28612, g9303)
--	g28914 = AND(g14092, g28643)
--	g28915 = AND(g28619, g9323)
--	g28919 = AND(g14107, g28644)
--	g28923 = AND(g28625, g9338)
--	g28931 = AND(g14153, g28645)
--	g28935 = AND(g14177, g28646)
--	g28936 = AND(g28619, g9384)
--	g28940 = AND(g14207, g28647)
--	g28944 = AND(g28625, g9404)
--	g28948 = AND(g14222, g28648)
--	g28949 = AND(g28630, g9419)
--	g28958 = AND(g14268, g28649)
--	g28962 = AND(g14292, g28650)
--	g28966 = AND(g28625, g9481)
--	g28970 = AND(g14322, g28651)
--	g28971 = AND(g28630, g9501)
--	g28986 = AND(g14390, g28652)
--	g28996 = AND(g14414, g28653)
--	g28997 = AND(g28630, g9623)
--	g29022 = AND(g14502, g28655)
--	g29130 = AND(g28397, g22221)
--	g29174 = AND(g29031, g20684)
--	g29175 = AND(g29009, g20687)
--	g29176 = AND(g29097, g20690)
--	g29180 = AND(g28982, g20714)
--	g29183 = AND(g29064, g20739)
--	g29186 = AND(g29063, g20769)
--	g29188 = AND(g29083, g20796)
--	g29196 = AND(g15022, g28741)
--	g29200 = AND(g15096, g28751)
--	g29203 = AND(g15118, g28755)
--	g29208 = AND(g15188, g28764)
--	g29211 = AND(g15210, g28768)
--	g29217 = AND(g15274, g28775)
--	g29220 = AND(g15296, g28779)
--	g29225 = AND(g15366, g28785)
--	g29229 = AND(g9293, g28791)
--	g29232 = AND(g9356, g28796)
--	g29233 = AND(g9374, g28799)
--	g29234 = AND(g9427, g28804)
--	g29235 = AND(g9453, g28807)
--	g29236 = AND(g9471, g28810)
--	g29238 = AND(g9569, g28814)
--	g29239 = AND(g9595, g28817)
--	g29240 = AND(g9613, g28820)
--	g29241 = AND(g9711, g28823)
--	g29242 = AND(g9737, g28826)
--	g29243 = AND(g9857, g28829)
--	g29248 = AND(g28855, g8836)
--	g29251 = AND(g28855, g8856)
--	g29252 = AND(g28859, g8863)
--	g29255 = AND(g28855, g8885)
--	g29256 = AND(g28859, g8894)
--	g29257 = AND(g28863, g8901)
--	g29259 = AND(g28859, g8925)
--	g29260 = AND(g28863, g8934)
--	g29261 = AND(g28867, g8941)
--	g29262 = AND(g28863, g8965)
--	g29263 = AND(g28867, g8974)
--	g29264 = AND(g28867, g8997)
--	g29284 = AND(g29001, g28871)
--	g29289 = AND(g29030, g28883)
--	g29294 = AND(g29053, g28900)
--	g29300 = AND(g29072, g28925)
--	g29302 = AND(g29026, g28928)
--	g29310 = AND(g28978, g28951)
--	g29312 = AND(g29049, g28955)
--	g29320 = AND(g29088, g28972)
--	g29321 = AND(g29008, g28979)
--	g29323 = AND(g29068, g28983)
--	g29329 = AND(g29096, g29002)
--	g29330 = AND(g29038, g29010)
--	g29332 = AND(g29080, g29019)
--	g29336 = AND(g29045, g29023)
--	g29337 = AND(g29103, g29032)
--	g29338 = AND(g29060, g29042)
--	g29341 = AND(g29062, g29046)
--	g29342 = AND(g29107, g29054)
--	g29344 = AND(g29076, g29065)
--	g29346 = AND(g29087, g29077)
--	g29411 = AND(g29090, g21932)
--	g29464 = AND(g29190, g8375)
--	g29465 = AND(g29191, g8424)
--	g29466 = AND(g8587, g29265)
--	g29467 = AND(g29340, g19467)
--	g29468 = AND(g29343, g19490)
--	g29469 = AND(g29345, g19511)
--	g29470 = AND(g29347, g19530)
--	g29471 = AND(g21461, g29266)
--	g29472 = AND(g21461, g29268)
--	g29473 = AND(g21508, g29269)
--	g29474 = AND(g21508, g29271)
--	g29475 = AND(g21544, g29272)
--	g29476 = AND(g21544, g29274)
--	g29477 = AND(g21580, g29275)
--	g29478 = AND(g21580, g29277)
--	g29479 = AND(g21461, g29280)
--	g29480 = AND(g21461, g29282)
--	g29481 = AND(g21508, g29283)
--	g29482 = AND(g21461, g29285)
--	g29483 = AND(g21508, g29286)
--	g29484 = AND(g21544, g29287)
--	g29485 = AND(g21508, g29290)
--	g29486 = AND(g21544, g29291)
--	g29487 = AND(g21580, g29292)
--	g29488 = AND(g21544, g29295)
--	g29489 = AND(g21580, g29296)
--	g29490 = AND(g21580, g29301)
--	g29502 = AND(g29350, g8912)
--	g29518 = AND(g28728, g29360)
--	g29520 = AND(g28731, g29361)
--	g29521 = AND(g28733, g29362)
--	g29522 = AND(g27735, g29363)
--	g29523 = AND(g28737, g29364)
--	g29524 = AND(g28739, g29365)
--	g29525 = AND(g29195, g29366)
--	g29526 = AND(g27741, g29367)
--	g29527 = AND(g28748, g29368)
--	g29528 = AND(g28750, g29369)
--	g29529 = AND(g29199, g29370)
--	g29531 = AND(g29202, g29371)
--	g29532 = AND(g27746, g29372)
--	g29533 = AND(g28762, g29373)
--	g29534 = AND(g29206, g29374)
--	g29536 = AND(g29207, g29375)
--	g29538 = AND(g29210, g29376)
--	g29539 = AND(g27754, g29377)
--	g29540 = AND(g26041, g29378)
--	g29541 = AND(g29214, g29379)
--	g29543 = AND(g29215, g29380)
--	g29545 = AND(g29216, g29381)
--	g29547 = AND(g29219, g29382)
--	g29548 = AND(g28784, g29383)
--	g29549 = AND(g26043, g29384)
--	g29550 = AND(g29222, g29385)
--	g29553 = AND(g29223, g29386)
--	g29555 = AND(g29224, g29387)
--	g29557 = AND(g28789, g29388)
--	g29558 = AND(g28790, g29389)
--	g29559 = AND(g26045, g29390)
--	g29560 = AND(g29227, g29391)
--	g29562 = AND(g29228, g29392)
--	g29564 = AND(g28794, g29393)
--	g29565 = AND(g28795, g29394)
--	g29566 = AND(g26047, g29395)
--	g29567 = AND(g29231, g29396)
--	g29572 = AND(g28802, g29397)
--	g29573 = AND(g28803, g29398)
--	g29575 = AND(g28813, g29402)
--	g29607 = AND(g29193, g11056)
--	g29610 = AND(g29349, g11123)
--	g29614 = AND(g29359, g11182)
--	g29615 = AND(g29245, g11185)
--	g29619 = AND(g29247, g11259)
--	g29622 = AND(g29250, g11327)
--	g29624 = AND(g29254, g11407)
--	g29625 = AND(g29189, g11472)
--	g29626 = AND(g29318, g11478)
--	g29790 = AND(g29491, g10918)
--	g29792 = AND(g29491, g10977)
--	g29793 = AND(g29491, g11063)
--	g29810 = AND(g29748, g22248)
--	g29811 = AND(g29703, g20644)
--	g29812 = AND(g29762, g12223)
--	g29813 = AND(g29760, g13869)
--	g29814 = AND(g29728, g22266)
--	g29815 = AND(g29727, g20662)
--	g29816 = AND(g29759, g13883)
--	g29817 = AND(g29709, g20694)
--	g29818 = AND(g29732, g22293)
--	g29819 = AND(g29751, g22294)
--	g29820 = AND(g29717, g20743)
--	g29821 = AND(g29731, g20746)
--	g29822 = AND(g29705, g22335)
--	g29827 = AND(g29741, g22356)
--	g29828 = AND(g29740, g20802)
--	g29833 = AND(g29725, g20813)
--	g29834 = AND(g29713, g22366)
--	g29839 = AND(g29747, g20827)
--	g29909 = AND(g29735, g19420, g19401)
--	g29910 = AND(g29779, g9961)
--	g29942 = AND(g29771, g28877)
--	g29944 = AND(g29782, g28889)
--	g29945 = AND(g29773, g28894)
--	g29946 = AND(g29778, g28906)
--	g29947 = AND(g29785, g28911)
--	g29948 = AND(g29775, g28916)
--	g29949 = AND(g29781, g28932)
--	g29950 = AND(g29788, g28937)
--	g29951 = AND(g29777, g28945)
--	g29952 = AND(g29784, g28959)
--	g29953 = AND(g29791, g28967)
--	g29954 = AND(g29770, g28975)
--	g29955 = AND(g29787, g28993)
--	g29956 = AND(g29780, g28998)
--	g29957 = AND(g29772, g29005)
--	g29958 = AND(g29783, g29027)
--	g29959 = AND(g29774, g29035)
--	g29960 = AND(g29786, g29050)
--	g29961 = AND(g29776, g29057)
--	g29962 = AND(g29789, g29069)
--	g29963 = AND(g29758, g13737)
--	g29964 = AND(g29757, g13786)
--	g29965 = AND(g29756, g11961)
--	g29966 = AND(g29755, g12004)
--	g29967 = AND(g29754, g12066)
--	g29968 = AND(g29765, g12119)
--	g29969 = AND(g29721, g22237)
--	g29970 = AND(g29764, g12178)
--	g29971 = AND(g29763, g13861)
--	g29980 = AND(g29881, g8324)
--	g29981 = AND(g29869, g8330)
--	g29982 = AND(g29893, g8336)
--	g29983 = AND(g29885, g8344)
--	g29984 = AND(g29873, g8351)
--	g29985 = AND(g29897, g8363)
--	g29986 = AND(g29877, g8366)
--	g29987 = AND(g29889, g8369)
--	g29988 = AND(g29881, g8382)
--	g29989 = AND(g29893, g8391)
--	g29990 = AND(g29885, g8397)
--	g29991 = AND(g29901, g8403)
--	g29992 = AND(g12441, g29909)
--	g29993 = AND(g29897, g8411)
--	g29994 = AND(g29889, g8418)
--	g29995 = AND(g29893, g8434)
--	g29996 = AND(g29901, g8443)
--	g29997 = AND(g29918, g22277)
--	g29998 = AND(g29922, g22278)
--	g29999 = AND(g29924, g22279)
--	g30000 = AND(g10767, g29930)
--	g30001 = AND(g29897, g8449)
--	g30002 = AND(g29905, g8455)
--	g30003 = AND(g29901, g8469)
--	g30004 = AND(g29926, g22295)
--	g30005 = AND(g29905, g8478)
--	g30006 = AND(g29928, g22310)
--	g30007 = AND(g29905, g8494)
--	g30008 = AND(g29919, g22334)
--	g30009 = AND(g29929, g22357)
--	g30077 = AND(g29823, g10963)
--	g30079 = AND(g29823, g10988)
--	g30080 = AND(g29829, g10996)
--	g30081 = AND(g29823, g11022)
--	g30082 = AND(g29829, g11036)
--	g30083 = AND(g29835, g11048)
--	g30085 = AND(g29829, g11092)
--	g30086 = AND(g29835, g11108)
--	g30087 = AND(g29840, g11120)
--	g30088 = AND(g29844, g11138)
--	g30089 = AND(g29835, g11160)
--	g30090 = AND(g29840, g11176)
--	g30091 = AND(g29844, g11202)
--	g30092 = AND(g29849, g11205)
--	g30093 = AND(g29853, g11222)
--	g30094 = AND(g29840, g11246)
--	g30095 = AND(g29857, g11265)
--	g30096 = AND(g29844, g11268)
--	g30097 = AND(g29849, g11271)
--	g30098 = AND(g29853, g11284)
--	g30099 = AND(g29861, g11287)
--	g30100 = AND(g29865, g11306)
--	g30101 = AND(g29857, g11341)
--	g30102 = AND(g29849, g11348)
--	g30103 = AND(g29869, g11358)
--	g30104 = AND(g29853, g11361)
--	g30105 = AND(g29861, g11364)
--	g30106 = AND(g29865, g11379)
--	g30107 = AND(g29873, g11382)
--	g30108 = AND(g29877, g11401)
--	g30109 = AND(g29857, g11411)
--	g30110 = AND(g29881, g11417)
--	g30111 = AND(g29869, g11425)
--	g30112 = AND(g29861, g11432)
--	g30113 = AND(g29885, g11444)
--	g30114 = AND(g29865, g11447)
--	g30115 = AND(g29873, g11450)
--	g30116 = AND(g29921, g22236)
--	g30117 = AND(g29877, g11465)
--	g30118 = AND(g29889, g11468)
--	g30123 = AND(g30070, g20641)
--	g30127 = AND(g30065, g20719)
--	g30128 = AND(g30062, g20722)
--	g30129 = AND(g30071, g20725)
--	g30131 = AND(g30059, g20749)
--	g30132 = AND(g30068, g20776)
--	g30133 = AND(g30067, g20799)
--	g30138 = AND(g30069, g20816)
--	g30216 = AND(g30036, g8921)
--	g30217 = AND(g30036, g8955)
--	g30218 = AND(g30040, g8961)
--	g30219 = AND(g30036, g8980)
--	g30220 = AND(g30040, g8987)
--	g30221 = AND(g30044, g8993)
--	g30222 = AND(g30040, g9010)
--	g30223 = AND(g30044, g9016)
--	g30224 = AND(g30048, g9022)
--	g30225 = AND(g30044, g9035)
--	g30226 = AND(g30048, g9041)
--	g30227 = AND(g30048, g9058)
--	g30327 = AND(g30187, g8321)
--	g30330 = AND(g30195, g8333)
--	g30333 = AND(g30191, g8341)
--	g30334 = AND(g30203, g8347)
--	g30337 = AND(g30199, g8354)
--	g30340 = AND(g30207, g8372)
--	g30345 = AND(g30195, g8388)
--	g30348 = AND(g30203, g8400)
--	g30351 = AND(g30199, g8408)
--	g30352 = AND(g30211, g8414)
--	g30355 = AND(g30207, g8421)
--	g30361 = AND(g30203, g8440)
--	g30364 = AND(g30211, g8452)
--	g30367 = AND(g30207, g8460)
--	g30372 = AND(g8594, g30228)
--	g30374 = AND(g30211, g8475)
--	g30387 = AND(g30229, g8888)
--	g30388 = AND(g30229, g8918)
--	g30389 = AND(g30233, g8928)
--	g30390 = AND(g30229, g8952)
--	g30391 = AND(g30233, g8958)
--	g30392 = AND(g30237, g8968)
--	g30393 = AND(g30233, g8984)
--	g30394 = AND(g30237, g8990)
--	g30395 = AND(g30241, g9000)
--	g30396 = AND(g30237, g9013)
--	g30397 = AND(g30241, g9019)
--	g30398 = AND(g30241, g9038)
--	g30407 = AND(g30134, g10991)
--	g30409 = AND(g30134, g11025)
--	g30410 = AND(g30139, g11028)
--	g30411 = AND(g30143, g11039)
--	g30436 = AND(g30134, g11079)
--	g30437 = AND(g30139, g11082)
--	g30438 = AND(g30147, g11085)
--	g30440 = AND(g30143, g11095)
--	g30441 = AND(g30151, g11098)
--	g30442 = AND(g30155, g11111)
--	g30444 = AND(g30139, g11132)
--	g30445 = AND(g30147, g11135)
--	g30447 = AND(g30143, g11145)
--	g30448 = AND(g30151, g11148)
--	g30449 = AND(g30159, g11151)
--	g30451 = AND(g30155, g11163)
--	g30452 = AND(g30163, g11166)
--	g30453 = AND(g30167, g11179)
--	g30454 = AND(g30147, g11199)
--	g30457 = AND(g30151, g11216)
--	g30458 = AND(g30159, g11219)
--	g30460 = AND(g30155, g11231)
--	g30461 = AND(g30163, g11234)
--	g30462 = AND(g30171, g11237)
--	g30464 = AND(g30167, g11249)
--	g30465 = AND(g30175, g11252)
--	g30467 = AND(g30179, g11274)
--	g30469 = AND(g30159, g11281)
--	g30472 = AND(g30163, g11300)
--	g30473 = AND(g30171, g11303)
--	g30475 = AND(g30167, g11315)
--	g30476 = AND(g30175, g11318)
--	g30477 = AND(g30183, g11321)
--	g30478 = AND(g30187, g11344)
--	g30481 = AND(g30179, g11351)
--	g30484 = AND(g30191, g11367)
--	g30486 = AND(g30171, g11376)
--	g30489 = AND(g30175, g11395)
--	g30490 = AND(g30183, g11398)
--	g30492 = AND(g30187, g11414)
--	g30495 = AND(g30179, g11422)
--	g30496 = AND(g30195, g11428)
--	g30499 = AND(g30191, g11435)
--	g30502 = AND(g30199, g11453)
--	g30504 = AND(g30183, g11462)
--	g30696 = AND(g30383, g10943)
--	g30697 = AND(g30383, g11011)
--	g30698 = AND(g30383, g11126)
--	g30728 = AND(g30605, g22252)
--	g30735 = AND(g30629, g22268)
--	g30736 = AND(g30584, g20669)
--	g30743 = AND(g30610, g22283)
--	g30744 = AND(g30609, g20697)
--	g30750 = AND(g30593, g20729)
--	g30754 = AND(g30614, g22313)
--	g30755 = AND(g30632, g22314)
--	g30757 = AND(g30601, g20780)
--	g30758 = AND(g30613, g20783)
--	g30759 = AND(g30588, g22360)
--	g30760 = AND(g30622, g22379)
--	g30761 = AND(g30621, g20822)
--	g30762 = AND(g30608, g20830)
--	g30763 = AND(g30597, g22386)
--	g30764 = AND(g30628, g20837)
--	g30766 = AND(g30617, g19457, g19431)
--	g30916 = AND(g30785, g22251)
--	g30917 = AND(g12446, g30766)
--	g30918 = AND(g30780, g22296)
--	g30919 = AND(g30786, g22297)
--	g30920 = AND(g30787, g22298)
--	g30921 = AND(g10773, g30791)
--	g30922 = AND(g30788, g22315)
--	g30923 = AND(g30789, g22338)
--	g30924 = AND(g30783, g22359)
--	g30925 = AND(g30790, g22380)
--	g30944 = AND(g30935, g20666)
--	g30945 = AND(g30931, g20754)
--	g30946 = AND(g30930, g20757)
--	g30947 = AND(g30936, g20760)
--	g30948 = AND(g30929, g20786)
--	g30949 = AND(g30933, g20806)
--	g30950 = AND(g30932, g20819)
--	g30951 = AND(g30934, g20833)
--	g30953 = AND(g8605, g30952)
--	
--	g9144 = OR(g2986, g5389)
--	g10778 = OR(g2929, g8022)
--	g12377 = OR(g7553, g11059)
--	g12407 = OR(g7573, g10779)
--	g12886 = OR(g9534, g3398)
--	g12926 = OR(g9676, g3554)
--	g12955 = OR(g9822, g3710)
--	g12984 = OR(g9968, g3866)
--	g16539 = OR(g15880, g14657)
--	g16571 = OR(g15913, g14691)
--	g16595 = OR(g15942, g14725)
--	g16615 = OR(g15971, g14753)
--	g17973 = OR(g11623, g15659)
--	g19181 = OR(g17729, g17979)
--	g19186 = OR(g18419, g17887)
--	g19187 = OR(g18419, g17729)
--	g19188 = OR(g17830, g18096)
--	g19191 = OR(g17807, g17887)
--	g19192 = OR(g18183, g18270)
--	g19193 = OR(g18492, g17998)
--	g19194 = OR(g18492, g17830)
--	g19195 = OR(g17942, g18212)
--	g19200 = OR(g18346, g18424)
--	g19201 = OR(g18183, g18424)
--	g19202 = OR(g17919, g17998)
--	g19203 = OR(g18290, g18363)
--	g19204 = OR(g18556, g18115)
--	g19205 = OR(g18556, g17942)
--	g19206 = OR(g18053, g18319)
--	g19209 = OR(g18079, g18346)
--	g19210 = OR(g18079, g18183)
--	g19211 = OR(g18441, g18497)
--	g19212 = OR(g18290, g18497)
--	g19213 = OR(g18030, g18115)
--	g19214 = OR(g18383, g18458)
--	g19215 = OR(g18606, g18231)
--	g19216 = OR(g18606, g18053)
--	g19221 = OR(g18270, g18346)
--	g19222 = OR(g18195, g18441)
--	g19223 = OR(g18195, g18290)
--	g19224 = OR(g18514, g18561)
--	g19225 = OR(g18383, g18561)
--	g19226 = OR(g18147, g18231)
--	g19227 = OR(g18478, g18531)
--	I25477 = OR(g17024, g17000, g16992)
--	g19230 = OR(g16985, g16965, I25477)
--	g19231 = OR(g18363, g18441)
--	g19232 = OR(g18302, g18514)
--	g19233 = OR(g18302, g18383)
--	g19234 = OR(g18578, g18611)
--	g19235 = OR(g18478, g18611)
--	I25495 = OR(g17158, g17137, g17115)
--	g19240 = OR(g17083, g17050, I25495)
--	g19242 = OR(g14244, g16501)
--	I25500 = OR(g17058, g17030, g17016)
--	g19243 = OR(g16995, g16986, I25500)
--	g19244 = OR(g18458, g18514)
--	g19245 = OR(g18395, g18578)
--	g19246 = OR(g18395, g18478)
--	g19250 = OR(g17729, g17807)
--	I25516 = OR(g17173, g17160, g17142)
--	g19253 = OR(g17121, g17085, I25516)
--	g19255 = OR(g14366, g16523)
--	I25521 = OR(g17093, g17064, g17046)
--	g19256 = OR(g17019, g16996, I25521)
--	g19257 = OR(g18531, g18578)
--	g19263 = OR(g17887, g17979)
--	g19264 = OR(g17830, g17919)
--	I25549 = OR(g17190, g17175, g17165)
--	g19266 = OR(g17148, g17123, I25549)
--	g19268 = OR(g14478, g16554)
--	I25554 = OR(g17131, g17099, g17080)
--	g19269 = OR(g17049, g17020, I25554)
--	g19275 = OR(g16867, g16515, g19001)
--	g19278 = OR(g17998, g18096)
--	g19279 = OR(g17942, g18030)
--	I25588 = OR(g17201, g17192, g17180)
--	g19281 = OR(g17171, g17150, I25588)
--	g19283 = OR(g14565, g16586)
--	g19294 = OR(g16895, g16546, g16507)
--	g19297 = OR(g18115, g18212)
--	g19298 = OR(g18053, g18147)
--	g19312 = OR(g16924, g16578, g16529)
--	g19315 = OR(g18231, g18319)
--	g19333 = OR(g16954, g16602, g16560)
--	g19450 = OR(g14837, g16682)
--	g19477 = OR(g14910, g16708)
--	g19500 = OR(g14991, g16739)
--	g19503 = OR(g16884, g16697, g16665)
--	g19521 = OR(g15080, g16781)
--	g19522 = OR(g16913, g16728, g16686)
--	g19532 = OR(g16943, g16770, g16712)
--	g19542 = OR(g16974, g16797, g16743)
--	I26429 = OR(g17979, g17887, g17807)
--	g19981 = OR(g17729, g18419, I26429)
--	I26455 = OR(g18424, g18346, g18270)
--	g20015 = OR(g18183, g18079, I26455)
--	I26461 = OR(g18096, g17998, g17919)
--	g20019 = OR(g17830, g18492, I26461)
--	I26491 = OR(g18497, g18441, g18363)
--	g20057 = OR(g18290, g18195, I26491)
--	I26497 = OR(g18212, g18115, g18030)
--	g20061 = OR(g17942, g18556, I26497)
--	I26532 = OR(g18561, g18514, g18458)
--	g20098 = OR(g18383, g18302, I26532)
--	I26538 = OR(g18319, g18231, g18147)
--	g20102 = OR(g18053, g18606, I26538)
--	I26571 = OR(g18611, g18578, g18531)
--	g20123 = OR(g18478, g18395, I26571)
--	g21120 = OR(g19484, g16515, g14071)
--	g21139 = OR(g19505, g16546, g14186)
--	g21159 = OR(g19524, g16578, g14301)
--	g21179 = OR(g19534, g16602, g14423)
--	g21244 = OR(g19578, g16697, g14776)
--	g21253 = OR(g19608, g16728, g14811)
--	g21261 = OR(g19641, g16770, g14863)
--	g21269 = OR(g19681, g16797, g14936)
--	g21501 = OR(g20522, g16867, g14071)
--	g21536 = OR(g20522, g19484, g19001)
--	g21540 = OR(g20542, g16895, g14186)
--	g21572 = OR(g20542, g19505, g16507)
--	g21576 = OR(g19067, g16924, g14301)
--	g21605 = OR(g19067, g19524, g16529)
--	g21609 = OR(g19084, g16954, g14423)
--	g21634 = OR(g19084, g19534, g16560)
--	g21774 = OR(g19121, g16884, g14776)
--	g21787 = OR(g19121, g19578, g16665)
--	I28305 = OR(g20197, g20177, g20145)
--	g21788 = OR(g20117, g20094, I28305)
--	g21789 = OR(g19128, g16913, g14811)
--	I28318 = OR(g19092, g19088, g19079)
--	g21799 = OR(g16505, g20538, g18994, I28318)
--	g21800 = OR(g18665, g20270, g20248, g18647)
--	g21801 = OR(g19128, g19608, g16686)
--	I28323 = OR(g20227, g20211, g20183)
--	g21802 = OR(g20147, g20119, I28323)
--	g21803 = OR(g19135, g16943, g14863)
--	g21806 = OR(g20116, g20093, g18547, g19097)
--	I28330 = OR(g19099, g19094, g19089)
--	g21807 = OR(g16527, g19063, g19007, I28330)
--	g21808 = OR(g18688, g20282, g20271, g18650)
--	g21809 = OR(g19135, g19641, g16712)
--	I28335 = OR(g20254, g20241, g20217)
--	g21810 = OR(g20185, g20149, I28335)
--	g21811 = OR(g19138, g16974, g14936)
--	g21813 = OR(g20146, g20118, g18597, g19104)
--	I28341 = OR(g19106, g19101, g19095)
--	g21814 = OR(g16558, g19080, g16513, I28341)
--	g21815 = OR(g18717, g20293, g20283, g18654)
--	g21816 = OR(g19138, g19681, g16743)
--	I28346 = OR(g20277, g20268, g20247)
--	g21817 = OR(g20219, g20187, I28346)
--	g21819 = OR(g20184, g20148, g18629, g19109)
--	I28351 = OR(g19111, g19108, g19102)
--	g21820 = OR(g16590, g19090, g16535, I28351)
--	g21821 = OR(g18753, g20309, g20294, g18668)
--	g21823 = OR(g20218, g20186, g18638, g19116)
--	I28365 = OR(g20280, g18652, g18649)
--	g21844 = OR(g20222, g18645, I28365)
--	I28369 = OR(g20291, g18666, g18653)
--	g21846 = OR(g20249, g18648, I28369)
--	I28374 = OR(g20307, g18689, g18667)
--	g21849 = OR(g20272, g18651, I28374)
--	I28380 = OR(g20326, g18718, g18690)
--	g21856 = OR(g20284, g18655, I28380)
--	g22175 = OR(g16075, g20842)
--	g22190 = OR(g16113, g20850)
--	g22199 = OR(g16164, g20858)
--	g22205 = OR(g16223, g20866)
--	g22811 = OR(g562, g559, g12451, g21851)
--	g23052 = OR(g21800, g21788, g21844)
--	g23071 = OR(g21808, g21802, g21846)
--	g23084 = OR(g21815, g21810, g21849)
--	g23089 = OR(g21806, g21799)
--	g23100 = OR(g21821, g21817, g21856)
--	g23107 = OR(g21813, g21807)
--	g23120 = OR(g21819, g21814)
--	g23129 = OR(g21823, g21820)
--	g23319 = OR(g14493, g22385)
--	g23688 = OR(g23106, g21906)
--	g23742 = OR(g23119, g21920)
--	g23797 = OR(g23128, g21938)
--	g23850 = OR(g23139, g20647)
--	g23919 = OR(g22666, g23140)
--	g24239 = OR(g19387, g22401)
--	g24244 = OR(g14144, g22317)
--	g24245 = OR(g19417, g22402)
--	g24252 = OR(g14259, g22342)
--	g24254 = OR(g19454, g22403)
--	g24257 = OR(g14381, g22365)
--	g24258 = OR(g19481, g22404)
--	g24633 = OR(g24094, g20842)
--	g24653 = OR(g24095, g20850)
--	g24672 = OR(g24097, g20858)
--	g24691 = OR(g24103, g20866)
--	g24890 = OR(g23639, g23144)
--	g24909 = OR(g23726, g23142)
--	g24925 = OR(g23772, g23141)
--	g24965 = OR(g23922, g23945)
--	g24978 = OR(g23954, g23974)
--	g24989 = OR(g23983, g24004)
--	g25000 = OR(g24013, g24038)
--	g25183 = OR(g24958, g24893)
--	g25186 = OR(g24969, g24916)
--	g25190 = OR(g24982, g24933)
--	g25195 = OR(g24993, g24945)
--	g25489 = OR(g24795, g16466)
--	g25490 = OR(g24759, g23146)
--	g25520 = OR(g24813, g23145)
--	g25566 = OR(g24843, g23143)
--	g26320 = OR(g25852, g25870)
--	g26367 = OR(g25873, g25882)
--	g26410 = OR(g25885, g25887)
--	g26451 = OR(g25890, g25892)
--	g26974 = OR(g26157, g23147)
--	g27113 = OR(g1248, g1245, g26534)
--	g28501 = OR(g27738, g25764)
--	g28512 = OR(g26481, g27738)
--	g28529 = OR(g27743, g25818)
--	g28540 = OR(g26497, g27743)
--	g28556 = OR(g27751, g25853)
--	g28567 = OR(g26512, g27751)
--	g28584 = OR(g27756, g25874)
--	g28595 = OR(g26520, g27756)
--	g29348 = OR(g1942, g1939, g29113)
--	g30305 = OR(g2636, g2633, g30072)
--	
--	I15167 = NAND(g2981, g2874)
--	I15168 = NAND(g2981, I15167)
--	I15169 = NAND(g2874, I15167)
--	g7855 = NAND(I15168, I15169)
--	I15183 = NAND(g2975, g2978)
--	I15184 = NAND(g2975, I15183)
--	I15185 = NAND(g2978, I15183)
--	g7875 = NAND(I15184, I15185)
--	I15190 = NAND(g2956, g2959)
--	I15191 = NAND(g2956, I15190)
--	I15192 = NAND(g2959, I15190)
--	g7876 = NAND(I15191, I15192)
--	I15204 = NAND(g2969, g2972)
--	I15205 = NAND(g2969, I15204)
--	I15206 = NAND(g2972, I15204)
--	g7895 = NAND(I15205, I15206)
--	I15211 = NAND(g2947, g2953)
--	I15212 = NAND(g2947, I15211)
--	I15213 = NAND(g2953, I15211)
--	g7896 = NAND(I15212, I15213)
--	I15237 = NAND(g2963, g2966)
--	I15238 = NAND(g2963, I15237)
--	I15239 = NAND(g2966, I15237)
--	g7922 = NAND(I15238, I15239)
--	I15244 = NAND(g2941, g2944)
--	I15245 = NAND(g2941, I15244)
--	I15246 = NAND(g2944, I15244)
--	g7923 = NAND(I15245, I15246)
--	I15276 = NAND(g2935, g2938)
--	I15277 = NAND(g2935, I15276)
--	I15278 = NAND(g2938, I15276)
--	g7970 = NAND(I15277, I15278)
--	g8381 = NAND(g8182, g8120, g8044, g7989)
--	g8533 = NAND(g3398, g3366)
--	g8547 = NAND(g3398, g3366)
--	g8550 = NAND(g3554, g3522)
--	g8560 = NAND(g3554, g3522)
--	g8563 = NAND(g3710, g3678)
--	g8571 = NAND(g3710, g3678)
--	g8574 = NAND(g3866, g3834)
--	g8577 = NAND(g3866, g3834)
--	I16879 = NAND(g4203, g3998)
--	I16880 = NAND(g4203, I16879)
--	I16881 = NAND(g3998, I16879)
--	g9883 = NAND(I16880, I16881)
--	I16965 = NAND(g4734, g4452)
--	I16966 = NAND(g4734, I16965)
--	I16967 = NAND(g4452, I16965)
--	g10003 = NAND(I16966, I16967)
--	g10038 = NAND(g7772, g3366)
--	I17059 = NAND(g6637, g6309)
--	I17060 = NAND(g6637, I17059)
--	I17061 = NAND(g6309, I17059)
--	g10095 = NAND(I17060, I17061)
--	g10147 = NAND(g7788, g3522)
--	I17149 = NAND(g7465, g7142)
--	I17150 = NAND(g7465, I17149)
--	I17151 = NAND(g7142, I17149)
--	g10185 = NAND(I17150, I17151)
--	g10252 = NAND(g7802, g3678)
--	g10354 = NAND(g7815, g3834)
--	g10649 = NAND(g3398, g6912)
--	g10676 = NAND(g3398, g6678)
--	g10677 = NAND(g3398, g6912)
--	g10679 = NAND(g3554, g7162)
--	g10703 = NAND(g3398, g6678)
--	g10705 = NAND(g3554, g6980)
--	g10706 = NAND(g3554, g7162)
--	g10708 = NAND(g3710, g7358)
--	g10723 = NAND(g3554, g6980)
--	g10725 = NAND(g3710, g7230)
--	g10726 = NAND(g3710, g7358)
--	g10728 = NAND(g3866, g7488)
--	g10744 = NAND(g3710, g7230)
--	g10746 = NAND(g3866, g7426)
--	g10747 = NAND(g3866, g7488)
--	g10763 = NAND(g3866, g7426)
--	I18106 = NAND(g7875, g7855)
--	I18107 = NAND(g7875, I18106)
--	I18108 = NAND(g7855, I18106)
--	g11188 = NAND(I18107, I18108)
--	I18113 = NAND(g3997, g8181)
--	I18114 = NAND(g3997, I18113)
--	I18115 = NAND(g8181, I18113)
--	g11189 = NAND(I18114, I18115)
--	I18190 = NAND(g7922, g7895)
--	I18191 = NAND(g7922, I18190)
--	I18192 = NAND(g7895, I18190)
--	g11262 = NAND(I18191, I18192)
--	I18197 = NAND(g7896, g7876)
--	I18198 = NAND(g7896, I18197)
--	I18199 = NAND(g7876, I18197)
--	g11263 = NAND(I18198, I18199)
--	I18204 = NAND(g7975, g4202)
--	I18205 = NAND(g7975, I18204)
--	I18206 = NAND(g4202, I18204)
--	g11264 = NAND(I18205, I18206)
--	I18280 = NAND(g7970, g7923)
--	I18281 = NAND(g7970, I18280)
--	I18282 = NAND(g7923, I18280)
--	g11330 = NAND(I18281, I18282)
--	I18287 = NAND(g8256, g8102)
--	I18288 = NAND(g8256, I18287)
--	I18289 = NAND(g8102, I18287)
--	g11331 = NAND(I18288, I18289)
--	I18368 = NAND(g4325, g4093)
--	I18369 = NAND(g4325, I18368)
--	I18370 = NAND(g4093, I18368)
--	g11410 = NAND(I18369, I18370)
--	g11617 = NAND(g8313, g2883)
--	I18799 = NAND(g11410, g11331)
--	I18800 = NAND(g11410, I18799)
--	I18801 = NAND(g11331, I18799)
--	g11621 = NAND(I18800, I18801)
--	g11661 = NAND(g9534, g3366)
--	g11662 = NAND(g9534, g3366)
--	g11672 = NAND(g9534, g3366)
--	g11673 = NAND(g9676, g3522)
--	g11674 = NAND(g9676, g3522)
--	g11683 = NAND(g9534, g3366)
--	g11684 = NAND(g9676, g3522)
--	g11685 = NAND(g9822, g3678)
--	g11686 = NAND(g9822, g3678)
--	g11691 = NAND(g9534, g3366)
--	g11692 = NAND(g9676, g3522)
--	g11693 = NAND(g9822, g3678)
--	g11694 = NAND(g9968, g3834)
--	g11695 = NAND(g9968, g3834)
--	g11696 = NAND(g9534, g3366)
--	g11698 = NAND(g9676, g3522)
--	g11699 = NAND(g9822, g3678)
--	g11700 = NAND(g9968, g3834)
--	g11701 = NAND(g9534, g3366)
--	g11702 = NAND(g9676, g3522)
--	g11704 = NAND(g9822, g3678)
--	g11705 = NAND(g9968, g3834)
--	g11707 = NAND(g9534, g3366)
--	g11708 = NAND(g9534, g3366)
--	g11709 = NAND(g9676, g3522)
--	g11710 = NAND(g9822, g3678)
--	g11712 = NAND(g9968, g3834)
--	g11713 = NAND(g10481, g9144)
--	g11716 = NAND(g9534, g3366)
--	g11717 = NAND(g9676, g3522)
--	g11718 = NAND(g9676, g3522)
--	g11719 = NAND(g9822, g3678)
--	g11720 = NAND(g9968, g3834)
--	g11721 = NAND(g9534, g3366)
--	g11722 = NAND(g9676, g3522)
--	g11723 = NAND(g9822, g3678)
--	g11724 = NAND(g9822, g3678)
--	g11725 = NAND(g9968, g3834)
--	g11726 = NAND(g9676, g3522)
--	g11727 = NAND(g9822, g3678)
--	g11728 = NAND(g9968, g3834)
--	g11729 = NAND(g9968, g3834)
--	g11730 = NAND(g9822, g3678)
--	g11731 = NAND(g9968, g3834)
--	g11733 = NAND(g9968, g3834)
--	g12433 = NAND(g2879, g10778)
--	g12486 = NAND(g8278, g6448)
--	g12503 = NAND(g8278, g5438)
--	g12506 = NAND(g8287, g6713)
--	g12520 = NAND(g8287, g5473)
--	g12523 = NAND(g8296, g7015)
--	g12535 = NAND(g8296, g5512)
--	g12538 = NAND(g8305, g7265)
--	g12544 = NAND(g8305, g5556)
--	I20031 = NAND(g10003, g9883)
--	I20032 = NAND(g10003, I20031)
--	I20033 = NAND(g9883, I20031)
--	g12988 = NAND(I20032, I20033)
--	I20048 = NAND(g10185, g10095)
--	I20049 = NAND(g10185, I20048)
--	I20050 = NAND(g10095, I20048)
--	g12999 = NAND(I20049, I20050)
--	g13020 = NAND(g9534, g6912)
--	g13021 = NAND(g9534, g6912)
--	g13026 = NAND(g9534, g6678)
--	g13027 = NAND(g9534, g6912)
--	g13028 = NAND(g9534, g6678)
--	g13029 = NAND(g9676, g7162)
--	g13030 = NAND(g9676, g7162)
--	g13034 = NAND(g9534, g6678)
--	g13035 = NAND(g9534, g6912)
--	g13037 = NAND(g9676, g6980)
--	g13038 = NAND(g9676, g7162)
--	g13039 = NAND(g9676, g6980)
--	g13040 = NAND(g9822, g7358)
--	g13041 = NAND(g9822, g7358)
--	g13044 = NAND(g9534, g6678)
--	g13045 = NAND(g9534, g6912)
--	g13047 = NAND(g9676, g6980)
--	g13048 = NAND(g9676, g7162)
--	g13050 = NAND(g9822, g7230)
--	g13051 = NAND(g9822, g7358)
--	g13052 = NAND(g9822, g7230)
--	g13053 = NAND(g9968, g7488)
--	g13054 = NAND(g9968, g7488)
--	g13058 = NAND(g9534, g6678)
--	g13059 = NAND(g9534, g6912)
--	g13061 = NAND(g9676, g6980)
--	g13062 = NAND(g9676, g7162)
--	g13064 = NAND(g9822, g7230)
--	g13065 = NAND(g9822, g7358)
--	g13067 = NAND(g9968, g7426)
--	g13068 = NAND(g9968, g7488)
--	g13069 = NAND(g9968, g7426)
--	g13071 = NAND(g9534, g6678)
--	g13072 = NAND(g9534, g6912)
--	g13074 = NAND(g9676, g6980)
--	g13075 = NAND(g9676, g7162)
--	g13077 = NAND(g9822, g7230)
--	g13078 = NAND(g9822, g7358)
--	g13080 = NAND(g9968, g7426)
--	g13081 = NAND(g9968, g7488)
--	g13087 = NAND(g9534, g6678)
--	g13088 = NAND(g9534, g6912)
--	g13089 = NAND(g9534, g6912)
--	g13090 = NAND(g9676, g6980)
--	g13091 = NAND(g9676, g7162)
--	g13093 = NAND(g9822, g7230)
--	g13094 = NAND(g9822, g7358)
--	g13096 = NAND(g9968, g7426)
--	g13097 = NAND(g9968, g7488)
--	g13098 = NAND(g9534, g6678)
--	g13099 = NAND(g9534, g6912)
--	g13100 = NAND(g9534, g6678)
--	g13102 = NAND(g9676, g6980)
--	g13103 = NAND(g9676, g7162)
--	g13104 = NAND(g9676, g7162)
--	g13105 = NAND(g9822, g7230)
--	g13106 = NAND(g9822, g7358)
--	g13108 = NAND(g9968, g7426)
--	g13109 = NAND(g9968, g7488)
--	g13112 = NAND(g9534, g6678)
--	g13113 = NAND(g9534, g6912)
--	g13114 = NAND(g9676, g6980)
--	g13115 = NAND(g9676, g7162)
--	g13116 = NAND(g9676, g6980)
--	g13118 = NAND(g9822, g7230)
--	g13119 = NAND(g9822, g7358)
--	g13120 = NAND(g9822, g7358)
--	g13121 = NAND(g9968, g7426)
--	g13122 = NAND(g9968, g7488)
--	g13123 = NAND(g9534, g6678)
--	g13125 = NAND(g9676, g6980)
--	g13126 = NAND(g9676, g7162)
--	g13127 = NAND(g9822, g7230)
--	g13128 = NAND(g9822, g7358)
--	g13129 = NAND(g9822, g7230)
--	g13131 = NAND(g9968, g7426)
--	g13132 = NAND(g9968, g7488)
--	g13133 = NAND(g9968, g7488)
--	g13134 = NAND(g9676, g6980)
--	g13136 = NAND(g9822, g7230)
--	g13137 = NAND(g9822, g7358)
--	g13138 = NAND(g9968, g7426)
--	g13139 = NAND(g9968, g7488)
--	g13140 = NAND(g9968, g7426)
--	g13142 = NAND(g9822, g7230)
--	g13144 = NAND(g9968, g7426)
--	g13145 = NAND(g9968, g7488)
--	g13146 = NAND(g9968, g7426)
--	g13147 = NAND(g8278, g3306)
--	g13150 = NAND(g8287, g3462)
--	g13156 = NAND(g8296, g3618)
--	g13165 = NAND(g8305, g3774)
--	g13245 = NAND(g10779, g7901)
--	g13305 = NAND(g8317, g2993)
--	I20429 = NAND(g11262, g11188)
--	I20430 = NAND(g11262, I20429)
--	I20431 = NAND(g11188, I20429)
--	g13348 = NAND(I20430, I20431)
--	I20465 = NAND(g11330, g11263)
--	I20466 = NAND(g11330, I20465)
--	I20467 = NAND(g11263, I20465)
--	g13370 = NAND(I20466, I20467)
--	I20504 = NAND(g11264, g11189)
--	I20505 = NAND(g11264, I20504)
--	I20506 = NAND(g11189, I20504)
--	g13399 = NAND(I20505, I20506)
--	g13476 = NAND(g12565, g3254)
--	g13478 = NAND(g12611, g3410)
--	g13482 = NAND(g12657, g3566)
--	g13494 = NAND(g12565, g3254)
--	g13495 = NAND(g12611, g3410)
--	g13497 = NAND(g12657, g3566)
--	g13501 = NAND(g12711, g3722)
--	I20743 = NAND(g11621, g13399)
--	I20744 = NAND(g11621, I20743)
--	I20745 = NAND(g13399, I20743)
--	g13507 = NAND(I20744, I20745)
--	g13510 = NAND(g12565, g3254)
--	g13511 = NAND(g12611, g3410)
--	g13512 = NAND(g12657, g3566)
--	g13514 = NAND(g12711, g3722)
--	g13518 = NAND(g12565, g3254)
--	g13524 = NAND(g12611, g3410)
--	g13525 = NAND(g12657, g3566)
--	g13526 = NAND(g12711, g3722)
--	g13528 = NAND(g12565, g3254)
--	g13529 = NAND(g12611, g3410)
--	g13535 = NAND(g12657, g3566)
--	g13536 = NAND(g12711, g3722)
--	g13537 = NAND(g12565, g3254)
--	g13538 = NAND(g12565, g3254)
--	g13539 = NAND(g12611, g3410)
--	g13540 = NAND(g12657, g3566)
--	g13546 = NAND(g12711, g3722)
--	g13547 = NAND(g12565, g3254)
--	g13548 = NAND(g12611, g3410)
--	g13549 = NAND(g12611, g3410)
--	g13550 = NAND(g12657, g3566)
--	g13551 = NAND(g12711, g3722)
--	g13557 = NAND(g12611, g3410)
--	g13558 = NAND(g12657, g3566)
--	g13559 = NAND(g12657, g3566)
--	g13560 = NAND(g12711, g3722)
--	g13561 = NAND(g12657, g3566)
--	g13562 = NAND(g12711, g3722)
--	g13563 = NAND(g12711, g3722)
--	g13564 = NAND(g12711, g3722)
--	g13599 = NAND(g12886, g3366)
--	g13611 = NAND(g12926, g3522)
--	g13621 = NAND(g12955, g3678)
--	g13633 = NAND(g12984, g3834)
--	g13893 = NAND(g8580, g12463)
--	g13915 = NAND(g8822, g12473, g12463)
--	g13934 = NAND(g8587, g12478)
--	g13957 = NAND(g10730, g12473)
--	g13971 = NAND(g8846, g12490, g12478)
--	g13990 = NAND(g8594, g12495)
--	g14027 = NAND(g10749, g12490)
--	g14041 = NAND(g8873, g12510, g12495)
--	g14060 = NAND(g8605, g12515)
--	g14118 = NAND(g10767, g12510)
--	g14132 = NAND(g8911, g12527, g12515)
--	g14233 = NAND(g10773, g12527)
--	g15454 = NAND(g9232, g9150, g12780)
--	g15540 = NAND(g9310, g9174, g12819)
--	g15618 = NAND(g9391, g9216, g12857)
--	g15660 = NAND(g13401, g12354)
--	g15664 = NAND(g12565, g6314)
--	g15694 = NAND(g9488, g9277, g12898)
--	g15718 = NAND(g13286, g12354)
--	g15719 = NAND(g13401, g12392)
--	g15720 = NAND(g12565, g6232)
--	g15721 = NAND(g12565, g6314)
--	g15723 = NAND(g12611, g6519)
--	g15756 = NAND(g13313, g12354)
--	g15757 = NAND(g11622, g12392)
--	g15758 = NAND(g12565, g6232)
--	g15759 = NAND(g12565, g6314)
--	g15760 = NAND(g12611, g6369)
--	g15761 = NAND(g12611, g6519)
--	g15763 = NAND(g12657, g6783)
--	g15782 = NAND(g13332, g12354)
--	g15783 = NAND(g11643, g12392)
--	g15784 = NAND(g12565, g6232)
--	g15785 = NAND(g12565, g6314)
--	g15786 = NAND(g12611, g6369)
--	g15787 = NAND(g12611, g6519)
--	g15788 = NAND(g12657, g6574)
--	g15789 = NAND(g12657, g6783)
--	g15791 = NAND(g12711, g7085)
--	g15803 = NAND(g13375, g12354)
--	g15804 = NAND(g11660, g12392)
--	g15805 = NAND(g12565, g6232)
--	g15806 = NAND(g12565, g6314)
--	g15807 = NAND(g12611, g6369)
--	g15808 = NAND(g12611, g6519)
--	g15809 = NAND(g12657, g6574)
--	g15810 = NAND(g12657, g6783)
--	g15811 = NAND(g12711, g6838)
--	g15812 = NAND(g12711, g7085)
--	I22062 = NAND(g12999, g12988)
--	I22063 = NAND(g12999, I22062)
--	I22064 = NAND(g12988, I22062)
--	g15814 = NAND(I22063, I22064)
--	g15818 = NAND(g13024, g12354)
--	g15819 = NAND(g13286, g12392)
--	g15820 = NAND(g12565, g6232)
--	g15821 = NAND(g12565, g6314)
--	g15822 = NAND(g12611, g6369)
--	g15823 = NAND(g12611, g6519)
--	g15824 = NAND(g12657, g6574)
--	g15825 = NAND(g12657, g6783)
--	g15826 = NAND(g12711, g6838)
--	g15827 = NAND(g12711, g7085)
--	g15830 = NAND(g13310, g12392)
--	g15831 = NAND(g13313, g12392)
--	g15832 = NAND(g12565, g6232)
--	g15833 = NAND(g12565, g6314)
--	g15834 = NAND(g12611, g6369)
--	g15835 = NAND(g12611, g6519)
--	g15836 = NAND(g12657, g6574)
--	g15837 = NAND(g12657, g6783)
--	g15838 = NAND(g12711, g6838)
--	g15839 = NAND(g12711, g7085)
--	g15841 = NAND(g13331, g12392)
--	g15842 = NAND(g13332, g12392)
--	g15843 = NAND(g12565, g6314)
--	g15844 = NAND(g12565, g6232)
--	g15845 = NAND(g12565, g6314)
--	g15846 = NAND(g12611, g6369)
--	g15847 = NAND(g12611, g6519)
--	g15848 = NAND(g12657, g6574)
--	g15849 = NAND(g12657, g6783)
--	g15850 = NAND(g12711, g6838)
--	g15851 = NAND(g12711, g7085)
--	g15853 = NAND(g13310, g12354)
--	g15854 = NAND(g13353, g12392)
--	g15855 = NAND(g13354, g12392)
--	g15856 = NAND(g12565, g6232)
--	g15857 = NAND(g12565, g6314)
--	g15858 = NAND(g12565, g6232)
--	g15866 = NAND(g12611, g6519)
--	g15867 = NAND(g12611, g6369)
--	g15868 = NAND(g12611, g6519)
--	g15869 = NAND(g12657, g6574)
--	g15870 = NAND(g12657, g6783)
--	g15871 = NAND(g12711, g6838)
--	g15872 = NAND(g12711, g7085)
--	g15877 = NAND(g13374, g12392)
--	g15878 = NAND(g13375, g12392)
--	g15879 = NAND(g12565, g6232)
--	g15887 = NAND(g12611, g6369)
--	g15888 = NAND(g12611, g6519)
--	g15889 = NAND(g12611, g6369)
--	g15897 = NAND(g12657, g6783)
--	g15898 = NAND(g12657, g6574)
--	g15899 = NAND(g12657, g6783)
--	g15900 = NAND(g12711, g6838)
--	g15901 = NAND(g12711, g7085)
--	g15903 = NAND(g13404, g12392)
--	g15912 = NAND(g12611, g6369)
--	g15920 = NAND(g12657, g6574)
--	g15921 = NAND(g12657, g6783)
--	g15922 = NAND(g12657, g6574)
--	g15930 = NAND(g12711, g7085)
--	g15931 = NAND(g12711, g6838)
--	g15932 = NAND(g12711, g7085)
--	g15941 = NAND(g12657, g6574)
--	g15949 = NAND(g12711, g6838)
--	g15950 = NAND(g12711, g7085)
--	g15951 = NAND(g12711, g6838)
--	g15970 = NAND(g12711, g6838)
--	g15990 = NAND(g12886, g6912)
--	g15992 = NAND(g12886, g6678)
--	g15993 = NAND(g12926, g7162)
--	g15995 = NAND(g12926, g6980)
--	g15996 = NAND(g12955, g7358)
--	g15999 = NAND(g12955, g7230)
--	g16000 = NAND(g12984, g7488)
--	g16006 = NAND(g12984, g7426)
--	g16085 = NAND(g12883, g633)
--	g16123 = NAND(g12923, g1319)
--	I22282 = NAND(g2962, g13348)
--	I22283 = NAND(g2962, I22282)
--	I22284 = NAND(g13348, I22282)
--	g16132 = NAND(I22283, I22284)
--	g16174 = NAND(g12952, g2013)
--	I22316 = NAND(g2934, g13370)
--	I22317 = NAND(g2934, I22316)
--	I22318 = NAND(g13370, I22316)
--	g16181 = NAND(I22317, I22318)
--	g16233 = NAND(g12981, g2707)
--	g16341 = NAND(g12377, g12407)
--	g16412 = NAND(g12565, g3254)
--	g16439 = NAND(g13082, g2912)
--	g16442 = NAND(g12565, g3254)
--	g16446 = NAND(g12611, g3410)
--	g16463 = NAND(g13004, g3018)
--	g16536 = NAND(g15873, g2896)
--	I22630 = NAND(g13507, g15978)
--	I22631 = NAND(g13507, I22630)
--	I22632 = NAND(g15978, I22630)
--	g16566 = NAND(I22631, I22632)
--	I22705 = NAND(g13348, g15661)
--	I22706 = NAND(g13348, I22705)
--	I22707 = NAND(g15661, I22705)
--	g16662 = NAND(I22706, I22707)
--	I22884 = NAND(g13370, g15661)
--	I22885 = NAND(g13370, I22884)
--	I22886 = NAND(g15661, I22884)
--	g16935 = NAND(I22885, I22886)
--	I22900 = NAND(g15022, g14000)
--	I22901 = NAND(g15022, I22900)
--	I22902 = NAND(g14000, I22900)
--	g16965 = NAND(I22901, I22902)
--	I22917 = NAND(g15096, g13945)
--	I22918 = NAND(g15096, I22917)
--	I22919 = NAND(g13945, I22917)
--	g16985 = NAND(I22918, I22919)
--	I22924 = NAND(g15118, g14091)
--	I22925 = NAND(g15118, I22924)
--	I22926 = NAND(g14091, I22924)
--	g16986 = NAND(I22925, I22926)
--	I22936 = NAND(g9150, g13906)
--	I22937 = NAND(g9150, I22936)
--	I22938 = NAND(g13906, I22936)
--	g16992 = NAND(I22937, I22938)
--	I22945 = NAND(g15188, g14015)
--	I22946 = NAND(g15188, I22945)
--	I22947 = NAND(g14015, I22945)
--	g16995 = NAND(I22946, I22947)
--	I22952 = NAND(g15210, g14206)
--	I22953 = NAND(g15210, I22952)
--	I22954 = NAND(g14206, I22952)
--	g16996 = NAND(I22953, I22954)
--	I22962 = NAND(g9161, g13885)
--	I22963 = NAND(g9161, I22962)
--	I22964 = NAND(g13885, I22962)
--	g17000 = NAND(I22963, I22964)
--	I22972 = NAND(g9174, g13962)
--	I22973 = NAND(g9174, I22972)
--	I22974 = NAND(g13962, I22972)
--	g17016 = NAND(I22973, I22974)
--	I22981 = NAND(g15274, g14106)
--	I22982 = NAND(g15274, I22981)
--	I22983 = NAND(g14106, I22981)
--	g17019 = NAND(I22982, I22983)
--	I22988 = NAND(g15296, g14321)
--	I22989 = NAND(g15296, I22988)
--	I22990 = NAND(g14321, I22988)
--	g17020 = NAND(I22989, I22990)
--	I22998 = NAND(g9187, g13872)
--	I22999 = NAND(g9187, I22998)
--	I23000 = NAND(g13872, I22998)
--	g17024 = NAND(I22999, I23000)
--	I23008 = NAND(g9203, g13926)
--	I23009 = NAND(g9203, I23008)
--	I23010 = NAND(g13926, I23008)
--	g17030 = NAND(I23009, I23010)
--	I23018 = NAND(g9216, g14032)
--	I23019 = NAND(g9216, I23018)
--	I23020 = NAND(g14032, I23018)
--	g17046 = NAND(I23019, I23020)
--	I23027 = NAND(g15366, g14221)
--	I23028 = NAND(g15366, I23027)
--	I23029 = NAND(g14221, I23027)
--	g17049 = NAND(I23028, I23029)
--	I23034 = NAND(g9232, g13864)
--	I23035 = NAND(g9232, I23034)
--	I23036 = NAND(g13864, I23034)
--	g17050 = NAND(I23035, I23036)
--	I23045 = NAND(g9248, g13894)
--	I23046 = NAND(g9248, I23045)
--	I23047 = NAND(g13894, I23045)
--	g17058 = NAND(I23046, I23047)
--	I23055 = NAND(g9264, g13982)
--	I23056 = NAND(g9264, I23055)
--	I23057 = NAND(g13982, I23055)
--	g17064 = NAND(I23056, I23057)
--	I23065 = NAND(g9277, g14123)
--	I23066 = NAND(g9277, I23065)
--	I23067 = NAND(g14123, I23065)
--	g17080 = NAND(I23066, I23067)
--	I23074 = NAND(g9293, g13856)
--	I23075 = NAND(g9293, I23074)
--	I23076 = NAND(g13856, I23074)
--	g17083 = NAND(I23075, I23076)
--	I23082 = NAND(g9310, g13879)
--	I23083 = NAND(g9310, I23082)
--	I23084 = NAND(g13879, I23082)
--	g17085 = NAND(I23083, I23084)
--	I23093 = NAND(g9326, g13935)
--	I23094 = NAND(g9326, I23093)
--	I23095 = NAND(g13935, I23093)
--	g17093 = NAND(I23094, I23095)
--	I23103 = NAND(g9342, g14052)
--	I23104 = NAND(g9342, I23103)
--	I23105 = NAND(g14052, I23103)
--	g17099 = NAND(I23104, I23105)
--	I23113 = NAND(g9356, g13848)
--	I23114 = NAND(g9356, I23113)
--	I23115 = NAND(g13848, I23113)
--	g17115 = NAND(I23114, I23115)
--	g17118 = NAND(g13915, g13893)
--	I23123 = NAND(g9374, g13866)
--	I23124 = NAND(g9374, I23123)
--	I23125 = NAND(g13866, I23123)
--	g17121 = NAND(I23124, I23125)
--	I23131 = NAND(g9391, g13901)
--	I23132 = NAND(g9391, I23131)
--	I23133 = NAND(g13901, I23131)
--	g17123 = NAND(I23132, I23133)
--	I23142 = NAND(g9407, g13991)
--	I23143 = NAND(g9407, I23142)
--	I23144 = NAND(g13991, I23142)
--	g17131 = NAND(I23143, I23144)
--	I23152 = NAND(g9427, g14061)
--	I23153 = NAND(g9427, I23152)
--	I23154 = NAND(g14061, I23152)
--	g17137 = NAND(I23153, I23154)
--	g17139 = NAND(g13957, g13915)
--	I23161 = NAND(g9453, g13857)
--	I23162 = NAND(g9453, I23161)
--	I23163 = NAND(g13857, I23161)
--	g17142 = NAND(I23162, I23163)
--	g17145 = NAND(g13971, g13934)
--	I23171 = NAND(g9471, g13881)
--	I23172 = NAND(g9471, I23171)
--	I23173 = NAND(g13881, I23171)
--	g17148 = NAND(I23172, I23173)
--	I23179 = NAND(g9488, g13942)
--	I23180 = NAND(g9488, I23179)
--	I23181 = NAND(g13942, I23179)
--	g17150 = NAND(I23180, I23181)
--	I23190 = NAND(g9507, g13999)
--	I23191 = NAND(g9507, I23190)
--	I23192 = NAND(g13999, I23190)
--	g17158 = NAND(I23191, I23192)
--	g17159 = NAND(g14642, g14657)
--	I23198 = NAND(g9569, g14176)
--	I23199 = NAND(g9569, I23198)
--	I23200 = NAND(g14176, I23198)
--	g17160 = NAND(I23199, I23200)
--	g17162 = NAND(g14027, g13971)
--	I23207 = NAND(g9595, g13867)
--	I23208 = NAND(g9595, I23207)
--	I23209 = NAND(g13867, I23207)
--	g17165 = NAND(I23208, I23209)
--	g17168 = NAND(g14041, g13990)
--	I23217 = NAND(g9613, g13903)
--	I23218 = NAND(g9613, I23217)
--	I23219 = NAND(g13903, I23217)
--	g17171 = NAND(I23218, I23219)
--	I23225 = NAND(g9649, g14090)
--	I23226 = NAND(g9649, I23225)
--	I23227 = NAND(g14090, I23225)
--	g17173 = NAND(I23226, I23227)
--	g17174 = NAND(g14669, g14691)
--	I23233 = NAND(g9711, g14291)
--	I23234 = NAND(g9711, I23233)
--	I23235 = NAND(g14291, I23233)
--	g17175 = NAND(I23234, I23235)
--	g17177 = NAND(g14118, g14041)
--	I23242 = NAND(g9737, g13882)
--	I23243 = NAND(g9737, I23242)
--	I23244 = NAND(g13882, I23242)
--	g17180 = NAND(I23243, I23244)
--	g17183 = NAND(g14132, g14060)
--	I23256 = NAND(g9795, g14205)
--	I23257 = NAND(g9795, I23256)
--	I23258 = NAND(g14205, I23256)
--	g17190 = NAND(I23257, I23258)
--	g17191 = NAND(g14703, g14725)
--	I23264 = NAND(g9857, g14413)
--	I23265 = NAND(g9857, I23264)
--	I23266 = NAND(g14413, I23264)
--	g17192 = NAND(I23265, I23266)
--	g17194 = NAND(g14233, g14132)
--	I23277 = NAND(g9941, g14320)
--	I23278 = NAND(g9941, I23277)
--	I23279 = NAND(g14320, I23277)
--	g17201 = NAND(I23278, I23279)
--	g17202 = NAND(g14737, g14753)
--	I23806 = NAND(g14062, g9150)
--	I23807 = NAND(g14062, I23806)
--	I23808 = NAND(g9150, I23806)
--	g17729 = NAND(I23807, I23808)
--	I23878 = NAND(g14001, g9187)
--	I23879 = NAND(g14001, I23878)
--	I23880 = NAND(g9187, I23878)
--	g17807 = NAND(I23879, I23880)
--	I23893 = NAND(g14177, g9174)
--	I23894 = NAND(g14177, I23893)
--	I23895 = NAND(g9174, I23893)
--	g17830 = NAND(I23894, I23895)
--	I23941 = NAND(g13946, g9293)
--	I23942 = NAND(g13946, I23941)
--	I23943 = NAND(g9293, I23941)
--	g17887 = NAND(I23942, I23943)
--	I23958 = NAND(g6513, g14171)
--	I23959 = NAND(g6513, I23958)
--	I23960 = NAND(g14171, I23958)
--	g17913 = NAND(I23959, I23960)
--	I23966 = NAND(g14092, g9248)
--	I23967 = NAND(g14092, I23966)
--	I23968 = NAND(g9248, I23966)
--	g17919 = NAND(I23967, I23968)
--	I23981 = NAND(g14292, g9216)
--	I23982 = NAND(g14292, I23981)
--	I23983 = NAND(g9216, I23981)
--	g17942 = NAND(I23982, I23983)
--	I24005 = NAND(g7548, g15814)
--	I24006 = NAND(g7548, I24005)
--	I24007 = NAND(g15814, I24005)
--	g17968 = NAND(I24006, I24007)
--	I24015 = NAND(g13907, g9427)
--	I24016 = NAND(g13907, I24015)
--	I24017 = NAND(g9427, I24015)
--	g17979 = NAND(I24016, I24017)
--	g17985 = NAND(g14641, g9636)
--	I24028 = NAND(g6201, g14086)
--	I24029 = NAND(g6201, I24028)
--	I24030 = NAND(g14086, I24028)
--	g17992 = NAND(I24029, I24030)
--	I24036 = NAND(g14016, g9374)
--	I24037 = NAND(g14016, I24036)
--	I24038 = NAND(g9374, I24036)
--	g17998 = NAND(I24037, I24038)
--	I24053 = NAND(g6777, g14286)
--	I24054 = NAND(g6777, I24053)
--	I24055 = NAND(g14286, I24053)
--	g18024 = NAND(I24054, I24055)
--	I24061 = NAND(g14207, g9326)
--	I24062 = NAND(g14207, I24061)
--	I24063 = NAND(g9326, I24061)
--	g18030 = NAND(I24062, I24063)
--	I24076 = NAND(g14414, g9277)
--	I24077 = NAND(g14414, I24076)
--	I24078 = NAND(g9277, I24076)
--	g18053 = NAND(I24077, I24078)
--	I24091 = NAND(g13886, g15096)
--	I24092 = NAND(g13886, I24091)
--	I24093 = NAND(g15096, I24091)
--	g18079 = NAND(I24092, I24093)
--	I24102 = NAND(g6363, g14011)
--	I24103 = NAND(g6363, I24102)
--	I24104 = NAND(g14011, I24102)
--	g18090 = NAND(I24103, I24104)
--	I24110 = NAND(g13963, g9569)
--	I24111 = NAND(g13963, I24110)
--	I24112 = NAND(g9569, I24110)
--	g18096 = NAND(I24111, I24112)
--	g18102 = NAND(g14668, g9782)
--	I24123 = NAND(g6290, g14201)
--	I24124 = NAND(g6290, I24123)
--	I24125 = NAND(g14201, I24123)
--	g18109 = NAND(I24124, I24125)
--	I24131 = NAND(g14107, g9471)
--	I24132 = NAND(g14107, I24131)
--	I24133 = NAND(g9471, I24131)
--	g18115 = NAND(I24132, I24133)
--	I24148 = NAND(g7079, g14408)
--	I24149 = NAND(g7079, I24148)
--	I24150 = NAND(g14408, I24148)
--	g18141 = NAND(I24149, I24150)
--	I24156 = NAND(g14322, g9407)
--	I24157 = NAND(g14322, I24156)
--	I24158 = NAND(g9407, I24156)
--	g18147 = NAND(I24157, I24158)
--	I24178 = NAND(g13873, g9161)
--	I24179 = NAND(g13873, I24178)
--	I24180 = NAND(g9161, I24178)
--	g18183 = NAND(I24179, I24180)
--	I24186 = NAND(g6177, g13958)
--	I24187 = NAND(g6177, I24186)
--	I24188 = NAND(g13958, I24186)
--	g18189 = NAND(I24187, I24188)
--	I24194 = NAND(g13927, g15188)
--	I24195 = NAND(g13927, I24194)
--	I24196 = NAND(g15188, I24194)
--	g18195 = NAND(I24195, I24196)
--	I24205 = NAND(g6568, g14102)
--	I24206 = NAND(g6568, I24205)
--	I24207 = NAND(g14102, I24205)
--	g18206 = NAND(I24206, I24207)
--	I24213 = NAND(g14033, g9711)
--	I24214 = NAND(g14033, I24213)
--	I24215 = NAND(g9711, I24213)
--	g18212 = NAND(I24214, I24215)
--	g18218 = NAND(g14702, g9928)
--	I24226 = NAND(g6427, g14316)
--	I24227 = NAND(g6427, I24226)
--	I24228 = NAND(g14316, I24226)
--	g18225 = NAND(I24227, I24228)
--	I24234 = NAND(g14222, g9613)
--	I24235 = NAND(g14222, I24234)
--	I24236 = NAND(g9613, I24234)
--	g18231 = NAND(I24235, I24236)
--	I24251 = NAND(g7329, g14520)
--	I24252 = NAND(g7329, I24251)
--	I24253 = NAND(g14520, I24251)
--	g18257 = NAND(I24252, I24253)
--	I24263 = NAND(g14342, g9232)
--	I24264 = NAND(g14342, I24263)
--	I24265 = NAND(g9232, I24263)
--	g18270 = NAND(I24264, I24265)
--	I24271 = NAND(g6180, g13922)
--	I24272 = NAND(g6180, I24271)
--	I24273 = NAND(g13922, I24271)
--	g18276 = NAND(I24272, I24273)
--	I24278 = NAND(g6284, g13918)
--	I24279 = NAND(g6284, I24278)
--	I24280 = NAND(g13918, I24278)
--	g18277 = NAND(I24279, I24280)
--	I24290 = NAND(g13895, g9203)
--	I24291 = NAND(g13895, I24290)
--	I24292 = NAND(g9203, I24290)
--	g18290 = NAND(I24291, I24292)
--	I24298 = NAND(g6209, g14028)
--	I24299 = NAND(g6209, I24298)
--	I24300 = NAND(g14028, I24298)
--	g18296 = NAND(I24299, I24300)
--	I24306 = NAND(g13983, g15274)
--	I24307 = NAND(g13983, I24306)
--	I24308 = NAND(g15274, I24306)
--	g18302 = NAND(I24307, I24308)
--	I24317 = NAND(g6832, g14217)
--	I24318 = NAND(g6832, I24317)
--	I24319 = NAND(g14217, I24317)
--	g18313 = NAND(I24318, I24319)
--	I24325 = NAND(g14124, g9857)
--	I24326 = NAND(g14124, I24325)
--	I24327 = NAND(g9857, I24325)
--	g18319 = NAND(I24326, I24327)
--	g18325 = NAND(g14736, g10082)
--	I24338 = NAND(g6632, g14438)
--	I24339 = NAND(g6632, I24338)
--	I24340 = NAND(g14438, I24338)
--	g18332 = NAND(I24339, I24340)
--	I24351 = NAND(g14238, g9356)
--	I24352 = NAND(g14238, I24351)
--	I24353 = NAND(g9356, I24351)
--	g18346 = NAND(I24352, I24353)
--	I24361 = NAND(g6157, g14525)
--	I24362 = NAND(g6157, I24361)
--	I24363 = NAND(g14525, I24361)
--	g18354 = NAND(I24362, I24363)
--	I24372 = NAND(g14454, g9310)
--	I24373 = NAND(g14454, I24372)
--	I24374 = NAND(g9310, I24372)
--	g18363 = NAND(I24373, I24374)
--	I24380 = NAND(g6212, g13978)
--	I24381 = NAND(g6212, I24380)
--	I24382 = NAND(g13978, I24380)
--	g18369 = NAND(I24381, I24382)
--	I24387 = NAND(g6421, g13974)
--	I24388 = NAND(g6421, I24387)
--	I24389 = NAND(g13974, I24387)
--	g18370 = NAND(I24388, I24389)
--	I24399 = NAND(g13936, g9264)
--	I24400 = NAND(g13936, I24399)
--	I24401 = NAND(g9264, I24399)
--	g18383 = NAND(I24400, I24401)
--	I24407 = NAND(g6298, g14119)
--	I24408 = NAND(g6298, I24407)
--	I24409 = NAND(g14119, I24407)
--	g18389 = NAND(I24408, I24409)
--	I24415 = NAND(g14053, g15366)
--	I24416 = NAND(g14053, I24415)
--	I24417 = NAND(g15366, I24415)
--	g18395 = NAND(I24416, I24417)
--	I24426 = NAND(g7134, g14332)
--	I24427 = NAND(g7134, I24426)
--	I24428 = NAND(g14332, I24426)
--	g18406 = NAND(I24427, I24428)
--	I24436 = NAND(g14153, g15022)
--	I24437 = NAND(g14153, I24436)
--	I24438 = NAND(g15022, I24436)
--	g18419 = NAND(I24437, I24438)
--	I24443 = NAND(g14148, g9507)
--	I24444 = NAND(g14148, I24443)
--	I24445 = NAND(g9507, I24443)
--	g18424 = NAND(I24444, I24445)
--	I24452 = NAND(g6142, g14450)
--	I24453 = NAND(g6142, I24452)
--	I24454 = NAND(g14450, I24452)
--	g18431 = NAND(I24453, I24454)
--	I24464 = NAND(g14360, g9453)
--	I24465 = NAND(g14360, I24464)
--	I24466 = NAND(g9453, I24464)
--	g18441 = NAND(I24465, I24466)
--	I24474 = NAND(g6184, g14580)
--	I24475 = NAND(g6184, I24474)
--	I24476 = NAND(g14580, I24474)
--	g18449 = NAND(I24475, I24476)
--	I24485 = NAND(g14541, g9391)
--	I24486 = NAND(g14541, I24485)
--	I24487 = NAND(g9391, I24485)
--	g18458 = NAND(I24486, I24487)
--	I24493 = NAND(g6301, g14048)
--	I24494 = NAND(g6301, I24493)
--	I24495 = NAND(g14048, I24493)
--	g18464 = NAND(I24494, I24495)
--	I24500 = NAND(g6626, g14044)
--	I24501 = NAND(g6626, I24500)
--	I24502 = NAND(g14044, I24500)
--	g18465 = NAND(I24501, I24502)
--	I24512 = NAND(g13992, g9342)
--	I24513 = NAND(g13992, I24512)
--	I24514 = NAND(g9342, I24512)
--	g18478 = NAND(I24513, I24514)
--	I24520 = NAND(g6435, g14234)
--	I24521 = NAND(g6435, I24520)
--	I24522 = NAND(g14234, I24520)
--	g18484 = NAND(I24521, I24522)
--	I24530 = NAND(g6707, g14355)
--	I24531 = NAND(g6707, I24530)
--	I24532 = NAND(g14355, I24530)
--	g18491 = NAND(I24531, I24532)
--	I24537 = NAND(g14268, g15118)
--	I24538 = NAND(g14268, I24537)
--	I24539 = NAND(g15118, I24537)
--	g18492 = NAND(I24538, I24539)
--	I24544 = NAND(g14263, g9649)
--	I24545 = NAND(g14263, I24544)
--	I24546 = NAND(g9649, I24544)
--	g18497 = NAND(I24545, I24546)
--	I24553 = NAND(g6163, g14537)
--	I24554 = NAND(g6163, I24553)
--	I24555 = NAND(g14537, I24553)
--	g18504 = NAND(I24554, I24555)
--	I24565 = NAND(g14472, g9595)
--	I24566 = NAND(g14472, I24565)
--	I24567 = NAND(g9595, I24565)
--	g18514 = NAND(I24566, I24567)
--	I24575 = NAND(g6216, g14614)
--	I24576 = NAND(g6216, I24575)
--	I24577 = NAND(g14614, I24575)
--	g18522 = NAND(I24576, I24577)
--	I24586 = NAND(g14596, g9488)
--	I24587 = NAND(g14596, I24586)
--	I24588 = NAND(g9488, I24586)
--	g18531 = NAND(I24587, I24588)
--	I24594 = NAND(g6438, g14139)
--	I24595 = NAND(g6438, I24594)
--	I24596 = NAND(g14139, I24594)
--	g18537 = NAND(I24595, I24596)
--	I24601 = NAND(g6890, g14135)
--	I24602 = NAND(g6890, I24601)
--	I24603 = NAND(g14135, I24601)
--	g18538 = NAND(I24602, I24603)
--	I24611 = NAND(g15814, g15978)
--	I24612 = NAND(g15814, I24611)
--	I24613 = NAND(g15978, I24611)
--	g18542 = NAND(I24612, I24613)
--	I24624 = NAND(g6136, g14252)
--	I24625 = NAND(g6136, I24624)
--	I24626 = NAND(g14252, I24624)
--	g18553 = NAND(I24625, I24626)
--	I24632 = NAND(g7009, g14467)
--	I24633 = NAND(g7009, I24632)
--	I24634 = NAND(g14467, I24632)
--	g18555 = NAND(I24633, I24634)
--	I24639 = NAND(g14390, g15210)
--	I24640 = NAND(g14390, I24639)
--	I24641 = NAND(g15210, I24639)
--	g18556 = NAND(I24640, I24641)
--	I24646 = NAND(g14385, g9795)
--	I24647 = NAND(g14385, I24646)
--	I24648 = NAND(g9795, I24646)
--	g18561 = NAND(I24647, I24648)
--	I24655 = NAND(g6190, g14592)
--	I24656 = NAND(g6190, I24655)
--	I24657 = NAND(g14592, I24655)
--	g18568 = NAND(I24656, I24657)
--	I24667 = NAND(g14559, g9737)
--	I24668 = NAND(g14559, I24667)
--	I24669 = NAND(g9737, I24667)
--	g18578 = NAND(I24668, I24669)
--	I24677 = NAND(g6305, g14637)
--	I24678 = NAND(g6305, I24677)
--	I24679 = NAND(g14637, I24677)
--	g18586 = NAND(I24678, I24679)
--	I24694 = NAND(g6146, g14374)
--	I24695 = NAND(g6146, I24694)
--	I24696 = NAND(g14374, I24694)
--	g18603 = NAND(I24695, I24696)
--	I24702 = NAND(g7259, g14554)
--	I24703 = NAND(g7259, I24702)
--	I24704 = NAND(g14554, I24702)
--	g18605 = NAND(I24703, I24704)
--	I24709 = NAND(g14502, g15296)
--	I24710 = NAND(g14502, I24709)
--	I24711 = NAND(g15296, I24709)
--	g18606 = NAND(I24710, I24711)
--	I24716 = NAND(g14497, g9941)
--	I24717 = NAND(g14497, I24716)
--	I24718 = NAND(g9941, I24716)
--	g18611 = NAND(I24717, I24718)
--	I24725 = NAND(g6222, g14626)
--	I24726 = NAND(g6222, I24725)
--	I24727 = NAND(g14626, I24725)
--	g18618 = NAND(I24726, I24727)
--	I24743 = NAND(g6167, g14486)
--	I24744 = NAND(g6167, I24743)
--	I24745 = NAND(g14486, I24743)
--	g18635 = NAND(I24744, I24745)
--	I24751 = NAND(g7455, g14609)
--	I24752 = NAND(g7455, I24751)
--	I24753 = NAND(g14609, I24751)
--	g18637 = NAND(I24752, I24753)
--	I24763 = NAND(g6194, g14573)
--	I24764 = NAND(g6194, I24763)
--	I24765 = NAND(g14573, I24763)
--	g18644 = NAND(I24764, I24765)
--	g18977 = NAND(g15797, g3006)
--	I25030 = NAND(g8029, g13507)
--	I25031 = NAND(g8029, I25030)
--	I25032 = NAND(g13507, I25030)
--	g18980 = NAND(I25031, I25032)
--	g19067 = NAND(g16554, g16578)
--	g19084 = NAND(g16586, g16602)
--	g19103 = NAND(g18590, g2924)
--	g19121 = NAND(g16682, g16697)
--	g19128 = NAND(g16708, g16728)
--	g19135 = NAND(g16739, g16770)
--	g19138 = NAND(g16781, g16797)
--	g19141 = NAND(g3088, g16825)
--	g19152 = NAND(g5378, g18884)
--	I25532 = NAND(g52, g18179)
--	I25533 = NAND(g52, I25532)
--	I25534 = NAND(g18179, I25532)
--	g19261 = NAND(I25533, I25534)
--	I25539 = NAND(g92, g18174)
--	I25540 = NAND(g92, I25539)
--	I25541 = NAND(g18174, I25539)
--	g19262 = NAND(I25540, I25541)
--	I25560 = NAND(g56, g17724)
--	I25561 = NAND(g56, I25560)
--	I25562 = NAND(g17724, I25560)
--	g19271 = NAND(I25561, I25562)
--	I25571 = NAND(g740, g18286)
--	I25572 = NAND(g740, I25571)
--	I25573 = NAND(g18286, I25571)
--	g19276 = NAND(I25572, I25573)
--	I25578 = NAND(g780, g18281)
--	I25579 = NAND(g780, I25578)
--	I25580 = NAND(g18281, I25578)
--	g19277 = NAND(I25579, I25580)
--	I25595 = NAND(g61, g18074)
--	I25596 = NAND(g61, I25595)
--	I25597 = NAND(g18074, I25595)
--	g19286 = NAND(I25596, I25597)
--	g19288 = NAND(g14685, g8580, g17057)
--	I25605 = NAND(g744, g17825)
--	I25606 = NAND(g744, I25605)
--	I25607 = NAND(g17825, I25605)
--	g19290 = NAND(I25606, I25607)
--	I25616 = NAND(g1426, g18379)
--	I25617 = NAND(g1426, I25616)
--	I25618 = NAND(g18379, I25616)
--	g19295 = NAND(I25617, I25618)
--	I25623 = NAND(g1466, g18374)
--	I25624 = NAND(g1466, I25623)
--	I25625 = NAND(g18374, I25623)
--	g19296 = NAND(I25624, I25625)
--	I25633 = NAND(g65, g17640)
--	I25634 = NAND(g65, I25633)
--	I25635 = NAND(g17640, I25633)
--	g19300 = NAND(I25634, I25635)
--	I25643 = NAND(g749, g18190)
--	I25644 = NAND(g749, I25643)
--	I25645 = NAND(g18190, I25643)
--	g19304 = NAND(I25644, I25645)
--	g19306 = NAND(g14719, g8587, g17092)
--	I25653 = NAND(g1430, g17937)
--	I25654 = NAND(g1430, I25653)
--	I25655 = NAND(g17937, I25653)
--	g19308 = NAND(I25654, I25655)
--	I25664 = NAND(g2120, g18474)
--	I25665 = NAND(g2120, I25664)
--	I25666 = NAND(g18474, I25664)
--	g19313 = NAND(I25665, I25666)
--	I25671 = NAND(g2160, g18469)
--	I25672 = NAND(g2160, I25671)
--	I25673 = NAND(g18469, I25671)
--	g19314 = NAND(I25672, I25673)
--	I25681 = NAND(g70, g17974)
--	I25682 = NAND(g70, I25681)
--	I25683 = NAND(g17974, I25681)
--	g19318 = NAND(I25682, I25683)
--	I25690 = NAND(g753, g17741)
--	I25691 = NAND(g753, I25690)
--	I25692 = NAND(g17741, I25690)
--	g19321 = NAND(I25691, I25692)
--	I25700 = NAND(g1435, g18297)
--	I25701 = NAND(g1435, I25700)
--	I25702 = NAND(g18297, I25700)
--	g19325 = NAND(I25701, I25702)
--	g19327 = NAND(g14747, g8594, g17130)
--	I25710 = NAND(g2124, g18048)
--	I25711 = NAND(g2124, I25710)
--	I25712 = NAND(g18048, I25710)
--	g19329 = NAND(I25711, I25712)
--	I25721 = NAND(g74, g18341)
--	I25722 = NAND(g74, I25721)
--	I25723 = NAND(g18341, I25721)
--	g19334 = NAND(I25722, I25723)
--	I25731 = NAND(g758, g18091)
--	I25732 = NAND(g758, I25731)
--	I25733 = NAND(g18091, I25731)
--	g19345 = NAND(I25732, I25733)
--	I25740 = NAND(g1439, g17842)
--	I25741 = NAND(g1439, I25740)
--	I25742 = NAND(g17842, I25740)
--	g19348 = NAND(I25741, I25742)
--	I25750 = NAND(g2129, g18390)
--	I25751 = NAND(g2129, I25750)
--	I25752 = NAND(g18390, I25750)
--	g19352 = NAND(I25751, I25752)
--	g19354 = NAND(g14768, g8605, g17157)
--	I25761 = NAND(g79, g17882)
--	I25762 = NAND(g79, I25761)
--	I25763 = NAND(g17882, I25761)
--	g19357 = NAND(I25762, I25763)
--	I25771 = NAND(g762, g18436)
--	I25772 = NAND(g762, I25771)
--	I25773 = NAND(g18436, I25771)
--	g19368 = NAND(I25772, I25773)
--	I25781 = NAND(g1444, g18207)
--	I25782 = NAND(g1444, I25781)
--	I25783 = NAND(g18207, I25781)
--	g19379 = NAND(I25782, I25783)
--	I25790 = NAND(g2133, g17954)
--	I25791 = NAND(g2133, I25790)
--	I25792 = NAND(g17954, I25790)
--	g19382 = NAND(I25791, I25792)
--	I25800 = NAND(g83, g18265)
--	I25801 = NAND(g83, I25800)
--	I25802 = NAND(g18265, I25800)
--	g19386 = NAND(I25801, I25802)
--	I25809 = NAND(g767, g17993)
--	I25810 = NAND(g767, I25809)
--	I25811 = NAND(g17993, I25809)
--	g19389 = NAND(I25810, I25811)
--	I25819 = NAND(g1448, g18509)
--	I25820 = NAND(g1448, I25819)
--	I25821 = NAND(g18509, I25819)
--	g19400 = NAND(I25820, I25821)
--	I25829 = NAND(g2138, g18314)
--	I25830 = NAND(g2138, I25829)
--	I25831 = NAND(g18314, I25829)
--	g19411 = NAND(I25830, I25831)
--	I25838 = NAND(g88, g17802)
--	I25839 = NAND(g88, I25838)
--	I25840 = NAND(g17802, I25838)
--	g19414 = NAND(I25839, I25840)
--	I25846 = NAND(g771, g18358)
--	I25847 = NAND(g771, I25846)
--	I25848 = NAND(g18358, I25846)
--	g19416 = NAND(I25847, I25848)
--	I25855 = NAND(g1453, g18110)
--	I25856 = NAND(g1453, I25855)
--	I25857 = NAND(g18110, I25855)
--	g19419 = NAND(I25856, I25857)
--	I25865 = NAND(g2142, g18573)
--	I25866 = NAND(g2142, I25865)
--	I25867 = NAND(g18573, I25865)
--	g19430 = NAND(I25866, I25867)
--	I25880 = NAND(g776, g17914)
--	I25881 = NAND(g776, I25880)
--	I25882 = NAND(g17914, I25880)
--	g19451 = NAND(I25881, I25882)
--	I25888 = NAND(g1457, g18453)
--	I25889 = NAND(g1457, I25888)
--	I25890 = NAND(g18453, I25888)
--	g19453 = NAND(I25889, I25890)
--	I25897 = NAND(g2147, g18226)
--	I25898 = NAND(g2147, I25897)
--	I25899 = NAND(g18226, I25897)
--	g19456 = NAND(I25898, I25899)
--	I25913 = NAND(g1462, g18025)
--	I25914 = NAND(g1462, I25913)
--	I25915 = NAND(g18025, I25913)
--	g19478 = NAND(I25914, I25915)
--	I25921 = NAND(g2151, g18526)
--	I25922 = NAND(g2151, I25921)
--	I25923 = NAND(g18526, I25921)
--	g19480 = NAND(I25922, I25923)
--	I25938 = NAND(g2156, g18142)
--	I25939 = NAND(g2156, I25938)
--	I25940 = NAND(g18142, I25938)
--	g19501 = NAND(I25939, I25940)
--	g19865 = NAND(g16607, g9636)
--	g19896 = NAND(g16625, g9782)
--	g19921 = NAND(g16639, g9928)
--	g19936 = NAND(g16650, g10082)
--	g19954 = NAND(g17186, g92)
--	g19984 = NAND(g17197, g780)
--	g20022 = NAND(g17204, g1466)
--	g20064 = NAND(g17209, g2160)
--	g20473 = NAND(g18085, g646)
--	g20481 = NAND(g18201, g1332)
--	g20487 = NAND(g18308, g2026)
--	g20493 = NAND(g18401, g2720)
--	g20497 = NAND(g5410, g18886)
--	g20522 = NAND(g16501, g16515)
--	g20537 = NAND(g18626, g3036)
--	g20542 = NAND(g16523, g16546)
--	g20633 = NAND(g20164, g3254)
--	g20648 = NAND(g20164, g3254)
--	g20658 = NAND(g20198, g3410)
--	g20672 = NAND(g20164, g3254)
--	g20683 = NAND(g20198, g3410)
--	g20693 = NAND(g20228, g3566)
--	g20700 = NAND(g20153, g2903)
--	g20703 = NAND(g20164, g3254)
--	g20707 = NAND(g20198, g3410)
--	g20718 = NAND(g20228, g3566)
--	g20728 = NAND(g20255, g3722)
--	g20738 = NAND(g20198, g3410)
--	g20742 = NAND(g20228, g3566)
--	g20753 = NAND(g20255, g3722)
--	g20775 = NAND(g20228, g3566)
--	g20779 = NAND(g20255, g3722)
--	g20805 = NAND(g20255, g3722)
--	g20825 = NAND(g19219, g15959)
--	g21659 = NAND(g20164, g6314)
--	I28189 = NAND(g14079, g19444)
--	I28190 = NAND(g14079, I28189)
--	I28191 = NAND(g19444, I28189)
--	g21660 = NAND(I28190, I28191)
--	g21685 = NAND(g20164, g6232)
--	g21686 = NAND(g20164, g6314)
--	g21688 = NAND(g20198, g6519)
--	I28217 = NAND(g14194, g19471)
--	I28218 = NAND(g14194, I28217)
--	I28219 = NAND(g19471, I28217)
--	g21689 = NAND(I28218, I28219)
--	g21714 = NAND(g20164, g6232)
--	g21715 = NAND(g20164, g6314)
--	g21720 = NAND(g14256, g15177, g19871, g19842)
--	g21721 = NAND(g20198, g6369)
--	g21722 = NAND(g20198, g6519)
--	g21724 = NAND(g20228, g6783)
--	I28247 = NAND(g14309, g19494)
--	I28248 = NAND(g14309, I28247)
--	I28249 = NAND(g19494, I28247)
--	g21725 = NAND(I28248, I28249)
--	g21736 = NAND(g20164, g6232)
--	g21737 = NAND(g20164, g6314)
--	g21740 = NAND(g20198, g6369)
--	g21741 = NAND(g20198, g6519)
--	g21746 = NAND(g14378, g15263, g19902, g19875)
--	g21747 = NAND(g20228, g6574)
--	g21748 = NAND(g20228, g6783)
--	g21750 = NAND(g20255, g7085)
--	I28271 = NAND(g14431, g19515)
--	I28272 = NAND(g14431, I28271)
--	I28273 = NAND(g19515, I28271)
--	g21751 = NAND(I28272, I28273)
--	g21759 = NAND(g20164, g6232)
--	g21760 = NAND(g20198, g6369)
--	g21761 = NAND(g20198, g6519)
--	g21764 = NAND(g20228, g6574)
--	g21765 = NAND(g20228, g6783)
--	g21770 = NAND(g14490, g15355, g19927, g19906)
--	g21771 = NAND(g20255, g6838)
--	g21772 = NAND(g20255, g7085)
--	g21775 = NAND(g20198, g6369)
--	g21776 = NAND(g20228, g6574)
--	g21777 = NAND(g20228, g6783)
--	g21780 = NAND(g20255, g6838)
--	g21781 = NAND(g20255, g7085)
--	g21786 = NAND(g14577, g15441, g19942, g19931)
--	g21790 = NAND(g20228, g6574)
--	g21791 = NAND(g20255, g6838)
--	g21792 = NAND(g20255, g7085)
--	g21804 = NAND(g20255, g6838)
--	g21848 = NAND(g17807, g19181, g19186)
--	g21850 = NAND(g17979, g19187, g19191)
--	g21855 = NAND(g17919, g19188, g19193)
--	g21857 = NAND(g18079, g19192, g19200)
--	g21858 = NAND(g18096, g19194, g19202)
--	g21859 = NAND(g18030, g19195, g19204)
--	g21860 = NAND(g18270, g19201, g19209)
--	g21862 = NAND(g18195, g19203, g19211)
--	g21863 = NAND(g18212, g19205, g19213)
--	g21864 = NAND(g18147, g19206, g19215)
--	g21865 = NAND(g18424, g19210, g19221)
--	g21866 = NAND(g18363, g19212, g19222)
--	g21868 = NAND(g18302, g19214, g19224)
--	g21869 = NAND(g18319, g19216, g19226)
--	g21870 = NAND(g18497, g19223, g19231)
--	g21871 = NAND(g18458, g19225, g19232)
--	g21873 = NAND(g18395, g19227, g19234)
--	g21874 = NAND(g18561, g19233, g19244)
--	g21875 = NAND(g18531, g19235, g19245)
--	g21877 = NAND(g18611, g19246, g19257)
--	g21879 = NAND(g18419, g19250, g19263)
--	g21881 = NAND(g18492, g19264, g19278)
--	g21885 = NAND(g18556, g19279, g19297)
--	g21888 = NAND(g18606, g19298, g19315)
--	g21903 = NAND(g20008, g3013)
--	g21976 = NAND(g19242, g21120, g19275)
--	g21983 = NAND(g19255, g21139, g19294)
--	g21989 = NAND(g21048, g18623)
--	g21991 = NAND(g21501, g21536)
--	g21996 = NAND(g19268, g21159, g19312)
--	g22002 = NAND(g21065, g21711)
--	g22005 = NAND(g21540, g21572)
--	g22009 = NAND(g19283, g21179, g19333)
--	g22016 = NAND(g21576, g21605)
--	g22021 = NAND(g21609, g21634)
--	g22050 = NAND(g19450, g21244, g19503)
--	g22069 = NAND(g19477, g21253, g19522)
--	g22083 = NAND(g21774, g21787)
--	g22093 = NAND(g19500, g21261, g19532)
--	g22108 = NAND(g21789, g21801)
--	g22118 = NAND(g19521, g21269, g19542)
--	g22134 = NAND(g21803, g21809)
--	g22157 = NAND(g21811, g21816)
--	I28726 = NAND(g21887, g13519)
--	I28727 = NAND(g21887, I28726)
--	I28728 = NAND(g13519, I28726)
--	g22188 = NAND(I28727, I28728)
--	I28741 = NAND(g21890, g13530)
--	I28742 = NAND(g21890, I28741)
--	I28743 = NAND(g13530, I28741)
--	g22197 = NAND(I28742, I28743)
--	I28753 = NAND(g21893, g13541)
--	I28754 = NAND(g21893, I28753)
--	I28755 = NAND(g13541, I28753)
--	g22203 = NAND(I28754, I28755)
--	I28765 = NAND(g21901, g13552)
--	I28766 = NAND(g21901, I28765)
--	I28767 = NAND(g13552, I28765)
--	g22209 = NAND(I28766, I28767)
--	g22317 = NAND(g21152, g21241, g21136)
--	g22339 = NAND(g14442, g21149, g10694)
--	g22342 = NAND(g21172, g21249, g21156)
--	g22362 = NAND(g14529, g21169, g10714)
--	g22365 = NAND(g21192, g21258, g21176)
--	g22381 = NAND(g21211, g14442, g10694)
--	g22382 = NAND(g14584, g21189, g10735)
--	g22385 = NAND(g21207, g21266, g21196)
--	g22396 = NAND(g21219, g14529, g10714)
--	g22397 = NAND(g14618, g21204, g10754)
--	g22399 = NAND(g21230, g14584, g10735)
--	g22400 = NAND(g21235, g14618, g10754)
--	g22608 = NAND(g20842, g20885)
--	g22644 = NAND(g20850, g20904)
--	g22668 = NAND(g16075, g21271)
--	g22680 = NAND(g20858, g20928)
--	g22708 = NAND(g16113, g21278)
--	g22720 = NAND(g20866, g20956)
--	g22739 = NAND(g16164, g21285)
--	g22771 = NAND(g16223, g21293)
--	g22809 = NAND(g21850, g21848, g21879)
--	g22844 = NAND(g21865, g21860, g21857)
--	g22845 = NAND(g19441, g20885)
--	g22846 = NAND(g8278, g21660)
--	g22850 = NAND(g21858, g21855, g21881)
--	g22876 = NAND(g21238, g83)
--	g22879 = NAND(g21870, g21866, g21862)
--	g22880 = NAND(g19468, g20904)
--	g22881 = NAND(g8287, g21689)
--	g22885 = NAND(g21863, g21859, g21885)
--	g22911 = NAND(g21246, g771)
--	g22914 = NAND(g21874, g21871, g21868)
--	g22915 = NAND(g19491, g20928)
--	g22916 = NAND(g8296, g21725)
--	g22920 = NAND(g21869, g21864, g21888)
--	g22936 = NAND(g21255, g1457)
--	g22939 = NAND(g21877, g21875, g21873)
--	g22940 = NAND(g19512, g20956)
--	g22941 = NAND(g8305, g21751)
--	g22942 = NAND(g21263, g2151)
--	g22992 = NAND(g21636, g672)
--	g23003 = NAND(g21667, g1358)
--	g23017 = NAND(g21696, g2052)
--	g23033 = NAND(g21732, g2746)
--	g23320 = NAND(g23066, g23051)
--	g23325 = NAND(g23080, g23070)
--	g23331 = NAND(g22999, g22174)
--	g23335 = NAND(g23096, g23083)
--	g23340 = NAND(g23013, g22189)
--	g23344 = NAND(g23113, g23099)
--	g23349 = NAND(g23029, g22198)
--	g23353 = NAND(g23046, g22204)
--	g23360 = NAND(g21980, g21975)
--	g23364 = NAND(g21987, g21981)
--	g23368 = NAND(g23135, g22288)
--	g23372 = NAND(g22000, g21988)
--	g23376 = NAND(g18435, g22812)
--	g23377 = NAND(g21968, g22308)
--	g23381 = NAND(g22013, g22001)
--	g23387 = NAND(g18508, g22852)
--	g23388 = NAND(g21971, g22336)
--	g23394 = NAND(g18572, g22887)
--	g23395 = NAND(g21973, g22361)
--	g23402 = NAND(g18622, g22922)
--	g23478 = NAND(g22809, g14442, g10694)
--	g23486 = NAND(g22844, g14442, g10694)
--	g23489 = NAND(g22850, g14529, g10714)
--	g23495 = NAND(g10694, g14442, g22316)
--	g23502 = NAND(g22879, g14529, g10714)
--	g23505 = NAND(g22885, g14584, g10735)
--	g23511 = NAND(g10714, g14529, g22341)
--	g23518 = NAND(g22914, g14584, g10735)
--	g23521 = NAND(g22920, g14618, g10754)
--	g23526 = NAND(g10735, g14584, g22364)
--	g23533 = NAND(g22939, g14618, g10754)
--	g23537 = NAND(g10754, g14618, g22384)
--	I30790 = NAND(g22846, g14079)
--	I30791 = NAND(g22846, I30790)
--	I30792 = NAND(g14079, I30790)
--	g23660 = NAND(I30791, I30792)
--	I30868 = NAND(g22881, g14194)
--	I30869 = NAND(g22881, I30868)
--	I30870 = NAND(g14194, I30868)
--	g23710 = NAND(I30869, I30870)
--	I30952 = NAND(g22916, g14309)
--	I30953 = NAND(g22916, I30952)
--	I30954 = NAND(g14309, I30952)
--	g23764 = NAND(I30953, I30954)
--	I31035 = NAND(g22941, g14431)
--	I31036 = NAND(g22941, I31035)
--	I31037 = NAND(g14431, I31035)
--	g23819 = NAND(I31036, I31037)
--	g23906 = NAND(g22812, g13958)
--	g23936 = NAND(g22812, g13922)
--	g23937 = NAND(g22812, g13918)
--	g23938 = NAND(g22852, g14028)
--	g23953 = NAND(g22812, g14525)
--	g23968 = NAND(g22852, g13978)
--	g23969 = NAND(g22852, g13974)
--	g23970 = NAND(g22887, g14119)
--	g23973 = NAND(g22812, g14450)
--	g23982 = NAND(g22852, g14580)
--	g23997 = NAND(g22887, g14048)
--	g23998 = NAND(g22887, g14044)
--	g23999 = NAND(g22922, g14234)
--	g24002 = NAND(g22812, g14355)
--	g24003 = NAND(g22852, g14537)
--	g24012 = NAND(g22887, g14614)
--	g24027 = NAND(g22922, g14139)
--	g24028 = NAND(g22922, g14135)
--	g24034 = NAND(g22812, g14252)
--	g24036 = NAND(g22852, g14467)
--	g24037 = NAND(g22887, g14592)
--	g24046 = NAND(g22922, g14637)
--	g24052 = NAND(g22812, g14171)
--	g24054 = NAND(g22852, g14374)
--	g24056 = NAND(g22887, g14554)
--	g24057 = NAND(g22922, g14626)
--	g24058 = NAND(g22812, g14086)
--	g24065 = NAND(g22852, g14286)
--	g24067 = NAND(g22887, g14486)
--	g24069 = NAND(g22922, g14609)
--	g24070 = NAND(g22812, g14011)
--	g24071 = NAND(g22852, g14201)
--	g24078 = NAND(g22887, g14408)
--	g24080 = NAND(g22922, g14573)
--	g24081 = NAND(g22852, g14102)
--	g24082 = NAND(g22887, g14316)
--	g24089 = NAND(g22922, g14520)
--	g24090 = NAND(g22887, g14217)
--	g24091 = NAND(g22922, g14438)
--	g24093 = NAND(g22922, g14332)
--	g24100 = NAND(g20885, g22175)
--	g24109 = NAND(g20904, g22190)
--	g24126 = NAND(g20928, g22199)
--	g24145 = NAND(g20956, g22205)
--	g24442 = NAND(g23644, g3306)
--	g24443 = NAND(g23644, g3306)
--	g24444 = NAND(g23694, g3462)
--	g24447 = NAND(g23644, g3306)
--	g24448 = NAND(g23923, g3338)
--	g24449 = NAND(g23694, g3462)
--	g24450 = NAND(g23748, g3618)
--	g24451 = NAND(g23644, g3306)
--	g24452 = NAND(g23923, g3338)
--	g24453 = NAND(g23694, g3462)
--	g24454 = NAND(g23955, g3494)
--	g24455 = NAND(g23748, g3618)
--	g24456 = NAND(g23803, g3774)
--	g24457 = NAND(g23923, g3338)
--	g24458 = NAND(g23694, g3462)
--	g24459 = NAND(g23955, g3494)
--	g24460 = NAND(g23748, g3618)
--	g24461 = NAND(g23984, g3650)
--	g24462 = NAND(g23803, g3774)
--	g24463 = NAND(g23923, g3338)
--	g24464 = NAND(g23955, g3494)
--	g24465 = NAND(g23748, g3618)
--	g24466 = NAND(g23984, g3650)
--	g24467 = NAND(g23803, g3774)
--	g24468 = NAND(g24014, g3806)
--	g24469 = NAND(g23955, g3494)
--	g24470 = NAND(g23984, g3650)
--	g24471 = NAND(g23803, g3774)
--	g24472 = NAND(g24014, g3806)
--	g24474 = NAND(g23984, g3650)
--	g24475 = NAND(g24014, g3806)
--	g24477 = NAND(g24014, g3806)
--	g24616 = NAND(g499, g23376)
--	g24627 = NAND(g1186, g23387)
--	g24641 = NAND(g1880, g23394)
--	g24660 = NAND(g2574, g23402)
--	I32265 = NAND(g17903, g23936)
--	I32266 = NAND(g17903, I32265)
--	I32267 = NAND(g23936, I32265)
--	g24753 = NAND(I32266, I32267)
--	I32284 = NAND(g17815, g23953)
--	I32285 = NAND(g17815, I32284)
--	I32286 = NAND(g23953, I32284)
--	g24766 = NAND(I32285, I32286)
--	I32295 = NAND(g18014, g23968)
--	I32296 = NAND(g18014, I32295)
--	I32297 = NAND(g23968, I32295)
--	g24771 = NAND(I32296, I32297)
--	I32308 = NAND(g17903, g23973)
--	I32309 = NAND(g17903, I32308)
--	I32310 = NAND(g23973, I32308)
--	g24778 = NAND(I32309, I32310)
--	I32323 = NAND(g17927, g23982)
--	I32324 = NAND(g17927, I32323)
--	I32325 = NAND(g23982, I32323)
--	g24787 = NAND(I32324, I32325)
--	I32333 = NAND(g18131, g23997)
--	I32334 = NAND(g18131, I32333)
--	I32335 = NAND(g23997, I32333)
--	g24791 = NAND(I32334, I32335)
--	I32345 = NAND(g17815, g24002)
--	I32346 = NAND(g17815, I32345)
--	I32347 = NAND(g24002, I32345)
--	g24797 = NAND(I32346, I32347)
--	I32355 = NAND(g18014, g24003)
--	I32356 = NAND(g18014, I32355)
--	I32357 = NAND(g24003, I32355)
--	g24801 = NAND(I32356, I32357)
--	I32368 = NAND(g18038, g24012)
--	I32369 = NAND(g18038, I32368)
--	I32370 = NAND(g24012, I32368)
--	g24808 = NAND(I32369, I32370)
--	I32378 = NAND(g18247, g24027)
--	I32379 = NAND(g18247, I32378)
--	I32380 = NAND(g24027, I32378)
--	g24812 = NAND(I32379, I32380)
--	g24814 = NAND(g24239, g24244)
--	I32391 = NAND(g17903, g24034)
--	I32392 = NAND(g17903, I32391)
--	I32393 = NAND(g24034, I32391)
--	g24817 = NAND(I32392, I32393)
--	I32400 = NAND(g17927, g24036)
--	I32401 = NAND(g17927, I32400)
--	I32402 = NAND(g24036, I32400)
--	g24820 = NAND(I32401, I32402)
--	I32409 = NAND(g18131, g24037)
--	I32410 = NAND(g18131, I32409)
--	I32411 = NAND(g24037, I32409)
--	g24823 = NAND(I32410, I32411)
--	I32422 = NAND(g18155, g24046)
--	I32423 = NAND(g18155, I32422)
--	I32424 = NAND(g24046, I32422)
--	g24830 = NAND(I32423, I32424)
--	I32430 = NAND(g17815, g24052)
--	I32431 = NAND(g17815, I32430)
--	I32432 = NAND(g24052, I32430)
--	g24832 = NAND(I32431, I32432)
--	g24833 = NAND(g24245, g24252)
--	I32443 = NAND(g18014, g24054)
--	I32444 = NAND(g18014, I32443)
--	I32445 = NAND(g24054, I32443)
--	g24837 = NAND(I32444, I32445)
--	I32451 = NAND(g18038, g24056)
--	I32452 = NAND(g18038, I32451)
--	I32453 = NAND(g24056, I32451)
--	g24839 = NAND(I32452, I32453)
--	I32460 = NAND(g18247, g24057)
--	I32461 = NAND(g18247, I32460)
--	I32462 = NAND(g24057, I32460)
--	g24842 = NAND(I32461, I32462)
--	I32468 = NAND(g17903, g24058)
--	I32469 = NAND(g17903, I32468)
--	I32470 = NAND(g24058, I32468)
--	g24844 = NAND(I32469, I32470)
--	I32478 = NAND(g17927, g24065)
--	I32479 = NAND(g17927, I32478)
--	I32480 = NAND(g24065, I32478)
--	g24848 = NAND(I32479, I32480)
--	g24849 = NAND(g24254, g24257)
--	I32490 = NAND(g18131, g24067)
--	I32491 = NAND(g18131, I32490)
--	I32492 = NAND(g24067, I32490)
--	g24852 = NAND(I32491, I32492)
--	I32498 = NAND(g18155, g24069)
--	I32499 = NAND(g18155, I32498)
--	I32500 = NAND(g24069, I32498)
--	g24854 = NAND(I32499, I32500)
--	I32509 = NAND(g17815, g24070)
--	I32510 = NAND(g17815, I32509)
--	I32511 = NAND(g24070, I32509)
--	g24857 = NAND(I32510, I32511)
--	I32518 = NAND(g18014, g24071)
--	I32519 = NAND(g18014, I32518)
--	I32520 = NAND(g24071, I32518)
--	g24860 = NAND(I32519, I32520)
--	I32526 = NAND(g18038, g24078)
--	I32527 = NAND(g18038, I32526)
--	I32528 = NAND(g24078, I32526)
--	g24862 = NAND(I32527, I32528)
--	g24863 = NAND(g24258, g23319)
--	I32538 = NAND(g18247, g24080)
--	I32539 = NAND(g18247, I32538)
--	I32540 = NAND(g24080, I32538)
--	g24866 = NAND(I32539, I32540)
--	I32546 = NAND(g17903, g23906)
--	I32547 = NAND(g17903, I32546)
--	I32548 = NAND(g23906, I32546)
--	g24868 = NAND(I32547, I32548)
--	I32559 = NAND(g17927, g24081)
--	I32560 = NAND(g17927, I32559)
--	I32561 = NAND(g24081, I32559)
--	g24873 = NAND(I32560, I32561)
--	I32567 = NAND(g18131, g24082)
--	I32568 = NAND(g18131, I32567)
--	I32569 = NAND(g24082, I32567)
--	g24875 = NAND(I32568, I32569)
--	I32575 = NAND(g18155, g24089)
--	I32576 = NAND(g18155, I32575)
--	I32577 = NAND(g24089, I32575)
--	g24877 = NAND(I32576, I32577)
--	I32586 = NAND(g17815, g23937)
--	I32587 = NAND(g17815, I32586)
--	I32588 = NAND(g23937, I32586)
--	g24880 = NAND(I32587, I32588)
--	I32595 = NAND(g18014, g23938)
--	I32596 = NAND(g18014, I32595)
--	I32597 = NAND(g23938, I32595)
--	g24883 = NAND(I32596, I32597)
--	I32607 = NAND(g18038, g24090)
--	I32608 = NAND(g18038, I32607)
--	I32609 = NAND(g24090, I32607)
--	g24887 = NAND(I32608, I32609)
--	I32615 = NAND(g18247, g24091)
--	I32616 = NAND(g18247, I32615)
--	I32617 = NAND(g24091, I32615)
--	g24889 = NAND(I32616, I32617)
--	I32624 = NAND(g17927, g23969)
--	I32625 = NAND(g17927, I32624)
--	I32626 = NAND(g23969, I32624)
--	g24897 = NAND(I32625, I32626)
--	I32633 = NAND(g18131, g23970)
--	I32634 = NAND(g18131, I32633)
--	I32635 = NAND(g23970, I32633)
--	g24900 = NAND(I32634, I32635)
--	I32645 = NAND(g18155, g24093)
--	I32646 = NAND(g18155, I32645)
--	I32647 = NAND(g24093, I32645)
--	g24904 = NAND(I32646, I32647)
--	I32659 = NAND(g18038, g23998)
--	I32660 = NAND(g18038, I32659)
--	I32661 = NAND(g23998, I32659)
--	g24920 = NAND(I32660, I32661)
--	I32668 = NAND(g18247, g23999)
--	I32669 = NAND(g18247, I32668)
--	I32670 = NAND(g23999, I32668)
--	g24923 = NAND(I32669, I32670)
--	I32677 = NAND(g23823, g14165)
--	I32678 = NAND(g23823, I32677)
--	I32679 = NAND(g14165, I32677)
--	g24928 = NAND(I32678, I32679)
--	I32686 = NAND(g18155, g24028)
--	I32687 = NAND(g18155, I32686)
--	I32688 = NAND(g24028, I32686)
--	g24937 = NAND(I32687, I32688)
--	I32695 = NAND(g23858, g14280)
--	I32696 = NAND(g23858, I32695)
--	I32697 = NAND(g14280, I32695)
--	g24940 = NAND(I32696, I32697)
--	I32708 = NAND(g23892, g14402)
--	I32709 = NAND(g23892, I32708)
--	I32710 = NAND(g14402, I32708)
--	g24951 = NAND(I32709, I32710)
--	I32724 = NAND(g23913, g14514)
--	I32725 = NAND(g23913, I32724)
--	I32726 = NAND(g14514, I32724)
--	g24963 = NAND(I32725, I32726)
--	g24975 = NAND(g23497, g74)
--	g24986 = NAND(g23513, g762)
--	g24997 = NAND(g23528, g1448)
--	g25004 = NAND(g23644, g6448)
--	g25005 = NAND(g23539, g2142)
--	g25008 = NAND(g23644, g5438)
--	g25009 = NAND(g23644, g6448)
--	g25010 = NAND(g23694, g6713)
--	g25011 = NAND(g23644, g5438)
--	g25012 = NAND(g23644, g6448)
--	g25013 = NAND(g23923, g6643)
--	g25014 = NAND(g23694, g5473)
--	g25015 = NAND(g23694, g6713)
--	g25016 = NAND(g23748, g7015)
--	g25017 = NAND(g23644, g5438)
--	g25018 = NAND(g23644, g6448)
--	g25019 = NAND(g23923, g6486)
--	g25020 = NAND(g23923, g6643)
--	g25021 = NAND(g23694, g5473)
--	g25022 = NAND(g23694, g6713)
--	g25023 = NAND(g23955, g6945)
--	g25024 = NAND(g23748, g5512)
--	g25025 = NAND(g23748, g7015)
--	g25026 = NAND(g23803, g7265)
--	g25028 = NAND(g23644, g5438)
--	g25029 = NAND(g23923, g6486)
--	g25030 = NAND(g23923, g6643)
--	g25031 = NAND(g23694, g5473)
--	g25032 = NAND(g23694, g6713)
--	g25033 = NAND(g23955, g6751)
--	g25034 = NAND(g23955, g6945)
--	g25035 = NAND(g23748, g5512)
--	g25036 = NAND(g23748, g7015)
--	g25037 = NAND(g23984, g7195)
--	g25038 = NAND(g23803, g5556)
--	g25039 = NAND(g23803, g7265)
--	g25040 = NAND(g23923, g6486)
--	g25041 = NAND(g23923, g6643)
--	g25043 = NAND(g23694, g5473)
--	g25044 = NAND(g23955, g6751)
--	g25045 = NAND(g23955, g6945)
--	g25046 = NAND(g23748, g5512)
--	g25047 = NAND(g23748, g7015)
--	g25048 = NAND(g23984, g7053)
--	g25049 = NAND(g23984, g7195)
--	g25050 = NAND(g23803, g5556)
--	g25051 = NAND(g23803, g7265)
--	g25052 = NAND(g24014, g7391)
--	g25053 = NAND(g23923, g6486)
--	g25054 = NAND(g23955, g6751)
--	g25055 = NAND(g23955, g6945)
--	g25057 = NAND(g23748, g5512)
--	g25058 = NAND(g23984, g7053)
--	g25059 = NAND(g23984, g7195)
--	g25060 = NAND(g23803, g5556)
--	g25061 = NAND(g23803, g7265)
--	g25062 = NAND(g24014, g7303)
--	g25063 = NAND(g24014, g7391)
--	g25064 = NAND(g23955, g6751)
--	g25065 = NAND(g23984, g7053)
--	g25066 = NAND(g23984, g7195)
--	g25068 = NAND(g23803, g5556)
--	g25069 = NAND(g24014, g7303)
--	g25070 = NAND(g24014, g7391)
--	g25071 = NAND(g23984, g7053)
--	g25072 = NAND(g24014, g7303)
--	g25073 = NAND(g24014, g7391)
--	g25074 = NAND(g24014, g7303)
--	g25088 = NAND(g23950, g679)
--	g25096 = NAND(g23979, g1365)
--	g25106 = NAND(g24009, g2059)
--	g25112 = NAND(g24043, g2753)
--	g25200 = NAND(g24965, g3306)
--	g25203 = NAND(g24978, g3462)
--	g25205 = NAND(g24989, g3618)
--	g25210 = NAND(g25000, g3774)
--	g25312 = NAND(g21211, g14442, g10694, g24590)
--	g25320 = NAND(g21219, g14529, g10714, g24595)
--	g25331 = NAND(g21230, g14584, g10735, g24603)
--	g25340 = NAND(g21235, g14618, g10754, g24610)
--	g25927 = NAND(g24965, g6448)
--	g25928 = NAND(g24965, g5438)
--	g25929 = NAND(g24978, g6713)
--	g25930 = NAND(g24978, g5473)
--	g25931 = NAND(g24989, g7015)
--	g25933 = NAND(g24989, g5512)
--	g25934 = NAND(g25000, g7265)
--	g25936 = NAND(g25000, g5556)
--	g25954 = NAND(g22806, g24517)
--	g25958 = NAND(g22847, g24530)
--	g25964 = NAND(g22882, g24543)
--	g25969 = NAND(g22917, g24555)
--	g26059 = NAND(g25422, g25379, g25274)
--	g26066 = NAND(g25431, g25395, g25283)
--	g26073 = NAND(g25438, g25405, g25291)
--	g26079 = NAND(g25445, g25413, g25301)
--	g26106 = NAND(g23644, g25354)
--	g26119 = NAND(g8278, g14657, g25422, g25379)
--	g26120 = NAND(g23694, g25369)
--	g26129 = NAND(g8287, g14691, g25431, g25395)
--	g26130 = NAND(g23748, g25386)
--	g26143 = NAND(g8296, g14725, g25438, g25405)
--	g26144 = NAND(g23803, g25402)
--	g26148 = NAND(g8305, g14753, g25445, g25413)
--	g26356 = NAND(g16539, g25183)
--	g26399 = NAND(g16571, g25186)
--	g26440 = NAND(g16595, g25190)
--	g26458 = NAND(g25343, g65)
--	g26472 = NAND(g16615, g25195)
--	g26482 = NAND(g25357, g753)
--	g26498 = NAND(g25372, g1439)
--	g26513 = NAND(g25389, g2133)
--	g26772 = NAND(g26320, g3306)
--	g26779 = NAND(g26367, g3462)
--	g26785 = NAND(g26410, g3618)
--	g26792 = NAND(g26451, g3774)
--	I35020 = NAND(g26110, g26099)
--	I35021 = NAND(g26110, I35020)
--	I35022 = NAND(g26099, I35020)
--	g26859 = NAND(I35021, I35022)
--	I35034 = NAND(g26087, g26154)
--	I35035 = NAND(g26087, I35034)
--	I35036 = NAND(g26154, I35034)
--	g26865 = NAND(I35035, I35036)
--	I35042 = NAND(g26151, g26145)
--	I35043 = NAND(g26151, I35042)
--	I35044 = NAND(g26145, I35042)
--	g26867 = NAND(I35043, I35044)
--	I35057 = NAND(g26137, g26126)
--	I35058 = NAND(g26137, I35057)
--	I35059 = NAND(g26126, I35057)
--	g26874 = NAND(I35058, I35059)
--	g26892 = NAND(g25699, g26283, g25569, g25631)
--	g26902 = NAND(g25631, g26283, g25569)
--	g26906 = NAND(g25772, g26327, g25648, g25708)
--	g26911 = NAND(g25569, g26283)
--	g26915 = NAND(g25708, g26327, g25648)
--	g26918 = NAND(g25826, g26374, g25725, g25781)
--	g26925 = NAND(g25648, g26327)
--	g26928 = NAND(g25781, g26374, g25725)
--	g26931 = NAND(g25861, g26417, g25798, g25835)
--	I35123 = NAND(g26107, g26096)
--	I35124 = NAND(g26107, I35123)
--	I35125 = NAND(g26096, I35123)
--	g26934 = NAND(I35124, I35125)
--	g26938 = NAND(g25725, g26374)
--	g26941 = NAND(g25835, g26417, g25798)
--	g26947 = NAND(g25798, g26417)
--	g27117 = NAND(g26320, g6448)
--	g27118 = NAND(g26320, g5438)
--	g27119 = NAND(g26367, g6713)
--	g27121 = NAND(g26367, g5473)
--	g27122 = NAND(g26410, g7015)
--	g27124 = NAND(g26410, g5512)
--	g27125 = NAND(g26451, g7265)
--	g27130 = NAND(g26451, g5556)
--	I35701 = NAND(g26867, g26874)
--	I35702 = NAND(g26867, I35701)
--	I35703 = NAND(g26874, I35701)
--	g27379 = NAND(I35702, I35703)
--	I35714 = NAND(g26859, g26865)
--	I35715 = NAND(g26859, I35714)
--	I35716 = NAND(g26865, I35714)
--	g27382 = NAND(I35715, I35716)
--	g27390 = NAND(g26989, g6448)
--	g27395 = NAND(g26989, g5438)
--	g27400 = NAND(g27012, g6713)
--	g27408 = NAND(g27012, g5473)
--	g27413 = NAND(g27038, g7015)
--	g27426 = NAND(g27038, g5512)
--	g27431 = NAND(g27066, g7265)
--	g27447 = NAND(g27066, g5556)
--	I35904 = NAND(g27051, g14831)
--	I35905 = NAND(g27051, I35904)
--	I35906 = NAND(g14831, I35904)
--	g27528 = NAND(I35905, I35906)
--	I35944 = NAND(g27078, g14904)
--	I35945 = NAND(g27078, I35944)
--	I35946 = NAND(g14904, I35944)
--	g27550 = NAND(I35945, I35946)
--	I35974 = NAND(g27094, g14985)
--	I35975 = NAND(g27094, I35974)
--	I35976 = NAND(g14985, I35974)
--	g27566 = NAND(I35975, I35976)
--	g27571 = NAND(g26869, g56)
--	I35992 = NAND(g27106, g15074)
--	I35993 = NAND(g27106, I35992)
--	I35994 = NAND(g15074, I35992)
--	g27576 = NAND(I35993, I35994)
--	g27580 = NAND(g26878, g744)
--	g27583 = NAND(g26887, g1430)
--	g27587 = NAND(g26897, g2124)
--	g27626 = NAND(g26989, g3306)
--	g27627 = NAND(g27012, g3462)
--	g27628 = NAND(g27038, g3618)
--	g27630 = NAND(g27066, g3774)
--	g27738 = NAND(g25367, g27415)
--	g27743 = NAND(g25384, g27436)
--	g27751 = NAND(g25400, g27455)
--	g27756 = NAND(g25410, g27471)
--	I36256 = NAND(g27527, g15859)
--	I36257 = NAND(g27527, I36256)
--	I36258 = NAND(g15859, I36256)
--	g27801 = NAND(I36257, I36258)
--	I36270 = NAND(g27549, g15890)
--	I36271 = NAND(g27549, I36270)
--	I36272 = NAND(g15890, I36270)
--	g27809 = NAND(I36271, I36272)
--	I36289 = NAND(g27565, g15923)
--	I36290 = NAND(g27565, I36289)
--	I36291 = NAND(g15923, I36289)
--	g27830 = NAND(I36290, I36291)
--	I36300 = NAND(g27382, g27379)
--	I36301 = NAND(g27382, I36300)
--	I36302 = NAND(g27379, I36300)
--	g27838 = NAND(I36301, I36302)
--	I36314 = NAND(g27575, g15952)
--	I36315 = NAND(g27575, I36314)
--	I36316 = NAND(g15952, I36314)
--	g27846 = NAND(I36315, I36316)
--	I36591 = NAND(g27529, g14885)
--	I36592 = NAND(g27529, I36591)
--	I36593 = NAND(g14885, I36591)
--	g28046 = NAND(I36592, I36593)
--	I36666 = NAND(g27551, g14966)
--	I36667 = NAND(g27551, I36666)
--	I36668 = NAND(g14966, I36666)
--	g28075 = NAND(I36667, I36668)
--	I36731 = NAND(g27567, g15055)
--	I36732 = NAND(g27567, I36731)
--	I36733 = NAND(g15055, I36731)
--	g28100 = NAND(I36732, I36733)
--	I36779 = NAND(g27577, g15151)
--	I36780 = NAND(g27577, I36779)
--	I36781 = NAND(g15151, I36779)
--	g28118 = NAND(I36780, I36781)
--	I37295 = NAND(g27827, g27814)
--	I37296 = NAND(g27827, I37295)
--	I37297 = NAND(g27814, I37295)
--	g28384 = NAND(I37296, I37297)
--	I37303 = NAND(g27802, g27900)
--	I37304 = NAND(g27802, I37303)
--	I37305 = NAND(g27900, I37303)
--	g28386 = NAND(I37304, I37305)
--	I37311 = NAND(g27897, g27883)
--	I37312 = NAND(g27897, I37311)
--	I37313 = NAND(g27883, I37311)
--	g28388 = NAND(I37312, I37313)
--	I37322 = NAND(g27865, g27855)
--	I37323 = NAND(g27865, I37322)
--	I37324 = NAND(g27855, I37322)
--	g28391 = NAND(I37323, I37324)
--	I37356 = NAND(g27824, g27811)
--	I37357 = NAND(g27824, I37356)
--	I37358 = NAND(g27811, I37356)
--	g28415 = NAND(I37357, I37358)
--	I37813 = NAND(g28388, g28391)
--	I37814 = NAND(g28388, I37813)
--	I37815 = NAND(g28391, I37813)
--	g28842 = NAND(I37814, I37815)
--	I37822 = NAND(g28384, g28386)
--	I37823 = NAND(g28384, I37822)
--	I37824 = NAND(g28386, I37822)
--	g28845 = NAND(I37823, I37824)
--	g28978 = NAND(g9150, g28512)
--	g29001 = NAND(g9161, g28512)
--	g29008 = NAND(g9174, g28540)
--	g29026 = NAND(g9187, g28512)
--	g29030 = NAND(g9203, g28540)
--	g29038 = NAND(g9216, g28567)
--	g29045 = NAND(g9232, g28512)
--	g29049 = NAND(g9248, g28540)
--	g29053 = NAND(g9264, g28567)
--	g29060 = NAND(g9277, g28595)
--	g29062 = NAND(g9310, g28540)
--	g29068 = NAND(g9326, g28567)
--	g29072 = NAND(g9342, g28595)
--	g29076 = NAND(g9391, g28567)
--	g29080 = NAND(g9407, g28595)
--	g29087 = NAND(g9488, g28595)
--	g29088 = NAND(g9507, g28512)
--	g29096 = NAND(g9649, g28540)
--	g29103 = NAND(g9795, g28567)
--	g29107 = NAND(g9941, g28595)
--	I38378 = NAND(g28845, g28842)
--	I38379 = NAND(g28845, I38378)
--	I38380 = NAND(g28842, I38378)
--	g29265 = NAND(I38379, I38380)
--	I38810 = NAND(g29303, g15904)
--	I38811 = NAND(g29303, I38810)
--	I38812 = NAND(g15904, I38810)
--	g29498 = NAND(I38811, I38812)
--	I38820 = NAND(g29313, g15933)
--	I38821 = NAND(g29313, I38820)
--	I38822 = NAND(g15933, I38820)
--	g29500 = NAND(I38821, I38822)
--	I38831 = NAND(g29324, g15962)
--	I38832 = NAND(g29324, I38831)
--	I38833 = NAND(g15962, I38831)
--	g29503 = NAND(I38832, I38833)
--	I38841 = NAND(g29333, g15981)
--	I38842 = NAND(g29333, I38841)
--	I38843 = NAND(g15981, I38841)
--	g29505 = NAND(I38842, I38843)
--	I39323 = NAND(g29721, g29713)
--	I39324 = NAND(g29721, I39323)
--	I39325 = NAND(g29713, I39323)
--	g29911 = NAND(I39324, I39325)
--	I39331 = NAND(g29705, g29751)
--	I39332 = NAND(g29705, I39331)
--	I39333 = NAND(g29751, I39331)
--	g29913 = NAND(I39332, I39333)
--	I39339 = NAND(g29748, g29741)
--	I39340 = NAND(g29748, I39339)
--	I39341 = NAND(g29741, I39339)
--	g29915 = NAND(I39340, I39341)
--	I39347 = NAND(g29732, g29728)
--	I39348 = NAND(g29732, I39347)
--	I39349 = NAND(g29728, I39347)
--	g29917 = NAND(I39348, I39349)
--	I39359 = NAND(g29766, g15880)
--	I39360 = NAND(g29766, I39359)
--	I39361 = NAND(g15880, I39359)
--	g29923 = NAND(I39360, I39361)
--	I39367 = NAND(g29767, g15913)
--	I39368 = NAND(g29767, I39367)
--	I39369 = NAND(g15913, I39367)
--	g29925 = NAND(I39368, I39369)
--	I39375 = NAND(g29768, g15942)
--	I39376 = NAND(g29768, I39375)
--	I39377 = NAND(g15942, I39375)
--	g29927 = NAND(I39376, I39377)
--	I39384 = NAND(g29718, g29710)
--	I39385 = NAND(g29718, I39384)
--	I39386 = NAND(g29710, I39384)
--	g29930 = NAND(I39385, I39386)
--	I39391 = NAND(g29769, g15971)
--	I39392 = NAND(g29769, I39391)
--	I39393 = NAND(g15971, I39391)
--	g29931 = NAND(I39392, I39393)
--	I39532 = NAND(g29915, g29917)
--	I39533 = NAND(g29915, I39532)
--	I39534 = NAND(g29917, I39532)
--	g30034 = NAND(I39533, I39534)
--	I39539 = NAND(g29911, g29913)
--	I39540 = NAND(g29911, I39539)
--	I39541 = NAND(g29913, I39539)
--	g30035 = NAND(I39540, I39541)
--	I39689 = NAND(g30035, g30034)
--	I39690 = NAND(g30035, I39689)
--	I39691 = NAND(g30034, I39689)
--	g30228 = NAND(I39690, I39691)
--	I40558 = NAND(g30605, g30597)
--	I40559 = NAND(g30605, I40558)
--	I40560 = NAND(g30597, I40558)
--	g30768 = NAND(I40559, I40560)
--	I40571 = NAND(g30588, g30632)
--	I40572 = NAND(g30588, I40571)
--	I40573 = NAND(g30632, I40571)
--	g30771 = NAND(I40572, I40573)
--	I40587 = NAND(g30629, g30622)
--	I40588 = NAND(g30629, I40587)
--	I40589 = NAND(g30622, I40587)
--	g30775 = NAND(I40588, I40589)
--	I40603 = NAND(g30614, g30610)
--	I40604 = NAND(g30614, I40603)
--	I40605 = NAND(g30610, I40603)
--	g30779 = NAND(I40604, I40605)
--	I40627 = NAND(g30602, g30594)
--	I40628 = NAND(g30602, I40627)
--	I40629 = NAND(g30594, I40627)
--	g30791 = NAND(I40628, I40629)
--	I41010 = NAND(g30775, g30779)
--	I41011 = NAND(g30775, I41010)
--	I41012 = NAND(g30779, I41010)
--	g30926 = NAND(I41011, I41012)
--	I41017 = NAND(g30768, g30771)
--	I41018 = NAND(g30768, I41017)
--	I41019 = NAND(g30771, I41017)
--	g30927 = NAND(I41018, I41019)
--	I41064 = NAND(g30927, g30926)
--	I41065 = NAND(g30927, I41064)
--	I41066 = NAND(g30926, I41064)
--	g30952 = NAND(I41065, I41066)
--	
--	g7528 = NOR(g3151, g3142, g3147)
--	g7575 = NOR(g2984, g2985)
--	g7795 = NOR(g2992, g2991)
--	g8430 = NOR(g3198, g8120, g3194, g3191)
--	g10784 = NOR(g5630, g5649, g5676)
--	g10789 = NOR(g5650, g5677, g5709)
--	g10793 = NOR(g5658, g5687, g5728)
--	g10797 = NOR(g5678, g5710, g5757)
--	g10801 = NOR(g5688, g5729, g5767)
--	g10805 = NOR(g5696, g5739, g5786)
--	g10810 = NOR(g5711, g5758, g5807)
--	g10814 = NOR(g5730, g5768, g5816)
--	g10818 = NOR(g5740, g5787, g5826)
--	g10822 = NOR(g5748, g5797, g5845)
--	g10831 = NOR(g5769, g5817, g5863)
--	g10835 = NOR(g5788, g5827, g5872)
--	g10839 = NOR(g5798, g5846, g5882)
--	g10851 = NOR(g5828, g5873, g5910)
--	g10855 = NOR(g5847, g5883, g5919)
--	g10872 = NOR(g5884, g5920, g5949)
--	g11600 = NOR(g9049, g9064, g9078)
--	g11622 = NOR(g8183, g11332, g7928, g11069)
--	g11624 = NOR(g9062, g9075, g9091)
--	g11627 = NOR(g9063, g9077, g9093)
--	g11630 = NOR(g9066, g9081, g9097)
--	g11643 = NOR(g11481, g8045, g7928, g11069)
--	g11644 = NOR(g9076, g9092, g9102)
--	g11647 = NOR(g9079, g9094, g9103)
--	g11650 = NOR(g9080, g9096, g9105)
--	g11653 = NOR(g9083, g9100, g9109)
--	g11660 = NOR(g8183, g8045, g7928, g11069)
--	g11663 = NOR(g9095, g9104, g9112)
--	g11666 = NOR(g9098, g9106, g9113)
--	g11669 = NOR(g9099, g9108, g9115)
--	g11675 = NOR(g9107, g9114, g9120)
--	g11678 = NOR(g9110, g9116, g9121)
--	g11681 = NOR(g9111, g9118, g9123)
--	g11687 = NOR(g9117, g9122, g9126)
--	g11690 = NOR(g9119, g9124, g9127)
--	g11697 = NOR(g9125, g9131, g9133)
--	g11703 = NOR(g9132, g9137, g9139)
--	g11711 = NOR(g9138, g9143, g9145)
--	g11744 = NOR(g9241, g9301, g9364)
--	g11759 = NOR(g9302, g9365, g9438)
--	g11760 = NOR(g9319, g9382, g9461)
--	g11767 = NOR(g9366, g9439, g9518)
--	g11768 = NOR(g9367, g9441, g9521)
--	g11772 = NOR(g9383, g9462, g9580)
--	g11773 = NOR(g9400, g9479, g9603)
--	g11780 = NOR(g9440, g9519, g9630)
--	g11781 = NOR(g9442, g9522, g9633)
--	g11784 = NOR(g9463, g9581, g9660)
--	g11785 = NOR(g9464, g9583, g9663)
--	g11789 = NOR(g9480, g9604, g9722)
--	g11790 = NOR(g9497, g9621, g9745)
--	g11799 = NOR(g9520, g9631, g9759)
--	g11800 = NOR(g9523, g9634, g9762)
--	g11806 = NOR(g9582, g9661, g9776)
--	g11807 = NOR(g9584, g9664, g9779)
--	g11810 = NOR(g9605, g9723, g9806)
--	g11811 = NOR(g9606, g9725, g9809)
--	g11815 = NOR(g9622, g9746, g9868)
--	g11822 = NOR(g9632, g9760, g9888)
--	g11823 = NOR(g9635, g9763, g9891)
--	g11828 = NOR(g9639, g9764, g9892)
--	g11830 = NOR(g9647, g9773, g9901)
--	g11831 = NOR(g9648, g9775, g9904)
--	g11832 = NOR(g9662, g9777, g9905)
--	g11833 = NOR(g9665, g9780, g9908)
--	g11839 = NOR(g9724, g9807, g9922)
--	g11840 = NOR(g9726, g9810, g9925)
--	g11843 = NOR(g9747, g9869, g9952)
--	g11844 = NOR(g9748, g9871, g9955)
--	g11855 = NOR(g9761, g9889, g10009)
--	g11860 = NOR(g9765, g9893, g10012)
--	g11861 = NOR(g9766, g9894, g10013)
--	g11863 = NOR(g9774, g9902, g10035)
--	g11864 = NOR(g9778, g9906, g10042)
--	g11865 = NOR(g9781, g9909, g10045)
--	g11870 = NOR(g9785, g9910, g10046)
--	g11872 = NOR(g9793, g9919, g10055)
--	g11873 = NOR(g9794, g9921, g10058)
--	g11874 = NOR(g9808, g9923, g10059)
--	g11875 = NOR(g9811, g9926, g10062)
--	g11881 = NOR(g9870, g9953, g10076)
--	g11882 = NOR(g9872, g9956, g10079)
--	g11889 = NOR(g9887, g10007, g10101)
--	g11890 = NOR(g9890, g10010, g10103)
--	g11896 = NOR(g9903, g10036, g10112)
--	g11897 = NOR(g9907, g10043, g10118)
--	g11902 = NOR(g9911, g10047, g10121)
--	g11903 = NOR(g9912, g10048, g10122)
--	g11905 = NOR(g9920, g10056, g10144)
--	g11906 = NOR(g9924, g10060, g10151)
--	g11907 = NOR(g9927, g10063, g10154)
--	g11912 = NOR(g9931, g10064, g10155)
--	g11914 = NOR(g9939, g10073, g10164)
--	g11915 = NOR(g9940, g10075, g10167)
--	g11916 = NOR(g9954, g10077, g10168)
--	g11917 = NOR(g9957, g10080, g10171)
--	g11928 = NOR(g10008, g10102, g10192)
--	g11934 = NOR(g10011, g10104, g10193)
--	g11935 = NOR(g10014, g10106, g10196)
--	g11938 = NOR(g10037, g10113, g10201)
--	g11939 = NOR(g10041, g10116, g10206)
--	g11940 = NOR(g10044, g10119, g10208)
--	g11946 = NOR(g10057, g10145, g10217)
--	g11947 = NOR(g10061, g10152, g10223)
--	g11952 = NOR(g10065, g10156, g10226)
--	g11953 = NOR(g10066, g10157, g10227)
--	g11955 = NOR(g10074, g10165, g10249)
--	g11956 = NOR(g10078, g10169, g10256)
--	g11957 = NOR(g10081, g10172, g10259)
--	g11962 = NOR(g10085, g10173, g10260)
--	g11964 = NOR(g10093, g10182, g10269)
--	g11965 = NOR(g10094, g10184, g10272)
--	g11974 = NOR(g10105, g10194, g10279)
--	g11975 = NOR(g10107, g10197, g10282)
--	g11979 = NOR(g10114, g10202, g10288)
--	g11980 = NOR(g10115, g10204, g10291)
--	g11981 = NOR(g10117, g10207, g10294)
--	g11987 = NOR(g10120, g10209, g10295)
--	g11988 = NOR(g10123, g10211, g10298)
--	g11991 = NOR(g10146, g10218, g10303)
--	g11992 = NOR(g10150, g10221, g10308)
--	g11993 = NOR(g10153, g10224, g10310)
--	g11999 = NOR(g10166, g10250, g10319)
--	g12000 = NOR(g10170, g10257, g10325)
--	g12005 = NOR(g10174, g10261, g10328)
--	g12006 = NOR(g10175, g10262, g10329)
--	g12008 = NOR(g10183, g10270, g10351)
--	g12026 = NOR(g10195, g10280, g10360)
--	g12033 = NOR(g10199, g10284, g10362)
--	g12034 = NOR(g10200, g10286, g10365)
--	g12035 = NOR(g10203, g10289, g10367)
--	g12036 = NOR(g10205, g10292, g10370)
--	g12043 = NOR(g10210, g10296, g10372)
--	g12044 = NOR(g10212, g10299, g10375)
--	g12048 = NOR(g10219, g10304, g10381)
--	g12049 = NOR(g10220, g10306, g10384)
--	g12050 = NOR(g10222, g10309, g10387)
--	g12056 = NOR(g10225, g10311, g10388)
--	g12057 = NOR(g10228, g10313, g10391)
--	g12060 = NOR(g10251, g10320, g10396)
--	g12061 = NOR(g10255, g10323, g10401)
--	g12062 = NOR(g10258, g10326, g10403)
--	g12068 = NOR(g10271, g10352, g10412)
--	g12079 = NOR(g10281, g10361, g10422)
--	g12080 = NOR(g10285, g10363, g10430)
--	g12081 = NOR(g10287, g10366, g10433)
--	g12082 = NOR(g10290, g10368, g10435)
--	g12083 = NOR(g10293, g10371, g10438)
--	g12090 = NOR(g10297, g10373, g10439)
--	g12097 = NOR(g10301, g10377, g10441)
--	g12098 = NOR(g10302, g10379, g10444)
--	g12099 = NOR(g10305, g10382, g10446)
--	g12100 = NOR(g10307, g10385, g10449)
--	g12107 = NOR(g10312, g10389, g10451)
--	g12108 = NOR(g10314, g10392, g10454)
--	g12112 = NOR(g10321, g10397, g10460)
--	g12113 = NOR(g10322, g10399, g10463)
--	g12114 = NOR(g10324, g10402, g10466)
--	g12120 = NOR(g10327, g10404, g10467)
--	g12121 = NOR(g10330, g10406, g10470)
--	g12124 = NOR(g10353, g10413, g10475)
--	g12145 = NOR(g10364, g10431, g10492)
--	g12146 = NOR(g10369, g10436, g10496)
--	g12151 = NOR(g10374, g10440, g10498)
--	g12152 = NOR(g10378, g10442, g10506)
--	g12153 = NOR(g10380, g10445, g10509)
--	g12154 = NOR(g10383, g10447, g10511)
--	g12155 = NOR(g10386, g10450, g10514)
--	g12162 = NOR(g10390, g10452, g10515)
--	g12169 = NOR(g10394, g10456, g10517)
--	g12170 = NOR(g10395, g10458, g10520)
--	g12171 = NOR(g10398, g10461, g10522)
--	g12172 = NOR(g10400, g10464, g10525)
--	g12179 = NOR(g10405, g10468, g10527)
--	g12180 = NOR(g10407, g10471, g10530)
--	g12184 = NOR(g10414, g10476, g10536)
--	g12185 = NOR(g10415, g10478, g10539)
--	g12192 = NOR(g10423, g10485, g10548)
--	g12193 = NOR(g10432, g10493, g10555)
--	g12194 = NOR(g10434, g10494, g10556)
--	g12195 = NOR(g10437, g10497, g10558)
--	g12207 = NOR(g10443, g10507, g10566)
--	g12208 = NOR(g10448, g10512, g10570)
--	g12213 = NOR(g10453, g10516, g10572)
--	g12214 = NOR(g10457, g10518, g10580)
--	g12215 = NOR(g10459, g10521, g10583)
--	g12216 = NOR(g10462, g10523, g10585)
--	g12217 = NOR(g10465, g10526, g10588)
--	g12224 = NOR(g10469, g10528, g10589)
--	g12231 = NOR(g10473, g10532, g10591)
--	g12232 = NOR(g10474, g10534, g10594)
--	g12233 = NOR(g10477, g10537, g10596)
--	g12234 = NOR(g10479, g10540, g10599)
--	g12245 = NOR(g10495, g10557, g10604)
--	g12247 = NOR(g10499, g10559, g10605)
--	g12248 = NOR(g10508, g10567, g10612)
--	g12249 = NOR(g10510, g10568, g10613)
--	g12250 = NOR(g10513, g10571, g10615)
--	g12262 = NOR(g10519, g10581, g10623)
--	g12263 = NOR(g10524, g10586, g10627)
--	g12268 = NOR(g10529, g10590, g10629)
--	g12269 = NOR(g10533, g10592, g10637)
--	g12270 = NOR(g10535, g10595, g10640)
--	g12271 = NOR(g10538, g10597, g10642)
--	g12272 = NOR(g10541, g10600, g10645)
--	g12288 = NOR(g10569, g10614, g10651)
--	g12290 = NOR(g10573, g10616, g10652)
--	g12291 = NOR(g10582, g10624, g10659)
--	g12292 = NOR(g10584, g10625, g10660)
--	g12293 = NOR(g10587, g10628, g10662)
--	g12305 = NOR(g10593, g10638, g10670)
--	g12306 = NOR(g10598, g10643, g10674)
--	g12324 = NOR(g10626, g10661, g10681)
--	g12326 = NOR(g10630, g10663, g10682)
--	g12327 = NOR(g10639, g10671, g10689)
--	g12328 = NOR(g10641, g10672, g10690)
--	g12329 = NOR(g10644, g10675, g10692)
--	g12339 = NOR(g10650, g10678, g10704)
--	g12352 = NOR(g10673, g10691, g10710)
--	g12369 = NOR(g10680, g10707, g10724)
--	g12388 = NOR(g10709, g10727, g10745)
--	g12418 = NOR(g10729, g10748, g10764)
--	g12431 = NOR(g8580, g10730)
--	g12436 = NOR(g8587, g10749)
--	g12441 = NOR(g8594, g10767)
--	g12446 = NOR(g8605, g10773)
--	g12451 = NOR(g499, g8983)
--	g12457 = NOR(g9009, g9033, g9048)
--	g12467 = NOR(g9034, g9056, g9065)
--	g12482 = NOR(g9057, g9073, g9082)
--	g12487 = NOR(g10108, g10198, g10283)
--	g12499 = NOR(g9074, g9090, g9101)
--	g12507 = NOR(g10213, g10300, g10376)
--	g12524 = NOR(g10315, g10393, g10455)
--	g12539 = NOR(g10408, g10472, g10531)
--	g12698 = NOR(g11347, g11420, g8327)
--	g12747 = NOR(g11421, g8328, g8385)
--	g12755 = NOR(g11431, g8339, g8394)
--	g12780 = NOR(g9187, g9161)
--	g12781 = NOR(g8329, g8386, g8431)
--	g12789 = NOR(g8340, g8395, g8437)
--	g12797 = NOR(g8350, g8406, g8446)
--	g12814 = NOR(g8387, g8432, g8463)
--	g12819 = NOR(g9248, g9203)
--	g12820 = NOR(g8396, g8438, g8466)
--	g12828 = NOR(g8407, g8447, g8472)
--	g12836 = NOR(g8417, g8458, g8481)
--	g12849 = NOR(g8433, g8464, g8485)
--	g12852 = NOR(g8439, g8467, g8488)
--	g12857 = NOR(g9326, g9264)
--	g12858 = NOR(g8448, g8473, g8491)
--	g12866 = NOR(g8459, g8482, g8497)
--	g12880 = NOR(g8465, g8486, g8502)
--	g12883 = NOR(g10038, g6284)
--	g12890 = NOR(g8468, g8489, g8505)
--	g12893 = NOR(g8474, g8492, g8508)
--	g12898 = NOR(g9407, g9342)
--	g12899 = NOR(g8483, g8498, g8511)
--	g12912 = NOR(g8484, g8500, g8515)
--	g12913 = NOR(g8487, g8503, g8518)
--	g12920 = NOR(g8490, g8506, g8521)
--	g12923 = NOR(g10147, g6421)
--	g12930 = NOR(g8493, g8509, g8524)
--	g12933 = NOR(g8499, g8512, g8527)
--	g12939 = NOR(g8501, g8516, g8531)
--	g12941 = NOR(g8504, g8519, g8534)
--	g12942 = NOR(g8507, g8522, g8537)
--	g12949 = NOR(g8510, g8525, g8540)
--	g12952 = NOR(g10252, g6626)
--	g12959 = NOR(g8513, g8528, g8543)
--	g12967 = NOR(g8517, g8532, g8546)
--	g12968 = NOR(g8520, g8535, g8548)
--	g12970 = NOR(g8523, g8538, g8551)
--	g12971 = NOR(g8526, g8541, g8554)
--	g12978 = NOR(g8529, g8544, g8557)
--	g12981 = NOR(g10354, g6890)
--	g12991 = NOR(g8536, g8549, g8559)
--	g12992 = NOR(g8539, g8552, g8561)
--	g12994 = NOR(g8542, g8555, g8564)
--	g12995 = NOR(g8545, g8558, g8567)
--	g13001 = NOR(g8553, g8562, g8570)
--	g13002 = NOR(g8556, g8565, g8572)
--	g13022 = NOR(g8566, g8573, g8576)
--	g13024 = NOR(g11481, g8045, g7928, g7880)
--	g13111 = NOR(g8601, g8612, g8621)
--	g13124 = NOR(g8613, g8625, g8631)
--	g13135 = NOR(g8626, g8635, g8650)
--	g13143 = NOR(g8636, g8654, g8666)
--	g13149 = NOR(g8676, g8687, g8703)
--	g13155 = NOR(g8688, g8705, g8722)
--	g13160 = NOR(g8704, g8717, g8751)
--	g13164 = NOR(g8706, g8724, g8760)
--	g13171 = NOR(g8723, g8755, g8774)
--	g13175 = NOR(g8725, g8762, g8783)
--	g13182 = NOR(g8761, g8778, g8797)
--	g13194 = NOR(g8784, g8801, g8816)
--	g13228 = NOR(g8841, g8861, g8892)
--	g13251 = NOR(g8868, g8899, g8932)
--	g13274 = NOR(g8906, g8939, g8972)
--	g13286 = NOR(g11481, g11332, g11190, g7880)
--	g13299 = NOR(g8946, g8979, g9004)
--	g13310 = NOR(g11481, g11332, g11190, g11069)
--	g13313 = NOR(g8183, g11332, g11190, g7880)
--	g13331 = NOR(g8183, g11332, g11190, g11069)
--	g13332 = NOR(g11481, g8045, g11190, g7880)
--	g13353 = NOR(g11481, g8045, g11190, g11069)
--	g13354 = NOR(g8183, g8045, g11190, g7880)
--	g13374 = NOR(g8183, g8045, g11190, g11069)
--	g13375 = NOR(g11481, g11332, g7928, g7880)
--	g13378 = NOR(g9026, g9047, g9061)
--	g13401 = NOR(g11481, g11332, g7928, g11069)
--	g13404 = NOR(g8183, g11332, g7928, g7880)
--	g15661 = NOR(g11737, g7345)
--	g15797 = NOR(g13305, g7143)
--	g15873 = NOR(g11617, g7562)
--	g15959 = NOR(g2814, g13082)
--	g15978 = NOR(g11737, g7152)
--	g16020 = NOR(g6200, g12457, g10952)
--	g16036 = NOR(g6289, g12467, g10952)
--	g16058 = NOR(g6426, g12482, g10952)
--	g16082 = NOR(g10952, g6140, g12487)
--	g16094 = NOR(g6631, g12499, g10952)
--	g16120 = NOR(g10952, g6161, g12507)
--	g16171 = NOR(g10952, g6188, g12524)
--	g16230 = NOR(g10952, g6220, g12539)
--	g16498 = NOR(g14158, g14347)
--	g16520 = NOR(g14273, g14459)
--	g16551 = NOR(g14395, g14546)
--	g16567 = NOR(g15904, g15880, g15859)
--	g16570 = NOR(g15904, g15880, g14630)
--	g16583 = NOR(g14507, g14601)
--	g16591 = NOR(g15933, g15913, g15890)
--	g16594 = NOR(g15933, g15913, g14650)
--	g16611 = NOR(g15962, g15942, g15923)
--	g16614 = NOR(g15962, g15942, g14677)
--	g16629 = NOR(g15981, g15971, g15952)
--	g16632 = NOR(g15981, g15971, g14711)
--	g16643 = NOR(g15904, g14642, g15859)
--	g16654 = NOR(g14690, g12477)
--	g16655 = NOR(g15933, g14669, g15890)
--	g16671 = NOR(g14724, g12494)
--	g16672 = NOR(g15962, g14703, g15923)
--	g16679 = NOR(g14797, g14895)
--	g16692 = NOR(g14752, g12514)
--	g16693 = NOR(g15981, g14737, g15952)
--	g16705 = NOR(g14849, g14976)
--	g16718 = NOR(g14773, g12531)
--	g16736 = NOR(g14922, g15065)
--	g16778 = NOR(g15003, g15161)
--	g16802 = NOR(g13469, g3897)
--	g16803 = NOR(g15593, g12908)
--	g16823 = NOR(g5362, g13469)
--	g16824 = NOR(g15658, g12938)
--	g16829 = NOR(g14956, g12564)
--	g16835 = NOR(g15717, g12966)
--	g16841 = NOR(g15021, g12607)
--	g16844 = NOR(g15754, g12989)
--	g16845 = NOR(g15755, g12990)
--	g16847 = NOR(g15095, g12650)
--	g16851 = NOR(g15781, g13000)
--	g16853 = NOR(g15801, g13009)
--	g16854 = NOR(g15802, g13010)
--	g16857 = NOR(g15817, g13023)
--	g16860 = NOR(g15828, g13031)
--	g16861 = NOR(g15829, g13032)
--	g16866 = NOR(g15840, g13042)
--	g16880 = NOR(g15852, g13056)
--	g17012 = NOR(g14657, g14642, g15859)
--	g17025 = NOR(g15904, g15880, g15859)
--	g17042 = NOR(g14691, g14669, g15890)
--	g17051 = NOR(g14657, g15880, g14630)
--	g17059 = NOR(g15933, g15913, g15890)
--	g17076 = NOR(g14725, g14703, g15923)
--	g17086 = NOR(g14691, g15913, g14650)
--	g17094 = NOR(g15962, g15942, g15923)
--	g17111 = NOR(g14753, g14737, g15952)
--	g17124 = NOR(g14725, g15942, g14677)
--	g17132 = NOR(g15981, g15971, g15952)
--	g17151 = NOR(g14753, g15971, g14711)
--	g17186 = NOR(g7949, g14144)
--	g17197 = NOR(g8000, g14259)
--	g17204 = NOR(g8075, g14381)
--	g17209 = NOR(g8160, g14493)
--	g17213 = NOR(g4326, g14442)
--	g17215 = NOR(g15904, g14642)
--	g17216 = NOR(g4495, g14529)
--	g17218 = NOR(g15933, g14669)
--	g17219 = NOR(g4671, g14584)
--	g17220 = NOR(g15962, g14703)
--	g17221 = NOR(g4848, g14618)
--	g17222 = NOR(g15998, g16003)
--	g17223 = NOR(g15981, g14737)
--	g17224 = NOR(g16004, g16009)
--	g17225 = NOR(g16008, g16015)
--	g17226 = NOR(g16010, g16017)
--	g17228 = NOR(g16016, g16029)
--	g17229 = NOR(g16019, g16032)
--	g17234 = NOR(g16028, g16045)
--	g17235 = NOR(g16030, g16047)
--	g17236 = NOR(g16033, g16051)
--	g17246 = NOR(g16046, g16066)
--	g17247 = NOR(g16050, g16070)
--	g17248 = NOR(g16052, g16072)
--	g17269 = NOR(g16067, g16100)
--	g17270 = NOR(g16071, g16104)
--	g17271 = NOR(g16073, g16106)
--	g17302 = NOR(g16103, g16135)
--	g17303 = NOR(g16105, g16137)
--	g17340 = NOR(g16136, g16183)
--	g17341 = NOR(g16138, g16185)
--	g17383 = NOR(g16184, g16238)
--	g17429 = NOR(g16239, g16288)
--	g17507 = NOR(g16298, g13318)
--	g17896 = NOR(g14352, g16020)
--	g18007 = NOR(g14464, g16036)
--	g18085 = NOR(g16085, g6363)
--	g18124 = NOR(g14551, g16058)
--	g18201 = NOR(g16123, g6568)
--	g18240 = NOR(g14606, g16094)
--	g18308 = NOR(g16174, g6832)
--	g18352 = NOR(g16082, g14249)
--	g18401 = NOR(g16233, g7134)
--	g18430 = NOR(g16020, g14352)
--	g18447 = NOR(g16120, g14371)
--	g18503 = NOR(g16036, g14464)
--	g18520 = NOR(g16171, g14483)
--	g18548 = NOR(g14249, g16082)
--	g18567 = NOR(g16058, g14551)
--	g18584 = NOR(g16230, g14570)
--	g18590 = NOR(g16439, g7522)
--	g18598 = NOR(g14371, g16120)
--	g18617 = NOR(g16094, g14606)
--	g18623 = NOR(g15902, g2814)
--	g18626 = NOR(g16463, g7549)
--	g18630 = NOR(g14483, g16171)
--	g18639 = NOR(g14570, g16230)
--	g18669 = NOR(g13623, g13634)
--	g18678 = NOR(g13625, g11771)
--	g18707 = NOR(g13636, g11788)
--	g18719 = NOR(g13643, g13656)
--	g18726 = NOR(g13645, g11805)
--	g18743 = NOR(g13648, g11814)
--	g18754 = NOR(g13655, g11816)
--	g18755 = NOR(g13871, g12274)
--	g18763 = NOR(g13671, g11838)
--	g18780 = NOR(g13674, g11847)
--	g18781 = NOR(g13675, g11851)
--	g18782 = NOR(g13676, g13705)
--	g18794 = NOR(g13701, g11880)
--	g18803 = NOR(g13704, g11885)
--	g18804 = NOR(g13905, g12331)
--	g18820 = NOR(g13738, g11922)
--	g18821 = NOR(g13740, g11926)
--	g18835 = NOR(g13788, g11966)
--	g18836 = NOR(g13789, g11967)
--	g18837 = NOR(g13998, g12376)
--	g18852 = NOR(g13815, g12012)
--	g18866 = NOR(g13834, g12069)
--	g18867 = NOR(g13835, g12070)
--	g18868 = NOR(g14143, g12419)
--	g18883 = NOR(g13846, g12128)
--	g18885 = NOR(g13847, g12129)
--	g18906 = NOR(g13855, g12186)
--	g18907 = NOR(g14336, g12429)
--	g18942 = NOR(g13870, g12273)
--	g18957 = NOR(g13884, g12307)
--	g18968 = NOR(g13904, g12330)
--	g18975 = NOR(g13944, g12353)
--	g19144 = NOR(g17268, g14884)
--	g19149 = NOR(g17339, g15020)
--	g19153 = NOR(g17381, g15093)
--	g19154 = NOR(g17382, g15094)
--	g19157 = NOR(g17428, g15171)
--	g19160 = NOR(g17446, g15178)
--	g19162 = NOR(g17485, g15243)
--	g19163 = NOR(g17486, g15244)
--	g19165 = NOR(g17526, g15264)
--	g19167 = NOR(g17556, g15320)
--	g19171 = NOR(g17616, g15356)
--	g19172 = NOR(g17635, g15388)
--	g19173 = NOR(g17636, g15389)
--	g19177 = NOR(g17713, g15442)
--	g19178 = NOR(g17718, g15452)
--	g19179 = NOR(g17719, g15453)
--	g19184 = NOR(g17798, g15520)
--	g19219 = NOR(g18165, g15753)
--	g20008 = NOR(g18977, g7338)
--	g20054 = NOR(g19001, g16867)
--	g20095 = NOR(g16507, g16895)
--	g20120 = NOR(g16529, g16924)
--	g20150 = NOR(g16560, g16954)
--	g20153 = NOR(g16536, g7583)
--	g20299 = NOR(g16665, g16884)
--	g20310 = NOR(g16850, g13654)
--	g20314 = NOR(g13646, g16855)
--	g20318 = NOR(g16686, g16913)
--	g20333 = NOR(g13672, g16859)
--	g20337 = NOR(g16712, g16943)
--	g20343 = NOR(g16856, g13703)
--	g20353 = NOR(g13702, g16864)
--	g20357 = NOR(g16743, g16974)
--	g20375 = NOR(g13739, g16879)
--	g20376 = NOR(g16865, g13787)
--	g20417 = NOR(g16907, g13833)
--	g20682 = NOR(g19160, g10024)
--	g20717 = NOR(g19165, g10133)
--	g20752 = NOR(g19171, g10238)
--	g20789 = NOR(g19177, g10340)
--	g20841 = NOR(g14767, g19552)
--	g20874 = NOR(g17301, g19594)
--	g20875 = NOR(g19584, g17352)
--	g20876 = NOR(g19585, g17353)
--	g20877 = NOR(g3919, g19830)
--	g20878 = NOR(g19600, g17395)
--	g20879 = NOR(g19601, g17396)
--	g20880 = NOR(g19602, g17397)
--	g20881 = NOR(g19603, g17398)
--	g20882 = NOR(g19614, g17408)
--	g20883 = NOR(g19615, g17409)
--	g20884 = NOR(g5394, g19830)
--	g20891 = NOR(g19626, g17447)
--	g20892 = NOR(g19627, g17448)
--	g20893 = NOR(g19628, g17449)
--	g20894 = NOR(g19629, g17450)
--	g20895 = NOR(g19633, g17461)
--	g20896 = NOR(g19634, g17462)
--	g20897 = NOR(g19635, g17463)
--	g20898 = NOR(g19636, g17464)
--	g20899 = NOR(g19647, g17474)
--	g20900 = NOR(g19648, g17475)
--	g20901 = NOR(g19660, g17508)
--	g20902 = NOR(g19661, g17509)
--	g20903 = NOR(g19662, g17510)
--	g20910 = NOR(g19666, g17527)
--	g20911 = NOR(g19667, g17528)
--	g20912 = NOR(g19668, g17529)
--	g20913 = NOR(g19669, g17530)
--	g20914 = NOR(g19673, g17541)
--	g20915 = NOR(g19674, g17542)
--	g20916 = NOR(g19675, g17543)
--	g20917 = NOR(g19676, g17544)
--	g20918 = NOR(g19687, g17554)
--	g20919 = NOR(g19688, g17555)
--	g20920 = NOR(g19691, g19726)
--	g20921 = NOR(g19697, g17576)
--	g20922 = NOR(g19698, g17577)
--	g20923 = NOR(g19699, g17578)
--	g20924 = NOR(g19700, g15257)
--	g20925 = NOR(g19708, g17598)
--	g20926 = NOR(g19709, g17599)
--	g20927 = NOR(g19710, g17600)
--	g20934 = NOR(g19714, g17617)
--	g20935 = NOR(g19715, g17618)
--	g20936 = NOR(g19716, g17619)
--	g20937 = NOR(g19717, g17620)
--	g20938 = NOR(g19721, g17631)
--	g20939 = NOR(g19722, g17632)
--	g20940 = NOR(g19723, g17633)
--	g20941 = NOR(g19724, g17634)
--	g20944 = NOR(g19731, g17652)
--	g20945 = NOR(g19732, g17653)
--	g20946 = NOR(g19733, g17654)
--	g20947 = NOR(g19734, g15335)
--	g20948 = NOR(g19735, g15336)
--	g20949 = NOR(g19741, g17673)
--	g20950 = NOR(g19742, g17674)
--	g20951 = NOR(g19743, g17675)
--	g20952 = NOR(g19744, g15349)
--	g20953 = NOR(g19752, g17695)
--	g20954 = NOR(g19753, g17696)
--	g20955 = NOR(g19754, g17697)
--	g20962 = NOR(g19758, g17714)
--	g20963 = NOR(g19759, g17715)
--	g20964 = NOR(g19760, g17716)
--	g20965 = NOR(g19761, g17717)
--	g20966 = NOR(g19765, g17734)
--	g20967 = NOR(g19766, g17735)
--	g20968 = NOR(g19767, g17736)
--	g20969 = NOR(g19768, g15402)
--	g20970 = NOR(g19769, g15403)
--	g20972 = NOR(g19774, g17752)
--	g20973 = NOR(g19775, g17753)
--	g20974 = NOR(g19776, g17754)
--	g20975 = NOR(g19777, g15421)
--	g20976 = NOR(g19778, g15422)
--	g20977 = NOR(g19784, g17773)
--	g20978 = NOR(g19785, g17774)
--	g20979 = NOR(g19786, g17775)
--	g20980 = NOR(g19787, g15435)
--	g20981 = NOR(g19795, g17795)
--	g20982 = NOR(g19796, g17796)
--	g20983 = NOR(g19797, g17797)
--	g20989 = NOR(g19802, g17812)
--	g20990 = NOR(g19803, g17813)
--	g20991 = NOR(g19804, g17814)
--	g20992 = NOR(g19805, g15470)
--	g20993 = NOR(g19807, g17835)
--	g20994 = NOR(g19808, g17836)
--	g20995 = NOR(g19809, g17837)
--	g20996 = NOR(g19810, g15486)
--	g20997 = NOR(g19811, g15487)
--	g20999 = NOR(g19816, g17853)
--	g21000 = NOR(g19817, g17854)
--	g21001 = NOR(g19818, g17855)
--	g21002 = NOR(g19819, g15505)
--	g21003 = NOR(g19820, g15506)
--	g21004 = NOR(g19826, g17874)
--	g21005 = NOR(g19827, g17875)
--	g21006 = NOR(g19828, g17876)
--	g21007 = NOR(g19829, g15519)
--	g21008 = NOR(g19836, g17877)
--	g21009 = NOR(g19839, g17900)
--	g21010 = NOR(g19840, g17901)
--	g21011 = NOR(g19841, g17902)
--	g21015 = NOR(g19846, g17924)
--	g21016 = NOR(g19847, g17925)
--	g21017 = NOR(g19848, g17926)
--	g21018 = NOR(g19849, g15556)
--	g21019 = NOR(g19851, g17947)
--	g21020 = NOR(g19852, g17948)
--	g21021 = NOR(g19853, g17949)
--	g21022 = NOR(g19854, g15572)
--	g21023 = NOR(g19855, g15573)
--	g21025 = NOR(g19860, g17965)
--	g21026 = NOR(g19861, g17966)
--	g21027 = NOR(g19862, g17967)
--	g21028 = NOR(g19863, g15591)
--	g21029 = NOR(g19864, g15592)
--	g21031 = NOR(g19869, g17989)
--	g21032 = NOR(g19870, g17990)
--	g21033 = NOR(g19872, g18011)
--	g21034 = NOR(g19873, g18012)
--	g21035 = NOR(g19874, g18013)
--	g21039 = NOR(g19879, g18035)
--	g21040 = NOR(g19880, g18036)
--	g21041 = NOR(g19881, g18037)
--	g21042 = NOR(g19882, g15634)
--	g21043 = NOR(g19884, g18058)
--	g21044 = NOR(g19885, g18059)
--	g21045 = NOR(g19886, g18060)
--	g21046 = NOR(g19887, g15650)
--	g21047 = NOR(g19888, g15651)
--	g21048 = NOR(g19889, g18062)
--	g21051 = NOR(g19895, g18088)
--	g21052 = NOR(g19900, g18106)
--	g21053 = NOR(g19901, g18107)
--	g21054 = NOR(g19903, g18128)
--	g21055 = NOR(g19904, g18129)
--	g21056 = NOR(g19905, g18130)
--	g21060 = NOR(g19910, g18152)
--	g21061 = NOR(g19911, g18153)
--	g21062 = NOR(g19912, g18154)
--	g21063 = NOR(g19913, g15710)
--	g21065 = NOR(g19914, g18169)
--	g21070 = NOR(g19920, g18204)
--	g21071 = NOR(g19925, g18222)
--	g21072 = NOR(g19926, g18223)
--	g21073 = NOR(g19928, g18244)
--	g21074 = NOR(g19929, g18245)
--	g21075 = NOR(g19930, g18246)
--	g21080 = NOR(g19935, g18311)
--	g21081 = NOR(g19940, g18329)
--	g21082 = NOR(g19941, g18330)
--	g21083 = NOR(g19943, g18333)
--	g21084 = NOR(g20011, g20048)
--	g21094 = NOR(g19952, g18404)
--	g21095 = NOR(g20012, g20049, g20084)
--	g21096 = NOR(g20013, g20051, g20087)
--	g21104 = NOR(g20050, g20085, g20106)
--	g21105 = NOR(g20052, g20088, g20109)
--	g21106 = NOR(g20053, g20090, g20112)
--	g21116 = NOR(g20086, g20107, g20131)
--	g21117 = NOR(g20089, g20110, g20133)
--	g21118 = NOR(g20091, g20113, g20136)
--	g21119 = NOR(g20092, g20115, g20139)
--	g21133 = NOR(g20108, g20132, g20156)
--	g21134 = NOR(g20111, g20134, g20157)
--	g21135 = NOR(g20114, g20137, g20160)
--	g21147 = NOR(g20135, g20158, g20188)
--	g21148 = NOR(g20138, g20161, g20190)
--	g21149 = NOR(g20015, g19981)
--	g21167 = NOR(g20159, g20189)
--	g21168 = NOR(g20162, g20191, g20220)
--	g21169 = NOR(g20057, g20019)
--	g21183 = NOR(g20192, g20221)
--	g21189 = NOR(g20098, g20061)
--	g21204 = NOR(g20123, g20102)
--	g21211 = NOR(g19240, g19230)
--	g21219 = NOR(g19253, g19243)
--	g21227 = NOR(g18414, g18485, g20295)
--	g21228 = NOR(g19388, g17118)
--	g21230 = NOR(g19266, g19256)
--	g21233 = NOR(g19418, g17145)
--	g21235 = NOR(g19281, g19269)
--	g21238 = NOR(g19954, g5890)
--	g21242 = NOR(g19455, g17168)
--	g21246 = NOR(g19984, g5929)
--	g21250 = NOR(g19482, g17183)
--	g21255 = NOR(g20022, g5963)
--	g21263 = NOR(g20064, g5992)
--	g21316 = NOR(g20460, g16111)
--	g21331 = NOR(g20472, g16153)
--	g21346 = NOR(g20480, g13247)
--	g21364 = NOR(g20486, g13266)
--	g21385 = NOR(g20492, g13289)
--	g21407 = NOR(g20499, g13316)
--	g21432 = NOR(g20502, g13335)
--	g21435 = NOR(g20503, g16385)
--	g21467 = NOR(g20506, g13355)
--	g21470 = NOR(g20512, g16417)
--	g21502 = NOR(g20525, g16445)
--	g21615 = NOR(g16567, g19957)
--	g21618 = NOR(g20016, g14079, g14165)
--	g21636 = NOR(g20473, g6513)
--	g21643 = NOR(g16591, g19987)
--	g21646 = NOR(g20058, g14194, g14280)
--	g21665 = NOR(g20507, g18352)
--	g21667 = NOR(g20481, g6777)
--	g21674 = NOR(g16611, g20025)
--	g21677 = NOR(g20099, g14309, g14402)
--	g21694 = NOR(g20526, g18447)
--	g21696 = NOR(g20487, g7079)
--	g21703 = NOR(g16629, g20067)
--	g21706 = NOR(g20124, g14431, g14514)
--	g21711 = NOR(g19830, g15780)
--	g21730 = NOR(g20545, g18520)
--	g21732 = NOR(g20493, g7329)
--	g21738 = NOR(g19444, g17893, g14079)
--	g21739 = NOR(g20507, g18430)
--	g21756 = NOR(g19070, g18584)
--	g21762 = NOR(g19471, g18004, g14194)
--	g21763 = NOR(g20526, g18503)
--	g21778 = NOR(g19494, g18121, g14309)
--	g21779 = NOR(g20545, g18567)
--	g21793 = NOR(g19515, g18237, g14431)
--	g21794 = NOR(g19070, g18617)
--	g21796 = NOR(g19830, g13004)
--	g21842 = NOR(g13609, g19150)
--	g21843 = NOR(g13619, g19155)
--	g21845 = NOR(g13631, g19161)
--	g21847 = NOR(g13642, g19166)
--	g21851 = NOR(g19252, g8842)
--	g21878 = NOR(g16964, g19228)
--	g21880 = NOR(g13854, g19236)
--	g21882 = NOR(g13862, g19248)
--	g21884 = NOR(g19260, g19284)
--	g21887 = NOR(g13519, g19289)
--	g21889 = NOR(g19285, g19316)
--	g21890 = NOR(g13530, g19307)
--	g21893 = NOR(g13541, g19328)
--	g21894 = NOR(g19317, g19356)
--	g21901 = NOR(g13552, g19355)
--	g21968 = NOR(g21234, g19476)
--	g21969 = NOR(g20895, g10133)
--	g21970 = NOR(g17182, g21226)
--	g21971 = NOR(g21243, g19499)
--	g21972 = NOR(g20914, g10238)
--	g21973 = NOR(g21251, g19520)
--	g21974 = NOR(g20938, g10340)
--	g21975 = NOR(g21245, g21259)
--	g21980 = NOR(g21252, g19531, g19540)
--	g21981 = NOR(g21254, g21267)
--	g21987 = NOR(g21260, g19541, g19544)
--	g21988 = NOR(g21262, g21276)
--	g22000 = NOR(g21268, g19545, g19547)
--	g22001 = NOR(g21270, g21283)
--	g22013 = NOR(g21277, g19548, g19551)
--	g22025 = NOR(g21284, g19549)
--	g22026 = NOR(g21083, g18407)
--	g22027 = NOR(g21290, g19553)
--	g22028 = NOR(g21291, g19554)
--	g22029 = NOR(g21292, g19555)
--	g22030 = NOR(g21298, g19557)
--	g22031 = NOR(g21299, g19558)
--	g22032 = NOR(g21300, g19559)
--	g22033 = NOR(g21301, g19560)
--	g22034 = NOR(g21302, g19561)
--	g22035 = NOR(g21303, g19562)
--	g22037 = NOR(g21304, g19564)
--	g22038 = NOR(g21305, g19565)
--	g22039 = NOR(g21306, g19566)
--	g22040 = NOR(g21307, g19567)
--	g22041 = NOR(g21308, g19568)
--	g22042 = NOR(g21309, g19569)
--	g22043 = NOR(g21310, g19570)
--	g22044 = NOR(g21311, g19571)
--	g22045 = NOR(g21312, g19572)
--	g22047 = NOR(g21313, g19574)
--	g22048 = NOR(g21314, g19575)
--	g22049 = NOR(g21315, g19576)
--	g22054 = NOR(g21319, g19586)
--	g22055 = NOR(g21320, g19587)
--	g22056 = NOR(g21321, g19588)
--	g22057 = NOR(g21322, g19589)
--	g22058 = NOR(g21323, g19590)
--	g22059 = NOR(g21324, g19591)
--	g22060 = NOR(g21325, g19592)
--	g22061 = NOR(g21326, g19593)
--	g22063 = NOR(g21328, g19597)
--	g22064 = NOR(g21329, g19598)
--	g22065 = NOR(g21330, g19599)
--	g22066 = NOR(g21334, g19604)
--	g22067 = NOR(g21335, g19605)
--	g22068 = NOR(g21336, g19606)
--	g22073 = NOR(g21337, g19616)
--	g22074 = NOR(g21338, g19617)
--	g22075 = NOR(g21339, g19618)
--	g22076 = NOR(g21340, g19619)
--	g22077 = NOR(g21341, g19620)
--	g22078 = NOR(g21342, g19621)
--	g22079 = NOR(g21343, g19623)
--	g22080 = NOR(g21344, g19624)
--	g22081 = NOR(g21345, g19625)
--	g22087 = NOR(g21349, g19630)
--	g22088 = NOR(g21350, g19631)
--	g22089 = NOR(g21351, g19632)
--	g22090 = NOR(g21352, g19637)
--	g22091 = NOR(g21353, g19638)
--	g22092 = NOR(g21354, g19639)
--	g22097 = NOR(g21355, g19649)
--	g22098 = NOR(g21356, g19650)
--	g22099 = NOR(g21357, g19651)
--	g22100 = NOR(g21360, g19653)
--	g22101 = NOR(g21361, g19654)
--	g22102 = NOR(g21362, g19655)
--	g22103 = NOR(g21363, g19656)
--	g22104 = NOR(g21367, g19663)
--	g22105 = NOR(g21368, g19664)
--	g22106 = NOR(g21369, g19665)
--	g22112 = NOR(g21370, g19670)
--	g22113 = NOR(g21371, g19671)
--	g22114 = NOR(g21372, g19672)
--	g22115 = NOR(g21373, g19677)
--	g22116 = NOR(g21374, g19678)
--	g22117 = NOR(g21375, g19679)
--	g22122 = NOR(g21378, g19692)
--	g22123 = NOR(g21379, g19693)
--	g22124 = NOR(g21380, g19694)
--	g22125 = NOR(g21381, g19695)
--	g22126 = NOR(g21389, g19701)
--	g22127 = NOR(g21390, g19702)
--	g22128 = NOR(g21391, g19703)
--	g22129 = NOR(g21392, g19704)
--	g22130 = NOR(g21393, g19711)
--	g22131 = NOR(g21394, g19712)
--	g22132 = NOR(g21395, g19713)
--	g22138 = NOR(g21396, g19718)
--	g22139 = NOR(g21397, g19719)
--	g22140 = NOR(g21398, g19720)
--	g22141 = NOR(g21401, g19727)
--	g22142 = NOR(g21402, g19728)
--	g22143 = NOR(g21403, g19729)
--	g22144 = NOR(g21410, g19730)
--	g22145 = NOR(g21411, g19736)
--	g22146 = NOR(g21412, g19737)
--	g22147 = NOR(g21413, g19738)
--	g22148 = NOR(g21414, g19739)
--	g22149 = NOR(g21419, g19745)
--	g22150 = NOR(g21420, g19746)
--	g22151 = NOR(g21421, g19747)
--	g22152 = NOR(g21422, g19748)
--	g22153 = NOR(g21423, g19755)
--	g22154 = NOR(g21424, g19756)
--	g22155 = NOR(g21425, g19757)
--	g22161 = NOR(g21428, g19764)
--	g22162 = NOR(g21438, g19770)
--	g22163 = NOR(g21439, g19771)
--	g22164 = NOR(g21440, g19772)
--	g22165 = NOR(g21444, g19773)
--	g22166 = NOR(g21445, g19779)
--	g22167 = NOR(g21446, g19780)
--	g22168 = NOR(g21447, g19781)
--	g22169 = NOR(g21448, g19782)
--	g22170 = NOR(g21453, g19788)
--	g22171 = NOR(g21454, g19789)
--	g22172 = NOR(g21455, g19790)
--	g22173 = NOR(g21456, g19791)
--	g22174 = NOR(g19868, g21593)
--	g22177 = NOR(g21476, g19806)
--	g22178 = NOR(g21480, g19812)
--	g22179 = NOR(g21481, g19813)
--	g22180 = NOR(g21482, g19814)
--	g22181 = NOR(g21486, g19815)
--	g22182 = NOR(g21487, g19821)
--	g22183 = NOR(g21488, g19822)
--	g22184 = NOR(g21489, g19823)
--	g22185 = NOR(g21490, g19824)
--	g22186 = NOR(g21497, g19837)
--	g22189 = NOR(g19899, g21622)
--	g22191 = NOR(g21517, g19850)
--	g22192 = NOR(g21521, g19856)
--	g22193 = NOR(g21522, g19857)
--	g22194 = NOR(g21523, g19858)
--	g22195 = NOR(g21527, g19859)
--	g22198 = NOR(g19924, g21650)
--	g22200 = NOR(g21553, g19883)
--	g22204 = NOR(g19939, g21681)
--	g22210 = NOR(g21610, g19932)
--	g22216 = NOR(g21635, g19944)
--	g22218 = NOR(g21639, g19949)
--	g22227 = NOR(g21658, g19953)
--	g22231 = NOR(g21666, g19971)
--	g22234 = NOR(g21670, g19976)
--	g22242 = NOR(g21687, g19983)
--	g22247 = NOR(g21695, g20001)
--	g22249 = NOR(g21699, g20006)
--	g22263 = NOR(g21723, g20021)
--	g22267 = NOR(g21731, g20039)
--	g22269 = NOR(g21735, g20044)
--	g22280 = NOR(g21749, g20063)
--	g22284 = NOR(g21757, g20081)
--	g22288 = NOR(g20144, g21805)
--	g22299 = NOR(g21773, g20104)
--	g22308 = NOR(g20182, g21812)
--	g22336 = NOR(g20216, g21818)
--	g22361 = NOR(g20246, g21822)
--	g22454 = NOR(g17012, g21891)
--	g22493 = NOR(g17042, g21899)
--	g22536 = NOR(g17076, g21911)
--	g22576 = NOR(g17111, g21925)
--	g22578 = NOR(g21892, g18982)
--	g22615 = NOR(g21900, g18990)
--	g22651 = NOR(g21912, g18997)
--	g22687 = NOR(g21926, g19010)
--	g22755 = NOR(g21271, g20842)
--	g22784 = NOR(g16075, g20885)
--	g22789 = NOR(g21278, g20850)
--	g22810 = NOR(g16075, g20842, g21271)
--	g22826 = NOR(g16113, g20904)
--	g22831 = NOR(g21285, g20858)
--	g22851 = NOR(g16113, g20850, g21278)
--	g22865 = NOR(g16164, g20928)
--	g22870 = NOR(g21293, g20866)
--	g22886 = NOR(g16164, g20858, g21285)
--	g22900 = NOR(g16223, g20956)
--	g22921 = NOR(g16223, g20866, g21293)
--	g22935 = NOR(g21903, g7466)
--	g22953 = NOR(g20700, g7595)
--	g22985 = NOR(g21618, g21049)
--	g22987 = NOR(g21646, g21068)
--	g22990 = NOR(g21677, g21078)
--	g22997 = NOR(g21706, g21092)
--	g22999 = NOR(g21085, g19241)
--	g23000 = NOR(g16909, g21067)
--	g23009 = NOR(g21738, g21107)
--	g23013 = NOR(g21097, g19254)
--	g23014 = NOR(g16939, g21077)
--	g23022 = NOR(g16968, g21086)
--	g23023 = NOR(g14256, g14175, g21123)
--	g23025 = NOR(g21762, g21124)
--	g23029 = NOR(g21111, g19267)
--	g23030 = NOR(g16970, g21091)
--	g23039 = NOR(g16989, g21098)
--	g23040 = NOR(g14378, g14290, g21142)
--	g23042 = NOR(g21778, g21143)
--	g23046 = NOR(g21128, g19282)
--	g23047 = NOR(g16991, g21103)
--	g23051 = NOR(g21121, g21153)
--	g23058 = NOR(g16999, g21112)
--	g23059 = NOR(g14490, g14412, g21162)
--	g23061 = NOR(g21793, g21163)
--	g23066 = NOR(g21138, g19303, g19320)
--	g23067 = NOR(g17015, g21122)
--	g23070 = NOR(g21140, g21173)
--	g23076 = NOR(g17023, g21129)
--	g23077 = NOR(g14577, g14524, g21182)
--	g23080 = NOR(g21158, g19324, g19347)
--	g23081 = NOR(g17045, g21141)
--	g23083 = NOR(g21160, g21193)
--	g23092 = NOR(g17055, g21154)
--	g23093 = NOR(g17056, g21155)
--	g23096 = NOR(g21178, g19351, g19381)
--	g23097 = NOR(g17079, g21161)
--	g23099 = NOR(g21180, g21208)
--	g23110 = NOR(g17090, g21174)
--	g23111 = NOR(g17091, g21175)
--	g23113 = NOR(g21198, g19385, g19413)
--	g23114 = NOR(g17114, g21181)
--	g23117 = NOR(g17117, g21188)
--	g23123 = NOR(g17128, g21194)
--	g23124 = NOR(g17129, g21195)
--	g23126 = NOR(g17144, g21203)
--	g23132 = NOR(g17155, g21209)
--	g23133 = NOR(g17156, g21210)
--	g23135 = NOR(g21229, g19449)
--	g23136 = NOR(g20878, g10024)
--	g23137 = NOR(g17167, g21218)
--	g23324 = NOR(g22144, g10024)
--	g23329 = NOR(g22165, g10133)
--	g23330 = NOR(g22186, g22777)
--	g23339 = NOR(g22181, g10238)
--	g23348 = NOR(g22195, g10340)
--	g23357 = NOR(g22210, g20127)
--	g23358 = NOR(g22227, g18407)
--	g23359 = NOR(g22216, g22907)
--	g23385 = NOR(g17393, g22517)
--	g23386 = NOR(g22483, g21388)
--	g23392 = NOR(g17460, g22557)
--	g23393 = NOR(g22526, g21418)
--	g23399 = NOR(g17506, g22581)
--	g23400 = NOR(g17540, g22597)
--	g23401 = NOR(g22566, g21452)
--	g23406 = NOR(g17597, g22618)
--	g23407 = NOR(g17630, g22634)
--	g23408 = NOR(g22606, g21494)
--	g23413 = NOR(g17694, g22654)
--	g23418 = NOR(g17794, g22690)
--	g23427 = NOR(g22699, g21589)
--	g23433 = NOR(g22726, g21611)
--	g23461 = NOR(g22841, g21707)
--	g23477 = NOR(g22906, g21758)
--	g23497 = NOR(g22876, g5606)
--	g23513 = NOR(g22911, g5631)
--	g23528 = NOR(g22936, g5659)
--	g23539 = NOR(g22942, g5697)
--	g23545 = NOR(g22984, g20285)
--	g23823 = NOR(g23009, g18490, g4456)
--	g23858 = NOR(g23025, g18554, g4632)
--	g23892 = NOR(g23042, g18604, g4809)
--	g23913 = NOR(g23061, g18636, g4985)
--	g23922 = NOR(g4456, g22985)
--	g23945 = NOR(g4456, g13565, g23009)
--	g23950 = NOR(g22992, g6707)
--	g23954 = NOR(g4632, g22987)
--	g23974 = NOR(g4632, g13573, g23025)
--	g23979 = NOR(g23003, g7009)
--	g23983 = NOR(g4809, g22990)
--	g24004 = NOR(g4809, g13582, g23042)
--	g24009 = NOR(g23017, g7259)
--	g24013 = NOR(g4985, g22997)
--	g24038 = NOR(g4985, g13602, g23061)
--	g24043 = NOR(g23033, g7455)
--	g24059 = NOR(g21990, g20809)
--	g24072 = NOR(g22004, g20826)
--	g24083 = NOR(g22015, g20836)
--	g24092 = NOR(g22020, g20840)
--	g24174 = NOR(g16894, g22206)
--	g24178 = NOR(g16908, g22211)
--	g24179 = NOR(g16923, g22214)
--	g24181 = NOR(g16938, g22220)
--	g24182 = NOR(g16953, g22223)
--	g24206 = NOR(g16966, g22228)
--	g24207 = NOR(g16967, g22229)
--	g24208 = NOR(g16969, g22235)
--	g24209 = NOR(g16984, g22238)
--	g24212 = NOR(g16987, g22244)
--	g24213 = NOR(g16988, g22245)
--	g24214 = NOR(g16990, g22250)
--	g24215 = NOR(g16993, g22254)
--	g24216 = NOR(g16994, g22255)
--	g24218 = NOR(g16997, g22264)
--	g24219 = NOR(g16998, g22265)
--	g24222 = NOR(g17017, g22272)
--	g24223 = NOR(g17018, g22273)
--	g24225 = NOR(g17021, g22281)
--	g24226 = NOR(g17022, g22282)
--	g24227 = NOR(g22270, g21137)
--	g24228 = NOR(g17028, g22285)
--	g24230 = NOR(g17047, g22291)
--	g24231 = NOR(g17048, g22292)
--	g24232 = NOR(g22637, g22665)
--	g24234 = NOR(g22289, g21157)
--	g24235 = NOR(g17062, g22305)
--	g24237 = NOR(g17081, g22311)
--	g24238 = NOR(g17082, g22312)
--	g24242 = NOR(g22309, g21177)
--	g24243 = NOR(g17097, g22333)
--	g24249 = NOR(g22337, g21197)
--	g24250 = NOR(g17135, g22358)
--	g24426 = NOR(g23386, g10024)
--	g24428 = NOR(g23544, g22398)
--	g24430 = NOR(g23393, g10133)
--	g24434 = NOR(g23401, g10238)
--	g24438 = NOR(g23408, g10340)
--	g24445 = NOR(g23427, g22777)
--	g24446 = NOR(g23433, g22907)
--	g24473 = NOR(g23461, g18407)
--	g24476 = NOR(g23477, g20127)
--	g24479 = NOR(g23593, g22516)
--	g24480 = NOR(g23617, g23659)
--	g24481 = NOR(g23618, g19696)
--	g24485 = NOR(g23625, g22556)
--	g24486 = NOR(g23643, g22577)
--	g24487 = NOR(g23666, g23709)
--	g24488 = NOR(g23667, g19740)
--	g24489 = NOR(g23674, g22596)
--	g24490 = NOR(g23686, g22607)
--	g24491 = NOR(g15247, g23735)
--	g24492 = NOR(g23689, g22610)
--	g24493 = NOR(g23693, g22614)
--	g24494 = NOR(g23716, g23763)
--	g24495 = NOR(g23717, g19783)
--	g24496 = NOR(g23724, g22633)
--	g24497 = NOR(g23734, g22638)
--	g24498 = NOR(g15324, g23777)
--	g24499 = NOR(g15325, g23778)
--	g24500 = NOR(g23740, g22643)
--	g24501 = NOR(g15339, g23790)
--	g24502 = NOR(g23743, g22646)
--	g24503 = NOR(g23747, g22650)
--	g24504 = NOR(g23770, g23818)
--	g24505 = NOR(g23771, g19825)
--	g24506 = NOR(g23776, g22667)
--	g24507 = NOR(g15391, g23824)
--	g24508 = NOR(g15392, g23825)
--	g24509 = NOR(g23789, g22674)
--	g24510 = NOR(g15410, g23830)
--	g24511 = NOR(g15411, g23831)
--	g24512 = NOR(g23795, g22679)
--	g24513 = NOR(g15425, g23843)
--	g24514 = NOR(g23798, g22682)
--	g24515 = NOR(g23802, g22686)
--	g24516 = NOR(g23820, g22700)
--	g24517 = NOR(g23822, g22701)
--	g24519 = NOR(g15459, g23855)
--	g24520 = NOR(g23829, g22707)
--	g24521 = NOR(g15475, g23859)
--	g24522 = NOR(g15476, g23860)
--	g24523 = NOR(g23842, g22714)
--	g24524 = NOR(g15494, g23865)
--	g24525 = NOR(g15495, g23866)
--	g24526 = NOR(g23848, g22719)
--	g24527 = NOR(g15509, g23878)
--	g24528 = NOR(g23851, g22722)
--	g24530 = NOR(g23857, g22732)
--	g24532 = NOR(g15545, g23889)
--	g24533 = NOR(g23864, g22738)
--	g24534 = NOR(g15561, g23893)
--	g24535 = NOR(g15562, g23894)
--	g24536 = NOR(g23877, g22745)
--	g24537 = NOR(g15580, g23899)
--	g24538 = NOR(g15581, g23900)
--	g24543 = NOR(g23891, g22764)
--	g24545 = NOR(g15623, g23910)
--	g24546 = NOR(g23898, g22770)
--	g24547 = NOR(g15639, g23914)
--	g24548 = NOR(g15640, g23915)
--	g24555 = NOR(g23912, g22798)
--	g24557 = NOR(g15699, g23942)
--	g24558 = NOR(g23917, g22804)
--	g24566 = NOR(g23944, g22842)
--	g24575 = NOR(g23972, g22874)
--	g24606 = NOR(g24183, g537)
--	g24613 = NOR(g23592, g22515)
--	g24622 = NOR(g23616, g22546)
--	g24623 = NOR(g24183, g529)
--	g24624 = NOR(g23624, g22555)
--	g24636 = NOR(g24183, g530)
--	g24637 = NOR(g23665, g22587)
--	g24638 = NOR(g23673, g22595)
--	g24652 = NOR(g24183, g531)
--	g24656 = NOR(g23715, g22624)
--	g24657 = NOR(g23723, g22632)
--	g24663 = NOR(g24183, g532)
--	g24675 = NOR(g23769, g22660)
--	g24681 = NOR(g24183, g533)
--	g24682 = NOR(g23688, g24183)
--	g24694 = NOR(g24183, g534)
--	g24708 = NOR(g23854, g22727)
--	g24711 = NOR(g24183, g536)
--	g24717 = NOR(g23886, g22754)
--	g24720 = NOR(g23888, g22759)
--	g24728 = NOR(g23907, g22788)
--	g24731 = NOR(g23909, g22793)
--	g24736 = NOR(g23939, g22830)
--	g24739 = NOR(g23941, g22835)
--	g24742 = NOR(g23971, g22869)
--	g24756 = NOR(g16089, g24211)
--	g24770 = NOR(g16119, g24217)
--	g24782 = NOR(g16160, g24221)
--	g24783 = NOR(g16161, g24224)
--	g24800 = NOR(g16211, g24229)
--	g24819 = NOR(g16262, g24236)
--	g24836 = NOR(g16309, g24241)
--	g24845 = NOR(g16350, g24246)
--	g24847 = NOR(g16356, g24247)
--	g24859 = NOR(g16390, g24253)
--	g24871 = NOR(g16422, g24256)
--	g25027 = NOR(g24227, g17001)
--	g25042 = NOR(g24234, g17031)
--	g25056 = NOR(g24242, g17065)
--	g25067 = NOR(g24249, g17100)
--	g25075 = NOR(g13880, g23483)
--	g25076 = NOR(g23409, g22187)
--	g25077 = NOR(g23414, g22196)
--	g25078 = NOR(g23419, g22201)
--	g25081 = NOR(g23423, g22202)
--	g25082 = NOR(g23428, g22207)
--	g25085 = NOR(g23432, g22208)
--	g25091 = NOR(g23434, g22215)
--	g25099 = NOR(g23440, g22224)
--	g25125 = NOR(g23510, g22340)
--	g25127 = NOR(g23525, g22363)
--	g25129 = NOR(g23536, g22383)
--	g25185 = NOR(g24492, g10024)
--	g25189 = NOR(g24502, g10133)
--	g25191 = NOR(g24516, g22777)
--	g25194 = NOR(g24514, g10238)
--	g25197 = NOR(g24528, g10340)
--	g25199 = NOR(g24558, g20127)
--	g25201 = NOR(g24575, g18407)
--	g25202 = NOR(g24566, g22907)
--	g25204 = NOR(g24745, g23547)
--	g25206 = NOR(g24746, g23550)
--	g25207 = NOR(g24747, g23551)
--	g25208 = NOR(g24748, g23552)
--	g25209 = NOR(g24749, g23554)
--	g25211 = NOR(g24750, g23558)
--	g25212 = NOR(g24751, g23559)
--	g25213 = NOR(g24752, g23560)
--	g25214 = NOR(g24754, g23563)
--	g25215 = NOR(g24755, g23564)
--	g25216 = NOR(g24757, g23565)
--	g25217 = NOR(g24758, g23567)
--	g25218 = NOR(g24760, g23571)
--	g25219 = NOR(g24761, g23572)
--	g25220 = NOR(g24762, g23573)
--	g25221 = NOR(g24767, g23577)
--	g25222 = NOR(g24768, g23578)
--	g25223 = NOR(g24769, g23579)
--	g25224 = NOR(g24772, g23582)
--	g25225 = NOR(g24773, g23583)
--	g25226 = NOR(g24774, g23584)
--	g25227 = NOR(g24775, g23586)
--	g25228 = NOR(g24776, g23590)
--	g25229 = NOR(g24777, g23591)
--	g25230 = NOR(g24779, g23598)
--	g25231 = NOR(g24780, g23599)
--	g25232 = NOR(g24781, g23600)
--	g25233 = NOR(g24788, g23604)
--	g25234 = NOR(g24789, g23605)
--	g25235 = NOR(g24790, g23606)
--	g25236 = NOR(g24792, g23609)
--	g25237 = NOR(g24793, g23610)
--	g25238 = NOR(g24794, g23611)
--	g25239 = NOR(g24796, g23615)
--	g25240 = NOR(g24798, g23622)
--	g25241 = NOR(g24799, g23623)
--	g25242 = NOR(g24802, g23630)
--	g25243 = NOR(g24803, g23631)
--	g25244 = NOR(g24804, g23632)
--	g25245 = NOR(g24809, g23636)
--	g25246 = NOR(g24810, g23637)
--	g25247 = NOR(g24811, g23638)
--	g25248 = NOR(g24818, g23664)
--	g25249 = NOR(g24821, g23671)
--	g25250 = NOR(g24822, g23672)
--	g25251 = NOR(g24824, g23679)
--	g25252 = NOR(g24825, g23680)
--	g25253 = NOR(g24826, g23681)
--	g25254 = NOR(g24831, g23687)
--	g25255 = NOR(g24838, g23714)
--	g25256 = NOR(g24840, g23721)
--	g25257 = NOR(g24841, g23722)
--	g25258 = NOR(g24846, g23741)
--	g25259 = NOR(g24853, g23768)
--	g25260 = NOR(g24858, g17737)
--	g25261 = NOR(g24861, g23796)
--	g25262 = NOR(g24869, g17824)
--	g25263 = NOR(g24874, g17838)
--	g25264 = NOR(g24876, g23849)
--	g25265 = NOR(g24878, g23852)
--	g25266 = NOR(g24881, g17912)
--	g25267 = NOR(g24884, g17936)
--	g25268 = NOR(g24888, g17950)
--	g25270 = NOR(g24898, g18023)
--	g25271 = NOR(g24901, g18047)
--	g25272 = NOR(g24905, g18061)
--	g25273 = NOR(g24907, g23904)
--	g25279 = NOR(g24921, g18140)
--	g25280 = NOR(g24924, g18164)
--	g25288 = NOR(g24938, g18256)
--	g25311 = NOR(g24964, g24029)
--	g25343 = NOR(g24975, g5623)
--	g25357 = NOR(g24986, g5651)
--	g25372 = NOR(g24997, g5689)
--	g25389 = NOR(g25005, g5741)
--	g25418 = NOR(g24482, g22319)
--	g25426 = NOR(g24183, g24616)
--	g25429 = NOR(g24482, g22319)
--	g25450 = NOR(g16018, g25086)
--	g25451 = NOR(g16048, g25102)
--	g25452 = NOR(g16101, g25117)
--	g25523 = NOR(g20842, g24429)
--	g25539 = NOR(g25088, g6157)
--	g25569 = NOR(g24708, g24490)
--	g25589 = NOR(g20850, g24433)
--	g25605 = NOR(g25096, g6184)
--	g25631 = NOR(g24717, g24497)
--	g25648 = NOR(g24720, g24500)
--	g25668 = NOR(g20858, g24437)
--	g25684 = NOR(g25106, g6216)
--	g25699 = NOR(g24613, g24506)
--	g25708 = NOR(g24728, g24509)
--	g25725 = NOR(g24731, g24512)
--	g25745 = NOR(g20866, g24440)
--	g25761 = NOR(g25112, g6305)
--	g25764 = NOR(g25076, g21615)
--	g25772 = NOR(g24624, g24520)
--	g25781 = NOR(g24736, g24523)
--	g25798 = NOR(g24739, g24526)
--	g25818 = NOR(g25077, g21643)
--	g25826 = NOR(g24638, g24533)
--	g25835 = NOR(g24742, g24536)
--	g25852 = NOR(g4456, g14831, g25078)
--	g25853 = NOR(g25081, g21674)
--	g25861 = NOR(g24657, g24546)
--	g25870 = NOR(g4456, g25078, g18429, g16075)
--	g25873 = NOR(g4632, g14904, g25082)
--	g25874 = NOR(g25085, g21703)
--	g25882 = NOR(g4632, g25082, g18502, g16113)
--	g25885 = NOR(g4809, g14985, g25091)
--	g25887 = NOR(g4809, g25091, g18566, g16164)
--	g25890 = NOR(g4985, g15074, g25099)
--	g25892 = NOR(g4985, g25099, g18616, g16223)
--	g25932 = NOR(g25125, g17001)
--	g25935 = NOR(g25127, g17031)
--	g25938 = NOR(g25129, g17065)
--	g25940 = NOR(g24428, g17100)
--	g25941 = NOR(g24529, g24540)
--	g25943 = NOR(g24541, g24550)
--	g25944 = NOR(g24542, g24552)
--	g25946 = NOR(g24553, g24561)
--	g25947 = NOR(g24554, g24563)
--	g25948 = NOR(g24564, g24571)
--	g25949 = NOR(g24565, g24573)
--	g25950 = NOR(g24574, g24580)
--	g25962 = NOR(g24591, g23496)
--	g25967 = NOR(g24596, g23512)
--	g25974 = NOR(g24604, g23527)
--	g25979 = NOR(g24611, g23538)
--	g26025 = NOR(g25392, g17193)
--	g26031 = NOR(g25273, g22777)
--	g26037 = NOR(g25311, g18407)
--	g26041 = NOR(g25475, g24855)
--	g26042 = NOR(g25505, g24867)
--	g26043 = NOR(g25506, g24870)
--	g26044 = NOR(g25552, g24882)
--	g26045 = NOR(g25553, g24885)
--	g26046 = NOR(g25618, g24899)
--	g26047 = NOR(g25619, g24902)
--	g26048 = NOR(g25628, g24906)
--	g26049 = NOR(g25629, g24908)
--	g26050 = NOR(g25697, g24922)
--	g26055 = NOR(g25881, g24974)
--	g26081 = NOR(g25470, g25482)
--	g26083 = NOR(g25426, g22319)
--	g26084 = NOR(g25487, g25513)
--	g26087 = NOR(g6068, g24183, g25319)
--	g26090 = NOR(g25518, g25560)
--	g26096 = NOR(g6068, g24183, g25394)
--	g26099 = NOR(g6068, g24183, g25313)
--	g26103 = NOR(g25565, g25626)
--	g26107 = NOR(g6068, g24183, g25383)
--	g26110 = NOR(g6068, g24183, g25305)
--	g26113 = NOR(g25426, g22319)
--	g26126 = NOR(g6068, g24183, g25368)
--	g26137 = NOR(g6068, g24183, g25355)
--	g26140 = NOR(g24183, g25430)
--	g26145 = NOR(g6068, g24183, g25347)
--	g26151 = NOR(g6068, g24183, g25335)
--	g26154 = NOR(g6068, g24183, g25329)
--	g26160 = NOR(g25951, g16162)
--	g26168 = NOR(g25953, g16212)
--	g26183 = NOR(g25957, g13270)
--	g26199 = NOR(g25961, g13291)
--	g26217 = NOR(g25963, g13320)
--	g26240 = NOR(g25968, g13340)
--	g26265 = NOR(g25972, g13360)
--	g26272 = NOR(g25973, g16423)
--	g26283 = NOR(g25954, g24486)
--	g26295 = NOR(g25977, g13385)
--	g26304 = NOR(g25978, g16451)
--	g26327 = NOR(g25958, g24493)
--	g26336 = NOR(g25981, g13481)
--	g26374 = NOR(g25964, g24503)
--	g26417 = NOR(g25969, g24515)
--	g26529 = NOR(g25962, g17001)
--	g26530 = NOR(g25967, g17031)
--	g26531 = NOR(g25974, g17065)
--	g26532 = NOR(g25979, g17100)
--	g26534 = NOR(g25321, g8869)
--	g26541 = NOR(g13755, g25269)
--	g26545 = NOR(g13790, g25277)
--	g26547 = NOR(g13796, g25278)
--	g26553 = NOR(g13816, g25282)
--	g26557 = NOR(g13818, g25286)
--	g26559 = NOR(g13824, g25287)
--	g26560 = NOR(g25281, g24559)
--	g26569 = NOR(g13837, g25290)
--	g26573 = NOR(g13839, g25294)
--	g26575 = NOR(g13845, g25295)
--	g26583 = NOR(g25289, g24569)
--	g26592 = NOR(g13851, g25300)
--	g26596 = NOR(g13853, g25304)
--	g26607 = NOR(g25299, g24578)
--	g26616 = NOR(g13860, g25310)
--	g26630 = NOR(g25309, g24585)
--	g26655 = NOR(g25328, g17084)
--	g26659 = NOR(g25334, g17116)
--	g26660 = NOR(g25208, g10024)
--	g26661 = NOR(g25337, g17122)
--	g26664 = NOR(g25346, g17138)
--	g26665 = NOR(g25348, g17143)
--	g26666 = NOR(g25216, g10133)
--	g26667 = NOR(g25351, g17149)
--	g26669 = NOR(g25360, g17161)
--	g26670 = NOR(g25362, g17166)
--	g26671 = NOR(g25226, g10238)
--	g26672 = NOR(g25365, g17172)
--	g26675 = NOR(g25375, g17176)
--	g26676 = NOR(g25377, g17181)
--	g26677 = NOR(g25238, g10340)
--	g26776 = NOR(g26042, g10024)
--	g26781 = NOR(g26044, g10133)
--	g26786 = NOR(g26049, g22777)
--	g26789 = NOR(g26046, g10238)
--	g26795 = NOR(g26050, g10340)
--	g26798 = NOR(g26055, g18407)
--	g26799 = NOR(g26158, g25453)
--	g26800 = NOR(g26163, g25457)
--	g26801 = NOR(g26171, g25461)
--	g26802 = NOR(g26188, g25466)
--	g26803 = NOR(g15105, g26213)
--	g26804 = NOR(g15172, g26235)
--	g26805 = NOR(g15173, g26236)
--	g26806 = NOR(g15197, g26244)
--	g26807 = NOR(g15245, g26261)
--	g26808 = NOR(g15246, g26262)
--	g26809 = NOR(g15258, g26270)
--	g26810 = NOR(g15259, g26271)
--	g26811 = NOR(g15283, g26279)
--	g26812 = NOR(g15321, g26291)
--	g26813 = NOR(g15337, g26302)
--	g26814 = NOR(g15338, g26303)
--	g26815 = NOR(g15350, g26311)
--	g26816 = NOR(g15351, g26312)
--	g26817 = NOR(g15375, g26317)
--	g26818 = NOR(g15407, g26335)
--	g26820 = NOR(g15423, g26346)
--	g26821 = NOR(g15424, g26347)
--	g26822 = NOR(g15436, g26352)
--	g26823 = NOR(g15437, g26353)
--	g26824 = NOR(g15491, g26382)
--	g26825 = NOR(g15507, g26390)
--	g26826 = NOR(g15508, g26391)
--	g26827 = NOR(g15577, g26425)
--	g26869 = NOR(g26458, g5642)
--	g26873 = NOR(g25483, g26260)
--	g26877 = NOR(g26140, g22319)
--	g26878 = NOR(g26482, g5680)
--	g26882 = NOR(g25514, g26301)
--	g26885 = NOR(g26140, g22319)
--	g26887 = NOR(g26498, g5732)
--	g26891 = NOR(g25561, g26345)
--	g26897 = NOR(g26513, g5790)
--	g26901 = NOR(g25627, g26389)
--	g26905 = NOR(g26096, g22319)
--	g26914 = NOR(g26107, g22319)
--	g26988 = NOR(g24893, g26023)
--	g26989 = NOR(g26663, g21913)
--	g27011 = NOR(g24916, g26026)
--	g27012 = NOR(g26668, g21931)
--	g27037 = NOR(g24933, g26028)
--	g27038 = NOR(g26674, g20640)
--	g27051 = NOR(g4456, g26081)
--	g27065 = NOR(g24945, g26029)
--	g27066 = NOR(g26024, g20665)
--	g27078 = NOR(g4632, g26084)
--	g27094 = NOR(g4809, g26090)
--	g27106 = NOR(g4985, g26103)
--	g27120 = NOR(g26560, g17001)
--	g27123 = NOR(g26583, g17031)
--	g27129 = NOR(g26607, g17065)
--	g27131 = NOR(g26630, g17100)
--	g27144 = NOR(g23451, g26052)
--	g27147 = NOR(g23458, g26054)
--	g27149 = NOR(g23462, g26060)
--	g27152 = NOR(g23467, g26062)
--	g27157 = NOR(g23471, g26067)
--	g27160 = NOR(g23476, g26069)
--	g27165 = NOR(g23484, g26074)
--	g27174 = NOR(g23494, g26080)
--	g27175 = NOR(g26075, g25342)
--	g27179 = NOR(g26082, g25356)
--	g27184 = NOR(g26085, g25371)
--	g27188 = NOR(g26091, g25388)
--	g27243 = NOR(g26802, g10340)
--	g27250 = NOR(g26955, g26166)
--	g27251 = NOR(g26958, g26186)
--	g27252 = NOR(g26963, g26207)
--	g27253 = NOR(g26965, g26212)
--	g27254 = NOR(g26968, g26231)
--	g27255 = NOR(g26969, g26233)
--	g27256 = NOR(g26970, g26234)
--	g27257 = NOR(g26971, g26243)
--	g27258 = NOR(g26977, g26257)
--	g27259 = NOR(g26978, g26258)
--	g27260 = NOR(g26979, g26259)
--	g27261 = NOR(g26980, g26263)
--	g27262 = NOR(g26981, g26268)
--	g27263 = NOR(g26982, g26269)
--	g27264 = NOR(g26984, g26278)
--	g27265 = NOR(g26993, g26288)
--	g27266 = NOR(g26994, g26289)
--	g27267 = NOR(g26995, g26290)
--	g27268 = NOR(g26996, g26292)
--	g27269 = NOR(g26997, g26293)
--	g27270 = NOR(g26998, g26298)
--	g27271 = NOR(g26999, g26299)
--	g27272 = NOR(g27000, g26300)
--	g27273 = NOR(g27001, g26307)
--	g27274 = NOR(g27002, g26309)
--	g27275 = NOR(g27003, g26310)
--	g27276 = NOR(g27004, g26316)
--	g27277 = NOR(g27005, g26318)
--	g27278 = NOR(g27006, g26319)
--	g27279 = NOR(g27007, g26324)
--	g27280 = NOR(g27008, g26325)
--	g27281 = NOR(g27009, g26326)
--	g27282 = NOR(g27016, g26332)
--	g27283 = NOR(g27017, g26333)
--	g27284 = NOR(g27018, g26334)
--	g27285 = NOR(g27019, g26339)
--	g27286 = NOR(g27020, g26340)
--	g27287 = NOR(g27021, g26342)
--	g27288 = NOR(g27022, g26343)
--	g27289 = NOR(g27023, g26344)
--	g27290 = NOR(g27024, g26348)
--	g27291 = NOR(g27025, g26350)
--	g27292 = NOR(g27026, g26351)
--	g27293 = NOR(g27027, g26357)
--	g27294 = NOR(g27028, g26361)
--	g27295 = NOR(g27029, g26362)
--	g27296 = NOR(g27030, g26363)
--	g27297 = NOR(g27031, g26365)
--	g27298 = NOR(g27032, g26366)
--	g27299 = NOR(g27033, g26371)
--	g27300 = NOR(g27034, g26372)
--	g27301 = NOR(g27035, g26373)
--	g27302 = NOR(g27042, g26379)
--	g27303 = NOR(g27043, g26380)
--	g27304 = NOR(g27044, g26381)
--	g27305 = NOR(g27045, g26383)
--	g27306 = NOR(g27046, g26384)
--	g27307 = NOR(g27047, g26386)
--	g27308 = NOR(g27048, g26387)
--	g27309 = NOR(g27049, g26388)
--	g27310 = NOR(g27050, g26392)
--	g27311 = NOR(g27053, g26396)
--	g27312 = NOR(g27054, g26397)
--	g27313 = NOR(g27055, g26400)
--	g27314 = NOR(g27056, g26404)
--	g27315 = NOR(g27057, g26405)
--	g27316 = NOR(g27058, g26406)
--	g27317 = NOR(g27059, g26408)
--	g27318 = NOR(g27060, g26409)
--	g27319 = NOR(g27061, g26414)
--	g27320 = NOR(g27062, g26415)
--	g27321 = NOR(g27063, g26416)
--	g27322 = NOR(g27070, g26422)
--	g27323 = NOR(g27071, g26423)
--	g27324 = NOR(g27072, g26424)
--	g27325 = NOR(g27073, g26426)
--	g27326 = NOR(g27074, g26427)
--	g27327 = NOR(g27077, g26432)
--	g27328 = NOR(g27080, g26437)
--	g27329 = NOR(g27081, g26438)
--	g27330 = NOR(g27082, g26441)
--	g27331 = NOR(g27083, g26445)
--	g27332 = NOR(g27084, g26446)
--	g27333 = NOR(g27085, g26447)
--	g27334 = NOR(g27086, g26449)
--	g27335 = NOR(g27087, g26450)
--	g27336 = NOR(g27088, g26455)
--	g27337 = NOR(g27089, g26456)
--	g27338 = NOR(g27090, g26457)
--	g27339 = NOR(g27093, g26464)
--	g27340 = NOR(g27096, g26469)
--	g27341 = NOR(g27097, g26470)
--	g27342 = NOR(g27098, g26473)
--	g27343 = NOR(g27099, g26477)
--	g27344 = NOR(g27100, g26478)
--	g27345 = NOR(g27101, g26479)
--	g27346 = NOR(g27105, g26488)
--	g27347 = NOR(g27108, g26493)
--	g27348 = NOR(g27109, g26494)
--	g27354 = NOR(g27112, g26504)
--	g27414 = NOR(g26770, g25187)
--	g27415 = NOR(g23104, g27181, g25128)
--	g27435 = NOR(g26777, g25193)
--	g27436 = NOR(g23118, g27187, g24427)
--	g27450 = NOR(g26902, g24613)
--	g27454 = NOR(g26783, g25196)
--	g27455 = NOR(g23127, g26758, g24431)
--	g27462 = NOR(g26892, g24622)
--	g27464 = NOR(g27178, g25975)
--	g27466 = NOR(g26915, g24624)
--	g27470 = NOR(g26790, g25198)
--	g27471 = NOR(g23138, g26764, g24435)
--	g27478 = NOR(g26754, g24432)
--	g27481 = NOR(g27182, g25980)
--	g27482 = NOR(g26906, g24637)
--	g27485 = NOR(g26928, g24638)
--	g27492 = NOR(g24958, g24633, g26771)
--	g27496 = NOR(g27185, g25178)
--	g27501 = NOR(g26763, g24436)
--	g27504 = NOR(g26918, g24656)
--	g27507 = NOR(g26941, g24657)
--	g27513 = NOR(g24969, g24653, g26778)
--	g27521 = NOR(g26766, g24439)
--	g27524 = NOR(g26931, g24675)
--	g27527 = NOR(g26759, g19087)
--	g27529 = NOR(g4456, g26873)
--	g27531 = NOR(g26760, g25181)
--	g27532 = NOR(g26761, g25182)
--	g27538 = NOR(g24982, g24672, g26784)
--	g27546 = NOR(g26769, g24441)
--	g27549 = NOR(g26765, g19093)
--	g27551 = NOR(g4632, g26882)
--	g27558 = NOR(g24993, g24691, g26791)
--	g27563 = NOR(g26922, g24708)
--	g27564 = NOR(g26767, g25184)
--	g27565 = NOR(g26768, g19100)
--	g27567 = NOR(g4809, g26891)
--	g27572 = NOR(g26911, g24717)
--	g27573 = NOR(g26773, g25188)
--	g27574 = NOR(g26935, g24720)
--	g27575 = NOR(g26774, g19107)
--	g27577 = NOR(g4985, g26901)
--	g27579 = NOR(g26775, g25192)
--	g27581 = NOR(g26925, g24728)
--	g27582 = NOR(g26944, g24731)
--	g27584 = NOR(g26938, g24736)
--	g27585 = NOR(g26950, g24739)
--	g27588 = NOR(g26947, g24742)
--	g27594 = NOR(g27175, g17001)
--	g27603 = NOR(g27179, g17031)
--	g27612 = NOR(g27184, g17065)
--	g27621 = NOR(g27188, g17100)
--	g27629 = NOR(g26829, g26051)
--	g27631 = NOR(g26833, g26053)
--	g27655 = NOR(g26842, g26061)
--	g27658 = NOR(g26851, g26068)
--	g27672 = NOR(g26799, g10024)
--	g27678 = NOR(g26800, g10133)
--	g27682 = NOR(g26801, g10238)
--	g27718 = NOR(g27251, g10133)
--	g27722 = NOR(g27252, g10238)
--	g27724 = NOR(g27254, g10340)
--	g27735 = NOR(g27394, g26961)
--	g27736 = NOR(g27396, g26962)
--	g27741 = NOR(g27407, g26966)
--	g27742 = NOR(g27409, g26967)
--	g27746 = NOR(g27425, g26972)
--	g27747 = NOR(g27427, g26973)
--	g27754 = NOR(g27446, g26985)
--	g27755 = NOR(g27448, g26986)
--	g27759 = NOR(g27495, g27052)
--	g27760 = NOR(g27509, g27076)
--	g27761 = NOR(g27516, g27079)
--	g27762 = NOR(g27530, g27091)
--	g27763 = NOR(g27534, g27092)
--	g27764 = NOR(g27541, g27095)
--	g27765 = NOR(g27552, g27103)
--	g27766 = NOR(g27554, g27104)
--	g27767 = NOR(g27561, g27107)
--	g27768 = NOR(g27568, g27110)
--	g27769 = NOR(g27570, g27111)
--	g27771 = NOR(g27578, g27115)
--	g27798 = NOR(g27632, g1223)
--	g27802 = NOR(g6087, g27632, g25330)
--	g27810 = NOR(g27632, g1215)
--	g27811 = NOR(g6087, g27632, g25404)
--	g27814 = NOR(g6087, g27632, g25322)
--	g27823 = NOR(g27632, g1216)
--	g27824 = NOR(g6087, g27632, g25399)
--	g27827 = NOR(g6087, g27632, g25314)
--	g27834 = NOR(g27478, g14630)
--	g27842 = NOR(g27632, g1217)
--	g27850 = NOR(g27501, g14650)
--	g27854 = NOR(g27632, g1218)
--	g27855 = NOR(g6087, g27632, g25385)
--	g27864 = NOR(g27632, g1219)
--	g27865 = NOR(g6087, g27632, g25370)
--	g27868 = NOR(g23742, g27632)
--	g27869 = NOR(g27632, g25437)
--	g27875 = NOR(g27521, g14677)
--	g27882 = NOR(g27632, g1220)
--	g27883 = NOR(g6087, g27632, g25361)
--	g27886 = NOR(g27632, g24627)
--	g27892 = NOR(g27546, g14711)
--	g27896 = NOR(g27632, g1222)
--	g27897 = NOR(g6087, g27632, g25349)
--	g27900 = NOR(g6087, g27632, g25338)
--	g27906 = NOR(g16127, g27656)
--	g27911 = NOR(g16170, g27657)
--	g27916 = NOR(g16219, g27659)
--	g27917 = NOR(g16220, g27660)
--	g27925 = NOR(g16276, g27661)
--	g27937 = NOR(g16321, g27666)
--	g27950 = NOR(g16367, g27673)
--	g27962 = NOR(g16394, g27679)
--	g27964 = NOR(g16400, g27680)
--	g27980 = NOR(g16428, g27681)
--	g27997 = NOR(g16456, g27242)
--	g28002 = NOR(g26032, g27246)
--	g28029 = NOR(g26033, g27247)
--	g28059 = NOR(g26034, g27248)
--	g28088 = NOR(g26036, g27249)
--	g28145 = NOR(g27629, g17001)
--	g28146 = NOR(g27631, g17031)
--	g28147 = NOR(g27655, g17065)
--	g28148 = NOR(g27658, g17100)
--	g28157 = NOR(g13902, g27370)
--	g28185 = NOR(g27356, g26845)
--	g28189 = NOR(g27359, g26853)
--	g28191 = NOR(g27365, g26860)
--	g28192 = NOR(g27372, g26866)
--	g28199 = NOR(g27250, g10024)
--	g28321 = NOR(g27742, g10133)
--	g28325 = NOR(g27747, g10238)
--	g28328 = NOR(g27755, g10340)
--	g28342 = NOR(g15460, g28008)
--	g28344 = NOR(g15526, g28027)
--	g28345 = NOR(g15527, g28028)
--	g28346 = NOR(g15546, g28035)
--	g28348 = NOR(g15594, g28050)
--	g28349 = NOR(g15595, g28051)
--	g28350 = NOR(g15604, g28057)
--	g28351 = NOR(g15605, g28058)
--	g28352 = NOR(g15624, g28065)
--	g28353 = NOR(g15666, g28073)
--	g28354 = NOR(g15670, g28079)
--	g28355 = NOR(g15671, g28080)
--	g28356 = NOR(g15680, g28086)
--	g28357 = NOR(g15681, g28087)
--	g28358 = NOR(g15700, g28094)
--	g28360 = NOR(g15725, g28098)
--	g28361 = NOR(g15729, g28104)
--	g28362 = NOR(g15730, g28105)
--	g28363 = NOR(g15739, g28111)
--	g28364 = NOR(g15740, g28112)
--	g28366 = NOR(g15765, g28116)
--	g28367 = NOR(g15769, g28122)
--	g28368 = NOR(g15770, g28123)
--	g28371 = NOR(g15793, g28127)
--	g28392 = NOR(g27886, g22344)
--	g28394 = NOR(g27869, g22344)
--	g28397 = NOR(g27869, g22344)
--	g28400 = NOR(g27886, g22344)
--	g28403 = NOR(g27811, g22344)
--	g28406 = NOR(g27824, g22344)
--	g28409 = NOR(g24676, g27801)
--	g28410 = NOR(g27748, g22344)
--	g28413 = NOR(g24695, g27809)
--	g28414 = NOR(g27748, g22344)
--	g28417 = NOR(g24712, g27830)
--	g28418 = NOR(g24723, g27846)
--	g28420 = NOR(g16031, g28171)
--	g28421 = NOR(g16068, g28176)
--	g28425 = NOR(g16133, g28188)
--	g28449 = NOR(g27727, g26780)
--	g28461 = NOR(g27729, g26787)
--	g28470 = NOR(g27671, g28193)
--	g28473 = NOR(g27730, g26794)
--	g28482 = NOR(g27731, g26797)
--	g28488 = NOR(g26755, g27719)
--	g28489 = NOR(g26756, g27720)
--	g28490 = NOR(g27240, g27721)
--	g28495 = NOR(g27244, g27723)
--	g28499 = NOR(g26027, g27725)
--	g28523 = NOR(g26035, g27732)
--	g28525 = NOR(g27245, g27726)
--	g28528 = NOR(g26030, g27728)
--	g28551 = NOR(g26038, g27733)
--	g28578 = NOR(g26039, g27734)
--	g28606 = NOR(g26040, g27737)
--	g28634 = NOR(g28185, g17001)
--	g28635 = NOR(g28189, g17031)
--	g28636 = NOR(g28191, g17065)
--	g28637 = NOR(g28192, g17100)
--	g28654 = NOR(g27770, g27355)
--	g28656 = NOR(g27772, g27358)
--	g28658 = NOR(g27773, g27364)
--	g28661 = NOR(g27775, g27371)
--	g28668 = NOR(g27736, g10024)
--	g28728 = NOR(g28422, g27904)
--	g28731 = NOR(g28423, g27908)
--	g28732 = NOR(g14894, g28426)
--	g28733 = NOR(g28424, g27909)
--	g28735 = NOR(g14957, g28430)
--	g28736 = NOR(g28427, g27913)
--	g28737 = NOR(g28428, g27914)
--	g28738 = NOR(g14975, g28433)
--	g28739 = NOR(g28429, g27915)
--	g28744 = NOR(g15030, g28439)
--	g28745 = NOR(g28431, g27922)
--	g28746 = NOR(g15046, g28441)
--	g28747 = NOR(g28434, g27923)
--	g28748 = NOR(g28435, g27924)
--	g28749 = NOR(g15064, g28444)
--	g28750 = NOR(g28436, g27926)
--	g28754 = NOR(g28440, g27931)
--	g28758 = NOR(g15126, g28451)
--	g28759 = NOR(g28442, g27935)
--	g28760 = NOR(g15142, g28453)
--	g28761 = NOR(g28445, g27936)
--	g28762 = NOR(g28446, g27938)
--	g28763 = NOR(g15160, g28456)
--	g28767 = NOR(g28452, g27945)
--	g28771 = NOR(g15218, g28463)
--	g28772 = NOR(g28454, g27949)
--	g28773 = NOR(g15234, g28465)
--	g28774 = NOR(g28457, g27951)
--	g28778 = NOR(g28464, g27963)
--	g28782 = NOR(g15304, g28475)
--	g28783 = NOR(g28466, g27968)
--	g28784 = NOR(g28468, g27970)
--	g28788 = NOR(g28476, g27984)
--	g28789 = NOR(g28477, g27985)
--	g28790 = NOR(g28478, g27991)
--	g28794 = NOR(g28484, g28009)
--	g28795 = NOR(g28485, g28015)
--	g28802 = NOR(g28492, g28036)
--	g28803 = NOR(g28493, g28042)
--	g28813 = NOR(g28497, g28066)
--	g28874 = NOR(g28657, g16221)
--	g28886 = NOR(g28659, g16277)
--	g28903 = NOR(g28660, g13295)
--	g28920 = NOR(g28662, g13322)
--	g28941 = NOR(g28663, g13343)
--	g28954 = NOR(g26673, g27241, g28323)
--	g28963 = NOR(g28664, g13365)
--	g28982 = NOR(g28665, g28670)
--	g28987 = NOR(g28666, g13390)
--	g28990 = NOR(g28667, g16457)
--	g29009 = NOR(g28669, g28320)
--	g29013 = NOR(g28671, g11607)
--	g29016 = NOR(g28672, g13487)
--	g29031 = NOR(g28319, g28324)
--	g29039 = NOR(g28322, g13500)
--	g29063 = NOR(g28326, g28329)
--	g29064 = NOR(g28327, g28330)
--	g29083 = NOR(g28331, g28333)
--	g29090 = NOR(g28332, g28334)
--	g29097 = NOR(g28335, g28336)
--	g29109 = NOR(g28654, g17001)
--	g29110 = NOR(g28656, g17031)
--	g29111 = NOR(g28658, g17065)
--	g29112 = NOR(g28661, g17100)
--	g29113 = NOR(g28381, g8907)
--	g29126 = NOR(g28373, g27774)
--	g29127 = NOR(g28376, g27779)
--	g29128 = NOR(g28380, g27783)
--	g29129 = NOR(g28385, g27790)
--	g29167 = NOR(g28841, g28396)
--	g29169 = NOR(g28843, g28398)
--	g29170 = NOR(g28844, g28399)
--	g29172 = NOR(g28846, g28401)
--	g29173 = NOR(g28847, g28402)
--	g29178 = NOR(g28848, g28404)
--	g29179 = NOR(g28849, g28405)
--	g29181 = NOR(g28850, g28407)
--	g29182 = NOR(g28851, g28408)
--	g29184 = NOR(g28852, g28411)
--	g29185 = NOR(g28853, g28412)
--	g29187 = NOR(g28854, g28416)
--	g29194 = NOR(g14958, g28881)
--	g29195 = NOR(g28880, g28438)
--	g29197 = NOR(g15031, g28893)
--	g29198 = NOR(g15047, g28898)
--	g29199 = NOR(g28892, g28448)
--	g29201 = NOR(g15104, g28910)
--	g29202 = NOR(g28897, g28450)
--	g29204 = NOR(g15127, g28915)
--	g29205 = NOR(g15143, g28923)
--	g29206 = NOR(g28909, g28459)
--	g29207 = NOR(g28914, g28460)
--	g29209 = NOR(g15196, g28936)
--	g29210 = NOR(g28919, g28462)
--	g29212 = NOR(g15219, g28944)
--	g29213 = NOR(g15235, g28949)
--	g29214 = NOR(g28931, g28469)
--	g29215 = NOR(g28935, g28471)
--	g29216 = NOR(g28940, g28472)
--	g29218 = NOR(g15282, g28966)
--	g29219 = NOR(g28948, g28474)
--	g29221 = NOR(g15305, g28971)
--	g29222 = NOR(g28958, g28479)
--	g29223 = NOR(g28962, g28480)
--	g29224 = NOR(g28970, g28481)
--	g29226 = NOR(g15374, g28997)
--	g29227 = NOR(g28986, g28486)
--	g29228 = NOR(g28996, g28487)
--	g29231 = NOR(g29022, g28494)
--	g29303 = NOR(g28716, g19112)
--	g29313 = NOR(g28717, g19117)
--	g29324 = NOR(g28718, g19124)
--	g29333 = NOR(g28719, g19131)
--	g29340 = NOR(g28337, g28722)
--	g29343 = NOR(g28338, g28724)
--	g29345 = NOR(g28339, g28726)
--	g29347 = NOR(g28340, g28729)
--	g29353 = NOR(g29126, g17001)
--	g29354 = NOR(g29127, g17031)
--	g29355 = NOR(g29128, g17065)
--	g29357 = NOR(g29129, g17100)
--	g29399 = NOR(g28834, g28378)
--	g29403 = NOR(g28836, g28383)
--	g29406 = NOR(g28838, g28387)
--	g29409 = NOR(g28840, g28389)
--	g29552 = NOR(g29130, g29411)
--	g29569 = NOR(g28708, g29174)
--	g29570 = NOR(g28709, g29175)
--	g29571 = NOR(g28710, g29176)
--	g29574 = NOR(g28712, g29180)
--	g29576 = NOR(g28713, g29183)
--	g29577 = NOR(g28714, g29186)
--	g29578 = NOR(g28715, g29188)
--	g29579 = NOR(g29399, g17001)
--	g29580 = NOR(g29403, g17031)
--	g29581 = NOR(g29406, g17065)
--	g29582 = NOR(g29409, g17100)
--	g29606 = NOR(g13878, g29248)
--	g29608 = NOR(g13892, g29251)
--	g29609 = NOR(g13900, g29252)
--	g29611 = NOR(g13913, g29255)
--	g29612 = NOR(g13933, g29256)
--	g29613 = NOR(g13941, g29257)
--	g29616 = NOR(g13969, g29259)
--	g29617 = NOR(g13989, g29260)
--	g29618 = NOR(g13997, g29261)
--	g29620 = NOR(g14039, g29262)
--	g29621 = NOR(g14059, g29263)
--	g29623 = NOR(g14130, g29264)
--	g29663 = NOR(g29518, g29284)
--	g29665 = NOR(g29521, g29289)
--	g29667 = NOR(g29524, g29294)
--	g29669 = NOR(g29528, g29300)
--	g29670 = NOR(g29529, g29302)
--	g29671 = NOR(g29534, g29310)
--	g29672 = NOR(g29536, g29312)
--	g29676 = NOR(g29540, g29320)
--	g29677 = NOR(g29543, g29321)
--	g29678 = NOR(g29545, g29323)
--	g29679 = NOR(g29549, g29329)
--	g29680 = NOR(g29553, g29330)
--	g29681 = NOR(g29555, g29332)
--	g29682 = NOR(g29557, g29336)
--	g29683 = NOR(g29559, g29337)
--	g29684 = NOR(g29562, g29338)
--	g29685 = NOR(g29564, g29341)
--	g29686 = NOR(g29566, g29342)
--	g29687 = NOR(g29572, g29344)
--	g29688 = NOR(g29575, g29346)
--	g29703 = NOR(g29583, g1917)
--	g29705 = NOR(g6104, g29583, g25339)
--	g29709 = NOR(g29583, g1909)
--	g29710 = NOR(g6104, g29583, g25412)
--	g29713 = NOR(g6104, g29583, g25332)
--	g29717 = NOR(g29583, g1910)
--	g29718 = NOR(g6104, g29583, g25409)
--	g29721 = NOR(g6104, g29583, g25323)
--	g29725 = NOR(g29583, g1911)
--	g29727 = NOR(g29583, g1912)
--	g29728 = NOR(g6104, g29583, g25401)
--	g29731 = NOR(g29583, g1913)
--	g29732 = NOR(g6104, g29583, g25387)
--	g29735 = NOR(g23797, g29583)
--	g29736 = NOR(g29583, g25444)
--	g29740 = NOR(g29583, g1914)
--	g29741 = NOR(g6104, g29583, g25376)
--	g29744 = NOR(g29583, g24641)
--	g29747 = NOR(g29583, g1916)
--	g29748 = NOR(g6104, g29583, g25363)
--	g29751 = NOR(g6104, g29583, g25352)
--	g29754 = NOR(g16178, g29607)
--	g29755 = NOR(g16229, g29610)
--	g29756 = NOR(g16284, g29614)
--	g29757 = NOR(g16285, g29615)
--	g29758 = NOR(g16335, g29619)
--	g29759 = NOR(g16379, g29622)
--	g29760 = NOR(g16411, g29624)
--	g29761 = NOR(g28707, g28711, g29466)
--	g29762 = NOR(g16432, g29625)
--	g29763 = NOR(g16438, g29626)
--	g29764 = NOR(g16462, g29464)
--	g29765 = NOR(g13492, g29465)
--	g29766 = NOR(g29467, g19142)
--	g29767 = NOR(g29468, g19143)
--	g29768 = NOR(g29469, g19146)
--	g29769 = NOR(g29470, g19148)
--	g29770 = NOR(g29471, g29196)
--	g29771 = NOR(g29472, g29200)
--	g29772 = NOR(g29473, g29203)
--	g29773 = NOR(g29474, g29208)
--	g29774 = NOR(g29475, g29211)
--	g29775 = NOR(g29476, g29217)
--	g29776 = NOR(g29477, g29220)
--	g29777 = NOR(g29478, g29225)
--	g29778 = NOR(g29479, g29229)
--	g29779 = NOR(g13943, g29502)
--	g29780 = NOR(g29480, g29232)
--	g29781 = NOR(g29481, g29233)
--	g29782 = NOR(g29482, g29234)
--	g29783 = NOR(g29483, g29235)
--	g29784 = NOR(g29484, g29236)
--	g29785 = NOR(g29485, g29238)
--	g29786 = NOR(g29486, g29239)
--	g29787 = NOR(g29487, g29240)
--	g29788 = NOR(g29488, g29241)
--	g29789 = NOR(g29489, g29242)
--	g29791 = NOR(g29490, g29243)
--	g29912 = NOR(g24676, g29716)
--	g29914 = NOR(g24695, g29724)
--	g29916 = NOR(g24712, g29726)
--	g29918 = NOR(g29744, g22367)
--	g29919 = NOR(g29736, g22367)
--	g29920 = NOR(g24723, g29739)
--	g29921 = NOR(g29736, g22367)
--	g29922 = NOR(g29744, g22367)
--	g29924 = NOR(g29710, g22367)
--	g29926 = NOR(g29718, g22367)
--	g29928 = NOR(g29673, g22367)
--	g29929 = NOR(g29673, g22367)
--	g29936 = NOR(g16049, g29790)
--	g29939 = NOR(g16102, g29792)
--	g29941 = NOR(g16182, g29793)
--	g30010 = NOR(g29520, g29942)
--	g30011 = NOR(g29522, g29944)
--	g30012 = NOR(g29523, g29945)
--	g30013 = NOR(g29525, g29946)
--	g30014 = NOR(g29526, g29947)
--	g30015 = NOR(g29527, g29948)
--	g30016 = NOR(g29531, g29949)
--	g30017 = NOR(g29532, g29950)
--	g30018 = NOR(g29533, g29951)
--	g30019 = NOR(g29538, g29952)
--	g30020 = NOR(g29539, g29953)
--	g30021 = NOR(g29541, g29954)
--	g30022 = NOR(g29547, g29955)
--	g30023 = NOR(g29548, g29956)
--	g30024 = NOR(g29550, g29957)
--	g30025 = NOR(g29558, g29958)
--	g30026 = NOR(g29560, g29959)
--	g30027 = NOR(g29565, g29960)
--	g30028 = NOR(g29567, g29961)
--	g30029 = NOR(g29573, g29962)
--	g30030 = NOR(g24676, g29923)
--	g30031 = NOR(g24695, g29925)
--	g30032 = NOR(g24712, g29927)
--	g30033 = NOR(g24723, g29931)
--	g30053 = NOR(g29963, g16286)
--	g30054 = NOR(g29964, g16336)
--	g30055 = NOR(g29965, g13326)
--	g30056 = NOR(g29966, g13345)
--	g30057 = NOR(g29967, g13368)
--	g30058 = NOR(g29968, g13395)
--	g30059 = NOR(g29969, g29811)
--	g30060 = NOR(g29970, g11612)
--	g30061 = NOR(g29971, g13493)
--	g30062 = NOR(g29810, g29815)
--	g30063 = NOR(g29812, g11637)
--	g30064 = NOR(g29813, g13506)
--	g30065 = NOR(g29814, g29817)
--	g30066 = NOR(g29816, g13517)
--	g30067 = NOR(g29818, g29820)
--	g30068 = NOR(g29819, g29821)
--	g30069 = NOR(g29822, g29828)
--	g30070 = NOR(g29827, g29833)
--	g30071 = NOR(g29834, g29839)
--	g30072 = NOR(g29910, g8947)
--	g30245 = NOR(g16074, g30077)
--	g30246 = NOR(g16107, g30079)
--	g30247 = NOR(g16112, g30080)
--	g30248 = NOR(g16139, g30081)
--	g30249 = NOR(g16158, g30082)
--	g30250 = NOR(g16163, g30083)
--	g30251 = NOR(g16198, g30085)
--	g30252 = NOR(g16217, g30086)
--	g30253 = NOR(g16222, g30087)
--	g30254 = NOR(g16242, g30088)
--	g30255 = NOR(g16263, g30089)
--	g30256 = NOR(g16282, g30090)
--	g30257 = NOR(g16290, g30091)
--	g30258 = NOR(g16291, g30092)
--	g30259 = NOR(g16301, g30093)
--	g30260 = NOR(g16322, g30094)
--	g30261 = NOR(g16342, g30095)
--	g30262 = NOR(g16343, g30096)
--	g30263 = NOR(g16344, g30097)
--	g30264 = NOR(g16348, g30098)
--	g30265 = NOR(g16349, g30099)
--	g30266 = NOR(g16359, g30100)
--	g30267 = NOR(g16380, g30101)
--	g30268 = NOR(g16382, g30102)
--	g30269 = NOR(g16386, g30103)
--	g30270 = NOR(g16387, g30104)
--	g30271 = NOR(g16388, g30105)
--	g30272 = NOR(g16392, g30106)
--	g30273 = NOR(g16393, g30107)
--	g30274 = NOR(g16403, g30108)
--	g30275 = NOR(g16413, g30109)
--	g30276 = NOR(g16415, g30110)
--	g30277 = NOR(g16418, g30111)
--	g30278 = NOR(g16420, g30112)
--	g30279 = NOR(g16424, g30113)
--	g30280 = NOR(g16425, g30114)
--	g30281 = NOR(g16426, g30115)
--	g30282 = NOR(g16430, g30117)
--	g30283 = NOR(g16431, g30118)
--	g30284 = NOR(g16444, g29980)
--	g30285 = NOR(g16447, g29981)
--	g30286 = NOR(g16449, g29982)
--	g30287 = NOR(g16452, g29983)
--	g30288 = NOR(g16454, g29984)
--	g30289 = NOR(g16458, g29985)
--	g30290 = NOR(g16459, g29986)
--	g30291 = NOR(g16460, g29987)
--	g30292 = NOR(g13477, g29988)
--	g30293 = NOR(g13480, g29989)
--	g30294 = NOR(g13483, g29990)
--	g30295 = NOR(g13485, g29991)
--	g30296 = NOR(g13488, g29993)
--	g30297 = NOR(g13490, g29994)
--	g30298 = NOR(g13496, g29995)
--	g30299 = NOR(g13499, g29996)
--	g30300 = NOR(g13502, g30001)
--	g30301 = NOR(g13504, g30002)
--	g30302 = NOR(g13513, g30003)
--	g30303 = NOR(g13516, g30005)
--	g30304 = NOR(g13527, g30007)
--	g30338 = NOR(g14297, g30225)
--	g30341 = NOR(g14328, g30226)
--	g30356 = NOR(g14419, g30227)
--	g30399 = NOR(g30116, g30123)
--	g30400 = NOR(g29997, g30127)
--	g30401 = NOR(g29998, g30128)
--	g30402 = NOR(g29999, g30129)
--	g30403 = NOR(g30004, g30131)
--	g30404 = NOR(g30006, g30132)
--	g30405 = NOR(g30008, g30133)
--	g30406 = NOR(g30009, g30138)
--	g30455 = NOR(g13953, g30216)
--	g30468 = NOR(g14007, g30217)
--	g30470 = NOR(g14023, g30218)
--	g30482 = NOR(g14067, g30219)
--	g30485 = NOR(g14098, g30220)
--	g30487 = NOR(g14114, g30221)
--	g30500 = NOR(g14182, g30222)
--	g30503 = NOR(g14213, g30223)
--	g30505 = NOR(g14229, g30224)
--	g30566 = NOR(g14327, g30398)
--	g30584 = NOR(g30412, g2611)
--	g30588 = NOR(g6119, g30412, g25353)
--	g30593 = NOR(g30412, g2603)
--	g30594 = NOR(g6119, g30412, g25419)
--	g30597 = NOR(g6119, g30412, g25341)
--	g30601 = NOR(g30412, g2604)
--	g30602 = NOR(g6119, g30412, g25417)
--	g30605 = NOR(g6119, g30412, g25333)
--	g30608 = NOR(g30412, g2605)
--	g30609 = NOR(g30412, g2606)
--	g30610 = NOR(g6119, g30412, g25411)
--	g30613 = NOR(g30412, g2607)
--	g30614 = NOR(g6119, g30412, g25403)
--	g30617 = NOR(g23850, g30412)
--	g30618 = NOR(g30412, g25449)
--	g30621 = NOR(g30412, g2608)
--	g30622 = NOR(g6119, g30412, g25393)
--	g30625 = NOR(g30412, g24660)
--	g30628 = NOR(g30412, g2610)
--	g30629 = NOR(g6119, g30412, g25378)
--	g30632 = NOR(g6119, g30412, g25366)
--	g30635 = NOR(g16108, g30407)
--	g30636 = NOR(g16140, g30409)
--	g30637 = NOR(g16141, g30410)
--	g30638 = NOR(g16159, g30411)
--	g30639 = NOR(g16186, g30436)
--	g30640 = NOR(g16187, g30437)
--	g30641 = NOR(g16188, g30438)
--	g30642 = NOR(g16199, g30440)
--	g30643 = NOR(g16200, g30441)
--	g30644 = NOR(g16218, g30442)
--	g30645 = NOR(g16240, g30444)
--	g30646 = NOR(g16241, g30445)
--	g30647 = NOR(g16251, g30447)
--	g30648 = NOR(g16252, g30448)
--	g30649 = NOR(g16253, g30449)
--	g30650 = NOR(g16264, g30451)
--	g30651 = NOR(g16265, g30452)
--	g30652 = NOR(g16283, g30453)
--	g30653 = NOR(g16289, g30454)
--	g30654 = NOR(g16299, g30457)
--	g30655 = NOR(g16300, g30458)
--	g30656 = NOR(g16310, g30460)
--	g30657 = NOR(g16311, g30461)
--	g30658 = NOR(g16312, g30462)
--	g30659 = NOR(g16323, g30464)
--	g30660 = NOR(g16324, g30465)
--	g30661 = NOR(g16345, g30467)
--	g30662 = NOR(g16347, g30469)
--	g30663 = NOR(g16357, g30472)
--	g30664 = NOR(g16358, g30473)
--	g30665 = NOR(g16368, g30475)
--	g30666 = NOR(g16369, g30476)
--	g30667 = NOR(g16370, g30477)
--	g30668 = NOR(g16381, g30478)
--	g30669 = NOR(g16383, g30481)
--	g30670 = NOR(g16389, g30484)
--	g30671 = NOR(g16391, g30486)
--	g30672 = NOR(g16401, g30489)
--	g30673 = NOR(g16402, g30490)
--	g30674 = NOR(g16414, g30492)
--	g30675 = NOR(g16416, g30495)
--	g30676 = NOR(g16419, g30496)
--	g30677 = NOR(g16421, g30499)
--	g30678 = NOR(g16427, g30502)
--	g30679 = NOR(g16429, g30504)
--	g30680 = NOR(g16443, g30327)
--	g30681 = NOR(g16448, g30330)
--	g30682 = NOR(g16450, g30333)
--	g30683 = NOR(g16453, g30334)
--	g30684 = NOR(g16455, g30337)
--	g30685 = NOR(g29992, g30000, g30372)
--	g30686 = NOR(g16461, g30340)
--	g30687 = NOR(g13479, g30345)
--	g30688 = NOR(g13484, g30348)
--	g30689 = NOR(g13486, g30351)
--	g30690 = NOR(g13489, g30352)
--	g30691 = NOR(g13491, g30355)
--	g30692 = NOR(g13498, g30361)
--	g30693 = NOR(g13503, g30364)
--	g30694 = NOR(g13505, g30367)
--	g30695 = NOR(g13515, g30374)
--	g30699 = NOR(g13914, g30387)
--	g30700 = NOR(g13952, g30388)
--	g30701 = NOR(g13970, g30389)
--	g30702 = NOR(g14006, g30390)
--	g30703 = NOR(g14022, g30391)
--	g30704 = NOR(g14040, g30392)
--	g30705 = NOR(g14097, g30393)
--	g30706 = NOR(g14113, g30394)
--	g30707 = NOR(g14131, g30395)
--	g30708 = NOR(g14212, g30396)
--	g30709 = NOR(g14228, g30397)
--	g30780 = NOR(g30625, g22387)
--	g30783 = NOR(g30618, g22387)
--	g30785 = NOR(g30618, g22387)
--	g30786 = NOR(g30625, g22387)
--	g30787 = NOR(g30594, g22387)
--	g30788 = NOR(g30602, g22387)
--	g30789 = NOR(g30575, g22387)
--	g30790 = NOR(g30575, g22387)
--	g30796 = NOR(g16069, g30696)
--	g30798 = NOR(g16134, g30697)
--	g30801 = NOR(g16237, g30698)
--	g30929 = NOR(g30728, g30736)
--	g30930 = NOR(g30735, g30744)
--	g30931 = NOR(g30743, g30750)
--	g30932 = NOR(g30754, g30757)
--	g30933 = NOR(g30755, g30758)
--	g30934 = NOR(g30759, g30761)
--	g30935 = NOR(g30760, g30762)
--	g30936 = NOR(g30763, g30764)
--	g30954 = NOR(g30916, g30944)
--	g30955 = NOR(g30918, g30945)
--	g30956 = NOR(g30919, g30946)
--	g30957 = NOR(g30920, g30947)
--	g30958 = NOR(g30922, g30948)
--	g30959 = NOR(g30923, g30949)
--	g30960 = NOR(g30924, g30950)
--	g30961 = NOR(g30925, g30951)
--	g30970 = NOR(g30917, g30921, g30953)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s38417 is
	port (
		CLK: in std_logic;
		G51: in std_logic;
		G563: in std_logic;
		G1249: in std_logic;
		G1943: in std_logic;
		G2637: in std_logic;
		G3212: in std_logic;
		G3213: in std_logic;
		G3214: in std_logic;
		G3215: in std_logic;
		G3216: in std_logic;
		G3217: in std_logic;
		G3218: in std_logic;
		G3219: in std_logic;
		G3220: in std_logic;
		G3221: in std_logic;
		G3222: in std_logic;
		G3223: in std_logic;
		G3224: in std_logic;
		G3225: in std_logic;
		G3226: in std_logic;
		G3227: in std_logic;
		G3228: in std_logic;
		G3229: in std_logic;
		G3230: in std_logic;
		G3231: in std_logic;
		G3232: in std_logic;
		G3233: in std_logic;
		G3234: in std_logic;
		G3993: out std_logic;
		G4088: out std_logic;
		G4090: out std_logic;
		G4200: out std_logic;
		G4321: out std_logic;
		G4323: out std_logic;
		G4450: out std_logic;
		G4590: out std_logic;
		G5388: out std_logic;
		G5437: out std_logic;
		G5472: out std_logic;
		G5511: out std_logic;
		G5549: out std_logic;
		G5555: out std_logic;
		G5595: out std_logic;
		G5612: out std_logic;
		G5629: out std_logic;
		G5637: out std_logic;
		G5648: out std_logic;
		G5657: out std_logic;
		G5686: out std_logic;
		G5695: out std_logic;
		G5738: out std_logic;
		G5747: out std_logic;
		G5796: out std_logic;
		G6225: out std_logic;
		G6231: out std_logic;
		G6313: out std_logic;
		G6368: out std_logic;
		G6442: out std_logic;
		G6447: out std_logic;
		G6485: out std_logic;
		G6518: out std_logic;
		G6573: out std_logic;
		G6642: out std_logic;
		G6677: out std_logic;
		G6712: out std_logic;
		G6750: out std_logic;
		G6782: out std_logic;
		G6837: out std_logic;
		G6895: out std_logic;
		G6911: out std_logic;
		G6944: out std_logic;
		G6979: out std_logic;
		G7014: out std_logic;
		G7052: out std_logic;
		G7084: out std_logic;
		G7161: out std_logic;
		G7194: out std_logic;
		G7229: out std_logic;
		G7264: out std_logic;
		G7302: out std_logic;
		G7334: out std_logic;
		G7357: out std_logic;
		G7390: out std_logic;
		G7425: out std_logic;
		G7487: out std_logic;
		G7519: out std_logic;
		G7909: out std_logic;
		G7956: out std_logic;
		G7961: out std_logic;
		G8007: out std_logic;
		G8012: out std_logic;
		G8021: out std_logic;
		G8023: out std_logic;
		G8030: out std_logic;
		G8082: out std_logic;
		G8087: out std_logic;
		G8096: out std_logic;
		G8106: out std_logic;
		G8167: out std_logic;
		G8175: out std_logic;
		G8249: out std_logic;
		G8251: out std_logic;
		G8258: out std_logic;
		G8259: out std_logic;
		G8260: out std_logic;
		G8261: out std_logic;
		G8262: out std_logic;
		G8263: out std_logic;
		G8264: out std_logic;
		G8265: out std_logic;
		G8266: out std_logic;
		G8267: out std_logic;
		G8268: out std_logic;
		G8269: out std_logic;
		G8270: out std_logic;
		G8271: out std_logic;
		G8272: out std_logic;
		G8273: out std_logic;
		G8274: out std_logic;
		G8275: out std_logic;
		G16297: out std_logic;
		G16355: out std_logic;
		G16399: out std_logic;
		G16437: out std_logic;
		G16496: out std_logic;
		G24734: out std_logic;
		G25420: out std_logic;
		G25435: out std_logic;
		G25442: out std_logic;
		G25489: out std_logic;
		G26104: out std_logic;
		G26135: out std_logic;
		G26149: out std_logic;
		G27380: out std_logic
	);
end entity;

architecture RTL of s38417 is
	attribute dont_touch: boolean;

	signal G1: std_logic; attribute dont_touch of G1: signal is true;
	signal G2: std_logic; attribute dont_touch of G2: signal is true;
	signal G5: std_logic; attribute dont_touch of G5: signal is true;
	signal G8: std_logic; attribute dont_touch of G8: signal is true;
	signal G11: std_logic; attribute dont_touch of G11: signal is true;
	signal G14: std_logic; attribute dont_touch of G14: signal is true;
	signal G17: std_logic; attribute dont_touch of G17: signal is true;
	signal G20: std_logic; attribute dont_touch of G20: signal is true;
	signal G23: std_logic; attribute dont_touch of G23: signal is true;
	signal G26: std_logic; attribute dont_touch of G26: signal is true;
	signal G27: std_logic; attribute dont_touch of G27: signal is true;
	signal G30: std_logic; attribute dont_touch of G30: signal is true;
	signal G33: std_logic; attribute dont_touch of G33: signal is true;
	signal G36: std_logic; attribute dont_touch of G36: signal is true;
	signal G39: std_logic; attribute dont_touch of G39: signal is true;
	signal G42: std_logic; attribute dont_touch of G42: signal is true;
	signal G45: std_logic; attribute dont_touch of G45: signal is true;
	signal G48: std_logic; attribute dont_touch of G48: signal is true;
	signal G52: std_logic; attribute dont_touch of G52: signal is true;
	signal G56: std_logic; attribute dont_touch of G56: signal is true;
	signal G61: std_logic; attribute dont_touch of G61: signal is true;
	signal G65: std_logic; attribute dont_touch of G65: signal is true;
	signal G70: std_logic; attribute dont_touch of G70: signal is true;
	signal G74: std_logic; attribute dont_touch of G74: signal is true;
	signal G79: std_logic; attribute dont_touch of G79: signal is true;
	signal G83: std_logic; attribute dont_touch of G83: signal is true;
	signal G88: std_logic; attribute dont_touch of G88: signal is true;
	signal G92: std_logic; attribute dont_touch of G92: signal is true;
	signal G97: std_logic; attribute dont_touch of G97: signal is true;
	signal G101: std_logic; attribute dont_touch of G101: signal is true;
	signal G105: std_logic; attribute dont_touch of G105: signal is true;
	signal G109: std_logic; attribute dont_touch of G109: signal is true;
	signal G113: std_logic; attribute dont_touch of G113: signal is true;
	signal G117: std_logic; attribute dont_touch of G117: signal is true;
	signal G121: std_logic; attribute dont_touch of G121: signal is true;
	signal G125: std_logic; attribute dont_touch of G125: signal is true;
	signal G129: std_logic; attribute dont_touch of G129: signal is true;
	signal G130: std_logic; attribute dont_touch of G130: signal is true;
	signal G131: std_logic; attribute dont_touch of G131: signal is true;
	signal G132: std_logic; attribute dont_touch of G132: signal is true;
	signal G133: std_logic; attribute dont_touch of G133: signal is true;
	signal G134: std_logic; attribute dont_touch of G134: signal is true;
	signal G135: std_logic; attribute dont_touch of G135: signal is true;
	signal G138: std_logic; attribute dont_touch of G138: signal is true;
	signal G141: std_logic; attribute dont_touch of G141: signal is true;
	signal G142: std_logic; attribute dont_touch of G142: signal is true;
	signal G143: std_logic; attribute dont_touch of G143: signal is true;
	signal G144: std_logic; attribute dont_touch of G144: signal is true;
	signal G145: std_logic; attribute dont_touch of G145: signal is true;
	signal G146: std_logic; attribute dont_touch of G146: signal is true;
	signal G147: std_logic; attribute dont_touch of G147: signal is true;
	signal G148: std_logic; attribute dont_touch of G148: signal is true;
	signal G149: std_logic; attribute dont_touch of G149: signal is true;
	signal G150: std_logic; attribute dont_touch of G150: signal is true;
	signal G151: std_logic; attribute dont_touch of G151: signal is true;
	signal G152: std_logic; attribute dont_touch of G152: signal is true;
	signal G153: std_logic; attribute dont_touch of G153: signal is true;
	signal G154: std_logic; attribute dont_touch of G154: signal is true;
	signal G155: std_logic; attribute dont_touch of G155: signal is true;
	signal G156: std_logic; attribute dont_touch of G156: signal is true;
	signal G157: std_logic; attribute dont_touch of G157: signal is true;
	signal G158: std_logic; attribute dont_touch of G158: signal is true;
	signal G159: std_logic; attribute dont_touch of G159: signal is true;
	signal G160: std_logic; attribute dont_touch of G160: signal is true;
	signal G161: std_logic; attribute dont_touch of G161: signal is true;
	signal G162: std_logic; attribute dont_touch of G162: signal is true;
	signal G163: std_logic; attribute dont_touch of G163: signal is true;
	signal G164: std_logic; attribute dont_touch of G164: signal is true;
	signal G165: std_logic; attribute dont_touch of G165: signal is true;
	signal G168: std_logic; attribute dont_touch of G168: signal is true;
	signal G169: std_logic; attribute dont_touch of G169: signal is true;
	signal G170: std_logic; attribute dont_touch of G170: signal is true;
	signal G171: std_logic; attribute dont_touch of G171: signal is true;
	signal G172: std_logic; attribute dont_touch of G172: signal is true;
	signal G173: std_logic; attribute dont_touch of G173: signal is true;
	signal G174: std_logic; attribute dont_touch of G174: signal is true;
	signal G175: std_logic; attribute dont_touch of G175: signal is true;
	signal G176: std_logic; attribute dont_touch of G176: signal is true;
	signal G177: std_logic; attribute dont_touch of G177: signal is true;
	signal G178: std_logic; attribute dont_touch of G178: signal is true;
	signal G179: std_logic; attribute dont_touch of G179: signal is true;
	signal G180: std_logic; attribute dont_touch of G180: signal is true;
	signal G181: std_logic; attribute dont_touch of G181: signal is true;
	signal G182: std_logic; attribute dont_touch of G182: signal is true;
	signal G185: std_logic; attribute dont_touch of G185: signal is true;
	signal G186: std_logic; attribute dont_touch of G186: signal is true;
	signal G189: std_logic; attribute dont_touch of G189: signal is true;
	signal G192: std_logic; attribute dont_touch of G192: signal is true;
	signal G195: std_logic; attribute dont_touch of G195: signal is true;
	signal G198: std_logic; attribute dont_touch of G198: signal is true;
	signal G201: std_logic; attribute dont_touch of G201: signal is true;
	signal G204: std_logic; attribute dont_touch of G204: signal is true;
	signal G207: std_logic; attribute dont_touch of G207: signal is true;
	signal G210: std_logic; attribute dont_touch of G210: signal is true;
	signal G213: std_logic; attribute dont_touch of G213: signal is true;
	signal G216: std_logic; attribute dont_touch of G216: signal is true;
	signal G219: std_logic; attribute dont_touch of G219: signal is true;
	signal G222: std_logic; attribute dont_touch of G222: signal is true;
	signal G225: std_logic; attribute dont_touch of G225: signal is true;
	signal G228: std_logic; attribute dont_touch of G228: signal is true;
	signal G231: std_logic; attribute dont_touch of G231: signal is true;
	signal G234: std_logic; attribute dont_touch of G234: signal is true;
	signal G237: std_logic; attribute dont_touch of G237: signal is true;
	signal G240: std_logic; attribute dont_touch of G240: signal is true;
	signal G243: std_logic; attribute dont_touch of G243: signal is true;
	signal G246: std_logic; attribute dont_touch of G246: signal is true;
	signal G249: std_logic; attribute dont_touch of G249: signal is true;
	signal G252: std_logic; attribute dont_touch of G252: signal is true;
	signal G255: std_logic; attribute dont_touch of G255: signal is true;
	signal G258: std_logic; attribute dont_touch of G258: signal is true;
	signal G261: std_logic; attribute dont_touch of G261: signal is true;
	signal G264: std_logic; attribute dont_touch of G264: signal is true;
	signal G267: std_logic; attribute dont_touch of G267: signal is true;
	signal G270: std_logic; attribute dont_touch of G270: signal is true;
	signal G273: std_logic; attribute dont_touch of G273: signal is true;
	signal G276: std_logic; attribute dont_touch of G276: signal is true;
	signal G279: std_logic; attribute dont_touch of G279: signal is true;
	signal G280: std_logic; attribute dont_touch of G280: signal is true;
	signal G281: std_logic; attribute dont_touch of G281: signal is true;
	signal G282: std_logic; attribute dont_touch of G282: signal is true;
	signal G283: std_logic; attribute dont_touch of G283: signal is true;
	signal G284: std_logic; attribute dont_touch of G284: signal is true;
	signal G285: std_logic; attribute dont_touch of G285: signal is true;
	signal G286: std_logic; attribute dont_touch of G286: signal is true;
	signal G287: std_logic; attribute dont_touch of G287: signal is true;
	signal G288: std_logic; attribute dont_touch of G288: signal is true;
	signal G289: std_logic; attribute dont_touch of G289: signal is true;
	signal G290: std_logic; attribute dont_touch of G290: signal is true;
	signal G291: std_logic; attribute dont_touch of G291: signal is true;
	signal G294: std_logic; attribute dont_touch of G294: signal is true;
	signal G295: std_logic; attribute dont_touch of G295: signal is true;
	signal G296: std_logic; attribute dont_touch of G296: signal is true;
	signal G297: std_logic; attribute dont_touch of G297: signal is true;
	signal G298: std_logic; attribute dont_touch of G298: signal is true;
	signal G299: std_logic; attribute dont_touch of G299: signal is true;
	signal G300: std_logic; attribute dont_touch of G300: signal is true;
	signal G301: std_logic; attribute dont_touch of G301: signal is true;
	signal G302: std_logic; attribute dont_touch of G302: signal is true;
	signal G303: std_logic; attribute dont_touch of G303: signal is true;
	signal G304: std_logic; attribute dont_touch of G304: signal is true;
	signal G305: std_logic; attribute dont_touch of G305: signal is true;
	signal G308: std_logic; attribute dont_touch of G308: signal is true;
	signal G309: std_logic; attribute dont_touch of G309: signal is true;
	signal G312: std_logic; attribute dont_touch of G312: signal is true;
	signal G313: std_logic; attribute dont_touch of G313: signal is true;
	signal G314: std_logic; attribute dont_touch of G314: signal is true;
	signal G315: std_logic; attribute dont_touch of G315: signal is true;
	signal G316: std_logic; attribute dont_touch of G316: signal is true;
	signal G317: std_logic; attribute dont_touch of G317: signal is true;
	signal G318: std_logic; attribute dont_touch of G318: signal is true;
	signal G319: std_logic; attribute dont_touch of G319: signal is true;
	signal G320: std_logic; attribute dont_touch of G320: signal is true;
	signal G321: std_logic; attribute dont_touch of G321: signal is true;
	signal G322: std_logic; attribute dont_touch of G322: signal is true;
	signal G323: std_logic; attribute dont_touch of G323: signal is true;
	signal G324: std_logic; attribute dont_touch of G324: signal is true;
	signal G325: std_logic; attribute dont_touch of G325: signal is true;
	signal G331: std_logic; attribute dont_touch of G331: signal is true;
	signal G337: std_logic; attribute dont_touch of G337: signal is true;
	signal G342: std_logic; attribute dont_touch of G342: signal is true;
	signal G343: std_logic; attribute dont_touch of G343: signal is true;
	signal G346: std_logic; attribute dont_touch of G346: signal is true;
	signal G349: std_logic; attribute dont_touch of G349: signal is true;
	signal G350: std_logic; attribute dont_touch of G350: signal is true;
	signal G351: std_logic; attribute dont_touch of G351: signal is true;
	signal G352: std_logic; attribute dont_touch of G352: signal is true;
	signal G353: std_logic; attribute dont_touch of G353: signal is true;
	signal G354: std_logic; attribute dont_touch of G354: signal is true;
	signal G357: std_logic; attribute dont_touch of G357: signal is true;
	signal G358: std_logic; attribute dont_touch of G358: signal is true;
	signal G361: std_logic; attribute dont_touch of G361: signal is true;
	signal G364: std_logic; attribute dont_touch of G364: signal is true;
	signal G365: std_logic; attribute dont_touch of G365: signal is true;
	signal G366: std_logic; attribute dont_touch of G366: signal is true;
	signal G367: std_logic; attribute dont_touch of G367: signal is true;
	signal G368: std_logic; attribute dont_touch of G368: signal is true;
	signal G369: std_logic; attribute dont_touch of G369: signal is true;
	signal G372: std_logic; attribute dont_touch of G372: signal is true;
	signal G373: std_logic; attribute dont_touch of G373: signal is true;
	signal G376: std_logic; attribute dont_touch of G376: signal is true;
	signal G379: std_logic; attribute dont_touch of G379: signal is true;
	signal G380: std_logic; attribute dont_touch of G380: signal is true;
	signal G381: std_logic; attribute dont_touch of G381: signal is true;
	signal G382: std_logic; attribute dont_touch of G382: signal is true;
	signal G383: std_logic; attribute dont_touch of G383: signal is true;
	signal G384: std_logic; attribute dont_touch of G384: signal is true;
	signal G387: std_logic; attribute dont_touch of G387: signal is true;
	signal G388: std_logic; attribute dont_touch of G388: signal is true;
	signal G391: std_logic; attribute dont_touch of G391: signal is true;
	signal G394: std_logic; attribute dont_touch of G394: signal is true;
	signal G395: std_logic; attribute dont_touch of G395: signal is true;
	signal G396: std_logic; attribute dont_touch of G396: signal is true;
	signal G397: std_logic; attribute dont_touch of G397: signal is true;
	signal G398: std_logic; attribute dont_touch of G398: signal is true;
	signal G401: std_logic; attribute dont_touch of G401: signal is true;
	signal G402: std_logic; attribute dont_touch of G402: signal is true;
	signal G403: std_logic; attribute dont_touch of G403: signal is true;
	signal G404: std_logic; attribute dont_touch of G404: signal is true;
	signal G405: std_logic; attribute dont_touch of G405: signal is true;
	signal G408: std_logic; attribute dont_touch of G408: signal is true;
	signal G411: std_logic; attribute dont_touch of G411: signal is true;
	signal G414: std_logic; attribute dont_touch of G414: signal is true;
	signal G417: std_logic; attribute dont_touch of G417: signal is true;
	signal G420: std_logic; attribute dont_touch of G420: signal is true;
	signal G423: std_logic; attribute dont_touch of G423: signal is true;
	signal G426: std_logic; attribute dont_touch of G426: signal is true;
	signal G427: std_logic; attribute dont_touch of G427: signal is true;
	signal G428: std_logic; attribute dont_touch of G428: signal is true;
	signal G429: std_logic; attribute dont_touch of G429: signal is true;
	signal G432: std_logic; attribute dont_touch of G432: signal is true;
	signal G435: std_logic; attribute dont_touch of G435: signal is true;
	signal G438: std_logic; attribute dont_touch of G438: signal is true;
	signal G441: std_logic; attribute dont_touch of G441: signal is true;
	signal G444: std_logic; attribute dont_touch of G444: signal is true;
	signal G447: std_logic; attribute dont_touch of G447: signal is true;
	signal G448: std_logic; attribute dont_touch of G448: signal is true;
	signal G449: std_logic; attribute dont_touch of G449: signal is true;
	signal G450: std_logic; attribute dont_touch of G450: signal is true;
	signal G451: std_logic; attribute dont_touch of G451: signal is true;
	signal G452: std_logic; attribute dont_touch of G452: signal is true;
	signal G453: std_logic; attribute dont_touch of G453: signal is true;
	signal G454: std_logic; attribute dont_touch of G454: signal is true;
	signal G455: std_logic; attribute dont_touch of G455: signal is true;
	signal G458: std_logic; attribute dont_touch of G458: signal is true;
	signal G461: std_logic; attribute dont_touch of G461: signal is true;
	signal G464: std_logic; attribute dont_touch of G464: signal is true;
	signal G465: std_logic; attribute dont_touch of G465: signal is true;
	signal G468: std_logic; attribute dont_touch of G468: signal is true;
	signal G471: std_logic; attribute dont_touch of G471: signal is true;
	signal G474: std_logic; attribute dont_touch of G474: signal is true;
	signal G477: std_logic; attribute dont_touch of G477: signal is true;
	signal G478: std_logic; attribute dont_touch of G478: signal is true;
	signal G479: std_logic; attribute dont_touch of G479: signal is true;
	signal G480: std_logic; attribute dont_touch of G480: signal is true;
	signal G481: std_logic; attribute dont_touch of G481: signal is true;
	signal G484: std_logic; attribute dont_touch of G484: signal is true;
	signal G485: std_logic; attribute dont_touch of G485: signal is true;
	signal G486: std_logic; attribute dont_touch of G486: signal is true;
	signal G487: std_logic; attribute dont_touch of G487: signal is true;
	signal G488: std_logic; attribute dont_touch of G488: signal is true;
	signal G489: std_logic; attribute dont_touch of G489: signal is true;
	signal G490: std_logic; attribute dont_touch of G490: signal is true;
	signal G493: std_logic; attribute dont_touch of G493: signal is true;
	signal G496: std_logic; attribute dont_touch of G496: signal is true;
	signal G499: std_logic; attribute dont_touch of G499: signal is true;
	signal G506: std_logic; attribute dont_touch of G506: signal is true;
	signal G507: std_logic; attribute dont_touch of G507: signal is true;
	signal G508: std_logic; attribute dont_touch of G508: signal is true;
	signal G509: std_logic; attribute dont_touch of G509: signal is true;
	signal G510: std_logic; attribute dont_touch of G510: signal is true;
	signal G513: std_logic; attribute dont_touch of G513: signal is true;
	signal G514: std_logic; attribute dont_touch of G514: signal is true;
	signal G515: std_logic; attribute dont_touch of G515: signal is true;
	signal G516: std_logic; attribute dont_touch of G516: signal is true;
	signal G517: std_logic; attribute dont_touch of G517: signal is true;
	signal G518: std_logic; attribute dont_touch of G518: signal is true;
	signal G519: std_logic; attribute dont_touch of G519: signal is true;
	signal G520: std_logic; attribute dont_touch of G520: signal is true;
	signal G523: std_logic; attribute dont_touch of G523: signal is true;
	signal G524: std_logic; attribute dont_touch of G524: signal is true;
	signal G525: std_logic; attribute dont_touch of G525: signal is true;
	signal G528: std_logic; attribute dont_touch of G528: signal is true;
	signal G529: std_logic; attribute dont_touch of G529: signal is true;
	signal G530: std_logic; attribute dont_touch of G530: signal is true;
	signal G531: std_logic; attribute dont_touch of G531: signal is true;
	signal G532: std_logic; attribute dont_touch of G532: signal is true;
	signal G533: std_logic; attribute dont_touch of G533: signal is true;
	signal G534: std_logic; attribute dont_touch of G534: signal is true;
	signal G535: std_logic; attribute dont_touch of G535: signal is true;
	signal G536: std_logic; attribute dont_touch of G536: signal is true;
	signal G537: std_logic; attribute dont_touch of G537: signal is true;
	signal G538: std_logic; attribute dont_touch of G538: signal is true;
	signal G541: std_logic; attribute dont_touch of G541: signal is true;
	signal G542: std_logic; attribute dont_touch of G542: signal is true;
	signal G543: std_logic; attribute dont_touch of G543: signal is true;
	signal G544: std_logic; attribute dont_touch of G544: signal is true;
	signal G545: std_logic; attribute dont_touch of G545: signal is true;
	signal G548: std_logic; attribute dont_touch of G548: signal is true;
	signal G549: std_logic; attribute dont_touch of G549: signal is true;
	signal G550: std_logic; attribute dont_touch of G550: signal is true;
	signal G551: std_logic; attribute dont_touch of G551: signal is true;
	signal G554: std_logic; attribute dont_touch of G554: signal is true;
	signal G557: std_logic; attribute dont_touch of G557: signal is true;
	signal G558: std_logic; attribute dont_touch of G558: signal is true;
	signal G559: std_logic; attribute dont_touch of G559: signal is true;
	signal G562: std_logic; attribute dont_touch of G562: signal is true;
	signal G564: std_logic; attribute dont_touch of G564: signal is true;
	signal G565: std_logic; attribute dont_touch of G565: signal is true;
	signal G566: std_logic; attribute dont_touch of G566: signal is true;
	signal G567: std_logic; attribute dont_touch of G567: signal is true;
	signal G568: std_logic; attribute dont_touch of G568: signal is true;
	signal G569: std_logic; attribute dont_touch of G569: signal is true;
	signal G570: std_logic; attribute dont_touch of G570: signal is true;
	signal G571: std_logic; attribute dont_touch of G571: signal is true;
	signal G572: std_logic; attribute dont_touch of G572: signal is true;
	signal G573: std_logic; attribute dont_touch of G573: signal is true;
	signal G574: std_logic; attribute dont_touch of G574: signal is true;
	signal G575: std_logic; attribute dont_touch of G575: signal is true;
	signal G576: std_logic; attribute dont_touch of G576: signal is true;
	signal G577: std_logic; attribute dont_touch of G577: signal is true;
	signal G578: std_logic; attribute dont_touch of G578: signal is true;
	signal G579: std_logic; attribute dont_touch of G579: signal is true;
	signal G580: std_logic; attribute dont_touch of G580: signal is true;
	signal G581: std_logic; attribute dont_touch of G581: signal is true;
	signal G582: std_logic; attribute dont_touch of G582: signal is true;
	signal G583: std_logic; attribute dont_touch of G583: signal is true;
	signal G584: std_logic; attribute dont_touch of G584: signal is true;
	signal G585: std_logic; attribute dont_touch of G585: signal is true;
	signal G586: std_logic; attribute dont_touch of G586: signal is true;
	signal G587: std_logic; attribute dont_touch of G587: signal is true;
	signal G590: std_logic; attribute dont_touch of G590: signal is true;
	signal G593: std_logic; attribute dont_touch of G593: signal is true;
	signal G596: std_logic; attribute dont_touch of G596: signal is true;
	signal G599: std_logic; attribute dont_touch of G599: signal is true;
	signal G602: std_logic; attribute dont_touch of G602: signal is true;
	signal G605: std_logic; attribute dont_touch of G605: signal is true;
	signal G608: std_logic; attribute dont_touch of G608: signal is true;
	signal G611: std_logic; attribute dont_touch of G611: signal is true;
	signal G614: std_logic; attribute dont_touch of G614: signal is true;
	signal G617: std_logic; attribute dont_touch of G617: signal is true;
	signal G620: std_logic; attribute dont_touch of G620: signal is true;
	signal G623: std_logic; attribute dont_touch of G623: signal is true;
	signal G626: std_logic; attribute dont_touch of G626: signal is true;
	signal G629: std_logic; attribute dont_touch of G629: signal is true;
	signal G630: std_logic; attribute dont_touch of G630: signal is true;
	signal G633: std_logic; attribute dont_touch of G633: signal is true;
	signal G640: std_logic; attribute dont_touch of G640: signal is true;
	signal G646: std_logic; attribute dont_touch of G646: signal is true;
	signal G653: std_logic; attribute dont_touch of G653: signal is true;
	signal G659: std_logic; attribute dont_touch of G659: signal is true;
	signal G660: std_logic; attribute dont_touch of G660: signal is true;
	signal G666: std_logic; attribute dont_touch of G666: signal is true;
	signal G672: std_logic; attribute dont_touch of G672: signal is true;
	signal G679: std_logic; attribute dont_touch of G679: signal is true;
	signal G686: std_logic; attribute dont_touch of G686: signal is true;
	signal G692: std_logic; attribute dont_touch of G692: signal is true;
	signal G698: std_logic; attribute dont_touch of G698: signal is true;
	signal G699: std_logic; attribute dont_touch of G699: signal is true;
	signal G700: std_logic; attribute dont_touch of G700: signal is true;
	signal G701: std_logic; attribute dont_touch of G701: signal is true;
	signal G702: std_logic; attribute dont_touch of G702: signal is true;
	signal G703: std_logic; attribute dont_touch of G703: signal is true;
	signal G704: std_logic; attribute dont_touch of G704: signal is true;
	signal G705: std_logic; attribute dont_touch of G705: signal is true;
	signal G706: std_logic; attribute dont_touch of G706: signal is true;
	signal G707: std_logic; attribute dont_touch of G707: signal is true;
	signal G708: std_logic; attribute dont_touch of G708: signal is true;
	signal G709: std_logic; attribute dont_touch of G709: signal is true;
	signal G710: std_logic; attribute dont_touch of G710: signal is true;
	signal G711: std_logic; attribute dont_touch of G711: signal is true;
	signal G712: std_logic; attribute dont_touch of G712: signal is true;
	signal G713: std_logic; attribute dont_touch of G713: signal is true;
	signal G714: std_logic; attribute dont_touch of G714: signal is true;
	signal G715: std_logic; attribute dont_touch of G715: signal is true;
	signal G716: std_logic; attribute dont_touch of G716: signal is true;
	signal G717: std_logic; attribute dont_touch of G717: signal is true;
	signal G718: std_logic; attribute dont_touch of G718: signal is true;
	signal G719: std_logic; attribute dont_touch of G719: signal is true;
	signal G720: std_logic; attribute dont_touch of G720: signal is true;
	signal G721: std_logic; attribute dont_touch of G721: signal is true;
	signal G722: std_logic; attribute dont_touch of G722: signal is true;
	signal G723: std_logic; attribute dont_touch of G723: signal is true;
	signal G724: std_logic; attribute dont_touch of G724: signal is true;
	signal G725: std_logic; attribute dont_touch of G725: signal is true;
	signal G726: std_logic; attribute dont_touch of G726: signal is true;
	signal G727: std_logic; attribute dont_touch of G727: signal is true;
	signal G728: std_logic; attribute dont_touch of G728: signal is true;
	signal G729: std_logic; attribute dont_touch of G729: signal is true;
	signal G730: std_logic; attribute dont_touch of G730: signal is true;
	signal G731: std_logic; attribute dont_touch of G731: signal is true;
	signal G732: std_logic; attribute dont_touch of G732: signal is true;
	signal G733: std_logic; attribute dont_touch of G733: signal is true;
	signal G734: std_logic; attribute dont_touch of G734: signal is true;
	signal G735: std_logic; attribute dont_touch of G735: signal is true;
	signal G736: std_logic; attribute dont_touch of G736: signal is true;
	signal G737: std_logic; attribute dont_touch of G737: signal is true;
	signal G738: std_logic; attribute dont_touch of G738: signal is true;
	signal G739: std_logic; attribute dont_touch of G739: signal is true;
	signal G740: std_logic; attribute dont_touch of G740: signal is true;
	signal G744: std_logic; attribute dont_touch of G744: signal is true;
	signal G749: std_logic; attribute dont_touch of G749: signal is true;
	signal G753: std_logic; attribute dont_touch of G753: signal is true;
	signal G758: std_logic; attribute dont_touch of G758: signal is true;
	signal G762: std_logic; attribute dont_touch of G762: signal is true;
	signal G767: std_logic; attribute dont_touch of G767: signal is true;
	signal G771: std_logic; attribute dont_touch of G771: signal is true;
	signal G776: std_logic; attribute dont_touch of G776: signal is true;
	signal G780: std_logic; attribute dont_touch of G780: signal is true;
	signal G785: std_logic; attribute dont_touch of G785: signal is true;
	signal G789: std_logic; attribute dont_touch of G789: signal is true;
	signal G793: std_logic; attribute dont_touch of G793: signal is true;
	signal G797: std_logic; attribute dont_touch of G797: signal is true;
	signal G801: std_logic; attribute dont_touch of G801: signal is true;
	signal G805: std_logic; attribute dont_touch of G805: signal is true;
	signal G809: std_logic; attribute dont_touch of G809: signal is true;
	signal G813: std_logic; attribute dont_touch of G813: signal is true;
	signal G817: std_logic; attribute dont_touch of G817: signal is true;
	signal G818: std_logic; attribute dont_touch of G818: signal is true;
	signal G819: std_logic; attribute dont_touch of G819: signal is true;
	signal G820: std_logic; attribute dont_touch of G820: signal is true;
	signal G821: std_logic; attribute dont_touch of G821: signal is true;
	signal G822: std_logic; attribute dont_touch of G822: signal is true;
	signal G823: std_logic; attribute dont_touch of G823: signal is true;
	signal G826: std_logic; attribute dont_touch of G826: signal is true;
	signal G829: std_logic; attribute dont_touch of G829: signal is true;
	signal G830: std_logic; attribute dont_touch of G830: signal is true;
	signal G831: std_logic; attribute dont_touch of G831: signal is true;
	signal G832: std_logic; attribute dont_touch of G832: signal is true;
	signal G833: std_logic; attribute dont_touch of G833: signal is true;
	signal G834: std_logic; attribute dont_touch of G834: signal is true;
	signal G835: std_logic; attribute dont_touch of G835: signal is true;
	signal G836: std_logic; attribute dont_touch of G836: signal is true;
	signal G837: std_logic; attribute dont_touch of G837: signal is true;
	signal G838: std_logic; attribute dont_touch of G838: signal is true;
	signal G839: std_logic; attribute dont_touch of G839: signal is true;
	signal G840: std_logic; attribute dont_touch of G840: signal is true;
	signal G841: std_logic; attribute dont_touch of G841: signal is true;
	signal G842: std_logic; attribute dont_touch of G842: signal is true;
	signal G843: std_logic; attribute dont_touch of G843: signal is true;
	signal G844: std_logic; attribute dont_touch of G844: signal is true;
	signal G845: std_logic; attribute dont_touch of G845: signal is true;
	signal G846: std_logic; attribute dont_touch of G846: signal is true;
	signal G847: std_logic; attribute dont_touch of G847: signal is true;
	signal G848: std_logic; attribute dont_touch of G848: signal is true;
	signal G849: std_logic; attribute dont_touch of G849: signal is true;
	signal G850: std_logic; attribute dont_touch of G850: signal is true;
	signal G851: std_logic; attribute dont_touch of G851: signal is true;
	signal G852: std_logic; attribute dont_touch of G852: signal is true;
	signal G853: std_logic; attribute dont_touch of G853: signal is true;
	signal G856: std_logic; attribute dont_touch of G856: signal is true;
	signal G857: std_logic; attribute dont_touch of G857: signal is true;
	signal G858: std_logic; attribute dont_touch of G858: signal is true;
	signal G859: std_logic; attribute dont_touch of G859: signal is true;
	signal G860: std_logic; attribute dont_touch of G860: signal is true;
	signal G861: std_logic; attribute dont_touch of G861: signal is true;
	signal G862: std_logic; attribute dont_touch of G862: signal is true;
	signal G863: std_logic; attribute dont_touch of G863: signal is true;
	signal G864: std_logic; attribute dont_touch of G864: signal is true;
	signal G865: std_logic; attribute dont_touch of G865: signal is true;
	signal G866: std_logic; attribute dont_touch of G866: signal is true;
	signal G867: std_logic; attribute dont_touch of G867: signal is true;
	signal G868: std_logic; attribute dont_touch of G868: signal is true;
	signal G869: std_logic; attribute dont_touch of G869: signal is true;
	signal G870: std_logic; attribute dont_touch of G870: signal is true;
	signal G873: std_logic; attribute dont_touch of G873: signal is true;
	signal G876: std_logic; attribute dont_touch of G876: signal is true;
	signal G879: std_logic; attribute dont_touch of G879: signal is true;
	signal G882: std_logic; attribute dont_touch of G882: signal is true;
	signal G885: std_logic; attribute dont_touch of G885: signal is true;
	signal G888: std_logic; attribute dont_touch of G888: signal is true;
	signal G891: std_logic; attribute dont_touch of G891: signal is true;
	signal G894: std_logic; attribute dont_touch of G894: signal is true;
	signal G897: std_logic; attribute dont_touch of G897: signal is true;
	signal G900: std_logic; attribute dont_touch of G900: signal is true;
	signal G903: std_logic; attribute dont_touch of G903: signal is true;
	signal G906: std_logic; attribute dont_touch of G906: signal is true;
	signal G909: std_logic; attribute dont_touch of G909: signal is true;
	signal G912: std_logic; attribute dont_touch of G912: signal is true;
	signal G915: std_logic; attribute dont_touch of G915: signal is true;
	signal G918: std_logic; attribute dont_touch of G918: signal is true;
	signal G921: std_logic; attribute dont_touch of G921: signal is true;
	signal G924: std_logic; attribute dont_touch of G924: signal is true;
	signal G927: std_logic; attribute dont_touch of G927: signal is true;
	signal G930: std_logic; attribute dont_touch of G930: signal is true;
	signal G933: std_logic; attribute dont_touch of G933: signal is true;
	signal G936: std_logic; attribute dont_touch of G936: signal is true;
	signal G939: std_logic; attribute dont_touch of G939: signal is true;
	signal G942: std_logic; attribute dont_touch of G942: signal is true;
	signal G945: std_logic; attribute dont_touch of G945: signal is true;
	signal G948: std_logic; attribute dont_touch of G948: signal is true;
	signal G951: std_logic; attribute dont_touch of G951: signal is true;
	signal G954: std_logic; attribute dont_touch of G954: signal is true;
	signal G957: std_logic; attribute dont_touch of G957: signal is true;
	signal G960: std_logic; attribute dont_touch of G960: signal is true;
	signal G963: std_logic; attribute dont_touch of G963: signal is true;
	signal G966: std_logic; attribute dont_touch of G966: signal is true;
	signal G967: std_logic; attribute dont_touch of G967: signal is true;
	signal G968: std_logic; attribute dont_touch of G968: signal is true;
	signal G969: std_logic; attribute dont_touch of G969: signal is true;
	signal G970: std_logic; attribute dont_touch of G970: signal is true;
	signal G971: std_logic; attribute dont_touch of G971: signal is true;
	signal G972: std_logic; attribute dont_touch of G972: signal is true;
	signal G973: std_logic; attribute dont_touch of G973: signal is true;
	signal G974: std_logic; attribute dont_touch of G974: signal is true;
	signal G975: std_logic; attribute dont_touch of G975: signal is true;
	signal G976: std_logic; attribute dont_touch of G976: signal is true;
	signal G977: std_logic; attribute dont_touch of G977: signal is true;
	signal G978: std_logic; attribute dont_touch of G978: signal is true;
	signal G981: std_logic; attribute dont_touch of G981: signal is true;
	signal G982: std_logic; attribute dont_touch of G982: signal is true;
	signal G983: std_logic; attribute dont_touch of G983: signal is true;
	signal G984: std_logic; attribute dont_touch of G984: signal is true;
	signal G985: std_logic; attribute dont_touch of G985: signal is true;
	signal G986: std_logic; attribute dont_touch of G986: signal is true;
	signal G987: std_logic; attribute dont_touch of G987: signal is true;
	signal G988: std_logic; attribute dont_touch of G988: signal is true;
	signal G989: std_logic; attribute dont_touch of G989: signal is true;
	signal G990: std_logic; attribute dont_touch of G990: signal is true;
	signal G991: std_logic; attribute dont_touch of G991: signal is true;
	signal G992: std_logic; attribute dont_touch of G992: signal is true;
	signal G995: std_logic; attribute dont_touch of G995: signal is true;
	signal G996: std_logic; attribute dont_touch of G996: signal is true;
	signal G999: std_logic; attribute dont_touch of G999: signal is true;
	signal G1000: std_logic; attribute dont_touch of G1000: signal is true;
	signal G1001: std_logic; attribute dont_touch of G1001: signal is true;
	signal G1002: std_logic; attribute dont_touch of G1002: signal is true;
	signal G1003: std_logic; attribute dont_touch of G1003: signal is true;
	signal G1004: std_logic; attribute dont_touch of G1004: signal is true;
	signal G1005: std_logic; attribute dont_touch of G1005: signal is true;
	signal G1006: std_logic; attribute dont_touch of G1006: signal is true;
	signal G1007: std_logic; attribute dont_touch of G1007: signal is true;
	signal G1008: std_logic; attribute dont_touch of G1008: signal is true;
	signal G1009: std_logic; attribute dont_touch of G1009: signal is true;
	signal G1010: std_logic; attribute dont_touch of G1010: signal is true;
	signal G1011: std_logic; attribute dont_touch of G1011: signal is true;
	signal G1012: std_logic; attribute dont_touch of G1012: signal is true;
	signal G1018: std_logic; attribute dont_touch of G1018: signal is true;
	signal G1024: std_logic; attribute dont_touch of G1024: signal is true;
	signal G1029: std_logic; attribute dont_touch of G1029: signal is true;
	signal G1030: std_logic; attribute dont_touch of G1030: signal is true;
	signal G1033: std_logic; attribute dont_touch of G1033: signal is true;
	signal G1036: std_logic; attribute dont_touch of G1036: signal is true;
	signal G1037: std_logic; attribute dont_touch of G1037: signal is true;
	signal G1038: std_logic; attribute dont_touch of G1038: signal is true;
	signal G1039: std_logic; attribute dont_touch of G1039: signal is true;
	signal G1040: std_logic; attribute dont_touch of G1040: signal is true;
	signal G1041: std_logic; attribute dont_touch of G1041: signal is true;
	signal G1044: std_logic; attribute dont_touch of G1044: signal is true;
	signal G1045: std_logic; attribute dont_touch of G1045: signal is true;
	signal G1048: std_logic; attribute dont_touch of G1048: signal is true;
	signal G1051: std_logic; attribute dont_touch of G1051: signal is true;
	signal G1052: std_logic; attribute dont_touch of G1052: signal is true;
	signal G1053: std_logic; attribute dont_touch of G1053: signal is true;
	signal G1054: std_logic; attribute dont_touch of G1054: signal is true;
	signal G1055: std_logic; attribute dont_touch of G1055: signal is true;
	signal G1056: std_logic; attribute dont_touch of G1056: signal is true;
	signal G1059: std_logic; attribute dont_touch of G1059: signal is true;
	signal G1060: std_logic; attribute dont_touch of G1060: signal is true;
	signal G1063: std_logic; attribute dont_touch of G1063: signal is true;
	signal G1066: std_logic; attribute dont_touch of G1066: signal is true;
	signal G1067: std_logic; attribute dont_touch of G1067: signal is true;
	signal G1068: std_logic; attribute dont_touch of G1068: signal is true;
	signal G1069: std_logic; attribute dont_touch of G1069: signal is true;
	signal G1070: std_logic; attribute dont_touch of G1070: signal is true;
	signal G1071: std_logic; attribute dont_touch of G1071: signal is true;
	signal G1074: std_logic; attribute dont_touch of G1074: signal is true;
	signal G1075: std_logic; attribute dont_touch of G1075: signal is true;
	signal G1078: std_logic; attribute dont_touch of G1078: signal is true;
	signal G1081: std_logic; attribute dont_touch of G1081: signal is true;
	signal G1082: std_logic; attribute dont_touch of G1082: signal is true;
	signal G1083: std_logic; attribute dont_touch of G1083: signal is true;
	signal G1084: std_logic; attribute dont_touch of G1084: signal is true;
	signal G1085: std_logic; attribute dont_touch of G1085: signal is true;
	signal G1088: std_logic; attribute dont_touch of G1088: signal is true;
	signal G1089: std_logic; attribute dont_touch of G1089: signal is true;
	signal G1090: std_logic; attribute dont_touch of G1090: signal is true;
	signal G1091: std_logic; attribute dont_touch of G1091: signal is true;
	signal G1092: std_logic; attribute dont_touch of G1092: signal is true;
	signal G1095: std_logic; attribute dont_touch of G1095: signal is true;
	signal G1098: std_logic; attribute dont_touch of G1098: signal is true;
	signal G1101: std_logic; attribute dont_touch of G1101: signal is true;
	signal G1104: std_logic; attribute dont_touch of G1104: signal is true;
	signal G1107: std_logic; attribute dont_touch of G1107: signal is true;
	signal G1110: std_logic; attribute dont_touch of G1110: signal is true;
	signal G1113: std_logic; attribute dont_touch of G1113: signal is true;
	signal G1114: std_logic; attribute dont_touch of G1114: signal is true;
	signal G1115: std_logic; attribute dont_touch of G1115: signal is true;
	signal G1116: std_logic; attribute dont_touch of G1116: signal is true;
	signal G1119: std_logic; attribute dont_touch of G1119: signal is true;
	signal G1122: std_logic; attribute dont_touch of G1122: signal is true;
	signal G1125: std_logic; attribute dont_touch of G1125: signal is true;
	signal G1128: std_logic; attribute dont_touch of G1128: signal is true;
	signal G1131: std_logic; attribute dont_touch of G1131: signal is true;
	signal G1134: std_logic; attribute dont_touch of G1134: signal is true;
	signal G1135: std_logic; attribute dont_touch of G1135: signal is true;
	signal G1136: std_logic; attribute dont_touch of G1136: signal is true;
	signal G1137: std_logic; attribute dont_touch of G1137: signal is true;
	signal G1138: std_logic; attribute dont_touch of G1138: signal is true;
	signal G1139: std_logic; attribute dont_touch of G1139: signal is true;
	signal G1140: std_logic; attribute dont_touch of G1140: signal is true;
	signal G1141: std_logic; attribute dont_touch of G1141: signal is true;
	signal G1142: std_logic; attribute dont_touch of G1142: signal is true;
	signal G1145: std_logic; attribute dont_touch of G1145: signal is true;
	signal G1148: std_logic; attribute dont_touch of G1148: signal is true;
	signal G1151: std_logic; attribute dont_touch of G1151: signal is true;
	signal G1152: std_logic; attribute dont_touch of G1152: signal is true;
	signal G1155: std_logic; attribute dont_touch of G1155: signal is true;
	signal G1158: std_logic; attribute dont_touch of G1158: signal is true;
	signal G1161: std_logic; attribute dont_touch of G1161: signal is true;
	signal G1164: std_logic; attribute dont_touch of G1164: signal is true;
	signal G1165: std_logic; attribute dont_touch of G1165: signal is true;
	signal G1166: std_logic; attribute dont_touch of G1166: signal is true;
	signal G1167: std_logic; attribute dont_touch of G1167: signal is true;
	signal G1168: std_logic; attribute dont_touch of G1168: signal is true;
	signal G1171: std_logic; attribute dont_touch of G1171: signal is true;
	signal G1172: std_logic; attribute dont_touch of G1172: signal is true;
	signal G1173: std_logic; attribute dont_touch of G1173: signal is true;
	signal G1174: std_logic; attribute dont_touch of G1174: signal is true;
	signal G1175: std_logic; attribute dont_touch of G1175: signal is true;
	signal G1176: std_logic; attribute dont_touch of G1176: signal is true;
	signal G1177: std_logic; attribute dont_touch of G1177: signal is true;
	signal G1180: std_logic; attribute dont_touch of G1180: signal is true;
	signal G1183: std_logic; attribute dont_touch of G1183: signal is true;
	signal G1186: std_logic; attribute dont_touch of G1186: signal is true;
	signal G1192: std_logic; attribute dont_touch of G1192: signal is true;
	signal G1193: std_logic; attribute dont_touch of G1193: signal is true;
	signal G1194: std_logic; attribute dont_touch of G1194: signal is true;
	signal G1195: std_logic; attribute dont_touch of G1195: signal is true;
	signal G1196: std_logic; attribute dont_touch of G1196: signal is true;
	signal G1199: std_logic; attribute dont_touch of G1199: signal is true;
	signal G1200: std_logic; attribute dont_touch of G1200: signal is true;
	signal G1201: std_logic; attribute dont_touch of G1201: signal is true;
	signal G1202: std_logic; attribute dont_touch of G1202: signal is true;
	signal G1203: std_logic; attribute dont_touch of G1203: signal is true;
	signal G1204: std_logic; attribute dont_touch of G1204: signal is true;
	signal G1205: std_logic; attribute dont_touch of G1205: signal is true;
	signal G1206: std_logic; attribute dont_touch of G1206: signal is true;
	signal G1209: std_logic; attribute dont_touch of G1209: signal is true;
	signal G1210: std_logic; attribute dont_touch of G1210: signal is true;
	signal G1211: std_logic; attribute dont_touch of G1211: signal is true;
	signal G1214: std_logic; attribute dont_touch of G1214: signal is true;
	signal G1215: std_logic; attribute dont_touch of G1215: signal is true;
	signal G1216: std_logic; attribute dont_touch of G1216: signal is true;
	signal G1217: std_logic; attribute dont_touch of G1217: signal is true;
	signal G1218: std_logic; attribute dont_touch of G1218: signal is true;
	signal G1219: std_logic; attribute dont_touch of G1219: signal is true;
	signal G1220: std_logic; attribute dont_touch of G1220: signal is true;
	signal G1221: std_logic; attribute dont_touch of G1221: signal is true;
	signal G1222: std_logic; attribute dont_touch of G1222: signal is true;
	signal G1223: std_logic; attribute dont_touch of G1223: signal is true;
	signal G1224: std_logic; attribute dont_touch of G1224: signal is true;
	signal G1227: std_logic; attribute dont_touch of G1227: signal is true;
	signal G1228: std_logic; attribute dont_touch of G1228: signal is true;
	signal G1229: std_logic; attribute dont_touch of G1229: signal is true;
	signal G1230: std_logic; attribute dont_touch of G1230: signal is true;
	signal G1231: std_logic; attribute dont_touch of G1231: signal is true;
	signal G1234: std_logic; attribute dont_touch of G1234: signal is true;
	signal G1235: std_logic; attribute dont_touch of G1235: signal is true;
	signal G1236: std_logic; attribute dont_touch of G1236: signal is true;
	signal G1237: std_logic; attribute dont_touch of G1237: signal is true;
	signal G1240: std_logic; attribute dont_touch of G1240: signal is true;
	signal G1243: std_logic; attribute dont_touch of G1243: signal is true;
	signal G1244: std_logic; attribute dont_touch of G1244: signal is true;
	signal G1245: std_logic; attribute dont_touch of G1245: signal is true;
	signal G1248: std_logic; attribute dont_touch of G1248: signal is true;
	signal G1250: std_logic; attribute dont_touch of G1250: signal is true;
	signal G1251: std_logic; attribute dont_touch of G1251: signal is true;
	signal G1252: std_logic; attribute dont_touch of G1252: signal is true;
	signal G1253: std_logic; attribute dont_touch of G1253: signal is true;
	signal G1254: std_logic; attribute dont_touch of G1254: signal is true;
	signal G1255: std_logic; attribute dont_touch of G1255: signal is true;
	signal G1256: std_logic; attribute dont_touch of G1256: signal is true;
	signal G1257: std_logic; attribute dont_touch of G1257: signal is true;
	signal G1258: std_logic; attribute dont_touch of G1258: signal is true;
	signal G1259: std_logic; attribute dont_touch of G1259: signal is true;
	signal G1260: std_logic; attribute dont_touch of G1260: signal is true;
	signal G1261: std_logic; attribute dont_touch of G1261: signal is true;
	signal G1262: std_logic; attribute dont_touch of G1262: signal is true;
	signal G1263: std_logic; attribute dont_touch of G1263: signal is true;
	signal G1264: std_logic; attribute dont_touch of G1264: signal is true;
	signal G1265: std_logic; attribute dont_touch of G1265: signal is true;
	signal G1266: std_logic; attribute dont_touch of G1266: signal is true;
	signal G1267: std_logic; attribute dont_touch of G1267: signal is true;
	signal G1268: std_logic; attribute dont_touch of G1268: signal is true;
	signal G1269: std_logic; attribute dont_touch of G1269: signal is true;
	signal G1270: std_logic; attribute dont_touch of G1270: signal is true;
	signal G1271: std_logic; attribute dont_touch of G1271: signal is true;
	signal G1272: std_logic; attribute dont_touch of G1272: signal is true;
	signal G1273: std_logic; attribute dont_touch of G1273: signal is true;
	signal G1276: std_logic; attribute dont_touch of G1276: signal is true;
	signal G1279: std_logic; attribute dont_touch of G1279: signal is true;
	signal G1282: std_logic; attribute dont_touch of G1282: signal is true;
	signal G1285: std_logic; attribute dont_touch of G1285: signal is true;
	signal G1288: std_logic; attribute dont_touch of G1288: signal is true;
	signal G1291: std_logic; attribute dont_touch of G1291: signal is true;
	signal G1294: std_logic; attribute dont_touch of G1294: signal is true;
	signal G1297: std_logic; attribute dont_touch of G1297: signal is true;
	signal G1300: std_logic; attribute dont_touch of G1300: signal is true;
	signal G1303: std_logic; attribute dont_touch of G1303: signal is true;
	signal G1306: std_logic; attribute dont_touch of G1306: signal is true;
	signal G1309: std_logic; attribute dont_touch of G1309: signal is true;
	signal G1312: std_logic; attribute dont_touch of G1312: signal is true;
	signal G1315: std_logic; attribute dont_touch of G1315: signal is true;
	signal G1316: std_logic; attribute dont_touch of G1316: signal is true;
	signal G1319: std_logic; attribute dont_touch of G1319: signal is true;
	signal G1326: std_logic; attribute dont_touch of G1326: signal is true;
	signal G1332: std_logic; attribute dont_touch of G1332: signal is true;
	signal G1339: std_logic; attribute dont_touch of G1339: signal is true;
	signal G1345: std_logic; attribute dont_touch of G1345: signal is true;
	signal G1346: std_logic; attribute dont_touch of G1346: signal is true;
	signal G1352: std_logic; attribute dont_touch of G1352: signal is true;
	signal G1358: std_logic; attribute dont_touch of G1358: signal is true;
	signal G1365: std_logic; attribute dont_touch of G1365: signal is true;
	signal G1372: std_logic; attribute dont_touch of G1372: signal is true;
	signal G1378: std_logic; attribute dont_touch of G1378: signal is true;
	signal G1384: std_logic; attribute dont_touch of G1384: signal is true;
	signal G1385: std_logic; attribute dont_touch of G1385: signal is true;
	signal G1386: std_logic; attribute dont_touch of G1386: signal is true;
	signal G1387: std_logic; attribute dont_touch of G1387: signal is true;
	signal G1388: std_logic; attribute dont_touch of G1388: signal is true;
	signal G1389: std_logic; attribute dont_touch of G1389: signal is true;
	signal G1390: std_logic; attribute dont_touch of G1390: signal is true;
	signal G1391: std_logic; attribute dont_touch of G1391: signal is true;
	signal G1392: std_logic; attribute dont_touch of G1392: signal is true;
	signal G1393: std_logic; attribute dont_touch of G1393: signal is true;
	signal G1394: std_logic; attribute dont_touch of G1394: signal is true;
	signal G1395: std_logic; attribute dont_touch of G1395: signal is true;
	signal G1396: std_logic; attribute dont_touch of G1396: signal is true;
	signal G1397: std_logic; attribute dont_touch of G1397: signal is true;
	signal G1398: std_logic; attribute dont_touch of G1398: signal is true;
	signal G1399: std_logic; attribute dont_touch of G1399: signal is true;
	signal G1400: std_logic; attribute dont_touch of G1400: signal is true;
	signal G1401: std_logic; attribute dont_touch of G1401: signal is true;
	signal G1402: std_logic; attribute dont_touch of G1402: signal is true;
	signal G1403: std_logic; attribute dont_touch of G1403: signal is true;
	signal G1404: std_logic; attribute dont_touch of G1404: signal is true;
	signal G1405: std_logic; attribute dont_touch of G1405: signal is true;
	signal G1406: std_logic; attribute dont_touch of G1406: signal is true;
	signal G1407: std_logic; attribute dont_touch of G1407: signal is true;
	signal G1408: std_logic; attribute dont_touch of G1408: signal is true;
	signal G1409: std_logic; attribute dont_touch of G1409: signal is true;
	signal G1410: std_logic; attribute dont_touch of G1410: signal is true;
	signal G1411: std_logic; attribute dont_touch of G1411: signal is true;
	signal G1412: std_logic; attribute dont_touch of G1412: signal is true;
	signal G1413: std_logic; attribute dont_touch of G1413: signal is true;
	signal G1414: std_logic; attribute dont_touch of G1414: signal is true;
	signal G1415: std_logic; attribute dont_touch of G1415: signal is true;
	signal G1416: std_logic; attribute dont_touch of G1416: signal is true;
	signal G1417: std_logic; attribute dont_touch of G1417: signal is true;
	signal G1418: std_logic; attribute dont_touch of G1418: signal is true;
	signal G1419: std_logic; attribute dont_touch of G1419: signal is true;
	signal G1420: std_logic; attribute dont_touch of G1420: signal is true;
	signal G1421: std_logic; attribute dont_touch of G1421: signal is true;
	signal G1422: std_logic; attribute dont_touch of G1422: signal is true;
	signal G1423: std_logic; attribute dont_touch of G1423: signal is true;
	signal G1424: std_logic; attribute dont_touch of G1424: signal is true;
	signal G1425: std_logic; attribute dont_touch of G1425: signal is true;
	signal G1426: std_logic; attribute dont_touch of G1426: signal is true;
	signal G1430: std_logic; attribute dont_touch of G1430: signal is true;
	signal G1435: std_logic; attribute dont_touch of G1435: signal is true;
	signal G1439: std_logic; attribute dont_touch of G1439: signal is true;
	signal G1444: std_logic; attribute dont_touch of G1444: signal is true;
	signal G1448: std_logic; attribute dont_touch of G1448: signal is true;
	signal G1453: std_logic; attribute dont_touch of G1453: signal is true;
	signal G1457: std_logic; attribute dont_touch of G1457: signal is true;
	signal G1462: std_logic; attribute dont_touch of G1462: signal is true;
	signal G1466: std_logic; attribute dont_touch of G1466: signal is true;
	signal G1471: std_logic; attribute dont_touch of G1471: signal is true;
	signal G1476: std_logic; attribute dont_touch of G1476: signal is true;
	signal G1481: std_logic; attribute dont_touch of G1481: signal is true;
	signal G1486: std_logic; attribute dont_touch of G1486: signal is true;
	signal G1491: std_logic; attribute dont_touch of G1491: signal is true;
	signal G1496: std_logic; attribute dont_touch of G1496: signal is true;
	signal G1501: std_logic; attribute dont_touch of G1501: signal is true;
	signal G1506: std_logic; attribute dont_touch of G1506: signal is true;
	signal G1511: std_logic; attribute dont_touch of G1511: signal is true;
	signal G1512: std_logic; attribute dont_touch of G1512: signal is true;
	signal G1513: std_logic; attribute dont_touch of G1513: signal is true;
	signal G1514: std_logic; attribute dont_touch of G1514: signal is true;
	signal G1515: std_logic; attribute dont_touch of G1515: signal is true;
	signal G1516: std_logic; attribute dont_touch of G1516: signal is true;
	signal G1517: std_logic; attribute dont_touch of G1517: signal is true;
	signal G1520: std_logic; attribute dont_touch of G1520: signal is true;
	signal G1523: std_logic; attribute dont_touch of G1523: signal is true;
	signal G1524: std_logic; attribute dont_touch of G1524: signal is true;
	signal G1525: std_logic; attribute dont_touch of G1525: signal is true;
	signal G1526: std_logic; attribute dont_touch of G1526: signal is true;
	signal G1527: std_logic; attribute dont_touch of G1527: signal is true;
	signal G1528: std_logic; attribute dont_touch of G1528: signal is true;
	signal G1529: std_logic; attribute dont_touch of G1529: signal is true;
	signal G1530: std_logic; attribute dont_touch of G1530: signal is true;
	signal G1531: std_logic; attribute dont_touch of G1531: signal is true;
	signal G1532: std_logic; attribute dont_touch of G1532: signal is true;
	signal G1533: std_logic; attribute dont_touch of G1533: signal is true;
	signal G1534: std_logic; attribute dont_touch of G1534: signal is true;
	signal G1535: std_logic; attribute dont_touch of G1535: signal is true;
	signal G1536: std_logic; attribute dont_touch of G1536: signal is true;
	signal G1537: std_logic; attribute dont_touch of G1537: signal is true;
	signal G1538: std_logic; attribute dont_touch of G1538: signal is true;
	signal G1539: std_logic; attribute dont_touch of G1539: signal is true;
	signal G1540: std_logic; attribute dont_touch of G1540: signal is true;
	signal G1541: std_logic; attribute dont_touch of G1541: signal is true;
	signal G1542: std_logic; attribute dont_touch of G1542: signal is true;
	signal G1543: std_logic; attribute dont_touch of G1543: signal is true;
	signal G1544: std_logic; attribute dont_touch of G1544: signal is true;
	signal G1545: std_logic; attribute dont_touch of G1545: signal is true;
	signal G1546: std_logic; attribute dont_touch of G1546: signal is true;
	signal G1547: std_logic; attribute dont_touch of G1547: signal is true;
	signal G1550: std_logic; attribute dont_touch of G1550: signal is true;
	signal G1551: std_logic; attribute dont_touch of G1551: signal is true;
	signal G1552: std_logic; attribute dont_touch of G1552: signal is true;
	signal G1553: std_logic; attribute dont_touch of G1553: signal is true;
	signal G1554: std_logic; attribute dont_touch of G1554: signal is true;
	signal G1555: std_logic; attribute dont_touch of G1555: signal is true;
	signal G1556: std_logic; attribute dont_touch of G1556: signal is true;
	signal G1557: std_logic; attribute dont_touch of G1557: signal is true;
	signal G1558: std_logic; attribute dont_touch of G1558: signal is true;
	signal G1559: std_logic; attribute dont_touch of G1559: signal is true;
	signal G1560: std_logic; attribute dont_touch of G1560: signal is true;
	signal G1561: std_logic; attribute dont_touch of G1561: signal is true;
	signal G1562: std_logic; attribute dont_touch of G1562: signal is true;
	signal G1563: std_logic; attribute dont_touch of G1563: signal is true;
	signal G1564: std_logic; attribute dont_touch of G1564: signal is true;
	signal G1567: std_logic; attribute dont_touch of G1567: signal is true;
	signal G1570: std_logic; attribute dont_touch of G1570: signal is true;
	signal G1573: std_logic; attribute dont_touch of G1573: signal is true;
	signal G1576: std_logic; attribute dont_touch of G1576: signal is true;
	signal G1579: std_logic; attribute dont_touch of G1579: signal is true;
	signal G1582: std_logic; attribute dont_touch of G1582: signal is true;
	signal G1585: std_logic; attribute dont_touch of G1585: signal is true;
	signal G1588: std_logic; attribute dont_touch of G1588: signal is true;
	signal G1591: std_logic; attribute dont_touch of G1591: signal is true;
	signal G1594: std_logic; attribute dont_touch of G1594: signal is true;
	signal G1597: std_logic; attribute dont_touch of G1597: signal is true;
	signal G1600: std_logic; attribute dont_touch of G1600: signal is true;
	signal G1603: std_logic; attribute dont_touch of G1603: signal is true;
	signal G1606: std_logic; attribute dont_touch of G1606: signal is true;
	signal G1609: std_logic; attribute dont_touch of G1609: signal is true;
	signal G1612: std_logic; attribute dont_touch of G1612: signal is true;
	signal G1615: std_logic; attribute dont_touch of G1615: signal is true;
	signal G1618: std_logic; attribute dont_touch of G1618: signal is true;
	signal G1621: std_logic; attribute dont_touch of G1621: signal is true;
	signal G1624: std_logic; attribute dont_touch of G1624: signal is true;
	signal G1627: std_logic; attribute dont_touch of G1627: signal is true;
	signal G1630: std_logic; attribute dont_touch of G1630: signal is true;
	signal G1633: std_logic; attribute dont_touch of G1633: signal is true;
	signal G1636: std_logic; attribute dont_touch of G1636: signal is true;
	signal G1639: std_logic; attribute dont_touch of G1639: signal is true;
	signal G1642: std_logic; attribute dont_touch of G1642: signal is true;
	signal G1645: std_logic; attribute dont_touch of G1645: signal is true;
	signal G1648: std_logic; attribute dont_touch of G1648: signal is true;
	signal G1651: std_logic; attribute dont_touch of G1651: signal is true;
	signal G1654: std_logic; attribute dont_touch of G1654: signal is true;
	signal G1657: std_logic; attribute dont_touch of G1657: signal is true;
	signal G1660: std_logic; attribute dont_touch of G1660: signal is true;
	signal G1661: std_logic; attribute dont_touch of G1661: signal is true;
	signal G1662: std_logic; attribute dont_touch of G1662: signal is true;
	signal G1663: std_logic; attribute dont_touch of G1663: signal is true;
	signal G1664: std_logic; attribute dont_touch of G1664: signal is true;
	signal G1665: std_logic; attribute dont_touch of G1665: signal is true;
	signal G1666: std_logic; attribute dont_touch of G1666: signal is true;
	signal G1667: std_logic; attribute dont_touch of G1667: signal is true;
	signal G1668: std_logic; attribute dont_touch of G1668: signal is true;
	signal G1669: std_logic; attribute dont_touch of G1669: signal is true;
	signal G1670: std_logic; attribute dont_touch of G1670: signal is true;
	signal G1671: std_logic; attribute dont_touch of G1671: signal is true;
	signal G1672: std_logic; attribute dont_touch of G1672: signal is true;
	signal G1675: std_logic; attribute dont_touch of G1675: signal is true;
	signal G1676: std_logic; attribute dont_touch of G1676: signal is true;
	signal G1677: std_logic; attribute dont_touch of G1677: signal is true;
	signal G1678: std_logic; attribute dont_touch of G1678: signal is true;
	signal G1679: std_logic; attribute dont_touch of G1679: signal is true;
	signal G1680: std_logic; attribute dont_touch of G1680: signal is true;
	signal G1681: std_logic; attribute dont_touch of G1681: signal is true;
	signal G1682: std_logic; attribute dont_touch of G1682: signal is true;
	signal G1683: std_logic; attribute dont_touch of G1683: signal is true;
	signal G1684: std_logic; attribute dont_touch of G1684: signal is true;
	signal G1685: std_logic; attribute dont_touch of G1685: signal is true;
	signal G1686: std_logic; attribute dont_touch of G1686: signal is true;
	signal G1689: std_logic; attribute dont_touch of G1689: signal is true;
	signal G1690: std_logic; attribute dont_touch of G1690: signal is true;
	signal G1693: std_logic; attribute dont_touch of G1693: signal is true;
	signal G1694: std_logic; attribute dont_touch of G1694: signal is true;
	signal G1695: std_logic; attribute dont_touch of G1695: signal is true;
	signal G1696: std_logic; attribute dont_touch of G1696: signal is true;
	signal G1697: std_logic; attribute dont_touch of G1697: signal is true;
	signal G1698: std_logic; attribute dont_touch of G1698: signal is true;
	signal G1699: std_logic; attribute dont_touch of G1699: signal is true;
	signal G1700: std_logic; attribute dont_touch of G1700: signal is true;
	signal G1701: std_logic; attribute dont_touch of G1701: signal is true;
	signal G1702: std_logic; attribute dont_touch of G1702: signal is true;
	signal G1703: std_logic; attribute dont_touch of G1703: signal is true;
	signal G1704: std_logic; attribute dont_touch of G1704: signal is true;
	signal G1705: std_logic; attribute dont_touch of G1705: signal is true;
	signal G1706: std_logic; attribute dont_touch of G1706: signal is true;
	signal G1712: std_logic; attribute dont_touch of G1712: signal is true;
	signal G1718: std_logic; attribute dont_touch of G1718: signal is true;
	signal G1723: std_logic; attribute dont_touch of G1723: signal is true;
	signal G1724: std_logic; attribute dont_touch of G1724: signal is true;
	signal G1727: std_logic; attribute dont_touch of G1727: signal is true;
	signal G1730: std_logic; attribute dont_touch of G1730: signal is true;
	signal G1731: std_logic; attribute dont_touch of G1731: signal is true;
	signal G1732: std_logic; attribute dont_touch of G1732: signal is true;
	signal G1733: std_logic; attribute dont_touch of G1733: signal is true;
	signal G1734: std_logic; attribute dont_touch of G1734: signal is true;
	signal G1735: std_logic; attribute dont_touch of G1735: signal is true;
	signal G1738: std_logic; attribute dont_touch of G1738: signal is true;
	signal G1739: std_logic; attribute dont_touch of G1739: signal is true;
	signal G1742: std_logic; attribute dont_touch of G1742: signal is true;
	signal G1745: std_logic; attribute dont_touch of G1745: signal is true;
	signal G1746: std_logic; attribute dont_touch of G1746: signal is true;
	signal G1747: std_logic; attribute dont_touch of G1747: signal is true;
	signal G1748: std_logic; attribute dont_touch of G1748: signal is true;
	signal G1749: std_logic; attribute dont_touch of G1749: signal is true;
	signal G1750: std_logic; attribute dont_touch of G1750: signal is true;
	signal G1753: std_logic; attribute dont_touch of G1753: signal is true;
	signal G1754: std_logic; attribute dont_touch of G1754: signal is true;
	signal G1757: std_logic; attribute dont_touch of G1757: signal is true;
	signal G1760: std_logic; attribute dont_touch of G1760: signal is true;
	signal G1761: std_logic; attribute dont_touch of G1761: signal is true;
	signal G1762: std_logic; attribute dont_touch of G1762: signal is true;
	signal G1763: std_logic; attribute dont_touch of G1763: signal is true;
	signal G1764: std_logic; attribute dont_touch of G1764: signal is true;
	signal G1765: std_logic; attribute dont_touch of G1765: signal is true;
	signal G1768: std_logic; attribute dont_touch of G1768: signal is true;
	signal G1769: std_logic; attribute dont_touch of G1769: signal is true;
	signal G1772: std_logic; attribute dont_touch of G1772: signal is true;
	signal G1775: std_logic; attribute dont_touch of G1775: signal is true;
	signal G1776: std_logic; attribute dont_touch of G1776: signal is true;
	signal G1777: std_logic; attribute dont_touch of G1777: signal is true;
	signal G1778: std_logic; attribute dont_touch of G1778: signal is true;
	signal G1779: std_logic; attribute dont_touch of G1779: signal is true;
	signal G1782: std_logic; attribute dont_touch of G1782: signal is true;
	signal G1783: std_logic; attribute dont_touch of G1783: signal is true;
	signal G1784: std_logic; attribute dont_touch of G1784: signal is true;
	signal G1785: std_logic; attribute dont_touch of G1785: signal is true;
	signal G1786: std_logic; attribute dont_touch of G1786: signal is true;
	signal G1789: std_logic; attribute dont_touch of G1789: signal is true;
	signal G1792: std_logic; attribute dont_touch of G1792: signal is true;
	signal G1795: std_logic; attribute dont_touch of G1795: signal is true;
	signal G1798: std_logic; attribute dont_touch of G1798: signal is true;
	signal G1801: std_logic; attribute dont_touch of G1801: signal is true;
	signal G1804: std_logic; attribute dont_touch of G1804: signal is true;
	signal G1807: std_logic; attribute dont_touch of G1807: signal is true;
	signal G1808: std_logic; attribute dont_touch of G1808: signal is true;
	signal G1809: std_logic; attribute dont_touch of G1809: signal is true;
	signal G1810: std_logic; attribute dont_touch of G1810: signal is true;
	signal G1813: std_logic; attribute dont_touch of G1813: signal is true;
	signal G1816: std_logic; attribute dont_touch of G1816: signal is true;
	signal G1819: std_logic; attribute dont_touch of G1819: signal is true;
	signal G1822: std_logic; attribute dont_touch of G1822: signal is true;
	signal G1825: std_logic; attribute dont_touch of G1825: signal is true;
	signal G1828: std_logic; attribute dont_touch of G1828: signal is true;
	signal G1829: std_logic; attribute dont_touch of G1829: signal is true;
	signal G1830: std_logic; attribute dont_touch of G1830: signal is true;
	signal G1831: std_logic; attribute dont_touch of G1831: signal is true;
	signal G1832: std_logic; attribute dont_touch of G1832: signal is true;
	signal G1833: std_logic; attribute dont_touch of G1833: signal is true;
	signal G1834: std_logic; attribute dont_touch of G1834: signal is true;
	signal G1835: std_logic; attribute dont_touch of G1835: signal is true;
	signal G1836: std_logic; attribute dont_touch of G1836: signal is true;
	signal G1839: std_logic; attribute dont_touch of G1839: signal is true;
	signal G1842: std_logic; attribute dont_touch of G1842: signal is true;
	signal G1845: std_logic; attribute dont_touch of G1845: signal is true;
	signal G1846: std_logic; attribute dont_touch of G1846: signal is true;
	signal G1849: std_logic; attribute dont_touch of G1849: signal is true;
	signal G1852: std_logic; attribute dont_touch of G1852: signal is true;
	signal G1855: std_logic; attribute dont_touch of G1855: signal is true;
	signal G1858: std_logic; attribute dont_touch of G1858: signal is true;
	signal G1859: std_logic; attribute dont_touch of G1859: signal is true;
	signal G1860: std_logic; attribute dont_touch of G1860: signal is true;
	signal G1861: std_logic; attribute dont_touch of G1861: signal is true;
	signal G1862: std_logic; attribute dont_touch of G1862: signal is true;
	signal G1865: std_logic; attribute dont_touch of G1865: signal is true;
	signal G1866: std_logic; attribute dont_touch of G1866: signal is true;
	signal G1867: std_logic; attribute dont_touch of G1867: signal is true;
	signal G1868: std_logic; attribute dont_touch of G1868: signal is true;
	signal G1869: std_logic; attribute dont_touch of G1869: signal is true;
	signal G1870: std_logic; attribute dont_touch of G1870: signal is true;
	signal G1871: std_logic; attribute dont_touch of G1871: signal is true;
	signal G1874: std_logic; attribute dont_touch of G1874: signal is true;
	signal G1877: std_logic; attribute dont_touch of G1877: signal is true;
	signal G1880: std_logic; attribute dont_touch of G1880: signal is true;
	signal G1886: std_logic; attribute dont_touch of G1886: signal is true;
	signal G1887: std_logic; attribute dont_touch of G1887: signal is true;
	signal G1888: std_logic; attribute dont_touch of G1888: signal is true;
	signal G1889: std_logic; attribute dont_touch of G1889: signal is true;
	signal G1890: std_logic; attribute dont_touch of G1890: signal is true;
	signal G1893: std_logic; attribute dont_touch of G1893: signal is true;
	signal G1894: std_logic; attribute dont_touch of G1894: signal is true;
	signal G1895: std_logic; attribute dont_touch of G1895: signal is true;
	signal G1896: std_logic; attribute dont_touch of G1896: signal is true;
	signal G1897: std_logic; attribute dont_touch of G1897: signal is true;
	signal G1898: std_logic; attribute dont_touch of G1898: signal is true;
	signal G1899: std_logic; attribute dont_touch of G1899: signal is true;
	signal G1900: std_logic; attribute dont_touch of G1900: signal is true;
	signal G1903: std_logic; attribute dont_touch of G1903: signal is true;
	signal G1904: std_logic; attribute dont_touch of G1904: signal is true;
	signal G1905: std_logic; attribute dont_touch of G1905: signal is true;
	signal G1908: std_logic; attribute dont_touch of G1908: signal is true;
	signal G1909: std_logic; attribute dont_touch of G1909: signal is true;
	signal G1910: std_logic; attribute dont_touch of G1910: signal is true;
	signal G1911: std_logic; attribute dont_touch of G1911: signal is true;
	signal G1912: std_logic; attribute dont_touch of G1912: signal is true;
	signal G1913: std_logic; attribute dont_touch of G1913: signal is true;
	signal G1914: std_logic; attribute dont_touch of G1914: signal is true;
	signal G1915: std_logic; attribute dont_touch of G1915: signal is true;
	signal G1916: std_logic; attribute dont_touch of G1916: signal is true;
	signal G1917: std_logic; attribute dont_touch of G1917: signal is true;
	signal G1918: std_logic; attribute dont_touch of G1918: signal is true;
	signal G1921: std_logic; attribute dont_touch of G1921: signal is true;
	signal G1922: std_logic; attribute dont_touch of G1922: signal is true;
	signal G1923: std_logic; attribute dont_touch of G1923: signal is true;
	signal G1924: std_logic; attribute dont_touch of G1924: signal is true;
	signal G1925: std_logic; attribute dont_touch of G1925: signal is true;
	signal G1928: std_logic; attribute dont_touch of G1928: signal is true;
	signal G1929: std_logic; attribute dont_touch of G1929: signal is true;
	signal G1930: std_logic; attribute dont_touch of G1930: signal is true;
	signal G1931: std_logic; attribute dont_touch of G1931: signal is true;
	signal G1934: std_logic; attribute dont_touch of G1934: signal is true;
	signal G1937: std_logic; attribute dont_touch of G1937: signal is true;
	signal G1938: std_logic; attribute dont_touch of G1938: signal is true;
	signal G1939: std_logic; attribute dont_touch of G1939: signal is true;
	signal G1942: std_logic; attribute dont_touch of G1942: signal is true;
	signal G1944: std_logic; attribute dont_touch of G1944: signal is true;
	signal G1945: std_logic; attribute dont_touch of G1945: signal is true;
	signal G1946: std_logic; attribute dont_touch of G1946: signal is true;
	signal G1947: std_logic; attribute dont_touch of G1947: signal is true;
	signal G1948: std_logic; attribute dont_touch of G1948: signal is true;
	signal G1949: std_logic; attribute dont_touch of G1949: signal is true;
	signal G1950: std_logic; attribute dont_touch of G1950: signal is true;
	signal G1951: std_logic; attribute dont_touch of G1951: signal is true;
	signal G1952: std_logic; attribute dont_touch of G1952: signal is true;
	signal G1953: std_logic; attribute dont_touch of G1953: signal is true;
	signal G1954: std_logic; attribute dont_touch of G1954: signal is true;
	signal G1955: std_logic; attribute dont_touch of G1955: signal is true;
	signal G1956: std_logic; attribute dont_touch of G1956: signal is true;
	signal G1957: std_logic; attribute dont_touch of G1957: signal is true;
	signal G1958: std_logic; attribute dont_touch of G1958: signal is true;
	signal G1959: std_logic; attribute dont_touch of G1959: signal is true;
	signal G1960: std_logic; attribute dont_touch of G1960: signal is true;
	signal G1961: std_logic; attribute dont_touch of G1961: signal is true;
	signal G1962: std_logic; attribute dont_touch of G1962: signal is true;
	signal G1963: std_logic; attribute dont_touch of G1963: signal is true;
	signal G1964: std_logic; attribute dont_touch of G1964: signal is true;
	signal G1965: std_logic; attribute dont_touch of G1965: signal is true;
	signal G1966: std_logic; attribute dont_touch of G1966: signal is true;
	signal G1967: std_logic; attribute dont_touch of G1967: signal is true;
	signal G1970: std_logic; attribute dont_touch of G1970: signal is true;
	signal G1973: std_logic; attribute dont_touch of G1973: signal is true;
	signal G1976: std_logic; attribute dont_touch of G1976: signal is true;
	signal G1979: std_logic; attribute dont_touch of G1979: signal is true;
	signal G1982: std_logic; attribute dont_touch of G1982: signal is true;
	signal G1985: std_logic; attribute dont_touch of G1985: signal is true;
	signal G1988: std_logic; attribute dont_touch of G1988: signal is true;
	signal G1991: std_logic; attribute dont_touch of G1991: signal is true;
	signal G1994: std_logic; attribute dont_touch of G1994: signal is true;
	signal G1997: std_logic; attribute dont_touch of G1997: signal is true;
	signal G2000: std_logic; attribute dont_touch of G2000: signal is true;
	signal G2003: std_logic; attribute dont_touch of G2003: signal is true;
	signal G2006: std_logic; attribute dont_touch of G2006: signal is true;
	signal G2009: std_logic; attribute dont_touch of G2009: signal is true;
	signal G2010: std_logic; attribute dont_touch of G2010: signal is true;
	signal G2013: std_logic; attribute dont_touch of G2013: signal is true;
	signal G2020: std_logic; attribute dont_touch of G2020: signal is true;
	signal G2026: std_logic; attribute dont_touch of G2026: signal is true;
	signal G2033: std_logic; attribute dont_touch of G2033: signal is true;
	signal G2039: std_logic; attribute dont_touch of G2039: signal is true;
	signal G2040: std_logic; attribute dont_touch of G2040: signal is true;
	signal G2046: std_logic; attribute dont_touch of G2046: signal is true;
	signal G2052: std_logic; attribute dont_touch of G2052: signal is true;
	signal G2059: std_logic; attribute dont_touch of G2059: signal is true;
	signal G2066: std_logic; attribute dont_touch of G2066: signal is true;
	signal G2072: std_logic; attribute dont_touch of G2072: signal is true;
	signal G2078: std_logic; attribute dont_touch of G2078: signal is true;
	signal G2079: std_logic; attribute dont_touch of G2079: signal is true;
	signal G2080: std_logic; attribute dont_touch of G2080: signal is true;
	signal G2081: std_logic; attribute dont_touch of G2081: signal is true;
	signal G2082: std_logic; attribute dont_touch of G2082: signal is true;
	signal G2083: std_logic; attribute dont_touch of G2083: signal is true;
	signal G2084: std_logic; attribute dont_touch of G2084: signal is true;
	signal G2085: std_logic; attribute dont_touch of G2085: signal is true;
	signal G2086: std_logic; attribute dont_touch of G2086: signal is true;
	signal G2087: std_logic; attribute dont_touch of G2087: signal is true;
	signal G2088: std_logic; attribute dont_touch of G2088: signal is true;
	signal G2089: std_logic; attribute dont_touch of G2089: signal is true;
	signal G2090: std_logic; attribute dont_touch of G2090: signal is true;
	signal G2091: std_logic; attribute dont_touch of G2091: signal is true;
	signal G2092: std_logic; attribute dont_touch of G2092: signal is true;
	signal G2093: std_logic; attribute dont_touch of G2093: signal is true;
	signal G2094: std_logic; attribute dont_touch of G2094: signal is true;
	signal G2095: std_logic; attribute dont_touch of G2095: signal is true;
	signal G2096: std_logic; attribute dont_touch of G2096: signal is true;
	signal G2097: std_logic; attribute dont_touch of G2097: signal is true;
	signal G2098: std_logic; attribute dont_touch of G2098: signal is true;
	signal G2099: std_logic; attribute dont_touch of G2099: signal is true;
	signal G2100: std_logic; attribute dont_touch of G2100: signal is true;
	signal G2101: std_logic; attribute dont_touch of G2101: signal is true;
	signal G2102: std_logic; attribute dont_touch of G2102: signal is true;
	signal G2103: std_logic; attribute dont_touch of G2103: signal is true;
	signal G2104: std_logic; attribute dont_touch of G2104: signal is true;
	signal G2105: std_logic; attribute dont_touch of G2105: signal is true;
	signal G2106: std_logic; attribute dont_touch of G2106: signal is true;
	signal G2107: std_logic; attribute dont_touch of G2107: signal is true;
	signal G2108: std_logic; attribute dont_touch of G2108: signal is true;
	signal G2109: std_logic; attribute dont_touch of G2109: signal is true;
	signal G2110: std_logic; attribute dont_touch of G2110: signal is true;
	signal G2111: std_logic; attribute dont_touch of G2111: signal is true;
	signal G2112: std_logic; attribute dont_touch of G2112: signal is true;
	signal G2113: std_logic; attribute dont_touch of G2113: signal is true;
	signal G2114: std_logic; attribute dont_touch of G2114: signal is true;
	signal G2115: std_logic; attribute dont_touch of G2115: signal is true;
	signal G2116: std_logic; attribute dont_touch of G2116: signal is true;
	signal G2117: std_logic; attribute dont_touch of G2117: signal is true;
	signal G2118: std_logic; attribute dont_touch of G2118: signal is true;
	signal G2119: std_logic; attribute dont_touch of G2119: signal is true;
	signal G2120: std_logic; attribute dont_touch of G2120: signal is true;
	signal G2124: std_logic; attribute dont_touch of G2124: signal is true;
	signal G2129: std_logic; attribute dont_touch of G2129: signal is true;
	signal G2133: std_logic; attribute dont_touch of G2133: signal is true;
	signal G2138: std_logic; attribute dont_touch of G2138: signal is true;
	signal G2142: std_logic; attribute dont_touch of G2142: signal is true;
	signal G2147: std_logic; attribute dont_touch of G2147: signal is true;
	signal G2151: std_logic; attribute dont_touch of G2151: signal is true;
	signal G2156: std_logic; attribute dont_touch of G2156: signal is true;
	signal G2160: std_logic; attribute dont_touch of G2160: signal is true;
	signal G2165: std_logic; attribute dont_touch of G2165: signal is true;
	signal G2170: std_logic; attribute dont_touch of G2170: signal is true;
	signal G2175: std_logic; attribute dont_touch of G2175: signal is true;
	signal G2180: std_logic; attribute dont_touch of G2180: signal is true;
	signal G2185: std_logic; attribute dont_touch of G2185: signal is true;
	signal G2190: std_logic; attribute dont_touch of G2190: signal is true;
	signal G2195: std_logic; attribute dont_touch of G2195: signal is true;
	signal G2200: std_logic; attribute dont_touch of G2200: signal is true;
	signal G2205: std_logic; attribute dont_touch of G2205: signal is true;
	signal G2206: std_logic; attribute dont_touch of G2206: signal is true;
	signal G2207: std_logic; attribute dont_touch of G2207: signal is true;
	signal G2208: std_logic; attribute dont_touch of G2208: signal is true;
	signal G2209: std_logic; attribute dont_touch of G2209: signal is true;
	signal G2210: std_logic; attribute dont_touch of G2210: signal is true;
	signal G2211: std_logic; attribute dont_touch of G2211: signal is true;
	signal G2214: std_logic; attribute dont_touch of G2214: signal is true;
	signal G2217: std_logic; attribute dont_touch of G2217: signal is true;
	signal G2218: std_logic; attribute dont_touch of G2218: signal is true;
	signal G2219: std_logic; attribute dont_touch of G2219: signal is true;
	signal G2220: std_logic; attribute dont_touch of G2220: signal is true;
	signal G2221: std_logic; attribute dont_touch of G2221: signal is true;
	signal G2222: std_logic; attribute dont_touch of G2222: signal is true;
	signal G2223: std_logic; attribute dont_touch of G2223: signal is true;
	signal G2224: std_logic; attribute dont_touch of G2224: signal is true;
	signal G2225: std_logic; attribute dont_touch of G2225: signal is true;
	signal G2226: std_logic; attribute dont_touch of G2226: signal is true;
	signal G2227: std_logic; attribute dont_touch of G2227: signal is true;
	signal G2228: std_logic; attribute dont_touch of G2228: signal is true;
	signal G2229: std_logic; attribute dont_touch of G2229: signal is true;
	signal G2230: std_logic; attribute dont_touch of G2230: signal is true;
	signal G2231: std_logic; attribute dont_touch of G2231: signal is true;
	signal G2232: std_logic; attribute dont_touch of G2232: signal is true;
	signal G2233: std_logic; attribute dont_touch of G2233: signal is true;
	signal G2234: std_logic; attribute dont_touch of G2234: signal is true;
	signal G2235: std_logic; attribute dont_touch of G2235: signal is true;
	signal G2236: std_logic; attribute dont_touch of G2236: signal is true;
	signal G2237: std_logic; attribute dont_touch of G2237: signal is true;
	signal G2238: std_logic; attribute dont_touch of G2238: signal is true;
	signal G2239: std_logic; attribute dont_touch of G2239: signal is true;
	signal G2240: std_logic; attribute dont_touch of G2240: signal is true;
	signal G2241: std_logic; attribute dont_touch of G2241: signal is true;
	signal G2244: std_logic; attribute dont_touch of G2244: signal is true;
	signal G2245: std_logic; attribute dont_touch of G2245: signal is true;
	signal G2246: std_logic; attribute dont_touch of G2246: signal is true;
	signal G2247: std_logic; attribute dont_touch of G2247: signal is true;
	signal G2248: std_logic; attribute dont_touch of G2248: signal is true;
	signal G2249: std_logic; attribute dont_touch of G2249: signal is true;
	signal G2250: std_logic; attribute dont_touch of G2250: signal is true;
	signal G2251: std_logic; attribute dont_touch of G2251: signal is true;
	signal G2252: std_logic; attribute dont_touch of G2252: signal is true;
	signal G2253: std_logic; attribute dont_touch of G2253: signal is true;
	signal G2254: std_logic; attribute dont_touch of G2254: signal is true;
	signal G2255: std_logic; attribute dont_touch of G2255: signal is true;
	signal G2256: std_logic; attribute dont_touch of G2256: signal is true;
	signal G2257: std_logic; attribute dont_touch of G2257: signal is true;
	signal G2258: std_logic; attribute dont_touch of G2258: signal is true;
	signal G2261: std_logic; attribute dont_touch of G2261: signal is true;
	signal G2264: std_logic; attribute dont_touch of G2264: signal is true;
	signal G2267: std_logic; attribute dont_touch of G2267: signal is true;
	signal G2270: std_logic; attribute dont_touch of G2270: signal is true;
	signal G2273: std_logic; attribute dont_touch of G2273: signal is true;
	signal G2276: std_logic; attribute dont_touch of G2276: signal is true;
	signal G2279: std_logic; attribute dont_touch of G2279: signal is true;
	signal G2282: std_logic; attribute dont_touch of G2282: signal is true;
	signal G2285: std_logic; attribute dont_touch of G2285: signal is true;
	signal G2288: std_logic; attribute dont_touch of G2288: signal is true;
	signal G2291: std_logic; attribute dont_touch of G2291: signal is true;
	signal G2294: std_logic; attribute dont_touch of G2294: signal is true;
	signal G2297: std_logic; attribute dont_touch of G2297: signal is true;
	signal G2300: std_logic; attribute dont_touch of G2300: signal is true;
	signal G2303: std_logic; attribute dont_touch of G2303: signal is true;
	signal G2306: std_logic; attribute dont_touch of G2306: signal is true;
	signal G2309: std_logic; attribute dont_touch of G2309: signal is true;
	signal G2312: std_logic; attribute dont_touch of G2312: signal is true;
	signal G2315: std_logic; attribute dont_touch of G2315: signal is true;
	signal G2318: std_logic; attribute dont_touch of G2318: signal is true;
	signal G2321: std_logic; attribute dont_touch of G2321: signal is true;
	signal G2324: std_logic; attribute dont_touch of G2324: signal is true;
	signal G2327: std_logic; attribute dont_touch of G2327: signal is true;
	signal G2330: std_logic; attribute dont_touch of G2330: signal is true;
	signal G2333: std_logic; attribute dont_touch of G2333: signal is true;
	signal G2336: std_logic; attribute dont_touch of G2336: signal is true;
	signal G2339: std_logic; attribute dont_touch of G2339: signal is true;
	signal G2342: std_logic; attribute dont_touch of G2342: signal is true;
	signal G2345: std_logic; attribute dont_touch of G2345: signal is true;
	signal G2348: std_logic; attribute dont_touch of G2348: signal is true;
	signal G2351: std_logic; attribute dont_touch of G2351: signal is true;
	signal G2354: std_logic; attribute dont_touch of G2354: signal is true;
	signal G2355: std_logic; attribute dont_touch of G2355: signal is true;
	signal G2356: std_logic; attribute dont_touch of G2356: signal is true;
	signal G2357: std_logic; attribute dont_touch of G2357: signal is true;
	signal G2358: std_logic; attribute dont_touch of G2358: signal is true;
	signal G2359: std_logic; attribute dont_touch of G2359: signal is true;
	signal G2360: std_logic; attribute dont_touch of G2360: signal is true;
	signal G2361: std_logic; attribute dont_touch of G2361: signal is true;
	signal G2362: std_logic; attribute dont_touch of G2362: signal is true;
	signal G2363: std_logic; attribute dont_touch of G2363: signal is true;
	signal G2364: std_logic; attribute dont_touch of G2364: signal is true;
	signal G2365: std_logic; attribute dont_touch of G2365: signal is true;
	signal G2366: std_logic; attribute dont_touch of G2366: signal is true;
	signal G2369: std_logic; attribute dont_touch of G2369: signal is true;
	signal G2370: std_logic; attribute dont_touch of G2370: signal is true;
	signal G2371: std_logic; attribute dont_touch of G2371: signal is true;
	signal G2372: std_logic; attribute dont_touch of G2372: signal is true;
	signal G2373: std_logic; attribute dont_touch of G2373: signal is true;
	signal G2374: std_logic; attribute dont_touch of G2374: signal is true;
	signal G2375: std_logic; attribute dont_touch of G2375: signal is true;
	signal G2376: std_logic; attribute dont_touch of G2376: signal is true;
	signal G2377: std_logic; attribute dont_touch of G2377: signal is true;
	signal G2378: std_logic; attribute dont_touch of G2378: signal is true;
	signal G2379: std_logic; attribute dont_touch of G2379: signal is true;
	signal G2380: std_logic; attribute dont_touch of G2380: signal is true;
	signal G2383: std_logic; attribute dont_touch of G2383: signal is true;
	signal G2384: std_logic; attribute dont_touch of G2384: signal is true;
	signal G2387: std_logic; attribute dont_touch of G2387: signal is true;
	signal G2388: std_logic; attribute dont_touch of G2388: signal is true;
	signal G2389: std_logic; attribute dont_touch of G2389: signal is true;
	signal G2390: std_logic; attribute dont_touch of G2390: signal is true;
	signal G2391: std_logic; attribute dont_touch of G2391: signal is true;
	signal G2392: std_logic; attribute dont_touch of G2392: signal is true;
	signal G2393: std_logic; attribute dont_touch of G2393: signal is true;
	signal G2394: std_logic; attribute dont_touch of G2394: signal is true;
	signal G2395: std_logic; attribute dont_touch of G2395: signal is true;
	signal G2396: std_logic; attribute dont_touch of G2396: signal is true;
	signal G2397: std_logic; attribute dont_touch of G2397: signal is true;
	signal G2398: std_logic; attribute dont_touch of G2398: signal is true;
	signal G2399: std_logic; attribute dont_touch of G2399: signal is true;
	signal G2400: std_logic; attribute dont_touch of G2400: signal is true;
	signal G2406: std_logic; attribute dont_touch of G2406: signal is true;
	signal G2412: std_logic; attribute dont_touch of G2412: signal is true;
	signal G2417: std_logic; attribute dont_touch of G2417: signal is true;
	signal G2418: std_logic; attribute dont_touch of G2418: signal is true;
	signal G2421: std_logic; attribute dont_touch of G2421: signal is true;
	signal G2424: std_logic; attribute dont_touch of G2424: signal is true;
	signal G2425: std_logic; attribute dont_touch of G2425: signal is true;
	signal G2426: std_logic; attribute dont_touch of G2426: signal is true;
	signal G2427: std_logic; attribute dont_touch of G2427: signal is true;
	signal G2428: std_logic; attribute dont_touch of G2428: signal is true;
	signal G2429: std_logic; attribute dont_touch of G2429: signal is true;
	signal G2432: std_logic; attribute dont_touch of G2432: signal is true;
	signal G2433: std_logic; attribute dont_touch of G2433: signal is true;
	signal G2436: std_logic; attribute dont_touch of G2436: signal is true;
	signal G2439: std_logic; attribute dont_touch of G2439: signal is true;
	signal G2440: std_logic; attribute dont_touch of G2440: signal is true;
	signal G2441: std_logic; attribute dont_touch of G2441: signal is true;
	signal G2442: std_logic; attribute dont_touch of G2442: signal is true;
	signal G2443: std_logic; attribute dont_touch of G2443: signal is true;
	signal G2444: std_logic; attribute dont_touch of G2444: signal is true;
	signal G2447: std_logic; attribute dont_touch of G2447: signal is true;
	signal G2448: std_logic; attribute dont_touch of G2448: signal is true;
	signal G2451: std_logic; attribute dont_touch of G2451: signal is true;
	signal G2454: std_logic; attribute dont_touch of G2454: signal is true;
	signal G2455: std_logic; attribute dont_touch of G2455: signal is true;
	signal G2456: std_logic; attribute dont_touch of G2456: signal is true;
	signal G2457: std_logic; attribute dont_touch of G2457: signal is true;
	signal G2458: std_logic; attribute dont_touch of G2458: signal is true;
	signal G2459: std_logic; attribute dont_touch of G2459: signal is true;
	signal G2462: std_logic; attribute dont_touch of G2462: signal is true;
	signal G2463: std_logic; attribute dont_touch of G2463: signal is true;
	signal G2466: std_logic; attribute dont_touch of G2466: signal is true;
	signal G2469: std_logic; attribute dont_touch of G2469: signal is true;
	signal G2470: std_logic; attribute dont_touch of G2470: signal is true;
	signal G2471: std_logic; attribute dont_touch of G2471: signal is true;
	signal G2472: std_logic; attribute dont_touch of G2472: signal is true;
	signal G2473: std_logic; attribute dont_touch of G2473: signal is true;
	signal G2476: std_logic; attribute dont_touch of G2476: signal is true;
	signal G2477: std_logic; attribute dont_touch of G2477: signal is true;
	signal G2478: std_logic; attribute dont_touch of G2478: signal is true;
	signal G2479: std_logic; attribute dont_touch of G2479: signal is true;
	signal G2480: std_logic; attribute dont_touch of G2480: signal is true;
	signal G2483: std_logic; attribute dont_touch of G2483: signal is true;
	signal G2486: std_logic; attribute dont_touch of G2486: signal is true;
	signal G2489: std_logic; attribute dont_touch of G2489: signal is true;
	signal G2492: std_logic; attribute dont_touch of G2492: signal is true;
	signal G2495: std_logic; attribute dont_touch of G2495: signal is true;
	signal G2498: std_logic; attribute dont_touch of G2498: signal is true;
	signal G2501: std_logic; attribute dont_touch of G2501: signal is true;
	signal G2502: std_logic; attribute dont_touch of G2502: signal is true;
	signal G2503: std_logic; attribute dont_touch of G2503: signal is true;
	signal G2504: std_logic; attribute dont_touch of G2504: signal is true;
	signal G2507: std_logic; attribute dont_touch of G2507: signal is true;
	signal G2510: std_logic; attribute dont_touch of G2510: signal is true;
	signal G2513: std_logic; attribute dont_touch of G2513: signal is true;
	signal G2516: std_logic; attribute dont_touch of G2516: signal is true;
	signal G2519: std_logic; attribute dont_touch of G2519: signal is true;
	signal G2522: std_logic; attribute dont_touch of G2522: signal is true;
	signal G2523: std_logic; attribute dont_touch of G2523: signal is true;
	signal G2524: std_logic; attribute dont_touch of G2524: signal is true;
	signal G2525: std_logic; attribute dont_touch of G2525: signal is true;
	signal G2526: std_logic; attribute dont_touch of G2526: signal is true;
	signal G2527: std_logic; attribute dont_touch of G2527: signal is true;
	signal G2528: std_logic; attribute dont_touch of G2528: signal is true;
	signal G2529: std_logic; attribute dont_touch of G2529: signal is true;
	signal G2530: std_logic; attribute dont_touch of G2530: signal is true;
	signal G2533: std_logic; attribute dont_touch of G2533: signal is true;
	signal G2536: std_logic; attribute dont_touch of G2536: signal is true;
	signal G2539: std_logic; attribute dont_touch of G2539: signal is true;
	signal G2540: std_logic; attribute dont_touch of G2540: signal is true;
	signal G2543: std_logic; attribute dont_touch of G2543: signal is true;
	signal G2546: std_logic; attribute dont_touch of G2546: signal is true;
	signal G2549: std_logic; attribute dont_touch of G2549: signal is true;
	signal G2552: std_logic; attribute dont_touch of G2552: signal is true;
	signal G2553: std_logic; attribute dont_touch of G2553: signal is true;
	signal G2554: std_logic; attribute dont_touch of G2554: signal is true;
	signal G2555: std_logic; attribute dont_touch of G2555: signal is true;
	signal G2556: std_logic; attribute dont_touch of G2556: signal is true;
	signal G2559: std_logic; attribute dont_touch of G2559: signal is true;
	signal G2560: std_logic; attribute dont_touch of G2560: signal is true;
	signal G2561: std_logic; attribute dont_touch of G2561: signal is true;
	signal G2562: std_logic; attribute dont_touch of G2562: signal is true;
	signal G2563: std_logic; attribute dont_touch of G2563: signal is true;
	signal G2564: std_logic; attribute dont_touch of G2564: signal is true;
	signal G2565: std_logic; attribute dont_touch of G2565: signal is true;
	signal G2568: std_logic; attribute dont_touch of G2568: signal is true;
	signal G2571: std_logic; attribute dont_touch of G2571: signal is true;
	signal G2574: std_logic; attribute dont_touch of G2574: signal is true;
	signal G2580: std_logic; attribute dont_touch of G2580: signal is true;
	signal G2581: std_logic; attribute dont_touch of G2581: signal is true;
	signal G2582: std_logic; attribute dont_touch of G2582: signal is true;
	signal G2583: std_logic; attribute dont_touch of G2583: signal is true;
	signal G2584: std_logic; attribute dont_touch of G2584: signal is true;
	signal G2587: std_logic; attribute dont_touch of G2587: signal is true;
	signal G2588: std_logic; attribute dont_touch of G2588: signal is true;
	signal G2589: std_logic; attribute dont_touch of G2589: signal is true;
	signal G2590: std_logic; attribute dont_touch of G2590: signal is true;
	signal G2591: std_logic; attribute dont_touch of G2591: signal is true;
	signal G2592: std_logic; attribute dont_touch of G2592: signal is true;
	signal G2593: std_logic; attribute dont_touch of G2593: signal is true;
	signal G2594: std_logic; attribute dont_touch of G2594: signal is true;
	signal G2597: std_logic; attribute dont_touch of G2597: signal is true;
	signal G2598: std_logic; attribute dont_touch of G2598: signal is true;
	signal G2599: std_logic; attribute dont_touch of G2599: signal is true;
	signal G2602: std_logic; attribute dont_touch of G2602: signal is true;
	signal G2603: std_logic; attribute dont_touch of G2603: signal is true;
	signal G2604: std_logic; attribute dont_touch of G2604: signal is true;
	signal G2605: std_logic; attribute dont_touch of G2605: signal is true;
	signal G2606: std_logic; attribute dont_touch of G2606: signal is true;
	signal G2607: std_logic; attribute dont_touch of G2607: signal is true;
	signal G2608: std_logic; attribute dont_touch of G2608: signal is true;
	signal G2609: std_logic; attribute dont_touch of G2609: signal is true;
	signal G2610: std_logic; attribute dont_touch of G2610: signal is true;
	signal G2611: std_logic; attribute dont_touch of G2611: signal is true;
	signal G2612: std_logic; attribute dont_touch of G2612: signal is true;
	signal G2615: std_logic; attribute dont_touch of G2615: signal is true;
	signal G2616: std_logic; attribute dont_touch of G2616: signal is true;
	signal G2617: std_logic; attribute dont_touch of G2617: signal is true;
	signal G2618: std_logic; attribute dont_touch of G2618: signal is true;
	signal G2619: std_logic; attribute dont_touch of G2619: signal is true;
	signal G2622: std_logic; attribute dont_touch of G2622: signal is true;
	signal G2623: std_logic; attribute dont_touch of G2623: signal is true;
	signal G2624: std_logic; attribute dont_touch of G2624: signal is true;
	signal G2625: std_logic; attribute dont_touch of G2625: signal is true;
	signal G2628: std_logic; attribute dont_touch of G2628: signal is true;
	signal G2631: std_logic; attribute dont_touch of G2631: signal is true;
	signal G2632: std_logic; attribute dont_touch of G2632: signal is true;
	signal G2633: std_logic; attribute dont_touch of G2633: signal is true;
	signal G2636: std_logic; attribute dont_touch of G2636: signal is true;
	signal G2638: std_logic; attribute dont_touch of G2638: signal is true;
	signal G2639: std_logic; attribute dont_touch of G2639: signal is true;
	signal G2640: std_logic; attribute dont_touch of G2640: signal is true;
	signal G2641: std_logic; attribute dont_touch of G2641: signal is true;
	signal G2642: std_logic; attribute dont_touch of G2642: signal is true;
	signal G2643: std_logic; attribute dont_touch of G2643: signal is true;
	signal G2644: std_logic; attribute dont_touch of G2644: signal is true;
	signal G2645: std_logic; attribute dont_touch of G2645: signal is true;
	signal G2646: std_logic; attribute dont_touch of G2646: signal is true;
	signal G2647: std_logic; attribute dont_touch of G2647: signal is true;
	signal G2648: std_logic; attribute dont_touch of G2648: signal is true;
	signal G2649: std_logic; attribute dont_touch of G2649: signal is true;
	signal G2650: std_logic; attribute dont_touch of G2650: signal is true;
	signal G2651: std_logic; attribute dont_touch of G2651: signal is true;
	signal G2652: std_logic; attribute dont_touch of G2652: signal is true;
	signal G2653: std_logic; attribute dont_touch of G2653: signal is true;
	signal G2654: std_logic; attribute dont_touch of G2654: signal is true;
	signal G2655: std_logic; attribute dont_touch of G2655: signal is true;
	signal G2656: std_logic; attribute dont_touch of G2656: signal is true;
	signal G2657: std_logic; attribute dont_touch of G2657: signal is true;
	signal G2658: std_logic; attribute dont_touch of G2658: signal is true;
	signal G2659: std_logic; attribute dont_touch of G2659: signal is true;
	signal G2660: std_logic; attribute dont_touch of G2660: signal is true;
	signal G2661: std_logic; attribute dont_touch of G2661: signal is true;
	signal G2664: std_logic; attribute dont_touch of G2664: signal is true;
	signal G2667: std_logic; attribute dont_touch of G2667: signal is true;
	signal G2670: std_logic; attribute dont_touch of G2670: signal is true;
	signal G2673: std_logic; attribute dont_touch of G2673: signal is true;
	signal G2676: std_logic; attribute dont_touch of G2676: signal is true;
	signal G2679: std_logic; attribute dont_touch of G2679: signal is true;
	signal G2682: std_logic; attribute dont_touch of G2682: signal is true;
	signal G2685: std_logic; attribute dont_touch of G2685: signal is true;
	signal G2688: std_logic; attribute dont_touch of G2688: signal is true;
	signal G2691: std_logic; attribute dont_touch of G2691: signal is true;
	signal G2694: std_logic; attribute dont_touch of G2694: signal is true;
	signal G2697: std_logic; attribute dont_touch of G2697: signal is true;
	signal G2700: std_logic; attribute dont_touch of G2700: signal is true;
	signal G2703: std_logic; attribute dont_touch of G2703: signal is true;
	signal G2704: std_logic; attribute dont_touch of G2704: signal is true;
	signal G2707: std_logic; attribute dont_touch of G2707: signal is true;
	signal G2714: std_logic; attribute dont_touch of G2714: signal is true;
	signal G2720: std_logic; attribute dont_touch of G2720: signal is true;
	signal G2727: std_logic; attribute dont_touch of G2727: signal is true;
	signal G2733: std_logic; attribute dont_touch of G2733: signal is true;
	signal G2734: std_logic; attribute dont_touch of G2734: signal is true;
	signal G2740: std_logic; attribute dont_touch of G2740: signal is true;
	signal G2746: std_logic; attribute dont_touch of G2746: signal is true;
	signal G2753: std_logic; attribute dont_touch of G2753: signal is true;
	signal G2760: std_logic; attribute dont_touch of G2760: signal is true;
	signal G2766: std_logic; attribute dont_touch of G2766: signal is true;
	signal G2772: std_logic; attribute dont_touch of G2772: signal is true;
	signal G2773: std_logic; attribute dont_touch of G2773: signal is true;
	signal G2774: std_logic; attribute dont_touch of G2774: signal is true;
	signal G2775: std_logic; attribute dont_touch of G2775: signal is true;
	signal G2776: std_logic; attribute dont_touch of G2776: signal is true;
	signal G2777: std_logic; attribute dont_touch of G2777: signal is true;
	signal G2778: std_logic; attribute dont_touch of G2778: signal is true;
	signal G2779: std_logic; attribute dont_touch of G2779: signal is true;
	signal G2780: std_logic; attribute dont_touch of G2780: signal is true;
	signal G2781: std_logic; attribute dont_touch of G2781: signal is true;
	signal G2782: std_logic; attribute dont_touch of G2782: signal is true;
	signal G2783: std_logic; attribute dont_touch of G2783: signal is true;
	signal G2784: std_logic; attribute dont_touch of G2784: signal is true;
	signal G2785: std_logic; attribute dont_touch of G2785: signal is true;
	signal G2786: std_logic; attribute dont_touch of G2786: signal is true;
	signal G2787: std_logic; attribute dont_touch of G2787: signal is true;
	signal G2788: std_logic; attribute dont_touch of G2788: signal is true;
	signal G2789: std_logic; attribute dont_touch of G2789: signal is true;
	signal G2790: std_logic; attribute dont_touch of G2790: signal is true;
	signal G2791: std_logic; attribute dont_touch of G2791: signal is true;
	signal G2792: std_logic; attribute dont_touch of G2792: signal is true;
	signal G2793: std_logic; attribute dont_touch of G2793: signal is true;
	signal G2794: std_logic; attribute dont_touch of G2794: signal is true;
	signal G2795: std_logic; attribute dont_touch of G2795: signal is true;
	signal G2796: std_logic; attribute dont_touch of G2796: signal is true;
	signal G2797: std_logic; attribute dont_touch of G2797: signal is true;
	signal G2798: std_logic; attribute dont_touch of G2798: signal is true;
	signal G2799: std_logic; attribute dont_touch of G2799: signal is true;
	signal G2800: std_logic; attribute dont_touch of G2800: signal is true;
	signal G2801: std_logic; attribute dont_touch of G2801: signal is true;
	signal G2802: std_logic; attribute dont_touch of G2802: signal is true;
	signal G2803: std_logic; attribute dont_touch of G2803: signal is true;
	signal G2804: std_logic; attribute dont_touch of G2804: signal is true;
	signal G2805: std_logic; attribute dont_touch of G2805: signal is true;
	signal G2806: std_logic; attribute dont_touch of G2806: signal is true;
	signal G2807: std_logic; attribute dont_touch of G2807: signal is true;
	signal G2808: std_logic; attribute dont_touch of G2808: signal is true;
	signal G2809: std_logic; attribute dont_touch of G2809: signal is true;
	signal G2810: std_logic; attribute dont_touch of G2810: signal is true;
	signal G2811: std_logic; attribute dont_touch of G2811: signal is true;
	signal G2812: std_logic; attribute dont_touch of G2812: signal is true;
	signal G2813: std_logic; attribute dont_touch of G2813: signal is true;
	signal G2814: std_logic; attribute dont_touch of G2814: signal is true;
	signal G2817: std_logic; attribute dont_touch of G2817: signal is true;
	signal G2818: std_logic; attribute dont_touch of G2818: signal is true;
	signal G2821: std_logic; attribute dont_touch of G2821: signal is true;
	signal G2824: std_logic; attribute dont_touch of G2824: signal is true;
	signal G2827: std_logic; attribute dont_touch of G2827: signal is true;
	signal G2830: std_logic; attribute dont_touch of G2830: signal is true;
	signal G2833: std_logic; attribute dont_touch of G2833: signal is true;
	signal G2836: std_logic; attribute dont_touch of G2836: signal is true;
	signal G2839: std_logic; attribute dont_touch of G2839: signal is true;
	signal G2842: std_logic; attribute dont_touch of G2842: signal is true;
	signal G2845: std_logic; attribute dont_touch of G2845: signal is true;
	signal G2848: std_logic; attribute dont_touch of G2848: signal is true;
	signal G2851: std_logic; attribute dont_touch of G2851: signal is true;
	signal G2854: std_logic; attribute dont_touch of G2854: signal is true;
	signal G2857: std_logic; attribute dont_touch of G2857: signal is true;
	signal G2858: std_logic; attribute dont_touch of G2858: signal is true;
	signal G2861: std_logic; attribute dont_touch of G2861: signal is true;
	signal G2864: std_logic; attribute dont_touch of G2864: signal is true;
	signal G2867: std_logic; attribute dont_touch of G2867: signal is true;
	signal G2870: std_logic; attribute dont_touch of G2870: signal is true;
	signal G2873: std_logic; attribute dont_touch of G2873: signal is true;
	signal G2874: std_logic; attribute dont_touch of G2874: signal is true;
	signal G2877: std_logic; attribute dont_touch of G2877: signal is true;
	signal G2878: std_logic; attribute dont_touch of G2878: signal is true;
	signal G2879: std_logic; attribute dont_touch of G2879: signal is true;
	signal G2883: std_logic; attribute dont_touch of G2883: signal is true;
	signal G2888: std_logic; attribute dont_touch of G2888: signal is true;
	signal G2892: std_logic; attribute dont_touch of G2892: signal is true;
	signal G2896: std_logic; attribute dont_touch of G2896: signal is true;
	signal G2900: std_logic; attribute dont_touch of G2900: signal is true;
	signal G2903: std_logic; attribute dont_touch of G2903: signal is true;
	signal G2908: std_logic; attribute dont_touch of G2908: signal is true;
	signal G2912: std_logic; attribute dont_touch of G2912: signal is true;
	signal G2917: std_logic; attribute dont_touch of G2917: signal is true;
	signal G2920: std_logic; attribute dont_touch of G2920: signal is true;
	signal G2924: std_logic; attribute dont_touch of G2924: signal is true;
	signal G2929: std_logic; attribute dont_touch of G2929: signal is true;
	signal G2930: std_logic; attribute dont_touch of G2930: signal is true;
	signal G2933: std_logic; attribute dont_touch of G2933: signal is true;
	signal G2934: std_logic; attribute dont_touch of G2934: signal is true;
	signal G2935: std_logic; attribute dont_touch of G2935: signal is true;
	signal G2938: std_logic; attribute dont_touch of G2938: signal is true;
	signal G2941: std_logic; attribute dont_touch of G2941: signal is true;
	signal G2944: std_logic; attribute dont_touch of G2944: signal is true;
	signal G2947: std_logic; attribute dont_touch of G2947: signal is true;
	signal G2950: std_logic; attribute dont_touch of G2950: signal is true;
	signal G2953: std_logic; attribute dont_touch of G2953: signal is true;
	signal G2956: std_logic; attribute dont_touch of G2956: signal is true;
	signal G2959: std_logic; attribute dont_touch of G2959: signal is true;
	signal G2962: std_logic; attribute dont_touch of G2962: signal is true;
	signal G2963: std_logic; attribute dont_touch of G2963: signal is true;
	signal G2966: std_logic; attribute dont_touch of G2966: signal is true;
	signal G2969: std_logic; attribute dont_touch of G2969: signal is true;
	signal G2972: std_logic; attribute dont_touch of G2972: signal is true;
	signal G2975: std_logic; attribute dont_touch of G2975: signal is true;
	signal G2978: std_logic; attribute dont_touch of G2978: signal is true;
	signal G2981: std_logic; attribute dont_touch of G2981: signal is true;
	signal G2984: std_logic; attribute dont_touch of G2984: signal is true;
	signal G2985: std_logic; attribute dont_touch of G2985: signal is true;
	signal G2986: std_logic; attribute dont_touch of G2986: signal is true;
	signal G2987: std_logic; attribute dont_touch of G2987: signal is true;
	signal G2990: std_logic; attribute dont_touch of G2990: signal is true;
	signal G2991: std_logic; attribute dont_touch of G2991: signal is true;
	signal G2992: std_logic; attribute dont_touch of G2992: signal is true;
	signal G2993: std_logic; attribute dont_touch of G2993: signal is true;
	signal G2997: std_logic; attribute dont_touch of G2997: signal is true;
	signal G2998: std_logic; attribute dont_touch of G2998: signal is true;
	signal G3002: std_logic; attribute dont_touch of G3002: signal is true;
	signal G3006: std_logic; attribute dont_touch of G3006: signal is true;
	signal G3010: std_logic; attribute dont_touch of G3010: signal is true;
	signal G3013: std_logic; attribute dont_touch of G3013: signal is true;
	signal G3018: std_logic; attribute dont_touch of G3018: signal is true;
	signal G3024: std_logic; attribute dont_touch of G3024: signal is true;
	signal G3028: std_logic; attribute dont_touch of G3028: signal is true;
	signal G3032: std_logic; attribute dont_touch of G3032: signal is true;
	signal G3036: std_logic; attribute dont_touch of G3036: signal is true;
	signal G3040: std_logic; attribute dont_touch of G3040: signal is true;
	signal G3043: std_logic; attribute dont_touch of G3043: signal is true;
	signal G3044: std_logic; attribute dont_touch of G3044: signal is true;
	signal G3045: std_logic; attribute dont_touch of G3045: signal is true;
	signal G3046: std_logic; attribute dont_touch of G3046: signal is true;
	signal G3047: std_logic; attribute dont_touch of G3047: signal is true;
	signal G3048: std_logic; attribute dont_touch of G3048: signal is true;
	signal G3049: std_logic; attribute dont_touch of G3049: signal is true;
	signal G3050: std_logic; attribute dont_touch of G3050: signal is true;
	signal G3051: std_logic; attribute dont_touch of G3051: signal is true;
	signal G3052: std_logic; attribute dont_touch of G3052: signal is true;
	signal G3053: std_logic; attribute dont_touch of G3053: signal is true;
	signal G3054: std_logic; attribute dont_touch of G3054: signal is true;
	signal G3055: std_logic; attribute dont_touch of G3055: signal is true;
	signal G3056: std_logic; attribute dont_touch of G3056: signal is true;
	signal G3057: std_logic; attribute dont_touch of G3057: signal is true;
	signal G3058: std_logic; attribute dont_touch of G3058: signal is true;
	signal G3059: std_logic; attribute dont_touch of G3059: signal is true;
	signal G3060: std_logic; attribute dont_touch of G3060: signal is true;
	signal G3061: std_logic; attribute dont_touch of G3061: signal is true;
	signal G3062: std_logic; attribute dont_touch of G3062: signal is true;
	signal G3063: std_logic; attribute dont_touch of G3063: signal is true;
	signal G3064: std_logic; attribute dont_touch of G3064: signal is true;
	signal G3065: std_logic; attribute dont_touch of G3065: signal is true;
	signal G3066: std_logic; attribute dont_touch of G3066: signal is true;
	signal G3067: std_logic; attribute dont_touch of G3067: signal is true;
	signal G3068: std_logic; attribute dont_touch of G3068: signal is true;
	signal G3069: std_logic; attribute dont_touch of G3069: signal is true;
	signal G3070: std_logic; attribute dont_touch of G3070: signal is true;
	signal G3071: std_logic; attribute dont_touch of G3071: signal is true;
	signal G3072: std_logic; attribute dont_touch of G3072: signal is true;
	signal G3073: std_logic; attribute dont_touch of G3073: signal is true;
	signal G3074: std_logic; attribute dont_touch of G3074: signal is true;
	signal G3075: std_logic; attribute dont_touch of G3075: signal is true;
	signal G3076: std_logic; attribute dont_touch of G3076: signal is true;
	signal G3077: std_logic; attribute dont_touch of G3077: signal is true;
	signal G3078: std_logic; attribute dont_touch of G3078: signal is true;
	signal G3079: std_logic; attribute dont_touch of G3079: signal is true;
	signal G3080: std_logic; attribute dont_touch of G3080: signal is true;
	signal G3083: std_logic; attribute dont_touch of G3083: signal is true;
	signal G3084: std_logic; attribute dont_touch of G3084: signal is true;
	signal G3085: std_logic; attribute dont_touch of G3085: signal is true;
	signal G3086: std_logic; attribute dont_touch of G3086: signal is true;
	signal G3087: std_logic; attribute dont_touch of G3087: signal is true;
	signal G3088: std_logic; attribute dont_touch of G3088: signal is true;
	signal G3091: std_logic; attribute dont_touch of G3091: signal is true;
	signal G3092: std_logic; attribute dont_touch of G3092: signal is true;
	signal G3093: std_logic; attribute dont_touch of G3093: signal is true;
	signal G3094: std_logic; attribute dont_touch of G3094: signal is true;
	signal G3095: std_logic; attribute dont_touch of G3095: signal is true;
	signal G3096: std_logic; attribute dont_touch of G3096: signal is true;
	signal G3097: std_logic; attribute dont_touch of G3097: signal is true;
	signal G3098: std_logic; attribute dont_touch of G3098: signal is true;
	signal G3099: std_logic; attribute dont_touch of G3099: signal is true;
	signal G3100: std_logic; attribute dont_touch of G3100: signal is true;
	signal G3101: std_logic; attribute dont_touch of G3101: signal is true;
	signal G3102: std_logic; attribute dont_touch of G3102: signal is true;
	signal G3103: std_logic; attribute dont_touch of G3103: signal is true;
	signal G3104: std_logic; attribute dont_touch of G3104: signal is true;
	signal G3105: std_logic; attribute dont_touch of G3105: signal is true;
	signal G3106: std_logic; attribute dont_touch of G3106: signal is true;
	signal G3107: std_logic; attribute dont_touch of G3107: signal is true;
	signal G3108: std_logic; attribute dont_touch of G3108: signal is true;
	signal G3109: std_logic; attribute dont_touch of G3109: signal is true;
	signal G3110: std_logic; attribute dont_touch of G3110: signal is true;
	signal G3111: std_logic; attribute dont_touch of G3111: signal is true;
	signal G3112: std_logic; attribute dont_touch of G3112: signal is true;
	signal G3113: std_logic; attribute dont_touch of G3113: signal is true;
	signal G3114: std_logic; attribute dont_touch of G3114: signal is true;
	signal G3117: std_logic; attribute dont_touch of G3117: signal is true;
	signal G3120: std_logic; attribute dont_touch of G3120: signal is true;
	signal G3123: std_logic; attribute dont_touch of G3123: signal is true;
	signal G3124: std_logic; attribute dont_touch of G3124: signal is true;
	signal G3125: std_logic; attribute dont_touch of G3125: signal is true;
	signal G3126: std_logic; attribute dont_touch of G3126: signal is true;
	signal G3127: std_logic; attribute dont_touch of G3127: signal is true;
	signal G3128: std_logic; attribute dont_touch of G3128: signal is true;
	signal G3129: std_logic; attribute dont_touch of G3129: signal is true;
	signal G3132: std_logic; attribute dont_touch of G3132: signal is true;
	signal G3133: std_logic; attribute dont_touch of G3133: signal is true;
	signal G3134: std_logic; attribute dont_touch of G3134: signal is true;
	signal G3135: std_logic; attribute dont_touch of G3135: signal is true;
	signal G3136: std_logic; attribute dont_touch of G3136: signal is true;
	signal G3139: std_logic; attribute dont_touch of G3139: signal is true;
	signal G3142: std_logic; attribute dont_touch of G3142: signal is true;
	signal G3147: std_logic; attribute dont_touch of G3147: signal is true;
	signal G3151: std_logic; attribute dont_touch of G3151: signal is true;
	signal G3155: std_logic; attribute dont_touch of G3155: signal is true;
	signal G3158: std_logic; attribute dont_touch of G3158: signal is true;
	signal G3161: std_logic; attribute dont_touch of G3161: signal is true;
	signal G3164: std_logic; attribute dont_touch of G3164: signal is true;
	signal G3167: std_logic; attribute dont_touch of G3167: signal is true;
	signal G3170: std_logic; attribute dont_touch of G3170: signal is true;
	signal G3173: std_logic; attribute dont_touch of G3173: signal is true;
	signal G3176: std_logic; attribute dont_touch of G3176: signal is true;
	signal G3179: std_logic; attribute dont_touch of G3179: signal is true;
	signal G3182: std_logic; attribute dont_touch of G3182: signal is true;
	signal G3185: std_logic; attribute dont_touch of G3185: signal is true;
	signal G3188: std_logic; attribute dont_touch of G3188: signal is true;
	signal G3191: std_logic; attribute dont_touch of G3191: signal is true;
	signal G3194: std_logic; attribute dont_touch of G3194: signal is true;
	signal G3197: std_logic; attribute dont_touch of G3197: signal is true;
	signal G3198: std_logic; attribute dont_touch of G3198: signal is true;
	signal G3201: std_logic; attribute dont_touch of G3201: signal is true;
	signal G3204: std_logic; attribute dont_touch of G3204: signal is true;
	signal G3207: std_logic; attribute dont_touch of G3207: signal is true;
	signal G3210: std_logic; attribute dont_touch of G3210: signal is true;
	signal G3211: std_logic; attribute dont_touch of G3211: signal is true;
	signal G3235: std_logic; attribute dont_touch of G3235: signal is true;
	signal G3236: std_logic; attribute dont_touch of G3236: signal is true;
	signal G3237: std_logic; attribute dont_touch of G3237: signal is true;
	signal G3238: std_logic; attribute dont_touch of G3238: signal is true;
	signal G3239: std_logic; attribute dont_touch of G3239: signal is true;
	signal G3240: std_logic; attribute dont_touch of G3240: signal is true;
	signal G3241: std_logic; attribute dont_touch of G3241: signal is true;
	signal G3242: std_logic; attribute dont_touch of G3242: signal is true;
	signal G3243: std_logic; attribute dont_touch of G3243: signal is true;
	signal G3244: std_logic; attribute dont_touch of G3244: signal is true;
	signal G3245: std_logic; attribute dont_touch of G3245: signal is true;
	signal G3246: std_logic; attribute dont_touch of G3246: signal is true;
	signal G3247: std_logic; attribute dont_touch of G3247: signal is true;
	signal G3248: std_logic; attribute dont_touch of G3248: signal is true;
	signal G3249: std_logic; attribute dont_touch of G3249: signal is true;
	signal G3250: std_logic; attribute dont_touch of G3250: signal is true;
	signal G3251: std_logic; attribute dont_touch of G3251: signal is true;
	signal G3252: std_logic; attribute dont_touch of G3252: signal is true;
	signal G3253: std_logic; attribute dont_touch of G3253: signal is true;
	signal G3254: std_logic; attribute dont_touch of G3254: signal is true;
	signal G3304: std_logic; attribute dont_touch of G3304: signal is true;
	signal G3305: std_logic; attribute dont_touch of G3305: signal is true;
	signal G3306: std_logic; attribute dont_touch of G3306: signal is true;
	signal G3337: std_logic; attribute dont_touch of G3337: signal is true;
	signal G3338: std_logic; attribute dont_touch of G3338: signal is true;
	signal G3365: std_logic; attribute dont_touch of G3365: signal is true;
	signal G3366: std_logic; attribute dont_touch of G3366: signal is true;
	signal G3398: std_logic; attribute dont_touch of G3398: signal is true;
	signal G3410: std_logic; attribute dont_touch of G3410: signal is true;
	signal G3460: std_logic; attribute dont_touch of G3460: signal is true;
	signal G3461: std_logic; attribute dont_touch of G3461: signal is true;
	signal G3462: std_logic; attribute dont_touch of G3462: signal is true;
	signal G3493: std_logic; attribute dont_touch of G3493: signal is true;
	signal G3494: std_logic; attribute dont_touch of G3494: signal is true;
	signal G3521: std_logic; attribute dont_touch of G3521: signal is true;
	signal G3522: std_logic; attribute dont_touch of G3522: signal is true;
	signal G3554: std_logic; attribute dont_touch of G3554: signal is true;
	signal G3566: std_logic; attribute dont_touch of G3566: signal is true;
	signal G3616: std_logic; attribute dont_touch of G3616: signal is true;
	signal G3617: std_logic; attribute dont_touch of G3617: signal is true;
	signal G3618: std_logic; attribute dont_touch of G3618: signal is true;
	signal G3649: std_logic; attribute dont_touch of G3649: signal is true;
	signal G3650: std_logic; attribute dont_touch of G3650: signal is true;
	signal G3677: std_logic; attribute dont_touch of G3677: signal is true;
	signal G3678: std_logic; attribute dont_touch of G3678: signal is true;
	signal G3710: std_logic; attribute dont_touch of G3710: signal is true;
	signal G3722: std_logic; attribute dont_touch of G3722: signal is true;
	signal G3772: std_logic; attribute dont_touch of G3772: signal is true;
	signal G3773: std_logic; attribute dont_touch of G3773: signal is true;
	signal G3774: std_logic; attribute dont_touch of G3774: signal is true;
	signal G3805: std_logic; attribute dont_touch of G3805: signal is true;
	signal G3806: std_logic; attribute dont_touch of G3806: signal is true;
	signal G3833: std_logic; attribute dont_touch of G3833: signal is true;
	signal G3834: std_logic; attribute dont_touch of G3834: signal is true;
	signal G3866: std_logic; attribute dont_touch of G3866: signal is true;
	signal G3878: std_logic; attribute dont_touch of G3878: signal is true;
	signal G3897: std_logic; attribute dont_touch of G3897: signal is true;
	signal G3900: std_logic; attribute dont_touch of G3900: signal is true;
	signal G3919: std_logic; attribute dont_touch of G3919: signal is true;
	signal G3922: std_logic; attribute dont_touch of G3922: signal is true;
	signal G3925: std_logic; attribute dont_touch of G3925: signal is true;
	signal G3928: std_logic; attribute dont_touch of G3928: signal is true;
	signal G3931: std_logic; attribute dont_touch of G3931: signal is true;
	signal G3934: std_logic; attribute dont_touch of G3934: signal is true;
	signal G3937: std_logic; attribute dont_touch of G3937: signal is true;
	signal G3940: std_logic; attribute dont_touch of G3940: signal is true;
	signal G3941: std_logic; attribute dont_touch of G3941: signal is true;
	signal G3942: std_logic; attribute dont_touch of G3942: signal is true;
	signal G3945: std_logic; attribute dont_touch of G3945: signal is true;
	signal G3948: std_logic; attribute dont_touch of G3948: signal is true;
	signal G3951: std_logic; attribute dont_touch of G3951: signal is true;
	signal G3954: std_logic; attribute dont_touch of G3954: signal is true;
	signal G3957: std_logic; attribute dont_touch of G3957: signal is true;
	signal G3960: std_logic; attribute dont_touch of G3960: signal is true;
	signal G3963: std_logic; attribute dont_touch of G3963: signal is true;
	signal G3966: std_logic; attribute dont_touch of G3966: signal is true;
	signal G3969: std_logic; attribute dont_touch of G3969: signal is true;
	signal G3972: std_logic; attribute dont_touch of G3972: signal is true;
	signal G3975: std_logic; attribute dont_touch of G3975: signal is true;
	signal G3978: std_logic; attribute dont_touch of G3978: signal is true;
	signal G3981: std_logic; attribute dont_touch of G3981: signal is true;
	signal G3984: std_logic; attribute dont_touch of G3984: signal is true;
	signal G3987: std_logic; attribute dont_touch of G3987: signal is true;
	signal G3990: std_logic; attribute dont_touch of G3990: signal is true;
	signal G3994: std_logic; attribute dont_touch of G3994: signal is true;
	signal G3995: std_logic; attribute dont_touch of G3995: signal is true;
	signal G3996: std_logic; attribute dont_touch of G3996: signal is true;
	signal G3997: std_logic; attribute dont_touch of G3997: signal is true;
	signal G3998: std_logic; attribute dont_touch of G3998: signal is true;
	signal G3999: std_logic; attribute dont_touch of G3999: signal is true;
	signal G4000: std_logic; attribute dont_touch of G4000: signal is true;
	signal G4003: std_logic; attribute dont_touch of G4003: signal is true;
	signal G4006: std_logic; attribute dont_touch of G4006: signal is true;
	signal G4009: std_logic; attribute dont_touch of G4009: signal is true;
	signal G4012: std_logic; attribute dont_touch of G4012: signal is true;
	signal G4015: std_logic; attribute dont_touch of G4015: signal is true;
	signal G4016: std_logic; attribute dont_touch of G4016: signal is true;
	signal G4017: std_logic; attribute dont_touch of G4017: signal is true;
	signal G4020: std_logic; attribute dont_touch of G4020: signal is true;
	signal G4023: std_logic; attribute dont_touch of G4023: signal is true;
	signal G4026: std_logic; attribute dont_touch of G4026: signal is true;
	signal G4029: std_logic; attribute dont_touch of G4029: signal is true;
	signal G4032: std_logic; attribute dont_touch of G4032: signal is true;
	signal G4035: std_logic; attribute dont_touch of G4035: signal is true;
	signal G4038: std_logic; attribute dont_touch of G4038: signal is true;
	signal G4041: std_logic; attribute dont_touch of G4041: signal is true;
	signal G4044: std_logic; attribute dont_touch of G4044: signal is true;
	signal G4047: std_logic; attribute dont_touch of G4047: signal is true;
	signal G4048: std_logic; attribute dont_touch of G4048: signal is true;
	signal G4049: std_logic; attribute dont_touch of G4049: signal is true;
	signal G4052: std_logic; attribute dont_touch of G4052: signal is true;
	signal G4055: std_logic; attribute dont_touch of G4055: signal is true;
	signal G4058: std_logic; attribute dont_touch of G4058: signal is true;
	signal G4061: std_logic; attribute dont_touch of G4061: signal is true;
	signal G4064: std_logic; attribute dont_touch of G4064: signal is true;
	signal G4067: std_logic; attribute dont_touch of G4067: signal is true;
	signal G4070: std_logic; attribute dont_touch of G4070: signal is true;
	signal G4073: std_logic; attribute dont_touch of G4073: signal is true;
	signal G4076: std_logic; attribute dont_touch of G4076: signal is true;
	signal G4079: std_logic; attribute dont_touch of G4079: signal is true;
	signal G4082: std_logic; attribute dont_touch of G4082: signal is true;
	signal G4085: std_logic; attribute dont_touch of G4085: signal is true;
	signal G4089: std_logic; attribute dont_touch of G4089: signal is true;
	signal G4091: std_logic; attribute dont_touch of G4091: signal is true;
	signal G4092: std_logic; attribute dont_touch of G4092: signal is true;
	signal G4093: std_logic; attribute dont_touch of G4093: signal is true;
	signal G4094: std_logic; attribute dont_touch of G4094: signal is true;
	signal G4095: std_logic; attribute dont_touch of G4095: signal is true;
	signal G4098: std_logic; attribute dont_touch of G4098: signal is true;
	signal G4101: std_logic; attribute dont_touch of G4101: signal is true;
	signal G4104: std_logic; attribute dont_touch of G4104: signal is true;
	signal G4107: std_logic; attribute dont_touch of G4107: signal is true;
	signal G4110: std_logic; attribute dont_touch of G4110: signal is true;
	signal G4111: std_logic; attribute dont_touch of G4111: signal is true;
	signal G4112: std_logic; attribute dont_touch of G4112: signal is true;
	signal G4115: std_logic; attribute dont_touch of G4115: signal is true;
	signal G4118: std_logic; attribute dont_touch of G4118: signal is true;
	signal G4121: std_logic; attribute dont_touch of G4121: signal is true;
	signal G4124: std_logic; attribute dont_touch of G4124: signal is true;
	signal G4127: std_logic; attribute dont_touch of G4127: signal is true;
	signal G4130: std_logic; attribute dont_touch of G4130: signal is true;
	signal G4133: std_logic; attribute dont_touch of G4133: signal is true;
	signal G4136: std_logic; attribute dont_touch of G4136: signal is true;
	signal G4139: std_logic; attribute dont_touch of G4139: signal is true;
	signal G4142: std_logic; attribute dont_touch of G4142: signal is true;
	signal G4143: std_logic; attribute dont_touch of G4143: signal is true;
	signal G4144: std_logic; attribute dont_touch of G4144: signal is true;
	signal G4147: std_logic; attribute dont_touch of G4147: signal is true;
	signal G4150: std_logic; attribute dont_touch of G4150: signal is true;
	signal G4153: std_logic; attribute dont_touch of G4153: signal is true;
	signal G4156: std_logic; attribute dont_touch of G4156: signal is true;
	signal G4159: std_logic; attribute dont_touch of G4159: signal is true;
	signal G4162: std_logic; attribute dont_touch of G4162: signal is true;
	signal G4165: std_logic; attribute dont_touch of G4165: signal is true;
	signal G4168: std_logic; attribute dont_touch of G4168: signal is true;
	signal G4171: std_logic; attribute dont_touch of G4171: signal is true;
	signal G4174: std_logic; attribute dont_touch of G4174: signal is true;
	signal G4175: std_logic; attribute dont_touch of G4175: signal is true;
	signal G4176: std_logic; attribute dont_touch of G4176: signal is true;
	signal G4179: std_logic; attribute dont_touch of G4179: signal is true;
	signal G4182: std_logic; attribute dont_touch of G4182: signal is true;
	signal G4185: std_logic; attribute dont_touch of G4185: signal is true;
	signal G4188: std_logic; attribute dont_touch of G4188: signal is true;
	signal G4191: std_logic; attribute dont_touch of G4191: signal is true;
	signal G4194: std_logic; attribute dont_touch of G4194: signal is true;
	signal G4197: std_logic; attribute dont_touch of G4197: signal is true;
	signal G4201: std_logic; attribute dont_touch of G4201: signal is true;
	signal G4202: std_logic; attribute dont_touch of G4202: signal is true;
	signal G4203: std_logic; attribute dont_touch of G4203: signal is true;
	signal G4204: std_logic; attribute dont_touch of G4204: signal is true;
	signal G4205: std_logic; attribute dont_touch of G4205: signal is true;
	signal G4208: std_logic; attribute dont_touch of G4208: signal is true;
	signal G4211: std_logic; attribute dont_touch of G4211: signal is true;
	signal G4214: std_logic; attribute dont_touch of G4214: signal is true;
	signal G4217: std_logic; attribute dont_touch of G4217: signal is true;
	signal G4220: std_logic; attribute dont_touch of G4220: signal is true;
	signal G4221: std_logic; attribute dont_touch of G4221: signal is true;
	signal G4224: std_logic; attribute dont_touch of G4224: signal is true;
	signal G4225: std_logic; attribute dont_touch of G4225: signal is true;
	signal G4228: std_logic; attribute dont_touch of G4228: signal is true;
	signal G4231: std_logic; attribute dont_touch of G4231: signal is true;
	signal G4234: std_logic; attribute dont_touch of G4234: signal is true;
	signal G4237: std_logic; attribute dont_touch of G4237: signal is true;
	signal G4240: std_logic; attribute dont_touch of G4240: signal is true;
	signal G4243: std_logic; attribute dont_touch of G4243: signal is true;
	signal G4246: std_logic; attribute dont_touch of G4246: signal is true;
	signal G4249: std_logic; attribute dont_touch of G4249: signal is true;
	signal G4250: std_logic; attribute dont_touch of G4250: signal is true;
	signal G4251: std_logic; attribute dont_touch of G4251: signal is true;
	signal G4254: std_logic; attribute dont_touch of G4254: signal is true;
	signal G4257: std_logic; attribute dont_touch of G4257: signal is true;
	signal G4260: std_logic; attribute dont_touch of G4260: signal is true;
	signal G4263: std_logic; attribute dont_touch of G4263: signal is true;
	signal G4266: std_logic; attribute dont_touch of G4266: signal is true;
	signal G4269: std_logic; attribute dont_touch of G4269: signal is true;
	signal G4272: std_logic; attribute dont_touch of G4272: signal is true;
	signal G4275: std_logic; attribute dont_touch of G4275: signal is true;
	signal G4278: std_logic; attribute dont_touch of G4278: signal is true;
	signal G4281: std_logic; attribute dont_touch of G4281: signal is true;
	signal G4282: std_logic; attribute dont_touch of G4282: signal is true;
	signal G4283: std_logic; attribute dont_touch of G4283: signal is true;
	signal G4286: std_logic; attribute dont_touch of G4286: signal is true;
	signal G4289: std_logic; attribute dont_touch of G4289: signal is true;
	signal G4292: std_logic; attribute dont_touch of G4292: signal is true;
	signal G4295: std_logic; attribute dont_touch of G4295: signal is true;
	signal G4298: std_logic; attribute dont_touch of G4298: signal is true;
	signal G4301: std_logic; attribute dont_touch of G4301: signal is true;
	signal G4304: std_logic; attribute dont_touch of G4304: signal is true;
	signal G4307: std_logic; attribute dont_touch of G4307: signal is true;
	signal G4310: std_logic; attribute dont_touch of G4310: signal is true;
	signal G4313: std_logic; attribute dont_touch of G4313: signal is true;
	signal G4314: std_logic; attribute dont_touch of G4314: signal is true;
	signal G4315: std_logic; attribute dont_touch of G4315: signal is true;
	signal G4318: std_logic; attribute dont_touch of G4318: signal is true;
	signal G4322: std_logic; attribute dont_touch of G4322: signal is true;
	signal G4324: std_logic; attribute dont_touch of G4324: signal is true;
	signal G4325: std_logic; attribute dont_touch of G4325: signal is true;
	signal G4326: std_logic; attribute dont_touch of G4326: signal is true;
	signal G4329: std_logic; attribute dont_touch of G4329: signal is true;
	signal G4332: std_logic; attribute dont_touch of G4332: signal is true;
	signal G4335: std_logic; attribute dont_touch of G4335: signal is true;
	signal G4338: std_logic; attribute dont_touch of G4338: signal is true;
	signal G4339: std_logic; attribute dont_touch of G4339: signal is true;
	signal G4340: std_logic; attribute dont_touch of G4340: signal is true;
	signal G4343: std_logic; attribute dont_touch of G4343: signal is true;
	signal G4346: std_logic; attribute dont_touch of G4346: signal is true;
	signal G4347: std_logic; attribute dont_touch of G4347: signal is true;
	signal G4348: std_logic; attribute dont_touch of G4348: signal is true;
	signal G4351: std_logic; attribute dont_touch of G4351: signal is true;
	signal G4354: std_logic; attribute dont_touch of G4354: signal is true;
	signal G4357: std_logic; attribute dont_touch of G4357: signal is true;
	signal G4360: std_logic; attribute dont_touch of G4360: signal is true;
	signal G4363: std_logic; attribute dont_touch of G4363: signal is true;
	signal G4366: std_logic; attribute dont_touch of G4366: signal is true;
	signal G4369: std_logic; attribute dont_touch of G4369: signal is true;
	signal G4372: std_logic; attribute dont_touch of G4372: signal is true;
	signal G4375: std_logic; attribute dont_touch of G4375: signal is true;
	signal G4376: std_logic; attribute dont_touch of G4376: signal is true;
	signal G4379: std_logic; attribute dont_touch of G4379: signal is true;
	signal G4380: std_logic; attribute dont_touch of G4380: signal is true;
	signal G4383: std_logic; attribute dont_touch of G4383: signal is true;
	signal G4386: std_logic; attribute dont_touch of G4386: signal is true;
	signal G4389: std_logic; attribute dont_touch of G4389: signal is true;
	signal G4392: std_logic; attribute dont_touch of G4392: signal is true;
	signal G4395: std_logic; attribute dont_touch of G4395: signal is true;
	signal G4398: std_logic; attribute dont_touch of G4398: signal is true;
	signal G4401: std_logic; attribute dont_touch of G4401: signal is true;
	signal G4404: std_logic; attribute dont_touch of G4404: signal is true;
	signal G4405: std_logic; attribute dont_touch of G4405: signal is true;
	signal G4406: std_logic; attribute dont_touch of G4406: signal is true;
	signal G4409: std_logic; attribute dont_touch of G4409: signal is true;
	signal G4412: std_logic; attribute dont_touch of G4412: signal is true;
	signal G4415: std_logic; attribute dont_touch of G4415: signal is true;
	signal G4418: std_logic; attribute dont_touch of G4418: signal is true;
	signal G4421: std_logic; attribute dont_touch of G4421: signal is true;
	signal G4424: std_logic; attribute dont_touch of G4424: signal is true;
	signal G4427: std_logic; attribute dont_touch of G4427: signal is true;
	signal G4430: std_logic; attribute dont_touch of G4430: signal is true;
	signal G4433: std_logic; attribute dont_touch of G4433: signal is true;
	signal G4436: std_logic; attribute dont_touch of G4436: signal is true;
	signal G4437: std_logic; attribute dont_touch of G4437: signal is true;
	signal G4438: std_logic; attribute dont_touch of G4438: signal is true;
	signal G4441: std_logic; attribute dont_touch of G4441: signal is true;
	signal G4444: std_logic; attribute dont_touch of G4444: signal is true;
	signal G4447: std_logic; attribute dont_touch of G4447: signal is true;
	signal G4451: std_logic; attribute dont_touch of G4451: signal is true;
	signal G4452: std_logic; attribute dont_touch of G4452: signal is true;
	signal G4453: std_logic; attribute dont_touch of G4453: signal is true;
	signal G4456: std_logic; attribute dont_touch of G4456: signal is true;
	signal G4465: std_logic; attribute dont_touch of G4465: signal is true;
	signal G4468: std_logic; attribute dont_touch of G4468: signal is true;
	signal G4471: std_logic; attribute dont_touch of G4471: signal is true;
	signal G4474: std_logic; attribute dont_touch of G4474: signal is true;
	signal G4475: std_logic; attribute dont_touch of G4475: signal is true;
	signal G4476: std_logic; attribute dont_touch of G4476: signal is true;
	signal G4479: std_logic; attribute dont_touch of G4479: signal is true;
	signal G4480: std_logic; attribute dont_touch of G4480: signal is true;
	signal G4483: std_logic; attribute dont_touch of G4483: signal is true;
	signal G4486: std_logic; attribute dont_touch of G4486: signal is true;
	signal G4489: std_logic; attribute dont_touch of G4489: signal is true;
	signal G4492: std_logic; attribute dont_touch of G4492: signal is true;
	signal G4495: std_logic; attribute dont_touch of G4495: signal is true;
	signal G4498: std_logic; attribute dont_touch of G4498: signal is true;
	signal G4501: std_logic; attribute dont_touch of G4501: signal is true;
	signal G4504: std_logic; attribute dont_touch of G4504: signal is true;
	signal G4507: std_logic; attribute dont_touch of G4507: signal is true;
	signal G4508: std_logic; attribute dont_touch of G4508: signal is true;
	signal G4509: std_logic; attribute dont_touch of G4509: signal is true;
	signal G4512: std_logic; attribute dont_touch of G4512: signal is true;
	signal G4515: std_logic; attribute dont_touch of G4515: signal is true;
	signal G4516: std_logic; attribute dont_touch of G4516: signal is true;
	signal G4517: std_logic; attribute dont_touch of G4517: signal is true;
	signal G4520: std_logic; attribute dont_touch of G4520: signal is true;
	signal G4523: std_logic; attribute dont_touch of G4523: signal is true;
	signal G4526: std_logic; attribute dont_touch of G4526: signal is true;
	signal G4529: std_logic; attribute dont_touch of G4529: signal is true;
	signal G4532: std_logic; attribute dont_touch of G4532: signal is true;
	signal G4535: std_logic; attribute dont_touch of G4535: signal is true;
	signal G4538: std_logic; attribute dont_touch of G4538: signal is true;
	signal G4541: std_logic; attribute dont_touch of G4541: signal is true;
	signal G4544: std_logic; attribute dont_touch of G4544: signal is true;
	signal G4545: std_logic; attribute dont_touch of G4545: signal is true;
	signal G4548: std_logic; attribute dont_touch of G4548: signal is true;
	signal G4549: std_logic; attribute dont_touch of G4549: signal is true;
	signal G4552: std_logic; attribute dont_touch of G4552: signal is true;
	signal G4555: std_logic; attribute dont_touch of G4555: signal is true;
	signal G4558: std_logic; attribute dont_touch of G4558: signal is true;
	signal G4561: std_logic; attribute dont_touch of G4561: signal is true;
	signal G4564: std_logic; attribute dont_touch of G4564: signal is true;
	signal G4567: std_logic; attribute dont_touch of G4567: signal is true;
	signal G4570: std_logic; attribute dont_touch of G4570: signal is true;
	signal G4573: std_logic; attribute dont_touch of G4573: signal is true;
	signal G4574: std_logic; attribute dont_touch of G4574: signal is true;
	signal G4575: std_logic; attribute dont_touch of G4575: signal is true;
	signal G4578: std_logic; attribute dont_touch of G4578: signal is true;
	signal G4581: std_logic; attribute dont_touch of G4581: signal is true;
	signal G4584: std_logic; attribute dont_touch of G4584: signal is true;
	signal G4587: std_logic; attribute dont_touch of G4587: signal is true;
	signal G4591: std_logic; attribute dont_touch of G4591: signal is true;
	signal G4592: std_logic; attribute dont_touch of G4592: signal is true;
	signal G4595: std_logic; attribute dont_touch of G4595: signal is true;
	signal G4598: std_logic; attribute dont_touch of G4598: signal is true;
	signal G4601: std_logic; attribute dont_touch of G4601: signal is true;
	signal G4602: std_logic; attribute dont_touch of G4602: signal is true;
	signal G4603: std_logic; attribute dont_touch of G4603: signal is true;
	signal G4606: std_logic; attribute dont_touch of G4606: signal is true;
	signal G4609: std_logic; attribute dont_touch of G4609: signal is true;
	signal G4610: std_logic; attribute dont_touch of G4610: signal is true;
	signal G4611: std_logic; attribute dont_touch of G4611: signal is true;
	signal G4614: std_logic; attribute dont_touch of G4614: signal is true;
	signal G4617: std_logic; attribute dont_touch of G4617: signal is true;
	signal G4620: std_logic; attribute dont_touch of G4620: signal is true;
	signal G4623: std_logic; attribute dont_touch of G4623: signal is true;
	signal G4626: std_logic; attribute dont_touch of G4626: signal is true;
	signal G4629: std_logic; attribute dont_touch of G4629: signal is true;
	signal G4632: std_logic; attribute dont_touch of G4632: signal is true;
	signal G4641: std_logic; attribute dont_touch of G4641: signal is true;
	signal G4644: std_logic; attribute dont_touch of G4644: signal is true;
	signal G4647: std_logic; attribute dont_touch of G4647: signal is true;
	signal G4650: std_logic; attribute dont_touch of G4650: signal is true;
	signal G4651: std_logic; attribute dont_touch of G4651: signal is true;
	signal G4652: std_logic; attribute dont_touch of G4652: signal is true;
	signal G4655: std_logic; attribute dont_touch of G4655: signal is true;
	signal G4656: std_logic; attribute dont_touch of G4656: signal is true;
	signal G4659: std_logic; attribute dont_touch of G4659: signal is true;
	signal G4662: std_logic; attribute dont_touch of G4662: signal is true;
	signal G4665: std_logic; attribute dont_touch of G4665: signal is true;
	signal G4668: std_logic; attribute dont_touch of G4668: signal is true;
	signal G4671: std_logic; attribute dont_touch of G4671: signal is true;
	signal G4674: std_logic; attribute dont_touch of G4674: signal is true;
	signal G4677: std_logic; attribute dont_touch of G4677: signal is true;
	signal G4680: std_logic; attribute dont_touch of G4680: signal is true;
	signal G4683: std_logic; attribute dont_touch of G4683: signal is true;
	signal G4684: std_logic; attribute dont_touch of G4684: signal is true;
	signal G4685: std_logic; attribute dont_touch of G4685: signal is true;
	signal G4688: std_logic; attribute dont_touch of G4688: signal is true;
	signal G4691: std_logic; attribute dont_touch of G4691: signal is true;
	signal G4692: std_logic; attribute dont_touch of G4692: signal is true;
	signal G4693: std_logic; attribute dont_touch of G4693: signal is true;
	signal G4696: std_logic; attribute dont_touch of G4696: signal is true;
	signal G4699: std_logic; attribute dont_touch of G4699: signal is true;
	signal G4702: std_logic; attribute dont_touch of G4702: signal is true;
	signal G4705: std_logic; attribute dont_touch of G4705: signal is true;
	signal G4708: std_logic; attribute dont_touch of G4708: signal is true;
	signal G4711: std_logic; attribute dont_touch of G4711: signal is true;
	signal G4714: std_logic; attribute dont_touch of G4714: signal is true;
	signal G4717: std_logic; attribute dont_touch of G4717: signal is true;
	signal G4720: std_logic; attribute dont_touch of G4720: signal is true;
	signal G4721: std_logic; attribute dont_touch of G4721: signal is true;
	signal G4724: std_logic; attribute dont_touch of G4724: signal is true;
	signal G4725: std_logic; attribute dont_touch of G4725: signal is true;
	signal G4728: std_logic; attribute dont_touch of G4728: signal is true;
	signal G4731: std_logic; attribute dont_touch of G4731: signal is true;
	signal G4734: std_logic; attribute dont_touch of G4734: signal is true;
	signal G4735: std_logic; attribute dont_touch of G4735: signal is true;
	signal G4736: std_logic; attribute dont_touch of G4736: signal is true;
	signal G4737: std_logic; attribute dont_touch of G4737: signal is true;
	signal G4740: std_logic; attribute dont_touch of G4740: signal is true;
	signal G4743: std_logic; attribute dont_touch of G4743: signal is true;
	signal G4746: std_logic; attribute dont_touch of G4746: signal is true;
	signal G4749: std_logic; attribute dont_touch of G4749: signal is true;
	signal G4752: std_logic; attribute dont_touch of G4752: signal is true;
	signal G4753: std_logic; attribute dont_touch of G4753: signal is true;
	signal G4754: std_logic; attribute dont_touch of G4754: signal is true;
	signal G4757: std_logic; attribute dont_touch of G4757: signal is true;
	signal G4760: std_logic; attribute dont_touch of G4760: signal is true;
	signal G4763: std_logic; attribute dont_touch of G4763: signal is true;
	signal G4766: std_logic; attribute dont_touch of G4766: signal is true;
	signal G4769: std_logic; attribute dont_touch of G4769: signal is true;
	signal G4772: std_logic; attribute dont_touch of G4772: signal is true;
	signal G4775: std_logic; attribute dont_touch of G4775: signal is true;
	signal G4778: std_logic; attribute dont_touch of G4778: signal is true;
	signal G4779: std_logic; attribute dont_touch of G4779: signal is true;
	signal G4780: std_logic; attribute dont_touch of G4780: signal is true;
	signal G4783: std_logic; attribute dont_touch of G4783: signal is true;
	signal G4786: std_logic; attribute dont_touch of G4786: signal is true;
	signal G4787: std_logic; attribute dont_touch of G4787: signal is true;
	signal G4788: std_logic; attribute dont_touch of G4788: signal is true;
	signal G4791: std_logic; attribute dont_touch of G4791: signal is true;
	signal G4794: std_logic; attribute dont_touch of G4794: signal is true;
	signal G4797: std_logic; attribute dont_touch of G4797: signal is true;
	signal G4800: std_logic; attribute dont_touch of G4800: signal is true;
	signal G4803: std_logic; attribute dont_touch of G4803: signal is true;
	signal G4806: std_logic; attribute dont_touch of G4806: signal is true;
	signal G4809: std_logic; attribute dont_touch of G4809: signal is true;
	signal G4818: std_logic; attribute dont_touch of G4818: signal is true;
	signal G4821: std_logic; attribute dont_touch of G4821: signal is true;
	signal G4824: std_logic; attribute dont_touch of G4824: signal is true;
	signal G4827: std_logic; attribute dont_touch of G4827: signal is true;
	signal G4828: std_logic; attribute dont_touch of G4828: signal is true;
	signal G4829: std_logic; attribute dont_touch of G4829: signal is true;
	signal G4832: std_logic; attribute dont_touch of G4832: signal is true;
	signal G4833: std_logic; attribute dont_touch of G4833: signal is true;
	signal G4836: std_logic; attribute dont_touch of G4836: signal is true;
	signal G4839: std_logic; attribute dont_touch of G4839: signal is true;
	signal G4842: std_logic; attribute dont_touch of G4842: signal is true;
	signal G4845: std_logic; attribute dont_touch of G4845: signal is true;
	signal G4848: std_logic; attribute dont_touch of G4848: signal is true;
	signal G4851: std_logic; attribute dont_touch of G4851: signal is true;
	signal G4854: std_logic; attribute dont_touch of G4854: signal is true;
	signal G4857: std_logic; attribute dont_touch of G4857: signal is true;
	signal G4860: std_logic; attribute dont_touch of G4860: signal is true;
	signal G4861: std_logic; attribute dont_touch of G4861: signal is true;
	signal G4862: std_logic; attribute dont_touch of G4862: signal is true;
	signal G4865: std_logic; attribute dont_touch of G4865: signal is true;
	signal G4868: std_logic; attribute dont_touch of G4868: signal is true;
	signal G4869: std_logic; attribute dont_touch of G4869: signal is true;
	signal G4870: std_logic; attribute dont_touch of G4870: signal is true;
	signal G4873: std_logic; attribute dont_touch of G4873: signal is true;
	signal G4876: std_logic; attribute dont_touch of G4876: signal is true;
	signal G4879: std_logic; attribute dont_touch of G4879: signal is true;
	signal G4882: std_logic; attribute dont_touch of G4882: signal is true;
	signal G4885: std_logic; attribute dont_touch of G4885: signal is true;
	signal G4888: std_logic; attribute dont_touch of G4888: signal is true;
	signal G4891: std_logic; attribute dont_touch of G4891: signal is true;
	signal G4894: std_logic; attribute dont_touch of G4894: signal is true;
	signal G4897: std_logic; attribute dont_touch of G4897: signal is true;
	signal G4898: std_logic; attribute dont_touch of G4898: signal is true;
	signal G4899: std_logic; attribute dont_touch of G4899: signal is true;
	signal G4902: std_logic; attribute dont_touch of G4902: signal is true;
	signal G4905: std_logic; attribute dont_touch of G4905: signal is true;
	signal G4908: std_logic; attribute dont_touch of G4908: signal is true;
	signal G4911: std_logic; attribute dont_touch of G4911: signal is true;
	signal G4912: std_logic; attribute dont_touch of G4912: signal is true;
	signal G4913: std_logic; attribute dont_touch of G4913: signal is true;
	signal G4916: std_logic; attribute dont_touch of G4916: signal is true;
	signal G4919: std_logic; attribute dont_touch of G4919: signal is true;
	signal G4922: std_logic; attribute dont_touch of G4922: signal is true;
	signal G4925: std_logic; attribute dont_touch of G4925: signal is true;
	signal G4928: std_logic; attribute dont_touch of G4928: signal is true;
	signal G4929: std_logic; attribute dont_touch of G4929: signal is true;
	signal G4930: std_logic; attribute dont_touch of G4930: signal is true;
	signal G4933: std_logic; attribute dont_touch of G4933: signal is true;
	signal G4936: std_logic; attribute dont_touch of G4936: signal is true;
	signal G4939: std_logic; attribute dont_touch of G4939: signal is true;
	signal G4942: std_logic; attribute dont_touch of G4942: signal is true;
	signal G4945: std_logic; attribute dont_touch of G4945: signal is true;
	signal G4948: std_logic; attribute dont_touch of G4948: signal is true;
	signal G4951: std_logic; attribute dont_touch of G4951: signal is true;
	signal G4954: std_logic; attribute dont_touch of G4954: signal is true;
	signal G4955: std_logic; attribute dont_touch of G4955: signal is true;
	signal G4956: std_logic; attribute dont_touch of G4956: signal is true;
	signal G4959: std_logic; attribute dont_touch of G4959: signal is true;
	signal G4962: std_logic; attribute dont_touch of G4962: signal is true;
	signal G4963: std_logic; attribute dont_touch of G4963: signal is true;
	signal G4964: std_logic; attribute dont_touch of G4964: signal is true;
	signal G4967: std_logic; attribute dont_touch of G4967: signal is true;
	signal G4970: std_logic; attribute dont_touch of G4970: signal is true;
	signal G4973: std_logic; attribute dont_touch of G4973: signal is true;
	signal G4976: std_logic; attribute dont_touch of G4976: signal is true;
	signal G4979: std_logic; attribute dont_touch of G4979: signal is true;
	signal G4982: std_logic; attribute dont_touch of G4982: signal is true;
	signal G4985: std_logic; attribute dont_touch of G4985: signal is true;
	signal G4994: std_logic; attribute dont_touch of G4994: signal is true;
	signal G4997: std_logic; attribute dont_touch of G4997: signal is true;
	signal G5000: std_logic; attribute dont_touch of G5000: signal is true;
	signal G5003: std_logic; attribute dont_touch of G5003: signal is true;
	signal G5004: std_logic; attribute dont_touch of G5004: signal is true;
	signal G5005: std_logic; attribute dont_touch of G5005: signal is true;
	signal G5008: std_logic; attribute dont_touch of G5008: signal is true;
	signal G5009: std_logic; attribute dont_touch of G5009: signal is true;
	signal G5012: std_logic; attribute dont_touch of G5012: signal is true;
	signal G5015: std_logic; attribute dont_touch of G5015: signal is true;
	signal G5018: std_logic; attribute dont_touch of G5018: signal is true;
	signal G5021: std_logic; attribute dont_touch of G5021: signal is true;
	signal G5024: std_logic; attribute dont_touch of G5024: signal is true;
	signal G5027: std_logic; attribute dont_touch of G5027: signal is true;
	signal G5030: std_logic; attribute dont_touch of G5030: signal is true;
	signal G5033: std_logic; attribute dont_touch of G5033: signal is true;
	signal G5034: std_logic; attribute dont_touch of G5034: signal is true;
	signal G5035: std_logic; attribute dont_touch of G5035: signal is true;
	signal G5038: std_logic; attribute dont_touch of G5038: signal is true;
	signal G5041: std_logic; attribute dont_touch of G5041: signal is true;
	signal G5044: std_logic; attribute dont_touch of G5044: signal is true;
	signal G5047: std_logic; attribute dont_touch of G5047: signal is true;
	signal G5050: std_logic; attribute dont_touch of G5050: signal is true;
	signal G5053: std_logic; attribute dont_touch of G5053: signal is true;
	signal G5056: std_logic; attribute dont_touch of G5056: signal is true;
	signal G5057: std_logic; attribute dont_touch of G5057: signal is true;
	signal G5058: std_logic; attribute dont_touch of G5058: signal is true;
	signal G5061: std_logic; attribute dont_touch of G5061: signal is true;
	signal G5064: std_logic; attribute dont_touch of G5064: signal is true;
	signal G5067: std_logic; attribute dont_touch of G5067: signal is true;
	signal G5070: std_logic; attribute dont_touch of G5070: signal is true;
	signal G5071: std_logic; attribute dont_touch of G5071: signal is true;
	signal G5072: std_logic; attribute dont_touch of G5072: signal is true;
	signal G5075: std_logic; attribute dont_touch of G5075: signal is true;
	signal G5078: std_logic; attribute dont_touch of G5078: signal is true;
	signal G5081: std_logic; attribute dont_touch of G5081: signal is true;
	signal G5084: std_logic; attribute dont_touch of G5084: signal is true;
	signal G5087: std_logic; attribute dont_touch of G5087: signal is true;
	signal G5088: std_logic; attribute dont_touch of G5088: signal is true;
	signal G5089: std_logic; attribute dont_touch of G5089: signal is true;
	signal G5092: std_logic; attribute dont_touch of G5092: signal is true;
	signal G5095: std_logic; attribute dont_touch of G5095: signal is true;
	signal G5098: std_logic; attribute dont_touch of G5098: signal is true;
	signal G5101: std_logic; attribute dont_touch of G5101: signal is true;
	signal G5104: std_logic; attribute dont_touch of G5104: signal is true;
	signal G5107: std_logic; attribute dont_touch of G5107: signal is true;
	signal G5110: std_logic; attribute dont_touch of G5110: signal is true;
	signal G5113: std_logic; attribute dont_touch of G5113: signal is true;
	signal G5114: std_logic; attribute dont_touch of G5114: signal is true;
	signal G5115: std_logic; attribute dont_touch of G5115: signal is true;
	signal G5118: std_logic; attribute dont_touch of G5118: signal is true;
	signal G5121: std_logic; attribute dont_touch of G5121: signal is true;
	signal G5122: std_logic; attribute dont_touch of G5122: signal is true;
	signal G5123: std_logic; attribute dont_touch of G5123: signal is true;
	signal G5126: std_logic; attribute dont_touch of G5126: signal is true;
	signal G5129: std_logic; attribute dont_touch of G5129: signal is true;
	signal G5132: std_logic; attribute dont_touch of G5132: signal is true;
	signal G5135: std_logic; attribute dont_touch of G5135: signal is true;
	signal G5138: std_logic; attribute dont_touch of G5138: signal is true;
	signal G5141: std_logic; attribute dont_touch of G5141: signal is true;
	signal G5142: std_logic; attribute dont_touch of G5142: signal is true;
	signal G5145: std_logic; attribute dont_touch of G5145: signal is true;
	signal G5148: std_logic; attribute dont_touch of G5148: signal is true;
	signal G5149: std_logic; attribute dont_touch of G5149: signal is true;
	signal G5150: std_logic; attribute dont_touch of G5150: signal is true;
	signal G5153: std_logic; attribute dont_touch of G5153: signal is true;
	signal G5156: std_logic; attribute dont_touch of G5156: signal is true;
	signal G5159: std_logic; attribute dont_touch of G5159: signal is true;
	signal G5162: std_logic; attribute dont_touch of G5162: signal is true;
	signal G5163: std_logic; attribute dont_touch of G5163: signal is true;
	signal G5164: std_logic; attribute dont_touch of G5164: signal is true;
	signal G5167: std_logic; attribute dont_touch of G5167: signal is true;
	signal G5170: std_logic; attribute dont_touch of G5170: signal is true;
	signal G5173: std_logic; attribute dont_touch of G5173: signal is true;
	signal G5176: std_logic; attribute dont_touch of G5176: signal is true;
	signal G5179: std_logic; attribute dont_touch of G5179: signal is true;
	signal G5182: std_logic; attribute dont_touch of G5182: signal is true;
	signal G5185: std_logic; attribute dont_touch of G5185: signal is true;
	signal G5186: std_logic; attribute dont_touch of G5186: signal is true;
	signal G5187: std_logic; attribute dont_touch of G5187: signal is true;
	signal G5190: std_logic; attribute dont_touch of G5190: signal is true;
	signal G5193: std_logic; attribute dont_touch of G5193: signal is true;
	signal G5196: std_logic; attribute dont_touch of G5196: signal is true;
	signal G5199: std_logic; attribute dont_touch of G5199: signal is true;
	signal G5200: std_logic; attribute dont_touch of G5200: signal is true;
	signal G5201: std_logic; attribute dont_touch of G5201: signal is true;
	signal G5204: std_logic; attribute dont_touch of G5204: signal is true;
	signal G5207: std_logic; attribute dont_touch of G5207: signal is true;
	signal G5210: std_logic; attribute dont_touch of G5210: signal is true;
	signal G5213: std_logic; attribute dont_touch of G5213: signal is true;
	signal G5216: std_logic; attribute dont_touch of G5216: signal is true;
	signal G5217: std_logic; attribute dont_touch of G5217: signal is true;
	signal G5218: std_logic; attribute dont_touch of G5218: signal is true;
	signal G5221: std_logic; attribute dont_touch of G5221: signal is true;
	signal G5224: std_logic; attribute dont_touch of G5224: signal is true;
	signal G5227: std_logic; attribute dont_touch of G5227: signal is true;
	signal G5230: std_logic; attribute dont_touch of G5230: signal is true;
	signal G5233: std_logic; attribute dont_touch of G5233: signal is true;
	signal G5234: std_logic; attribute dont_touch of G5234: signal is true;
	signal G5235: std_logic; attribute dont_touch of G5235: signal is true;
	signal G5238: std_logic; attribute dont_touch of G5238: signal is true;
	signal G5241: std_logic; attribute dont_touch of G5241: signal is true;
	signal G5242: std_logic; attribute dont_touch of G5242: signal is true;
	signal G5243: std_logic; attribute dont_touch of G5243: signal is true;
	signal G5246: std_logic; attribute dont_touch of G5246: signal is true;
	signal G5249: std_logic; attribute dont_touch of G5249: signal is true;
	signal G5252: std_logic; attribute dont_touch of G5252: signal is true;
	signal G5255: std_logic; attribute dont_touch of G5255: signal is true;
	signal G5256: std_logic; attribute dont_touch of G5256: signal is true;
	signal G5257: std_logic; attribute dont_touch of G5257: signal is true;
	signal G5260: std_logic; attribute dont_touch of G5260: signal is true;
	signal G5263: std_logic; attribute dont_touch of G5263: signal is true;
	signal G5266: std_logic; attribute dont_touch of G5266: signal is true;
	signal G5269: std_logic; attribute dont_touch of G5269: signal is true;
	signal G5272: std_logic; attribute dont_touch of G5272: signal is true;
	signal G5275: std_logic; attribute dont_touch of G5275: signal is true;
	signal G5278: std_logic; attribute dont_touch of G5278: signal is true;
	signal G5279: std_logic; attribute dont_touch of G5279: signal is true;
	signal G5280: std_logic; attribute dont_touch of G5280: signal is true;
	signal G5283: std_logic; attribute dont_touch of G5283: signal is true;
	signal G5286: std_logic; attribute dont_touch of G5286: signal is true;
	signal G5289: std_logic; attribute dont_touch of G5289: signal is true;
	signal G5292: std_logic; attribute dont_touch of G5292: signal is true;
	signal G5293: std_logic; attribute dont_touch of G5293: signal is true;
	signal G5296: std_logic; attribute dont_touch of G5296: signal is true;
	signal G5297: std_logic; attribute dont_touch of G5297: signal is true;
	signal G5298: std_logic; attribute dont_touch of G5298: signal is true;
	signal G5301: std_logic; attribute dont_touch of G5301: signal is true;
	signal G5304: std_logic; attribute dont_touch of G5304: signal is true;
	signal G5305: std_logic; attribute dont_touch of G5305: signal is true;
	signal G5306: std_logic; attribute dont_touch of G5306: signal is true;
	signal G5309: std_logic; attribute dont_touch of G5309: signal is true;
	signal G5312: std_logic; attribute dont_touch of G5312: signal is true;
	signal G5315: std_logic; attribute dont_touch of G5315: signal is true;
	signal G5318: std_logic; attribute dont_touch of G5318: signal is true;
	signal G5319: std_logic; attribute dont_touch of G5319: signal is true;
	signal G5320: std_logic; attribute dont_touch of G5320: signal is true;
	signal G5323: std_logic; attribute dont_touch of G5323: signal is true;
	signal G5326: std_logic; attribute dont_touch of G5326: signal is true;
	signal G5327: std_logic; attribute dont_touch of G5327: signal is true;
	signal G5330: std_logic; attribute dont_touch of G5330: signal is true;
	signal G5333: std_logic; attribute dont_touch of G5333: signal is true;
	signal G5334: std_logic; attribute dont_touch of G5334: signal is true;
	signal G5335: std_logic; attribute dont_touch of G5335: signal is true;
	signal G5338: std_logic; attribute dont_touch of G5338: signal is true;
	signal G5341: std_logic; attribute dont_touch of G5341: signal is true;
	signal G5342: std_logic; attribute dont_touch of G5342: signal is true;
	signal G5343: std_logic; attribute dont_touch of G5343: signal is true;
	signal G5346: std_logic; attribute dont_touch of G5346: signal is true;
	signal G5349: std_logic; attribute dont_touch of G5349: signal is true;
	signal G5352: std_logic; attribute dont_touch of G5352: signal is true;
	signal G5355: std_logic; attribute dont_touch of G5355: signal is true;
	signal G5358: std_logic; attribute dont_touch of G5358: signal is true;
	signal G5361: std_logic; attribute dont_touch of G5361: signal is true;
	signal G5362: std_logic; attribute dont_touch of G5362: signal is true;
	signal G5363: std_logic; attribute dont_touch of G5363: signal is true;
	signal G5366: std_logic; attribute dont_touch of G5366: signal is true;
	signal G5369: std_logic; attribute dont_touch of G5369: signal is true;
	signal G5372: std_logic; attribute dont_touch of G5372: signal is true;
	signal G5375: std_logic; attribute dont_touch of G5375: signal is true;
	signal G5378: std_logic; attribute dont_touch of G5378: signal is true;
	signal G5379: std_logic; attribute dont_touch of G5379: signal is true;
	signal G5382: std_logic; attribute dont_touch of G5382: signal is true;
	signal G5385: std_logic; attribute dont_touch of G5385: signal is true;
	signal G5389: std_logic; attribute dont_touch of G5389: signal is true;
	signal G5390: std_logic; attribute dont_touch of G5390: signal is true;
	signal G5391: std_logic; attribute dont_touch of G5391: signal is true;
	signal G5394: std_logic; attribute dont_touch of G5394: signal is true;
	signal G5395: std_logic; attribute dont_touch of G5395: signal is true;
	signal G5396: std_logic; attribute dont_touch of G5396: signal is true;
	signal G5397: std_logic; attribute dont_touch of G5397: signal is true;
	signal G5398: std_logic; attribute dont_touch of G5398: signal is true;
	signal G5399: std_logic; attribute dont_touch of G5399: signal is true;
	signal G5400: std_logic; attribute dont_touch of G5400: signal is true;
	signal G5401: std_logic; attribute dont_touch of G5401: signal is true;
	signal G5402: std_logic; attribute dont_touch of G5402: signal is true;
	signal G5403: std_logic; attribute dont_touch of G5403: signal is true;
	signal G5404: std_logic; attribute dont_touch of G5404: signal is true;
	signal G5405: std_logic; attribute dont_touch of G5405: signal is true;
	signal G5406: std_logic; attribute dont_touch of G5406: signal is true;
	signal G5407: std_logic; attribute dont_touch of G5407: signal is true;
	signal G5408: std_logic; attribute dont_touch of G5408: signal is true;
	signal G5409: std_logic; attribute dont_touch of G5409: signal is true;
	signal G5410: std_logic; attribute dont_touch of G5410: signal is true;
	signal G5411: std_logic; attribute dont_touch of G5411: signal is true;
	signal G5412: std_logic; attribute dont_touch of G5412: signal is true;
	signal G5413: std_logic; attribute dont_touch of G5413: signal is true;
	signal G5414: std_logic; attribute dont_touch of G5414: signal is true;
	signal G5415: std_logic; attribute dont_touch of G5415: signal is true;
	signal G5416: std_logic; attribute dont_touch of G5416: signal is true;
	signal G5417: std_logic; attribute dont_touch of G5417: signal is true;
	signal G5418: std_logic; attribute dont_touch of G5418: signal is true;
	signal G5419: std_logic; attribute dont_touch of G5419: signal is true;
	signal G5420: std_logic; attribute dont_touch of G5420: signal is true;
	signal G5421: std_logic; attribute dont_touch of G5421: signal is true;
	signal G5422: std_logic; attribute dont_touch of G5422: signal is true;
	signal G5423: std_logic; attribute dont_touch of G5423: signal is true;
	signal G5424: std_logic; attribute dont_touch of G5424: signal is true;
	signal G5425: std_logic; attribute dont_touch of G5425: signal is true;
	signal G5426: std_logic; attribute dont_touch of G5426: signal is true;
	signal G5427: std_logic; attribute dont_touch of G5427: signal is true;
	signal G5428: std_logic; attribute dont_touch of G5428: signal is true;
	signal G5431: std_logic; attribute dont_touch of G5431: signal is true;
	signal G5434: std_logic; attribute dont_touch of G5434: signal is true;
	signal G5438: std_logic; attribute dont_touch of G5438: signal is true;
	signal G5469: std_logic; attribute dont_touch of G5469: signal is true;
	signal G5473: std_logic; attribute dont_touch of G5473: signal is true;
	signal G5504: std_logic; attribute dont_touch of G5504: signal is true;
	signal G5507: std_logic; attribute dont_touch of G5507: signal is true;
	signal G5508: std_logic; attribute dont_touch of G5508: signal is true;
	signal G5512: std_logic; attribute dont_touch of G5512: signal is true;
	signal G5543: std_logic; attribute dont_touch of G5543: signal is true;
	signal G5546: std_logic; attribute dont_touch of G5546: signal is true;
	signal G5547: std_logic; attribute dont_touch of G5547: signal is true;
	signal G5548: std_logic; attribute dont_touch of G5548: signal is true;
	signal G5550: std_logic; attribute dont_touch of G5550: signal is true;
	signal G5551: std_logic; attribute dont_touch of G5551: signal is true;
	signal G5552: std_logic; attribute dont_touch of G5552: signal is true;
	signal G5556: std_logic; attribute dont_touch of G5556: signal is true;
	signal G5587: std_logic; attribute dont_touch of G5587: signal is true;
	signal G5590: std_logic; attribute dont_touch of G5590: signal is true;
	signal G5591: std_logic; attribute dont_touch of G5591: signal is true;
	signal G5592: std_logic; attribute dont_touch of G5592: signal is true;
	signal G5593: std_logic; attribute dont_touch of G5593: signal is true;
	signal G5594: std_logic; attribute dont_touch of G5594: signal is true;
	signal G5596: std_logic; attribute dont_touch of G5596: signal is true;
	signal G5597: std_logic; attribute dont_touch of G5597: signal is true;
	signal G5598: std_logic; attribute dont_touch of G5598: signal is true;
	signal G5601: std_logic; attribute dont_touch of G5601: signal is true;
	signal G5604: std_logic; attribute dont_touch of G5604: signal is true;
	signal G5605: std_logic; attribute dont_touch of G5605: signal is true;
	signal G5606: std_logic; attribute dont_touch of G5606: signal is true;
	signal G5609: std_logic; attribute dont_touch of G5609: signal is true;
	signal G5610: std_logic; attribute dont_touch of G5610: signal is true;
	signal G5611: std_logic; attribute dont_touch of G5611: signal is true;
	signal G5613: std_logic; attribute dont_touch of G5613: signal is true;
	signal G5614: std_logic; attribute dont_touch of G5614: signal is true;
	signal G5615: std_logic; attribute dont_touch of G5615: signal is true;
	signal G5618: std_logic; attribute dont_touch of G5618: signal is true;
	signal G5621: std_logic; attribute dont_touch of G5621: signal is true;
	signal G5622: std_logic; attribute dont_touch of G5622: signal is true;
	signal G5623: std_logic; attribute dont_touch of G5623: signal is true;
	signal G5626: std_logic; attribute dont_touch of G5626: signal is true;
	signal G5627: std_logic; attribute dont_touch of G5627: signal is true;
	signal G5628: std_logic; attribute dont_touch of G5628: signal is true;
	signal G5630: std_logic; attribute dont_touch of G5630: signal is true;
	signal G5631: std_logic; attribute dont_touch of G5631: signal is true;
	signal G5634: std_logic; attribute dont_touch of G5634: signal is true;
	signal G5635: std_logic; attribute dont_touch of G5635: signal is true;
	signal G5636: std_logic; attribute dont_touch of G5636: signal is true;
	signal G5638: std_logic; attribute dont_touch of G5638: signal is true;
	signal G5639: std_logic; attribute dont_touch of G5639: signal is true;
	signal G5640: std_logic; attribute dont_touch of G5640: signal is true;
	signal G5641: std_logic; attribute dont_touch of G5641: signal is true;
	signal G5642: std_logic; attribute dont_touch of G5642: signal is true;
	signal G5645: std_logic; attribute dont_touch of G5645: signal is true;
	signal G5646: std_logic; attribute dont_touch of G5646: signal is true;
	signal G5647: std_logic; attribute dont_touch of G5647: signal is true;
	signal G5649: std_logic; attribute dont_touch of G5649: signal is true;
	signal G5650: std_logic; attribute dont_touch of G5650: signal is true;
	signal G5651: std_logic; attribute dont_touch of G5651: signal is true;
	signal G5654: std_logic; attribute dont_touch of G5654: signal is true;
	signal G5655: std_logic; attribute dont_touch of G5655: signal is true;
	signal G5656: std_logic; attribute dont_touch of G5656: signal is true;
	signal G5658: std_logic; attribute dont_touch of G5658: signal is true;
	signal G5659: std_logic; attribute dont_touch of G5659: signal is true;
	signal G5662: std_logic; attribute dont_touch of G5662: signal is true;
	signal G5663: std_logic; attribute dont_touch of G5663: signal is true;
	signal G5664: std_logic; attribute dont_touch of G5664: signal is true;
	signal G5665: std_logic; attribute dont_touch of G5665: signal is true;
	signal G5666: std_logic; attribute dont_touch of G5666: signal is true;
	signal G5667: std_logic; attribute dont_touch of G5667: signal is true;
	signal G5668: std_logic; attribute dont_touch of G5668: signal is true;
	signal G5675: std_logic; attribute dont_touch of G5675: signal is true;
	signal G5676: std_logic; attribute dont_touch of G5676: signal is true;
	signal G5677: std_logic; attribute dont_touch of G5677: signal is true;
	signal G5678: std_logic; attribute dont_touch of G5678: signal is true;
	signal G5679: std_logic; attribute dont_touch of G5679: signal is true;
	signal G5680: std_logic; attribute dont_touch of G5680: signal is true;
	signal G5683: std_logic; attribute dont_touch of G5683: signal is true;
	signal G5684: std_logic; attribute dont_touch of G5684: signal is true;
	signal G5685: std_logic; attribute dont_touch of G5685: signal is true;
	signal G5687: std_logic; attribute dont_touch of G5687: signal is true;
	signal G5688: std_logic; attribute dont_touch of G5688: signal is true;
	signal G5689: std_logic; attribute dont_touch of G5689: signal is true;
	signal G5692: std_logic; attribute dont_touch of G5692: signal is true;
	signal G5693: std_logic; attribute dont_touch of G5693: signal is true;
	signal G5694: std_logic; attribute dont_touch of G5694: signal is true;
	signal G5696: std_logic; attribute dont_touch of G5696: signal is true;
	signal G5697: std_logic; attribute dont_touch of G5697: signal is true;
	signal G5700: std_logic; attribute dont_touch of G5700: signal is true;
	signal G5701: std_logic; attribute dont_touch of G5701: signal is true;
	signal G5702: std_logic; attribute dont_touch of G5702: signal is true;
	signal G5703: std_logic; attribute dont_touch of G5703: signal is true;
	signal G5704: std_logic; attribute dont_touch of G5704: signal is true;
	signal G5705: std_logic; attribute dont_touch of G5705: signal is true;
	signal G5706: std_logic; attribute dont_touch of G5706: signal is true;
	signal G5707: std_logic; attribute dont_touch of G5707: signal is true;
	signal G5708: std_logic; attribute dont_touch of G5708: signal is true;
	signal G5709: std_logic; attribute dont_touch of G5709: signal is true;
	signal G5710: std_logic; attribute dont_touch of G5710: signal is true;
	signal G5711: std_logic; attribute dont_touch of G5711: signal is true;
	signal G5712: std_logic; attribute dont_touch of G5712: signal is true;
	signal G5713: std_logic; attribute dont_touch of G5713: signal is true;
	signal G5714: std_logic; attribute dont_touch of G5714: signal is true;
	signal G5715: std_logic; attribute dont_touch of G5715: signal is true;
	signal G5716: std_logic; attribute dont_touch of G5716: signal is true;
	signal G5717: std_logic; attribute dont_touch of G5717: signal is true;
	signal G5718: std_logic; attribute dont_touch of G5718: signal is true;
	signal G5719: std_logic; attribute dont_touch of G5719: signal is true;
	signal G5720: std_logic; attribute dont_touch of G5720: signal is true;
	signal G5727: std_logic; attribute dont_touch of G5727: signal is true;
	signal G5728: std_logic; attribute dont_touch of G5728: signal is true;
	signal G5729: std_logic; attribute dont_touch of G5729: signal is true;
	signal G5730: std_logic; attribute dont_touch of G5730: signal is true;
	signal G5731: std_logic; attribute dont_touch of G5731: signal is true;
	signal G5732: std_logic; attribute dont_touch of G5732: signal is true;
	signal G5735: std_logic; attribute dont_touch of G5735: signal is true;
	signal G5736: std_logic; attribute dont_touch of G5736: signal is true;
	signal G5737: std_logic; attribute dont_touch of G5737: signal is true;
	signal G5739: std_logic; attribute dont_touch of G5739: signal is true;
	signal G5740: std_logic; attribute dont_touch of G5740: signal is true;
	signal G5741: std_logic; attribute dont_touch of G5741: signal is true;
	signal G5744: std_logic; attribute dont_touch of G5744: signal is true;
	signal G5745: std_logic; attribute dont_touch of G5745: signal is true;
	signal G5746: std_logic; attribute dont_touch of G5746: signal is true;
	signal G5748: std_logic; attribute dont_touch of G5748: signal is true;
	signal G5749: std_logic; attribute dont_touch of G5749: signal is true;
	signal G5750: std_logic; attribute dont_touch of G5750: signal is true;
	signal G5751: std_logic; attribute dont_touch of G5751: signal is true;
	signal G5752: std_logic; attribute dont_touch of G5752: signal is true;
	signal G5753: std_logic; attribute dont_touch of G5753: signal is true;
	signal G5754: std_logic; attribute dont_touch of G5754: signal is true;
	signal G5755: std_logic; attribute dont_touch of G5755: signal is true;
	signal G5756: std_logic; attribute dont_touch of G5756: signal is true;
	signal G5757: std_logic; attribute dont_touch of G5757: signal is true;
	signal G5758: std_logic; attribute dont_touch of G5758: signal is true;
	signal G5759: std_logic; attribute dont_touch of G5759: signal is true;
	signal G5760: std_logic; attribute dont_touch of G5760: signal is true;
	signal G5761: std_logic; attribute dont_touch of G5761: signal is true;
	signal G5762: std_logic; attribute dont_touch of G5762: signal is true;
	signal G5763: std_logic; attribute dont_touch of G5763: signal is true;
	signal G5764: std_logic; attribute dont_touch of G5764: signal is true;
	signal G5765: std_logic; attribute dont_touch of G5765: signal is true;
	signal G5766: std_logic; attribute dont_touch of G5766: signal is true;
	signal G5767: std_logic; attribute dont_touch of G5767: signal is true;
	signal G5768: std_logic; attribute dont_touch of G5768: signal is true;
	signal G5769: std_logic; attribute dont_touch of G5769: signal is true;
	signal G5770: std_logic; attribute dont_touch of G5770: signal is true;
	signal G5771: std_logic; attribute dont_touch of G5771: signal is true;
	signal G5772: std_logic; attribute dont_touch of G5772: signal is true;
	signal G5773: std_logic; attribute dont_touch of G5773: signal is true;
	signal G5774: std_logic; attribute dont_touch of G5774: signal is true;
	signal G5775: std_logic; attribute dont_touch of G5775: signal is true;
	signal G5776: std_logic; attribute dont_touch of G5776: signal is true;
	signal G5777: std_logic; attribute dont_touch of G5777: signal is true;
	signal G5778: std_logic; attribute dont_touch of G5778: signal is true;
	signal G5785: std_logic; attribute dont_touch of G5785: signal is true;
	signal G5786: std_logic; attribute dont_touch of G5786: signal is true;
	signal G5787: std_logic; attribute dont_touch of G5787: signal is true;
	signal G5788: std_logic; attribute dont_touch of G5788: signal is true;
	signal G5789: std_logic; attribute dont_touch of G5789: signal is true;
	signal G5790: std_logic; attribute dont_touch of G5790: signal is true;
	signal G5793: std_logic; attribute dont_touch of G5793: signal is true;
	signal G5794: std_logic; attribute dont_touch of G5794: signal is true;
	signal G5795: std_logic; attribute dont_touch of G5795: signal is true;
	signal G5797: std_logic; attribute dont_touch of G5797: signal is true;
	signal G5798: std_logic; attribute dont_touch of G5798: signal is true;
	signal G5799: std_logic; attribute dont_touch of G5799: signal is true;
	signal G5800: std_logic; attribute dont_touch of G5800: signal is true;
	signal G5801: std_logic; attribute dont_touch of G5801: signal is true;
	signal G5802: std_logic; attribute dont_touch of G5802: signal is true;
	signal G5803: std_logic; attribute dont_touch of G5803: signal is true;
	signal G5804: std_logic; attribute dont_touch of G5804: signal is true;
	signal G5805: std_logic; attribute dont_touch of G5805: signal is true;
	signal G5806: std_logic; attribute dont_touch of G5806: signal is true;
	signal G5807: std_logic; attribute dont_touch of G5807: signal is true;
	signal G5808: std_logic; attribute dont_touch of G5808: signal is true;
	signal G5809: std_logic; attribute dont_touch of G5809: signal is true;
	signal G5810: std_logic; attribute dont_touch of G5810: signal is true;
	signal G5811: std_logic; attribute dont_touch of G5811: signal is true;
	signal G5812: std_logic; attribute dont_touch of G5812: signal is true;
	signal G5813: std_logic; attribute dont_touch of G5813: signal is true;
	signal G5814: std_logic; attribute dont_touch of G5814: signal is true;
	signal G5815: std_logic; attribute dont_touch of G5815: signal is true;
	signal G5816: std_logic; attribute dont_touch of G5816: signal is true;
	signal G5817: std_logic; attribute dont_touch of G5817: signal is true;
	signal G5818: std_logic; attribute dont_touch of G5818: signal is true;
	signal G5819: std_logic; attribute dont_touch of G5819: signal is true;
	signal G5820: std_logic; attribute dont_touch of G5820: signal is true;
	signal G5821: std_logic; attribute dont_touch of G5821: signal is true;
	signal G5822: std_logic; attribute dont_touch of G5822: signal is true;
	signal G5823: std_logic; attribute dont_touch of G5823: signal is true;
	signal G5824: std_logic; attribute dont_touch of G5824: signal is true;
	signal G5825: std_logic; attribute dont_touch of G5825: signal is true;
	signal G5826: std_logic; attribute dont_touch of G5826: signal is true;
	signal G5827: std_logic; attribute dont_touch of G5827: signal is true;
	signal G5828: std_logic; attribute dont_touch of G5828: signal is true;
	signal G5829: std_logic; attribute dont_touch of G5829: signal is true;
	signal G5830: std_logic; attribute dont_touch of G5830: signal is true;
	signal G5831: std_logic; attribute dont_touch of G5831: signal is true;
	signal G5832: std_logic; attribute dont_touch of G5832: signal is true;
	signal G5833: std_logic; attribute dont_touch of G5833: signal is true;
	signal G5834: std_logic; attribute dont_touch of G5834: signal is true;
	signal G5835: std_logic; attribute dont_touch of G5835: signal is true;
	signal G5836: std_logic; attribute dont_touch of G5836: signal is true;
	signal G5837: std_logic; attribute dont_touch of G5837: signal is true;
	signal G5844: std_logic; attribute dont_touch of G5844: signal is true;
	signal G5845: std_logic; attribute dont_touch of G5845: signal is true;
	signal G5846: std_logic; attribute dont_touch of G5846: signal is true;
	signal G5847: std_logic; attribute dont_touch of G5847: signal is true;
	signal G5848: std_logic; attribute dont_touch of G5848: signal is true;
	signal G5849: std_logic; attribute dont_touch of G5849: signal is true;
	signal G5850: std_logic; attribute dont_touch of G5850: signal is true;
	signal G5851: std_logic; attribute dont_touch of G5851: signal is true;
	signal G5852: std_logic; attribute dont_touch of G5852: signal is true;
	signal G5853: std_logic; attribute dont_touch of G5853: signal is true;
	signal G5854: std_logic; attribute dont_touch of G5854: signal is true;
	signal G5855: std_logic; attribute dont_touch of G5855: signal is true;
	signal G5856: std_logic; attribute dont_touch of G5856: signal is true;
	signal G5857: std_logic; attribute dont_touch of G5857: signal is true;
	signal G5858: std_logic; attribute dont_touch of G5858: signal is true;
	signal G5859: std_logic; attribute dont_touch of G5859: signal is true;
	signal G5860: std_logic; attribute dont_touch of G5860: signal is true;
	signal G5861: std_logic; attribute dont_touch of G5861: signal is true;
	signal G5862: std_logic; attribute dont_touch of G5862: signal is true;
	signal G5863: std_logic; attribute dont_touch of G5863: signal is true;
	signal G5864: std_logic; attribute dont_touch of G5864: signal is true;
	signal G5865: std_logic; attribute dont_touch of G5865: signal is true;
	signal G5866: std_logic; attribute dont_touch of G5866: signal is true;
	signal G5867: std_logic; attribute dont_touch of G5867: signal is true;
	signal G5868: std_logic; attribute dont_touch of G5868: signal is true;
	signal G5869: std_logic; attribute dont_touch of G5869: signal is true;
	signal G5870: std_logic; attribute dont_touch of G5870: signal is true;
	signal G5871: std_logic; attribute dont_touch of G5871: signal is true;
	signal G5872: std_logic; attribute dont_touch of G5872: signal is true;
	signal G5873: std_logic; attribute dont_touch of G5873: signal is true;
	signal G5874: std_logic; attribute dont_touch of G5874: signal is true;
	signal G5875: std_logic; attribute dont_touch of G5875: signal is true;
	signal G5876: std_logic; attribute dont_touch of G5876: signal is true;
	signal G5877: std_logic; attribute dont_touch of G5877: signal is true;
	signal G5878: std_logic; attribute dont_touch of G5878: signal is true;
	signal G5879: std_logic; attribute dont_touch of G5879: signal is true;
	signal G5880: std_logic; attribute dont_touch of G5880: signal is true;
	signal G5881: std_logic; attribute dont_touch of G5881: signal is true;
	signal G5882: std_logic; attribute dont_touch of G5882: signal is true;
	signal G5883: std_logic; attribute dont_touch of G5883: signal is true;
	signal G5884: std_logic; attribute dont_touch of G5884: signal is true;
	signal G5885: std_logic; attribute dont_touch of G5885: signal is true;
	signal G5886: std_logic; attribute dont_touch of G5886: signal is true;
	signal G5887: std_logic; attribute dont_touch of G5887: signal is true;
	signal G5888: std_logic; attribute dont_touch of G5888: signal is true;
	signal G5889: std_logic; attribute dont_touch of G5889: signal is true;
	signal G5890: std_logic; attribute dont_touch of G5890: signal is true;
	signal G5893: std_logic; attribute dont_touch of G5893: signal is true;
	signal G5894: std_logic; attribute dont_touch of G5894: signal is true;
	signal G5895: std_logic; attribute dont_touch of G5895: signal is true;
	signal G5896: std_logic; attribute dont_touch of G5896: signal is true;
	signal G5897: std_logic; attribute dont_touch of G5897: signal is true;
	signal G5898: std_logic; attribute dont_touch of G5898: signal is true;
	signal G5899: std_logic; attribute dont_touch of G5899: signal is true;
	signal G5900: std_logic; attribute dont_touch of G5900: signal is true;
	signal G5901: std_logic; attribute dont_touch of G5901: signal is true;
	signal G5902: std_logic; attribute dont_touch of G5902: signal is true;
	signal G5903: std_logic; attribute dont_touch of G5903: signal is true;
	signal G5904: std_logic; attribute dont_touch of G5904: signal is true;
	signal G5905: std_logic; attribute dont_touch of G5905: signal is true;
	signal G5906: std_logic; attribute dont_touch of G5906: signal is true;
	signal G5907: std_logic; attribute dont_touch of G5907: signal is true;
	signal G5908: std_logic; attribute dont_touch of G5908: signal is true;
	signal G5909: std_logic; attribute dont_touch of G5909: signal is true;
	signal G5910: std_logic; attribute dont_touch of G5910: signal is true;
	signal G5911: std_logic; attribute dont_touch of G5911: signal is true;
	signal G5912: std_logic; attribute dont_touch of G5912: signal is true;
	signal G5913: std_logic; attribute dont_touch of G5913: signal is true;
	signal G5914: std_logic; attribute dont_touch of G5914: signal is true;
	signal G5915: std_logic; attribute dont_touch of G5915: signal is true;
	signal G5916: std_logic; attribute dont_touch of G5916: signal is true;
	signal G5917: std_logic; attribute dont_touch of G5917: signal is true;
	signal G5918: std_logic; attribute dont_touch of G5918: signal is true;
	signal G5919: std_logic; attribute dont_touch of G5919: signal is true;
	signal G5920: std_logic; attribute dont_touch of G5920: signal is true;
	signal G5921: std_logic; attribute dont_touch of G5921: signal is true;
	signal G5922: std_logic; attribute dont_touch of G5922: signal is true;
	signal G5923: std_logic; attribute dont_touch of G5923: signal is true;
	signal G5924: std_logic; attribute dont_touch of G5924: signal is true;
	signal G5925: std_logic; attribute dont_touch of G5925: signal is true;
	signal G5926: std_logic; attribute dont_touch of G5926: signal is true;
	signal G5927: std_logic; attribute dont_touch of G5927: signal is true;
	signal G5928: std_logic; attribute dont_touch of G5928: signal is true;
	signal G5929: std_logic; attribute dont_touch of G5929: signal is true;
	signal G5932: std_logic; attribute dont_touch of G5932: signal is true;
	signal G5933: std_logic; attribute dont_touch of G5933: signal is true;
	signal G5934: std_logic; attribute dont_touch of G5934: signal is true;
	signal G5935: std_logic; attribute dont_touch of G5935: signal is true;
	signal G5936: std_logic; attribute dont_touch of G5936: signal is true;
	signal G5937: std_logic; attribute dont_touch of G5937: signal is true;
	signal G5938: std_logic; attribute dont_touch of G5938: signal is true;
	signal G5939: std_logic; attribute dont_touch of G5939: signal is true;
	signal G5940: std_logic; attribute dont_touch of G5940: signal is true;
	signal G5941: std_logic; attribute dont_touch of G5941: signal is true;
	signal G5942: std_logic; attribute dont_touch of G5942: signal is true;
	signal G5943: std_logic; attribute dont_touch of G5943: signal is true;
	signal G5944: std_logic; attribute dont_touch of G5944: signal is true;
	signal G5945: std_logic; attribute dont_touch of G5945: signal is true;
	signal G5946: std_logic; attribute dont_touch of G5946: signal is true;
	signal G5947: std_logic; attribute dont_touch of G5947: signal is true;
	signal G5948: std_logic; attribute dont_touch of G5948: signal is true;
	signal G5949: std_logic; attribute dont_touch of G5949: signal is true;
	signal G5950: std_logic; attribute dont_touch of G5950: signal is true;
	signal G5951: std_logic; attribute dont_touch of G5951: signal is true;
	signal G5952: std_logic; attribute dont_touch of G5952: signal is true;
	signal G5953: std_logic; attribute dont_touch of G5953: signal is true;
	signal G5954: std_logic; attribute dont_touch of G5954: signal is true;
	signal G5955: std_logic; attribute dont_touch of G5955: signal is true;
	signal G5956: std_logic; attribute dont_touch of G5956: signal is true;
	signal G5957: std_logic; attribute dont_touch of G5957: signal is true;
	signal G5958: std_logic; attribute dont_touch of G5958: signal is true;
	signal G5959: std_logic; attribute dont_touch of G5959: signal is true;
	signal G5960: std_logic; attribute dont_touch of G5960: signal is true;
	signal G5961: std_logic; attribute dont_touch of G5961: signal is true;
	signal G5962: std_logic; attribute dont_touch of G5962: signal is true;
	signal G5963: std_logic; attribute dont_touch of G5963: signal is true;
	signal G5966: std_logic; attribute dont_touch of G5966: signal is true;
	signal G5967: std_logic; attribute dont_touch of G5967: signal is true;
	signal G5968: std_logic; attribute dont_touch of G5968: signal is true;
	signal G5969: std_logic; attribute dont_touch of G5969: signal is true;
	signal G5970: std_logic; attribute dont_touch of G5970: signal is true;
	signal G5971: std_logic; attribute dont_touch of G5971: signal is true;
	signal G5972: std_logic; attribute dont_touch of G5972: signal is true;
	signal G5973: std_logic; attribute dont_touch of G5973: signal is true;
	signal G5974: std_logic; attribute dont_touch of G5974: signal is true;
	signal G5975: std_logic; attribute dont_touch of G5975: signal is true;
	signal G5976: std_logic; attribute dont_touch of G5976: signal is true;
	signal G5977: std_logic; attribute dont_touch of G5977: signal is true;
	signal G5978: std_logic; attribute dont_touch of G5978: signal is true;
	signal G5979: std_logic; attribute dont_touch of G5979: signal is true;
	signal G5980: std_logic; attribute dont_touch of G5980: signal is true;
	signal G5981: std_logic; attribute dont_touch of G5981: signal is true;
	signal G5982: std_logic; attribute dont_touch of G5982: signal is true;
	signal G5983: std_logic; attribute dont_touch of G5983: signal is true;
	signal G5984: std_logic; attribute dont_touch of G5984: signal is true;
	signal G5985: std_logic; attribute dont_touch of G5985: signal is true;
	signal G5986: std_logic; attribute dont_touch of G5986: signal is true;
	signal G5987: std_logic; attribute dont_touch of G5987: signal is true;
	signal G5988: std_logic; attribute dont_touch of G5988: signal is true;
	signal G5989: std_logic; attribute dont_touch of G5989: signal is true;
	signal G5990: std_logic; attribute dont_touch of G5990: signal is true;
	signal G5991: std_logic; attribute dont_touch of G5991: signal is true;
	signal G5992: std_logic; attribute dont_touch of G5992: signal is true;
	signal G5995: std_logic; attribute dont_touch of G5995: signal is true;
	signal G5996: std_logic; attribute dont_touch of G5996: signal is true;
	signal G5997: std_logic; attribute dont_touch of G5997: signal is true;
	signal G5998: std_logic; attribute dont_touch of G5998: signal is true;
	signal G5999: std_logic; attribute dont_touch of G5999: signal is true;
	signal G6000: std_logic; attribute dont_touch of G6000: signal is true;
	signal G6014: std_logic; attribute dont_touch of G6014: signal is true;
	signal G6015: std_logic; attribute dont_touch of G6015: signal is true;
	signal G6016: std_logic; attribute dont_touch of G6016: signal is true;
	signal G6017: std_logic; attribute dont_touch of G6017: signal is true;
	signal G6018: std_logic; attribute dont_touch of G6018: signal is true;
	signal G6019: std_logic; attribute dont_touch of G6019: signal is true;
	signal G6020: std_logic; attribute dont_touch of G6020: signal is true;
	signal G6021: std_logic; attribute dont_touch of G6021: signal is true;
	signal G6022: std_logic; attribute dont_touch of G6022: signal is true;
	signal G6023: std_logic; attribute dont_touch of G6023: signal is true;
	signal G6024: std_logic; attribute dont_touch of G6024: signal is true;
	signal G6025: std_logic; attribute dont_touch of G6025: signal is true;
	signal G6026: std_logic; attribute dont_touch of G6026: signal is true;
	signal G6027: std_logic; attribute dont_touch of G6027: signal is true;
	signal G6028: std_logic; attribute dont_touch of G6028: signal is true;
	signal G6029: std_logic; attribute dont_touch of G6029: signal is true;
	signal G6030: std_logic; attribute dont_touch of G6030: signal is true;
	signal G6031: std_logic; attribute dont_touch of G6031: signal is true;
	signal G6032: std_logic; attribute dont_touch of G6032: signal is true;
	signal G6033: std_logic; attribute dont_touch of G6033: signal is true;
	signal G6034: std_logic; attribute dont_touch of G6034: signal is true;
	signal G6035: std_logic; attribute dont_touch of G6035: signal is true;
	signal G6036: std_logic; attribute dont_touch of G6036: signal is true;
	signal G6037: std_logic; attribute dont_touch of G6037: signal is true;
	signal G6038: std_logic; attribute dont_touch of G6038: signal is true;
	signal G6039: std_logic; attribute dont_touch of G6039: signal is true;
	signal G6040: std_logic; attribute dont_touch of G6040: signal is true;
	signal G6041: std_logic; attribute dont_touch of G6041: signal is true;
	signal G6042: std_logic; attribute dont_touch of G6042: signal is true;
	signal G6043: std_logic; attribute dont_touch of G6043: signal is true;
	signal G6044: std_logic; attribute dont_touch of G6044: signal is true;
	signal G6045: std_logic; attribute dont_touch of G6045: signal is true;
	signal G6046: std_logic; attribute dont_touch of G6046: signal is true;
	signal G6047: std_logic; attribute dont_touch of G6047: signal is true;
	signal G6048: std_logic; attribute dont_touch of G6048: signal is true;
	signal G6051: std_logic; attribute dont_touch of G6051: signal is true;
	signal G6052: std_logic; attribute dont_touch of G6052: signal is true;
	signal G6053: std_logic; attribute dont_touch of G6053: signal is true;
	signal G6054: std_logic; attribute dont_touch of G6054: signal is true;
	signal G6055: std_logic; attribute dont_touch of G6055: signal is true;
	signal G6056: std_logic; attribute dont_touch of G6056: signal is true;
	signal G6057: std_logic; attribute dont_touch of G6057: signal is true;
	signal G6058: std_logic; attribute dont_touch of G6058: signal is true;
	signal G6059: std_logic; attribute dont_touch of G6059: signal is true;
	signal G6060: std_logic; attribute dont_touch of G6060: signal is true;
	signal G6061: std_logic; attribute dont_touch of G6061: signal is true;
	signal G6062: std_logic; attribute dont_touch of G6062: signal is true;
	signal G6063: std_logic; attribute dont_touch of G6063: signal is true;
	signal G6064: std_logic; attribute dont_touch of G6064: signal is true;
	signal G6065: std_logic; attribute dont_touch of G6065: signal is true;
	signal G6066: std_logic; attribute dont_touch of G6066: signal is true;
	signal G6067: std_logic; attribute dont_touch of G6067: signal is true;
	signal G6068: std_logic; attribute dont_touch of G6068: signal is true;
	signal G6079: std_logic; attribute dont_touch of G6079: signal is true;
	signal G6080: std_logic; attribute dont_touch of G6080: signal is true;
	signal G6081: std_logic; attribute dont_touch of G6081: signal is true;
	signal G6082: std_logic; attribute dont_touch of G6082: signal is true;
	signal G6083: std_logic; attribute dont_touch of G6083: signal is true;
	signal G6084: std_logic; attribute dont_touch of G6084: signal is true;
	signal G6085: std_logic; attribute dont_touch of G6085: signal is true;
	signal G6086: std_logic; attribute dont_touch of G6086: signal is true;
	signal G6087: std_logic; attribute dont_touch of G6087: signal is true;
	signal G6098: std_logic; attribute dont_touch of G6098: signal is true;
	signal G6099: std_logic; attribute dont_touch of G6099: signal is true;
	signal G6100: std_logic; attribute dont_touch of G6100: signal is true;
	signal G6101: std_logic; attribute dont_touch of G6101: signal is true;
	signal G6102: std_logic; attribute dont_touch of G6102: signal is true;
	signal G6103: std_logic; attribute dont_touch of G6103: signal is true;
	signal G6104: std_logic; attribute dont_touch of G6104: signal is true;
	signal G6115: std_logic; attribute dont_touch of G6115: signal is true;
	signal G6116: std_logic; attribute dont_touch of G6116: signal is true;
	signal G6117: std_logic; attribute dont_touch of G6117: signal is true;
	signal G6118: std_logic; attribute dont_touch of G6118: signal is true;
	signal G6119: std_logic; attribute dont_touch of G6119: signal is true;
	signal G6130: std_logic; attribute dont_touch of G6130: signal is true;
	signal G6131: std_logic; attribute dont_touch of G6131: signal is true;
	signal G6134: std_logic; attribute dont_touch of G6134: signal is true;
	signal G6135: std_logic; attribute dont_touch of G6135: signal is true;
	signal G6136: std_logic; attribute dont_touch of G6136: signal is true;
	signal G6139: std_logic; attribute dont_touch of G6139: signal is true;
	signal G6140: std_logic; attribute dont_touch of G6140: signal is true;
	signal G6141: std_logic; attribute dont_touch of G6141: signal is true;
	signal G6142: std_logic; attribute dont_touch of G6142: signal is true;
	signal G6145: std_logic; attribute dont_touch of G6145: signal is true;
	signal G6146: std_logic; attribute dont_touch of G6146: signal is true;
	signal G6149: std_logic; attribute dont_touch of G6149: signal is true;
	signal G6153: std_logic; attribute dont_touch of G6153: signal is true;
	signal G6156: std_logic; attribute dont_touch of G6156: signal is true;
	signal G6157: std_logic; attribute dont_touch of G6157: signal is true;
	signal G6161: std_logic; attribute dont_touch of G6161: signal is true;
	signal G6162: std_logic; attribute dont_touch of G6162: signal is true;
	signal G6163: std_logic; attribute dont_touch of G6163: signal is true;
	signal G6166: std_logic; attribute dont_touch of G6166: signal is true;
	signal G6167: std_logic; attribute dont_touch of G6167: signal is true;
	signal G6170: std_logic; attribute dont_touch of G6170: signal is true;
	signal G6173: std_logic; attribute dont_touch of G6173: signal is true;
	signal G6177: std_logic; attribute dont_touch of G6177: signal is true;
	signal G6180: std_logic; attribute dont_touch of G6180: signal is true;
	signal G6183: std_logic; attribute dont_touch of G6183: signal is true;
	signal G6184: std_logic; attribute dont_touch of G6184: signal is true;
	signal G6188: std_logic; attribute dont_touch of G6188: signal is true;
	signal G6189: std_logic; attribute dont_touch of G6189: signal is true;
	signal G6190: std_logic; attribute dont_touch of G6190: signal is true;
	signal G6193: std_logic; attribute dont_touch of G6193: signal is true;
	signal G6194: std_logic; attribute dont_touch of G6194: signal is true;
	signal G6197: std_logic; attribute dont_touch of G6197: signal is true;
	signal G6200: std_logic; attribute dont_touch of G6200: signal is true;
	signal G6201: std_logic; attribute dont_touch of G6201: signal is true;
	signal G6204: std_logic; attribute dont_touch of G6204: signal is true;
	signal G6205: std_logic; attribute dont_touch of G6205: signal is true;
	signal G6209: std_logic; attribute dont_touch of G6209: signal is true;
	signal G6212: std_logic; attribute dont_touch of G6212: signal is true;
	signal G6215: std_logic; attribute dont_touch of G6215: signal is true;
	signal G6216: std_logic; attribute dont_touch of G6216: signal is true;
	signal G6220: std_logic; attribute dont_touch of G6220: signal is true;
	signal G6221: std_logic; attribute dont_touch of G6221: signal is true;
	signal G6222: std_logic; attribute dont_touch of G6222: signal is true;
	signal G6226: std_logic; attribute dont_touch of G6226: signal is true;
	signal G6227: std_logic; attribute dont_touch of G6227: signal is true;
	signal G6230: std_logic; attribute dont_touch of G6230: signal is true;
	signal G6232: std_logic; attribute dont_touch of G6232: signal is true;
	signal G6281: std_logic; attribute dont_touch of G6281: signal is true;
	signal G6284: std_logic; attribute dont_touch of G6284: signal is true;
	signal G6288: std_logic; attribute dont_touch of G6288: signal is true;
	signal G6289: std_logic; attribute dont_touch of G6289: signal is true;
	signal G6290: std_logic; attribute dont_touch of G6290: signal is true;
	signal G6293: std_logic; attribute dont_touch of G6293: signal is true;
	signal G6294: std_logic; attribute dont_touch of G6294: signal is true;
	signal G6298: std_logic; attribute dont_touch of G6298: signal is true;
	signal G6301: std_logic; attribute dont_touch of G6301: signal is true;
	signal G6304: std_logic; attribute dont_touch of G6304: signal is true;
	signal G6305: std_logic; attribute dont_touch of G6305: signal is true;
	signal G6309: std_logic; attribute dont_touch of G6309: signal is true;
	signal G6310: std_logic; attribute dont_touch of G6310: signal is true;
	signal G6314: std_logic; attribute dont_touch of G6314: signal is true;
	signal G6363: std_logic; attribute dont_touch of G6363: signal is true;
	signal G6367: std_logic; attribute dont_touch of G6367: signal is true;
	signal G6369: std_logic; attribute dont_touch of G6369: signal is true;
	signal G6418: std_logic; attribute dont_touch of G6418: signal is true;
	signal G6421: std_logic; attribute dont_touch of G6421: signal is true;
	signal G6425: std_logic; attribute dont_touch of G6425: signal is true;
	signal G6426: std_logic; attribute dont_touch of G6426: signal is true;
	signal G6427: std_logic; attribute dont_touch of G6427: signal is true;
	signal G6430: std_logic; attribute dont_touch of G6430: signal is true;
	signal G6431: std_logic; attribute dont_touch of G6431: signal is true;
	signal G6435: std_logic; attribute dont_touch of G6435: signal is true;
	signal G6438: std_logic; attribute dont_touch of G6438: signal is true;
	signal G6441: std_logic; attribute dont_touch of G6441: signal is true;
	signal G6443: std_logic; attribute dont_touch of G6443: signal is true;
	signal G6444: std_logic; attribute dont_touch of G6444: signal is true;
	signal G6448: std_logic; attribute dont_touch of G6448: signal is true;
	signal G6486: std_logic; attribute dont_touch of G6486: signal is true;
	signal G6512: std_logic; attribute dont_touch of G6512: signal is true;
	signal G6513: std_logic; attribute dont_touch of G6513: signal is true;
	signal G6517: std_logic; attribute dont_touch of G6517: signal is true;
	signal G6519: std_logic; attribute dont_touch of G6519: signal is true;
	signal G6568: std_logic; attribute dont_touch of G6568: signal is true;
	signal G6572: std_logic; attribute dont_touch of G6572: signal is true;
	signal G6574: std_logic; attribute dont_touch of G6574: signal is true;
	signal G6623: std_logic; attribute dont_touch of G6623: signal is true;
	signal G6626: std_logic; attribute dont_touch of G6626: signal is true;
	signal G6630: std_logic; attribute dont_touch of G6630: signal is true;
	signal G6631: std_logic; attribute dont_touch of G6631: signal is true;
	signal G6632: std_logic; attribute dont_touch of G6632: signal is true;
	signal G6635: std_logic; attribute dont_touch of G6635: signal is true;
	signal G6636: std_logic; attribute dont_touch of G6636: signal is true;
	signal G6637: std_logic; attribute dont_touch of G6637: signal is true;
	signal G6638: std_logic; attribute dont_touch of G6638: signal is true;
	signal G6641: std_logic; attribute dont_touch of G6641: signal is true;
	signal G6643: std_logic; attribute dont_touch of G6643: signal is true;
	signal G6672: std_logic; attribute dont_touch of G6672: signal is true;
	signal G6675: std_logic; attribute dont_touch of G6675: signal is true;
	signal G6676: std_logic; attribute dont_touch of G6676: signal is true;
	signal G6678: std_logic; attribute dont_touch of G6678: signal is true;
	signal G6707: std_logic; attribute dont_touch of G6707: signal is true;
	signal G6711: std_logic; attribute dont_touch of G6711: signal is true;
	signal G6713: std_logic; attribute dont_touch of G6713: signal is true;
	signal G6751: std_logic; attribute dont_touch of G6751: signal is true;
	signal G6776: std_logic; attribute dont_touch of G6776: signal is true;
	signal G6777: std_logic; attribute dont_touch of G6777: signal is true;
	signal G6781: std_logic; attribute dont_touch of G6781: signal is true;
	signal G6783: std_logic; attribute dont_touch of G6783: signal is true;
	signal G6832: std_logic; attribute dont_touch of G6832: signal is true;
	signal G6836: std_logic; attribute dont_touch of G6836: signal is true;
	signal G6838: std_logic; attribute dont_touch of G6838: signal is true;
	signal G6887: std_logic; attribute dont_touch of G6887: signal is true;
	signal G6890: std_logic; attribute dont_touch of G6890: signal is true;
	signal G6894: std_logic; attribute dont_touch of G6894: signal is true;
	signal G6896: std_logic; attribute dont_touch of G6896: signal is true;
	signal G6897: std_logic; attribute dont_touch of G6897: signal is true;
	signal G6898: std_logic; attribute dont_touch of G6898: signal is true;
	signal G6901: std_logic; attribute dont_touch of G6901: signal is true;
	signal G6905: std_logic; attribute dont_touch of G6905: signal is true;
	signal G6908: std_logic; attribute dont_touch of G6908: signal is true;
	signal G6912: std_logic; attribute dont_touch of G6912: signal is true;
	signal G6942: std_logic; attribute dont_touch of G6942: signal is true;
	signal G6943: std_logic; attribute dont_touch of G6943: signal is true;
	signal G6945: std_logic; attribute dont_touch of G6945: signal is true;
	signal G6974: std_logic; attribute dont_touch of G6974: signal is true;
	signal G6977: std_logic; attribute dont_touch of G6977: signal is true;
	signal G6978: std_logic; attribute dont_touch of G6978: signal is true;
	signal G6980: std_logic; attribute dont_touch of G6980: signal is true;
	signal G7009: std_logic; attribute dont_touch of G7009: signal is true;
	signal G7013: std_logic; attribute dont_touch of G7013: signal is true;
	signal G7015: std_logic; attribute dont_touch of G7015: signal is true;
	signal G7053: std_logic; attribute dont_touch of G7053: signal is true;
	signal G7078: std_logic; attribute dont_touch of G7078: signal is true;
	signal G7079: std_logic; attribute dont_touch of G7079: signal is true;
	signal G7083: std_logic; attribute dont_touch of G7083: signal is true;
	signal G7085: std_logic; attribute dont_touch of G7085: signal is true;
	signal G7134: std_logic; attribute dont_touch of G7134: signal is true;
	signal G7138: std_logic; attribute dont_touch of G7138: signal is true;
	signal G7139: std_logic; attribute dont_touch of G7139: signal is true;
	signal G7140: std_logic; attribute dont_touch of G7140: signal is true;
	signal G7141: std_logic; attribute dont_touch of G7141: signal is true;
	signal G7142: std_logic; attribute dont_touch of G7142: signal is true;
	signal G7143: std_logic; attribute dont_touch of G7143: signal is true;
	signal G7146: std_logic; attribute dont_touch of G7146: signal is true;
	signal G7149: std_logic; attribute dont_touch of G7149: signal is true;
	signal G7152: std_logic; attribute dont_touch of G7152: signal is true;
	signal G7153: std_logic; attribute dont_touch of G7153: signal is true;
	signal G7156: std_logic; attribute dont_touch of G7156: signal is true;
	signal G7157: std_logic; attribute dont_touch of G7157: signal is true;
	signal G7158: std_logic; attribute dont_touch of G7158: signal is true;
	signal G7162: std_logic; attribute dont_touch of G7162: signal is true;
	signal G7192: std_logic; attribute dont_touch of G7192: signal is true;
	signal G7193: std_logic; attribute dont_touch of G7193: signal is true;
	signal G7195: std_logic; attribute dont_touch of G7195: signal is true;
	signal G7224: std_logic; attribute dont_touch of G7224: signal is true;
	signal G7227: std_logic; attribute dont_touch of G7227: signal is true;
	signal G7228: std_logic; attribute dont_touch of G7228: signal is true;
	signal G7230: std_logic; attribute dont_touch of G7230: signal is true;
	signal G7259: std_logic; attribute dont_touch of G7259: signal is true;
	signal G7263: std_logic; attribute dont_touch of G7263: signal is true;
	signal G7265: std_logic; attribute dont_touch of G7265: signal is true;
	signal G7303: std_logic; attribute dont_touch of G7303: signal is true;
	signal G7328: std_logic; attribute dont_touch of G7328: signal is true;
	signal G7329: std_logic; attribute dont_touch of G7329: signal is true;
	signal G7333: std_logic; attribute dont_touch of G7333: signal is true;
	signal G7335: std_logic; attribute dont_touch of G7335: signal is true;
	signal G7336: std_logic; attribute dont_touch of G7336: signal is true;
	signal G7337: std_logic; attribute dont_touch of G7337: signal is true;
	signal G7338: std_logic; attribute dont_touch of G7338: signal is true;
	signal G7342: std_logic; attribute dont_touch of G7342: signal is true;
	signal G7345: std_logic; attribute dont_touch of G7345: signal is true;
	signal G7346: std_logic; attribute dont_touch of G7346: signal is true;
	signal G7347: std_logic; attribute dont_touch of G7347: signal is true;
	signal G7348: std_logic; attribute dont_touch of G7348: signal is true;
	signal G7349: std_logic; attribute dont_touch of G7349: signal is true;
	signal G7352: std_logic; attribute dont_touch of G7352: signal is true;
	signal G7353: std_logic; attribute dont_touch of G7353: signal is true;
	signal G7354: std_logic; attribute dont_touch of G7354: signal is true;
	signal G7358: std_logic; attribute dont_touch of G7358: signal is true;
	signal G7388: std_logic; attribute dont_touch of G7388: signal is true;
	signal G7389: std_logic; attribute dont_touch of G7389: signal is true;
	signal G7391: std_logic; attribute dont_touch of G7391: signal is true;
	signal G7420: std_logic; attribute dont_touch of G7420: signal is true;
	signal G7423: std_logic; attribute dont_touch of G7423: signal is true;
	signal G7424: std_logic; attribute dont_touch of G7424: signal is true;
	signal G7426: std_logic; attribute dont_touch of G7426: signal is true;
	signal G7455: std_logic; attribute dont_touch of G7455: signal is true;
	signal G7459: std_logic; attribute dont_touch of G7459: signal is true;
	signal G7460: std_logic; attribute dont_touch of G7460: signal is true;
	signal G7461: std_logic; attribute dont_touch of G7461: signal is true;
	signal G7462: std_logic; attribute dont_touch of G7462: signal is true;
	signal G7465: std_logic; attribute dont_touch of G7465: signal is true;
	signal G7466: std_logic; attribute dont_touch of G7466: signal is true;
	signal G7471: std_logic; attribute dont_touch of G7471: signal is true;
	signal G7475: std_logic; attribute dont_touch of G7475: signal is true;
	signal G7476: std_logic; attribute dont_touch of G7476: signal is true;
	signal G7477: std_logic; attribute dont_touch of G7477: signal is true;
	signal G7478: std_logic; attribute dont_touch of G7478: signal is true;
	signal G7479: std_logic; attribute dont_touch of G7479: signal is true;
	signal G7482: std_logic; attribute dont_touch of G7482: signal is true;
	signal G7483: std_logic; attribute dont_touch of G7483: signal is true;
	signal G7484: std_logic; attribute dont_touch of G7484: signal is true;
	signal G7488: std_logic; attribute dont_touch of G7488: signal is true;
	signal G7518: std_logic; attribute dont_touch of G7518: signal is true;
	signal G7520: std_logic; attribute dont_touch of G7520: signal is true;
	signal G7521: std_logic; attribute dont_touch of G7521: signal is true;
	signal G7522: std_logic; attribute dont_touch of G7522: signal is true;
	signal G7527: std_logic; attribute dont_touch of G7527: signal is true;
	signal G7528: std_logic; attribute dont_touch of G7528: signal is true;
	signal G7529: std_logic; attribute dont_touch of G7529: signal is true;
	signal G7530: std_logic; attribute dont_touch of G7530: signal is true;
	signal G7531: std_logic; attribute dont_touch of G7531: signal is true;
	signal G7532: std_logic; attribute dont_touch of G7532: signal is true;
	signal G7533: std_logic; attribute dont_touch of G7533: signal is true;
	signal G7534: std_logic; attribute dont_touch of G7534: signal is true;
	signal G7535: std_logic; attribute dont_touch of G7535: signal is true;
	signal G7538: std_logic; attribute dont_touch of G7538: signal is true;
	signal G7539: std_logic; attribute dont_touch of G7539: signal is true;
	signal G7540: std_logic; attribute dont_touch of G7540: signal is true;
	signal G7541: std_logic; attribute dont_touch of G7541: signal is true;
	signal G7542: std_logic; attribute dont_touch of G7542: signal is true;
	signal G7545: std_logic; attribute dont_touch of G7545: signal is true;
	signal G7548: std_logic; attribute dont_touch of G7548: signal is true;
	signal G7549: std_logic; attribute dont_touch of G7549: signal is true;
	signal G7553: std_logic; attribute dont_touch of G7553: signal is true;
	signal G7554: std_logic; attribute dont_touch of G7554: signal is true;
	signal G7555: std_logic; attribute dont_touch of G7555: signal is true;
	signal G7556: std_logic; attribute dont_touch of G7556: signal is true;
	signal G7557: std_logic; attribute dont_touch of G7557: signal is true;
	signal G7558: std_logic; attribute dont_touch of G7558: signal is true;
	signal G7559: std_logic; attribute dont_touch of G7559: signal is true;
	signal G7560: std_logic; attribute dont_touch of G7560: signal is true;
	signal G7561: std_logic; attribute dont_touch of G7561: signal is true;
	signal G7562: std_logic; attribute dont_touch of G7562: signal is true;
	signal G7566: std_logic; attribute dont_touch of G7566: signal is true;
	signal G7570: std_logic; attribute dont_touch of G7570: signal is true;
	signal G7573: std_logic; attribute dont_touch of G7573: signal is true;
	signal G7574: std_logic; attribute dont_touch of G7574: signal is true;
	signal G7575: std_logic; attribute dont_touch of G7575: signal is true;
	signal G7576: std_logic; attribute dont_touch of G7576: signal is true;
	signal G7577: std_logic; attribute dont_touch of G7577: signal is true;
	signal G7578: std_logic; attribute dont_touch of G7578: signal is true;
	signal G7579: std_logic; attribute dont_touch of G7579: signal is true;
	signal G7580: std_logic; attribute dont_touch of G7580: signal is true;
	signal G7581: std_logic; attribute dont_touch of G7581: signal is true;
	signal G7582: std_logic; attribute dont_touch of G7582: signal is true;
	signal G7583: std_logic; attribute dont_touch of G7583: signal is true;
	signal G7587: std_logic; attribute dont_touch of G7587: signal is true;
	signal G7590: std_logic; attribute dont_touch of G7590: signal is true;
	signal G7591: std_logic; attribute dont_touch of G7591: signal is true;
	signal G7592: std_logic; attribute dont_touch of G7592: signal is true;
	signal G7593: std_logic; attribute dont_touch of G7593: signal is true;
	signal G7594: std_logic; attribute dont_touch of G7594: signal is true;
	signal G7595: std_logic; attribute dont_touch of G7595: signal is true;
	signal G7600: std_logic; attribute dont_touch of G7600: signal is true;
	signal G7603: std_logic; attribute dont_touch of G7603: signal is true;
	signal G7604: std_logic; attribute dont_touch of G7604: signal is true;
	signal G7605: std_logic; attribute dont_touch of G7605: signal is true;
	signal G7606: std_logic; attribute dont_touch of G7606: signal is true;
	signal G7607: std_logic; attribute dont_touch of G7607: signal is true;
	signal G7610: std_logic; attribute dont_touch of G7610: signal is true;
	signal G7613: std_logic; attribute dont_touch of G7613: signal is true;
	signal G7614: std_logic; attribute dont_touch of G7614: signal is true;
	signal G7615: std_logic; attribute dont_touch of G7615: signal is true;
	signal G7616: std_logic; attribute dont_touch of G7616: signal is true;
	signal G7619: std_logic; attribute dont_touch of G7619: signal is true;
	signal G7622: std_logic; attribute dont_touch of G7622: signal is true;
	signal G7623: std_logic; attribute dont_touch of G7623: signal is true;
	signal G7626: std_logic; attribute dont_touch of G7626: signal is true;
	signal G7629: std_logic; attribute dont_touch of G7629: signal is true;
	signal G7632: std_logic; attribute dont_touch of G7632: signal is true;
	signal G7635: std_logic; attribute dont_touch of G7635: signal is true;
	signal G7638: std_logic; attribute dont_touch of G7638: signal is true;
	signal G7639: std_logic; attribute dont_touch of G7639: signal is true;
	signal G7642: std_logic; attribute dont_touch of G7642: signal is true;
	signal G7643: std_logic; attribute dont_touch of G7643: signal is true;
	signal G7646: std_logic; attribute dont_touch of G7646: signal is true;
	signal G7649: std_logic; attribute dont_touch of G7649: signal is true;
	signal G7652: std_logic; attribute dont_touch of G7652: signal is true;
	signal G7655: std_logic; attribute dont_touch of G7655: signal is true;
	signal G7658: std_logic; attribute dont_touch of G7658: signal is true;
	signal G7661: std_logic; attribute dont_touch of G7661: signal is true;
	signal G7664: std_logic; attribute dont_touch of G7664: signal is true;
	signal G7667: std_logic; attribute dont_touch of G7667: signal is true;
	signal G7670: std_logic; attribute dont_touch of G7670: signal is true;
	signal G7673: std_logic; attribute dont_touch of G7673: signal is true;
	signal G7676: std_logic; attribute dont_touch of G7676: signal is true;
	signal G7679: std_logic; attribute dont_touch of G7679: signal is true;
	signal G7682: std_logic; attribute dont_touch of G7682: signal is true;
	signal G7685: std_logic; attribute dont_touch of G7685: signal is true;
	signal G7688: std_logic; attribute dont_touch of G7688: signal is true;
	signal G7691: std_logic; attribute dont_touch of G7691: signal is true;
	signal G7694: std_logic; attribute dont_touch of G7694: signal is true;
	signal G7697: std_logic; attribute dont_touch of G7697: signal is true;
	signal G7700: std_logic; attribute dont_touch of G7700: signal is true;
	signal G7703: std_logic; attribute dont_touch of G7703: signal is true;
	signal G7706: std_logic; attribute dont_touch of G7706: signal is true;
	signal G7709: std_logic; attribute dont_touch of G7709: signal is true;
	signal G7712: std_logic; attribute dont_touch of G7712: signal is true;
	signal G7715: std_logic; attribute dont_touch of G7715: signal is true;
	signal G7718: std_logic; attribute dont_touch of G7718: signal is true;
	signal G7721: std_logic; attribute dont_touch of G7721: signal is true;
	signal G7724: std_logic; attribute dont_touch of G7724: signal is true;
	signal G7727: std_logic; attribute dont_touch of G7727: signal is true;
	signal G7730: std_logic; attribute dont_touch of G7730: signal is true;
	signal G7733: std_logic; attribute dont_touch of G7733: signal is true;
	signal G7736: std_logic; attribute dont_touch of G7736: signal is true;
	signal G7739: std_logic; attribute dont_touch of G7739: signal is true;
	signal G7742: std_logic; attribute dont_touch of G7742: signal is true;
	signal G7745: std_logic; attribute dont_touch of G7745: signal is true;
	signal G7748: std_logic; attribute dont_touch of G7748: signal is true;
	signal G7751: std_logic; attribute dont_touch of G7751: signal is true;
	signal G7754: std_logic; attribute dont_touch of G7754: signal is true;
	signal G7757: std_logic; attribute dont_touch of G7757: signal is true;
	signal G7760: std_logic; attribute dont_touch of G7760: signal is true;
	signal G7763: std_logic; attribute dont_touch of G7763: signal is true;
	signal G7766: std_logic; attribute dont_touch of G7766: signal is true;
	signal G7769: std_logic; attribute dont_touch of G7769: signal is true;
	signal G7772: std_logic; attribute dont_touch of G7772: signal is true;
	signal G7776: std_logic; attribute dont_touch of G7776: signal is true;
	signal G7779: std_logic; attribute dont_touch of G7779: signal is true;
	signal G7782: std_logic; attribute dont_touch of G7782: signal is true;
	signal G7785: std_logic; attribute dont_touch of G7785: signal is true;
	signal G7788: std_logic; attribute dont_touch of G7788: signal is true;
	signal G7792: std_logic; attribute dont_touch of G7792: signal is true;
	signal G7795: std_logic; attribute dont_touch of G7795: signal is true;
	signal G7796: std_logic; attribute dont_touch of G7796: signal is true;
	signal G7799: std_logic; attribute dont_touch of G7799: signal is true;
	signal G7802: std_logic; attribute dont_touch of G7802: signal is true;
	signal G7806: std_logic; attribute dont_touch of G7806: signal is true;
	signal G7809: std_logic; attribute dont_touch of G7809: signal is true;
	signal G7812: std_logic; attribute dont_touch of G7812: signal is true;
	signal G7815: std_logic; attribute dont_touch of G7815: signal is true;
	signal G7819: std_logic; attribute dont_touch of G7819: signal is true;
	signal G7822: std_logic; attribute dont_touch of G7822: signal is true;
	signal G7823: std_logic; attribute dont_touch of G7823: signal is true;
	signal G7826: std_logic; attribute dont_touch of G7826: signal is true;
	signal G7827: std_logic; attribute dont_touch of G7827: signal is true;
	signal G7830: std_logic; attribute dont_touch of G7830: signal is true;
	signal G7833: std_logic; attribute dont_touch of G7833: signal is true;
	signal G7834: std_logic; attribute dont_touch of G7834: signal is true;
	signal G7837: std_logic; attribute dont_touch of G7837: signal is true;
	signal G7838: std_logic; attribute dont_touch of G7838: signal is true;
	signal G7841: std_logic; attribute dont_touch of G7841: signal is true;
	signal G7842: std_logic; attribute dont_touch of G7842: signal is true;
	signal G7845: std_logic; attribute dont_touch of G7845: signal is true;
	signal G7848: std_logic; attribute dont_touch of G7848: signal is true;
	signal G7849: std_logic; attribute dont_touch of G7849: signal is true;
	signal G7852: std_logic; attribute dont_touch of G7852: signal is true;
	signal G7855: std_logic; attribute dont_touch of G7855: signal is true;
	signal G7856: std_logic; attribute dont_touch of G7856: signal is true;
	signal G7857: std_logic; attribute dont_touch of G7857: signal is true;
	signal G7858: std_logic; attribute dont_touch of G7858: signal is true;
	signal G7861: std_logic; attribute dont_touch of G7861: signal is true;
	signal G7862: std_logic; attribute dont_touch of G7862: signal is true;
	signal G7865: std_logic; attribute dont_touch of G7865: signal is true;
	signal G7868: std_logic; attribute dont_touch of G7868: signal is true;
	signal G7869: std_logic; attribute dont_touch of G7869: signal is true;
	signal G7872: std_logic; attribute dont_touch of G7872: signal is true;
	signal G7875: std_logic; attribute dont_touch of G7875: signal is true;
	signal G7876: std_logic; attribute dont_touch of G7876: signal is true;
	signal G7877: std_logic; attribute dont_touch of G7877: signal is true;
	signal G7878: std_logic; attribute dont_touch of G7878: signal is true;
	signal G7879: std_logic; attribute dont_touch of G7879: signal is true;
	signal G7880: std_logic; attribute dont_touch of G7880: signal is true;
	signal G7888: std_logic; attribute dont_touch of G7888: signal is true;
	signal G7891: std_logic; attribute dont_touch of G7891: signal is true;
	signal G7892: std_logic; attribute dont_touch of G7892: signal is true;
	signal G7895: std_logic; attribute dont_touch of G7895: signal is true;
	signal G7896: std_logic; attribute dont_touch of G7896: signal is true;
	signal G7897: std_logic; attribute dont_touch of G7897: signal is true;
	signal G7898: std_logic; attribute dont_touch of G7898: signal is true;
	signal G7899: std_logic; attribute dont_touch of G7899: signal is true;
	signal G7900: std_logic; attribute dont_touch of G7900: signal is true;
	signal G7901: std_logic; attribute dont_touch of G7901: signal is true;
	signal G7906: std_logic; attribute dont_touch of G7906: signal is true;
	signal G7910: std_logic; attribute dont_touch of G7910: signal is true;
	signal G7911: std_logic; attribute dont_touch of G7911: signal is true;
	signal G7912: std_logic; attribute dont_touch of G7912: signal is true;
	signal G7915: std_logic; attribute dont_touch of G7915: signal is true;
	signal G7916: std_logic; attribute dont_touch of G7916: signal is true;
	signal G7919: std_logic; attribute dont_touch of G7919: signal is true;
	signal G7922: std_logic; attribute dont_touch of G7922: signal is true;
	signal G7923: std_logic; attribute dont_touch of G7923: signal is true;
	signal G7924: std_logic; attribute dont_touch of G7924: signal is true;
	signal G7925: std_logic; attribute dont_touch of G7925: signal is true;
	signal G7926: std_logic; attribute dont_touch of G7926: signal is true;
	signal G7927: std_logic; attribute dont_touch of G7927: signal is true;
	signal G7928: std_logic; attribute dont_touch of G7928: signal is true;
	signal G7936: std_logic; attribute dont_touch of G7936: signal is true;
	signal G7949: std_logic; attribute dont_touch of G7949: signal is true;
	signal G7950: std_logic; attribute dont_touch of G7950: signal is true;
	signal G7953: std_logic; attribute dont_touch of G7953: signal is true;
	signal G7957: std_logic; attribute dont_touch of G7957: signal is true;
	signal G7958: std_logic; attribute dont_touch of G7958: signal is true;
	signal G7962: std_logic; attribute dont_touch of G7962: signal is true;
	signal G7963: std_logic; attribute dont_touch of G7963: signal is true;
	signal G7964: std_logic; attribute dont_touch of G7964: signal is true;
	signal G7967: std_logic; attribute dont_touch of G7967: signal is true;
	signal G7970: std_logic; attribute dont_touch of G7970: signal is true;
	signal G7971: std_logic; attribute dont_touch of G7971: signal is true;
	signal G7972: std_logic; attribute dont_touch of G7972: signal is true;
	signal G7973: std_logic; attribute dont_touch of G7973: signal is true;
	signal G7974: std_logic; attribute dont_touch of G7974: signal is true;
	signal G7975: std_logic; attribute dont_touch of G7975: signal is true;
	signal G7976: std_logic; attribute dont_touch of G7976: signal is true;
	signal G7989: std_logic; attribute dont_touch of G7989: signal is true;
	signal G7990: std_logic; attribute dont_touch of G7990: signal is true;
	signal G7993: std_logic; attribute dont_touch of G7993: signal is true;
	signal G7996: std_logic; attribute dont_touch of G7996: signal is true;
	signal G7999: std_logic; attribute dont_touch of G7999: signal is true;
	signal G8000: std_logic; attribute dont_touch of G8000: signal is true;
	signal G8001: std_logic; attribute dont_touch of G8001: signal is true;
	signal G8004: std_logic; attribute dont_touch of G8004: signal is true;
	signal G8008: std_logic; attribute dont_touch of G8008: signal is true;
	signal G8009: std_logic; attribute dont_touch of G8009: signal is true;
	signal G8013: std_logic; attribute dont_touch of G8013: signal is true;
	signal G8014: std_logic; attribute dont_touch of G8014: signal is true;
	signal G8015: std_logic; attribute dont_touch of G8015: signal is true;
	signal G8018: std_logic; attribute dont_touch of G8018: signal is true;
	signal G8022: std_logic; attribute dont_touch of G8022: signal is true;
	signal G8024: std_logic; attribute dont_touch of G8024: signal is true;
	signal G8025: std_logic; attribute dont_touch of G8025: signal is true;
	signal G8026: std_logic; attribute dont_touch of G8026: signal is true;
	signal G8027: std_logic; attribute dont_touch of G8027: signal is true;
	signal G8028: std_logic; attribute dont_touch of G8028: signal is true;
	signal G8029: std_logic; attribute dont_touch of G8029: signal is true;
	signal G8031: std_logic; attribute dont_touch of G8031: signal is true;
	signal G8044: std_logic; attribute dont_touch of G8044: signal is true;
	signal G8045: std_logic; attribute dont_touch of G8045: signal is true;
	signal G8053: std_logic; attribute dont_touch of G8053: signal is true;
	signal G8056: std_logic; attribute dont_touch of G8056: signal is true;
	signal G8059: std_logic; attribute dont_touch of G8059: signal is true;
	signal G8062: std_logic; attribute dont_touch of G8062: signal is true;
	signal G8065: std_logic; attribute dont_touch of G8065: signal is true;
	signal G8068: std_logic; attribute dont_touch of G8068: signal is true;
	signal G8071: std_logic; attribute dont_touch of G8071: signal is true;
	signal G8074: std_logic; attribute dont_touch of G8074: signal is true;
	signal G8075: std_logic; attribute dont_touch of G8075: signal is true;
	signal G8076: std_logic; attribute dont_touch of G8076: signal is true;
	signal G8079: std_logic; attribute dont_touch of G8079: signal is true;
	signal G8083: std_logic; attribute dont_touch of G8083: signal is true;
	signal G8084: std_logic; attribute dont_touch of G8084: signal is true;
	signal G8088: std_logic; attribute dont_touch of G8088: signal is true;
	signal G8089: std_logic; attribute dont_touch of G8089: signal is true;
	signal G8090: std_logic; attribute dont_touch of G8090: signal is true;
	signal G8093: std_logic; attribute dont_touch of G8093: signal is true;
	signal G8097: std_logic; attribute dont_touch of G8097: signal is true;
	signal G8098: std_logic; attribute dont_touch of G8098: signal is true;
	signal G8099: std_logic; attribute dont_touch of G8099: signal is true;
	signal G8100: std_logic; attribute dont_touch of G8100: signal is true;
	signal G8101: std_logic; attribute dont_touch of G8101: signal is true;
	signal G8102: std_logic; attribute dont_touch of G8102: signal is true;
	signal G8103: std_logic; attribute dont_touch of G8103: signal is true;
	signal G8107: std_logic; attribute dont_touch of G8107: signal is true;
	signal G8120: std_logic; attribute dont_touch of G8120: signal is true;
	signal G8123: std_logic; attribute dont_touch of G8123: signal is true;
	signal G8126: std_logic; attribute dont_touch of G8126: signal is true;
	signal G8129: std_logic; attribute dont_touch of G8129: signal is true;
	signal G8132: std_logic; attribute dont_touch of G8132: signal is true;
	signal G8135: std_logic; attribute dont_touch of G8135: signal is true;
	signal G8138: std_logic; attribute dont_touch of G8138: signal is true;
	signal G8141: std_logic; attribute dont_touch of G8141: signal is true;
	signal G8144: std_logic; attribute dont_touch of G8144: signal is true;
	signal G8147: std_logic; attribute dont_touch of G8147: signal is true;
	signal G8150: std_logic; attribute dont_touch of G8150: signal is true;
	signal G8153: std_logic; attribute dont_touch of G8153: signal is true;
	signal G8156: std_logic; attribute dont_touch of G8156: signal is true;
	signal G8159: std_logic; attribute dont_touch of G8159: signal is true;
	signal G8160: std_logic; attribute dont_touch of G8160: signal is true;
	signal G8161: std_logic; attribute dont_touch of G8161: signal is true;
	signal G8164: std_logic; attribute dont_touch of G8164: signal is true;
	signal G8168: std_logic; attribute dont_touch of G8168: signal is true;
	signal G8169: std_logic; attribute dont_touch of G8169: signal is true;
	signal G8172: std_logic; attribute dont_touch of G8172: signal is true;
	signal G8176: std_logic; attribute dont_touch of G8176: signal is true;
	signal G8177: std_logic; attribute dont_touch of G8177: signal is true;
	signal G8178: std_logic; attribute dont_touch of G8178: signal is true;
	signal G8179: std_logic; attribute dont_touch of G8179: signal is true;
	signal G8180: std_logic; attribute dont_touch of G8180: signal is true;
	signal G8181: std_logic; attribute dont_touch of G8181: signal is true;
	signal G8182: std_logic; attribute dont_touch of G8182: signal is true;
	signal G8183: std_logic; attribute dont_touch of G8183: signal is true;
	signal G8191: std_logic; attribute dont_touch of G8191: signal is true;
	signal G8194: std_logic; attribute dont_touch of G8194: signal is true;
	signal G8197: std_logic; attribute dont_touch of G8197: signal is true;
	signal G8200: std_logic; attribute dont_touch of G8200: signal is true;
	signal G8203: std_logic; attribute dont_touch of G8203: signal is true;
	signal G8206: std_logic; attribute dont_touch of G8206: signal is true;
	signal G8209: std_logic; attribute dont_touch of G8209: signal is true;
	signal G8212: std_logic; attribute dont_touch of G8212: signal is true;
	signal G8215: std_logic; attribute dont_touch of G8215: signal is true;
	signal G8218: std_logic; attribute dont_touch of G8218: signal is true;
	signal G8221: std_logic; attribute dont_touch of G8221: signal is true;
	signal G8224: std_logic; attribute dont_touch of G8224: signal is true;
	signal G8227: std_logic; attribute dont_touch of G8227: signal is true;
	signal G8230: std_logic; attribute dont_touch of G8230: signal is true;
	signal G8233: std_logic; attribute dont_touch of G8233: signal is true;
	signal G8236: std_logic; attribute dont_touch of G8236: signal is true;
	signal G8239: std_logic; attribute dont_touch of G8239: signal is true;
	signal G8242: std_logic; attribute dont_touch of G8242: signal is true;
	signal G8245: std_logic; attribute dont_touch of G8245: signal is true;
	signal G8246: std_logic; attribute dont_touch of G8246: signal is true;
	signal G8250: std_logic; attribute dont_touch of G8250: signal is true;
	signal G8252: std_logic; attribute dont_touch of G8252: signal is true;
	signal G8253: std_logic; attribute dont_touch of G8253: signal is true;
	signal G8254: std_logic; attribute dont_touch of G8254: signal is true;
	signal G8255: std_logic; attribute dont_touch of G8255: signal is true;
	signal G8256: std_logic; attribute dont_touch of G8256: signal is true;
	signal G8257: std_logic; attribute dont_touch of G8257: signal is true;
	signal G8276: std_logic; attribute dont_touch of G8276: signal is true;
	signal G8277: std_logic; attribute dont_touch of G8277: signal is true;
	signal G8278: std_logic; attribute dont_touch of G8278: signal is true;
	signal G8284: std_logic; attribute dont_touch of G8284: signal is true;
	signal G8285: std_logic; attribute dont_touch of G8285: signal is true;
	signal G8286: std_logic; attribute dont_touch of G8286: signal is true;
	signal G8287: std_logic; attribute dont_touch of G8287: signal is true;
	signal G8293: std_logic; attribute dont_touch of G8293: signal is true;
	signal G8294: std_logic; attribute dont_touch of G8294: signal is true;
	signal G8295: std_logic; attribute dont_touch of G8295: signal is true;
	signal G8296: std_logic; attribute dont_touch of G8296: signal is true;
	signal G8302: std_logic; attribute dont_touch of G8302: signal is true;
	signal G8303: std_logic; attribute dont_touch of G8303: signal is true;
	signal G8304: std_logic; attribute dont_touch of G8304: signal is true;
	signal G8305: std_logic; attribute dont_touch of G8305: signal is true;
	signal G8311: std_logic; attribute dont_touch of G8311: signal is true;
	signal G8312: std_logic; attribute dont_touch of G8312: signal is true;
	signal G8313: std_logic; attribute dont_touch of G8313: signal is true;
	signal G8317: std_logic; attribute dont_touch of G8317: signal is true;
	signal G8321: std_logic; attribute dont_touch of G8321: signal is true;
	signal G8324: std_logic; attribute dont_touch of G8324: signal is true;
	signal G8327: std_logic; attribute dont_touch of G8327: signal is true;
	signal G8328: std_logic; attribute dont_touch of G8328: signal is true;
	signal G8329: std_logic; attribute dont_touch of G8329: signal is true;
	signal G8330: std_logic; attribute dont_touch of G8330: signal is true;
	signal G8333: std_logic; attribute dont_touch of G8333: signal is true;
	signal G8336: std_logic; attribute dont_touch of G8336: signal is true;
	signal G8339: std_logic; attribute dont_touch of G8339: signal is true;
	signal G8340: std_logic; attribute dont_touch of G8340: signal is true;
	signal G8341: std_logic; attribute dont_touch of G8341: signal is true;
	signal G8344: std_logic; attribute dont_touch of G8344: signal is true;
	signal G8347: std_logic; attribute dont_touch of G8347: signal is true;
	signal G8350: std_logic; attribute dont_touch of G8350: signal is true;
	signal G8351: std_logic; attribute dont_touch of G8351: signal is true;
	signal G8354: std_logic; attribute dont_touch of G8354: signal is true;
	signal G8357: std_logic; attribute dont_touch of G8357: signal is true;
	signal G8360: std_logic; attribute dont_touch of G8360: signal is true;
	signal G8363: std_logic; attribute dont_touch of G8363: signal is true;
	signal G8366: std_logic; attribute dont_touch of G8366: signal is true;
	signal G8369: std_logic; attribute dont_touch of G8369: signal is true;
	signal G8372: std_logic; attribute dont_touch of G8372: signal is true;
	signal G8375: std_logic; attribute dont_touch of G8375: signal is true;
	signal G8378: std_logic; attribute dont_touch of G8378: signal is true;
	signal G8381: std_logic; attribute dont_touch of G8381: signal is true;
	signal G8382: std_logic; attribute dont_touch of G8382: signal is true;
	signal G8385: std_logic; attribute dont_touch of G8385: signal is true;
	signal G8386: std_logic; attribute dont_touch of G8386: signal is true;
	signal G8387: std_logic; attribute dont_touch of G8387: signal is true;
	signal G8388: std_logic; attribute dont_touch of G8388: signal is true;
	signal G8391: std_logic; attribute dont_touch of G8391: signal is true;
	signal G8394: std_logic; attribute dont_touch of G8394: signal is true;
	signal G8395: std_logic; attribute dont_touch of G8395: signal is true;
	signal G8396: std_logic; attribute dont_touch of G8396: signal is true;
	signal G8397: std_logic; attribute dont_touch of G8397: signal is true;
	signal G8400: std_logic; attribute dont_touch of G8400: signal is true;
	signal G8403: std_logic; attribute dont_touch of G8403: signal is true;
	signal G8406: std_logic; attribute dont_touch of G8406: signal is true;
	signal G8407: std_logic; attribute dont_touch of G8407: signal is true;
	signal G8408: std_logic; attribute dont_touch of G8408: signal is true;
	signal G8411: std_logic; attribute dont_touch of G8411: signal is true;
	signal G8414: std_logic; attribute dont_touch of G8414: signal is true;
	signal G8417: std_logic; attribute dont_touch of G8417: signal is true;
	signal G8418: std_logic; attribute dont_touch of G8418: signal is true;
	signal G8421: std_logic; attribute dont_touch of G8421: signal is true;
	signal G8424: std_logic; attribute dont_touch of G8424: signal is true;
	signal G8427: std_logic; attribute dont_touch of G8427: signal is true;
	signal G8430: std_logic; attribute dont_touch of G8430: signal is true;
	signal G8431: std_logic; attribute dont_touch of G8431: signal is true;
	signal G8432: std_logic; attribute dont_touch of G8432: signal is true;
	signal G8433: std_logic; attribute dont_touch of G8433: signal is true;
	signal G8434: std_logic; attribute dont_touch of G8434: signal is true;
	signal G8437: std_logic; attribute dont_touch of G8437: signal is true;
	signal G8438: std_logic; attribute dont_touch of G8438: signal is true;
	signal G8439: std_logic; attribute dont_touch of G8439: signal is true;
	signal G8440: std_logic; attribute dont_touch of G8440: signal is true;
	signal G8443: std_logic; attribute dont_touch of G8443: signal is true;
	signal G8446: std_logic; attribute dont_touch of G8446: signal is true;
	signal G8447: std_logic; attribute dont_touch of G8447: signal is true;
	signal G8448: std_logic; attribute dont_touch of G8448: signal is true;
	signal G8449: std_logic; attribute dont_touch of G8449: signal is true;
	signal G8452: std_logic; attribute dont_touch of G8452: signal is true;
	signal G8455: std_logic; attribute dont_touch of G8455: signal is true;
	signal G8458: std_logic; attribute dont_touch of G8458: signal is true;
	signal G8459: std_logic; attribute dont_touch of G8459: signal is true;
	signal G8460: std_logic; attribute dont_touch of G8460: signal is true;
	signal G8463: std_logic; attribute dont_touch of G8463: signal is true;
	signal G8464: std_logic; attribute dont_touch of G8464: signal is true;
	signal G8465: std_logic; attribute dont_touch of G8465: signal is true;
	signal G8466: std_logic; attribute dont_touch of G8466: signal is true;
	signal G8467: std_logic; attribute dont_touch of G8467: signal is true;
	signal G8468: std_logic; attribute dont_touch of G8468: signal is true;
	signal G8469: std_logic; attribute dont_touch of G8469: signal is true;
	signal G8472: std_logic; attribute dont_touch of G8472: signal is true;
	signal G8473: std_logic; attribute dont_touch of G8473: signal is true;
	signal G8474: std_logic; attribute dont_touch of G8474: signal is true;
	signal G8475: std_logic; attribute dont_touch of G8475: signal is true;
	signal G8478: std_logic; attribute dont_touch of G8478: signal is true;
	signal G8481: std_logic; attribute dont_touch of G8481: signal is true;
	signal G8482: std_logic; attribute dont_touch of G8482: signal is true;
	signal G8483: std_logic; attribute dont_touch of G8483: signal is true;
	signal G8484: std_logic; attribute dont_touch of G8484: signal is true;
	signal G8485: std_logic; attribute dont_touch of G8485: signal is true;
	signal G8486: std_logic; attribute dont_touch of G8486: signal is true;
	signal G8487: std_logic; attribute dont_touch of G8487: signal is true;
	signal G8488: std_logic; attribute dont_touch of G8488: signal is true;
	signal G8489: std_logic; attribute dont_touch of G8489: signal is true;
	signal G8490: std_logic; attribute dont_touch of G8490: signal is true;
	signal G8491: std_logic; attribute dont_touch of G8491: signal is true;
	signal G8492: std_logic; attribute dont_touch of G8492: signal is true;
	signal G8493: std_logic; attribute dont_touch of G8493: signal is true;
	signal G8494: std_logic; attribute dont_touch of G8494: signal is true;
	signal G8497: std_logic; attribute dont_touch of G8497: signal is true;
	signal G8498: std_logic; attribute dont_touch of G8498: signal is true;
	signal G8499: std_logic; attribute dont_touch of G8499: signal is true;
	signal G8500: std_logic; attribute dont_touch of G8500: signal is true;
	signal G8501: std_logic; attribute dont_touch of G8501: signal is true;
	signal G8502: std_logic; attribute dont_touch of G8502: signal is true;
	signal G8503: std_logic; attribute dont_touch of G8503: signal is true;
	signal G8504: std_logic; attribute dont_touch of G8504: signal is true;
	signal G8505: std_logic; attribute dont_touch of G8505: signal is true;
	signal G8506: std_logic; attribute dont_touch of G8506: signal is true;
	signal G8507: std_logic; attribute dont_touch of G8507: signal is true;
	signal G8508: std_logic; attribute dont_touch of G8508: signal is true;
	signal G8509: std_logic; attribute dont_touch of G8509: signal is true;
	signal G8510: std_logic; attribute dont_touch of G8510: signal is true;
	signal G8511: std_logic; attribute dont_touch of G8511: signal is true;
	signal G8512: std_logic; attribute dont_touch of G8512: signal is true;
	signal G8513: std_logic; attribute dont_touch of G8513: signal is true;
	signal G8514: std_logic; attribute dont_touch of G8514: signal is true;
	signal G8515: std_logic; attribute dont_touch of G8515: signal is true;
	signal G8516: std_logic; attribute dont_touch of G8516: signal is true;
	signal G8517: std_logic; attribute dont_touch of G8517: signal is true;
	signal G8518: std_logic; attribute dont_touch of G8518: signal is true;
	signal G8519: std_logic; attribute dont_touch of G8519: signal is true;
	signal G8520: std_logic; attribute dont_touch of G8520: signal is true;
	signal G8521: std_logic; attribute dont_touch of G8521: signal is true;
	signal G8522: std_logic; attribute dont_touch of G8522: signal is true;
	signal G8523: std_logic; attribute dont_touch of G8523: signal is true;
	signal G8524: std_logic; attribute dont_touch of G8524: signal is true;
	signal G8525: std_logic; attribute dont_touch of G8525: signal is true;
	signal G8526: std_logic; attribute dont_touch of G8526: signal is true;
	signal G8527: std_logic; attribute dont_touch of G8527: signal is true;
	signal G8528: std_logic; attribute dont_touch of G8528: signal is true;
	signal G8529: std_logic; attribute dont_touch of G8529: signal is true;
	signal G8530: std_logic; attribute dont_touch of G8530: signal is true;
	signal G8531: std_logic; attribute dont_touch of G8531: signal is true;
	signal G8532: std_logic; attribute dont_touch of G8532: signal is true;
	signal G8533: std_logic; attribute dont_touch of G8533: signal is true;
	signal G8534: std_logic; attribute dont_touch of G8534: signal is true;
	signal G8535: std_logic; attribute dont_touch of G8535: signal is true;
	signal G8536: std_logic; attribute dont_touch of G8536: signal is true;
	signal G8537: std_logic; attribute dont_touch of G8537: signal is true;
	signal G8538: std_logic; attribute dont_touch of G8538: signal is true;
	signal G8539: std_logic; attribute dont_touch of G8539: signal is true;
	signal G8540: std_logic; attribute dont_touch of G8540: signal is true;
	signal G8541: std_logic; attribute dont_touch of G8541: signal is true;
	signal G8542: std_logic; attribute dont_touch of G8542: signal is true;
	signal G8543: std_logic; attribute dont_touch of G8543: signal is true;
	signal G8544: std_logic; attribute dont_touch of G8544: signal is true;
	signal G8545: std_logic; attribute dont_touch of G8545: signal is true;
	signal G8546: std_logic; attribute dont_touch of G8546: signal is true;
	signal G8547: std_logic; attribute dont_touch of G8547: signal is true;
	signal G8548: std_logic; attribute dont_touch of G8548: signal is true;
	signal G8549: std_logic; attribute dont_touch of G8549: signal is true;
	signal G8550: std_logic; attribute dont_touch of G8550: signal is true;
	signal G8551: std_logic; attribute dont_touch of G8551: signal is true;
	signal G8552: std_logic; attribute dont_touch of G8552: signal is true;
	signal G8553: std_logic; attribute dont_touch of G8553: signal is true;
	signal G8554: std_logic; attribute dont_touch of G8554: signal is true;
	signal G8555: std_logic; attribute dont_touch of G8555: signal is true;
	signal G8556: std_logic; attribute dont_touch of G8556: signal is true;
	signal G8557: std_logic; attribute dont_touch of G8557: signal is true;
	signal G8558: std_logic; attribute dont_touch of G8558: signal is true;
	signal G8559: std_logic; attribute dont_touch of G8559: signal is true;
	signal G8560: std_logic; attribute dont_touch of G8560: signal is true;
	signal G8561: std_logic; attribute dont_touch of G8561: signal is true;
	signal G8562: std_logic; attribute dont_touch of G8562: signal is true;
	signal G8563: std_logic; attribute dont_touch of G8563: signal is true;
	signal G8564: std_logic; attribute dont_touch of G8564: signal is true;
	signal G8565: std_logic; attribute dont_touch of G8565: signal is true;
	signal G8566: std_logic; attribute dont_touch of G8566: signal is true;
	signal G8567: std_logic; attribute dont_touch of G8567: signal is true;
	signal G8568: std_logic; attribute dont_touch of G8568: signal is true;
	signal G8569: std_logic; attribute dont_touch of G8569: signal is true;
	signal G8570: std_logic; attribute dont_touch of G8570: signal is true;
	signal G8571: std_logic; attribute dont_touch of G8571: signal is true;
	signal G8572: std_logic; attribute dont_touch of G8572: signal is true;
	signal G8573: std_logic; attribute dont_touch of G8573: signal is true;
	signal G8574: std_logic; attribute dont_touch of G8574: signal is true;
	signal G8575: std_logic; attribute dont_touch of G8575: signal is true;
	signal G8576: std_logic; attribute dont_touch of G8576: signal is true;
	signal G8577: std_logic; attribute dont_touch of G8577: signal is true;
	signal G8578: std_logic; attribute dont_touch of G8578: signal is true;
	signal G8579: std_logic; attribute dont_touch of G8579: signal is true;
	signal G8580: std_logic; attribute dont_touch of G8580: signal is true;
	signal G8587: std_logic; attribute dont_touch of G8587: signal is true;
	signal G8594: std_logic; attribute dont_touch of G8594: signal is true;
	signal G8601: std_logic; attribute dont_touch of G8601: signal is true;
	signal G8602: std_logic; attribute dont_touch of G8602: signal is true;
	signal G8605: std_logic; attribute dont_touch of G8605: signal is true;
	signal G8612: std_logic; attribute dont_touch of G8612: signal is true;
	signal G8613: std_logic; attribute dont_touch of G8613: signal is true;
	signal G8614: std_logic; attribute dont_touch of G8614: signal is true;
	signal G8617: std_logic; attribute dont_touch of G8617: signal is true;
	signal G8620: std_logic; attribute dont_touch of G8620: signal is true;
	signal G8621: std_logic; attribute dont_touch of G8621: signal is true;
	signal G8622: std_logic; attribute dont_touch of G8622: signal is true;
	signal G8625: std_logic; attribute dont_touch of G8625: signal is true;
	signal G8626: std_logic; attribute dont_touch of G8626: signal is true;
	signal G8627: std_logic; attribute dont_touch of G8627: signal is true;
	signal G8630: std_logic; attribute dont_touch of G8630: signal is true;
	signal G8631: std_logic; attribute dont_touch of G8631: signal is true;
	signal G8632: std_logic; attribute dont_touch of G8632: signal is true;
	signal G8635: std_logic; attribute dont_touch of G8635: signal is true;
	signal G8636: std_logic; attribute dont_touch of G8636: signal is true;
	signal G8637: std_logic; attribute dont_touch of G8637: signal is true;
	signal G8640: std_logic; attribute dont_touch of G8640: signal is true;
	signal G8643: std_logic; attribute dont_touch of G8643: signal is true;
	signal G8646: std_logic; attribute dont_touch of G8646: signal is true;
	signal G8649: std_logic; attribute dont_touch of G8649: signal is true;
	signal G8650: std_logic; attribute dont_touch of G8650: signal is true;
	signal G8651: std_logic; attribute dont_touch of G8651: signal is true;
	signal G8654: std_logic; attribute dont_touch of G8654: signal is true;
	signal G8655: std_logic; attribute dont_touch of G8655: signal is true;
	signal G8658: std_logic; attribute dont_touch of G8658: signal is true;
	signal G8659: std_logic; attribute dont_touch of G8659: signal is true;
	signal G8662: std_logic; attribute dont_touch of G8662: signal is true;
	signal G8665: std_logic; attribute dont_touch of G8665: signal is true;
	signal G8666: std_logic; attribute dont_touch of G8666: signal is true;
	signal G8667: std_logic; attribute dont_touch of G8667: signal is true;
	signal G8670: std_logic; attribute dont_touch of G8670: signal is true;
	signal G8673: std_logic; attribute dont_touch of G8673: signal is true;
	signal G8676: std_logic; attribute dont_touch of G8676: signal is true;
	signal G8677: std_logic; attribute dont_touch of G8677: signal is true;
	signal G8678: std_logic; attribute dont_touch of G8678: signal is true;
	signal G8681: std_logic; attribute dont_touch of G8681: signal is true;
	signal G8684: std_logic; attribute dont_touch of G8684: signal is true;
	signal G8687: std_logic; attribute dont_touch of G8687: signal is true;
	signal G8688: std_logic; attribute dont_touch of G8688: signal is true;
	signal G8689: std_logic; attribute dont_touch of G8689: signal is true;
	signal G8690: std_logic; attribute dont_touch of G8690: signal is true;
	signal G8693: std_logic; attribute dont_touch of G8693: signal is true;
	signal G8696: std_logic; attribute dont_touch of G8696: signal is true;
	signal G8699: std_logic; attribute dont_touch of G8699: signal is true;
	signal G8700: std_logic; attribute dont_touch of G8700: signal is true;
	signal G8703: std_logic; attribute dont_touch of G8703: signal is true;
	signal G8704: std_logic; attribute dont_touch of G8704: signal is true;
	signal G8705: std_logic; attribute dont_touch of G8705: signal is true;
	signal G8706: std_logic; attribute dont_touch of G8706: signal is true;
	signal G8707: std_logic; attribute dont_touch of G8707: signal is true;
	signal G8708: std_logic; attribute dont_touch of G8708: signal is true;
	signal G8711: std_logic; attribute dont_touch of G8711: signal is true;
	signal G8714: std_logic; attribute dont_touch of G8714: signal is true;
	signal G8717: std_logic; attribute dont_touch of G8717: signal is true;
	signal G8718: std_logic; attribute dont_touch of G8718: signal is true;
	signal G8719: std_logic; attribute dont_touch of G8719: signal is true;
	signal G8722: std_logic; attribute dont_touch of G8722: signal is true;
	signal G8723: std_logic; attribute dont_touch of G8723: signal is true;
	signal G8724: std_logic; attribute dont_touch of G8724: signal is true;
	signal G8725: std_logic; attribute dont_touch of G8725: signal is true;
	signal G8726: std_logic; attribute dont_touch of G8726: signal is true;
	signal G8745: std_logic; attribute dont_touch of G8745: signal is true;
	signal G8748: std_logic; attribute dont_touch of G8748: signal is true;
	signal G8751: std_logic; attribute dont_touch of G8751: signal is true;
	signal G8752: std_logic; attribute dont_touch of G8752: signal is true;
	signal G8755: std_logic; attribute dont_touch of G8755: signal is true;
	signal G8756: std_logic; attribute dont_touch of G8756: signal is true;
	signal G8757: std_logic; attribute dont_touch of G8757: signal is true;
	signal G8760: std_logic; attribute dont_touch of G8760: signal is true;
	signal G8761: std_logic; attribute dont_touch of G8761: signal is true;
	signal G8762: std_logic; attribute dont_touch of G8762: signal is true;
	signal G8763: std_logic; attribute dont_touch of G8763: signal is true;
	signal G8766: std_logic; attribute dont_touch of G8766: signal is true;
	signal G8769: std_logic; attribute dont_touch of G8769: signal is true;
	signal G8770: std_logic; attribute dont_touch of G8770: signal is true;
	signal G8771: std_logic; attribute dont_touch of G8771: signal is true;
	signal G8774: std_logic; attribute dont_touch of G8774: signal is true;
	signal G8775: std_logic; attribute dont_touch of G8775: signal is true;
	signal G8778: std_logic; attribute dont_touch of G8778: signal is true;
	signal G8779: std_logic; attribute dont_touch of G8779: signal is true;
	signal G8780: std_logic; attribute dont_touch of G8780: signal is true;
	signal G8783: std_logic; attribute dont_touch of G8783: signal is true;
	signal G8784: std_logic; attribute dont_touch of G8784: signal is true;
	signal G8785: std_logic; attribute dont_touch of G8785: signal is true;
	signal G8788: std_logic; attribute dont_touch of G8788: signal is true;
	signal G8791: std_logic; attribute dont_touch of G8791: signal is true;
	signal G8792: std_logic; attribute dont_touch of G8792: signal is true;
	signal G8793: std_logic; attribute dont_touch of G8793: signal is true;
	signal G8794: std_logic; attribute dont_touch of G8794: signal is true;
	signal G8797: std_logic; attribute dont_touch of G8797: signal is true;
	signal G8798: std_logic; attribute dont_touch of G8798: signal is true;
	signal G8801: std_logic; attribute dont_touch of G8801: signal is true;
	signal G8802: std_logic; attribute dont_touch of G8802: signal is true;
	signal G8805: std_logic; attribute dont_touch of G8805: signal is true;
	signal G8808: std_logic; attribute dont_touch of G8808: signal is true;
	signal G8809: std_logic; attribute dont_touch of G8809: signal is true;
	signal G8810: std_logic; attribute dont_touch of G8810: signal is true;
	signal G8811: std_logic; attribute dont_touch of G8811: signal is true;
	signal G8812: std_logic; attribute dont_touch of G8812: signal is true;
	signal G8813: std_logic; attribute dont_touch of G8813: signal is true;
	signal G8816: std_logic; attribute dont_touch of G8816: signal is true;
	signal G8817: std_logic; attribute dont_touch of G8817: signal is true;
	signal G8820: std_logic; attribute dont_touch of G8820: signal is true;
	signal G8821: std_logic; attribute dont_touch of G8821: signal is true;
	signal G8822: std_logic; attribute dont_touch of G8822: signal is true;
	signal G8823: std_logic; attribute dont_touch of G8823: signal is true;
	signal G8824: std_logic; attribute dont_touch of G8824: signal is true;
	signal G8825: std_logic; attribute dont_touch of G8825: signal is true;
	signal G8826: std_logic; attribute dont_touch of G8826: signal is true;
	signal G8827: std_logic; attribute dont_touch of G8827: signal is true;
	signal G8828: std_logic; attribute dont_touch of G8828: signal is true;
	signal G8829: std_logic; attribute dont_touch of G8829: signal is true;
	signal G8832: std_logic; attribute dont_touch of G8832: signal is true;
	signal G8835: std_logic; attribute dont_touch of G8835: signal is true;
	signal G8836: std_logic; attribute dont_touch of G8836: signal is true;
	signal G8839: std_logic; attribute dont_touch of G8839: signal is true;
	signal G8840: std_logic; attribute dont_touch of G8840: signal is true;
	signal G8841: std_logic; attribute dont_touch of G8841: signal is true;
	signal G8842: std_logic; attribute dont_touch of G8842: signal is true;
	signal G8843: std_logic; attribute dont_touch of G8843: signal is true;
	signal G8844: std_logic; attribute dont_touch of G8844: signal is true;
	signal G8845: std_logic; attribute dont_touch of G8845: signal is true;
	signal G8846: std_logic; attribute dont_touch of G8846: signal is true;
	signal G8847: std_logic; attribute dont_touch of G8847: signal is true;
	signal G8850: std_logic; attribute dont_touch of G8850: signal is true;
	signal G8851: std_logic; attribute dont_touch of G8851: signal is true;
	signal G8852: std_logic; attribute dont_touch of G8852: signal is true;
	signal G8853: std_logic; attribute dont_touch of G8853: signal is true;
	signal G8856: std_logic; attribute dont_touch of G8856: signal is true;
	signal G8859: std_logic; attribute dont_touch of G8859: signal is true;
	signal G8860: std_logic; attribute dont_touch of G8860: signal is true;
	signal G8861: std_logic; attribute dont_touch of G8861: signal is true;
	signal G8862: std_logic; attribute dont_touch of G8862: signal is true;
	signal G8863: std_logic; attribute dont_touch of G8863: signal is true;
	signal G8866: std_logic; attribute dont_touch of G8866: signal is true;
	signal G8867: std_logic; attribute dont_touch of G8867: signal is true;
	signal G8868: std_logic; attribute dont_touch of G8868: signal is true;
	signal G8869: std_logic; attribute dont_touch of G8869: signal is true;
	signal G8870: std_logic; attribute dont_touch of G8870: signal is true;
	signal G8871: std_logic; attribute dont_touch of G8871: signal is true;
	signal G8872: std_logic; attribute dont_touch of G8872: signal is true;
	signal G8873: std_logic; attribute dont_touch of G8873: signal is true;
	signal G8874: std_logic; attribute dont_touch of G8874: signal is true;
	signal G8877: std_logic; attribute dont_touch of G8877: signal is true;
	signal G8878: std_logic; attribute dont_touch of G8878: signal is true;
	signal G8879: std_logic; attribute dont_touch of G8879: signal is true;
	signal G8882: std_logic; attribute dont_touch of G8882: signal is true;
	signal G8885: std_logic; attribute dont_touch of G8885: signal is true;
	signal G8888: std_logic; attribute dont_touch of G8888: signal is true;
	signal G8891: std_logic; attribute dont_touch of G8891: signal is true;
	signal G8892: std_logic; attribute dont_touch of G8892: signal is true;
	signal G8893: std_logic; attribute dont_touch of G8893: signal is true;
	signal G8894: std_logic; attribute dont_touch of G8894: signal is true;
	signal G8897: std_logic; attribute dont_touch of G8897: signal is true;
	signal G8898: std_logic; attribute dont_touch of G8898: signal is true;
	signal G8899: std_logic; attribute dont_touch of G8899: signal is true;
	signal G8900: std_logic; attribute dont_touch of G8900: signal is true;
	signal G8901: std_logic; attribute dont_touch of G8901: signal is true;
	signal G8904: std_logic; attribute dont_touch of G8904: signal is true;
	signal G8905: std_logic; attribute dont_touch of G8905: signal is true;
	signal G8906: std_logic; attribute dont_touch of G8906: signal is true;
	signal G8907: std_logic; attribute dont_touch of G8907: signal is true;
	signal G8908: std_logic; attribute dont_touch of G8908: signal is true;
	signal G8909: std_logic; attribute dont_touch of G8909: signal is true;
	signal G8910: std_logic; attribute dont_touch of G8910: signal is true;
	signal G8911: std_logic; attribute dont_touch of G8911: signal is true;
	signal G8912: std_logic; attribute dont_touch of G8912: signal is true;
	signal G8915: std_logic; attribute dont_touch of G8915: signal is true;
	signal G8918: std_logic; attribute dont_touch of G8918: signal is true;
	signal G8921: std_logic; attribute dont_touch of G8921: signal is true;
	signal G8924: std_logic; attribute dont_touch of G8924: signal is true;
	signal G8925: std_logic; attribute dont_touch of G8925: signal is true;
	signal G8928: std_logic; attribute dont_touch of G8928: signal is true;
	signal G8931: std_logic; attribute dont_touch of G8931: signal is true;
	signal G8932: std_logic; attribute dont_touch of G8932: signal is true;
	signal G8933: std_logic; attribute dont_touch of G8933: signal is true;
	signal G8934: std_logic; attribute dont_touch of G8934: signal is true;
	signal G8937: std_logic; attribute dont_touch of G8937: signal is true;
	signal G8938: std_logic; attribute dont_touch of G8938: signal is true;
	signal G8939: std_logic; attribute dont_touch of G8939: signal is true;
	signal G8940: std_logic; attribute dont_touch of G8940: signal is true;
	signal G8941: std_logic; attribute dont_touch of G8941: signal is true;
	signal G8944: std_logic; attribute dont_touch of G8944: signal is true;
	signal G8945: std_logic; attribute dont_touch of G8945: signal is true;
	signal G8946: std_logic; attribute dont_touch of G8946: signal is true;
	signal G8947: std_logic; attribute dont_touch of G8947: signal is true;
	signal G8948: std_logic; attribute dont_touch of G8948: signal is true;
	signal G8949: std_logic; attribute dont_touch of G8949: signal is true;
	signal G8952: std_logic; attribute dont_touch of G8952: signal is true;
	signal G8955: std_logic; attribute dont_touch of G8955: signal is true;
	signal G8958: std_logic; attribute dont_touch of G8958: signal is true;
	signal G8961: std_logic; attribute dont_touch of G8961: signal is true;
	signal G8964: std_logic; attribute dont_touch of G8964: signal is true;
	signal G8965: std_logic; attribute dont_touch of G8965: signal is true;
	signal G8968: std_logic; attribute dont_touch of G8968: signal is true;
	signal G8971: std_logic; attribute dont_touch of G8971: signal is true;
	signal G8972: std_logic; attribute dont_touch of G8972: signal is true;
	signal G8973: std_logic; attribute dont_touch of G8973: signal is true;
	signal G8974: std_logic; attribute dont_touch of G8974: signal is true;
	signal G8977: std_logic; attribute dont_touch of G8977: signal is true;
	signal G8978: std_logic; attribute dont_touch of G8978: signal is true;
	signal G8979: std_logic; attribute dont_touch of G8979: signal is true;
	signal G8980: std_logic; attribute dont_touch of G8980: signal is true;
	signal G8983: std_logic; attribute dont_touch of G8983: signal is true;
	signal G8984: std_logic; attribute dont_touch of G8984: signal is true;
	signal G8987: std_logic; attribute dont_touch of G8987: signal is true;
	signal G8990: std_logic; attribute dont_touch of G8990: signal is true;
	signal G8993: std_logic; attribute dont_touch of G8993: signal is true;
	signal G8996: std_logic; attribute dont_touch of G8996: signal is true;
	signal G8997: std_logic; attribute dont_touch of G8997: signal is true;
	signal G9000: std_logic; attribute dont_touch of G9000: signal is true;
	signal G9003: std_logic; attribute dont_touch of G9003: signal is true;
	signal G9004: std_logic; attribute dont_touch of G9004: signal is true;
	signal G9005: std_logic; attribute dont_touch of G9005: signal is true;
	signal G9006: std_logic; attribute dont_touch of G9006: signal is true;
	signal G9009: std_logic; attribute dont_touch of G9009: signal is true;
	signal G9010: std_logic; attribute dont_touch of G9010: signal is true;
	signal G9013: std_logic; attribute dont_touch of G9013: signal is true;
	signal G9016: std_logic; attribute dont_touch of G9016: signal is true;
	signal G9019: std_logic; attribute dont_touch of G9019: signal is true;
	signal G9022: std_logic; attribute dont_touch of G9022: signal is true;
	signal G9025: std_logic; attribute dont_touch of G9025: signal is true;
	signal G9026: std_logic; attribute dont_touch of G9026: signal is true;
	signal G9027: std_logic; attribute dont_touch of G9027: signal is true;
	signal G9033: std_logic; attribute dont_touch of G9033: signal is true;
	signal G9034: std_logic; attribute dont_touch of G9034: signal is true;
	signal G9035: std_logic; attribute dont_touch of G9035: signal is true;
	signal G9038: std_logic; attribute dont_touch of G9038: signal is true;
	signal G9041: std_logic; attribute dont_touch of G9041: signal is true;
	signal G9044: std_logic; attribute dont_touch of G9044: signal is true;
	signal G9047: std_logic; attribute dont_touch of G9047: signal is true;
	signal G9048: std_logic; attribute dont_touch of G9048: signal is true;
	signal G9049: std_logic; attribute dont_touch of G9049: signal is true;
	signal G9050: std_logic; attribute dont_touch of G9050: signal is true;
	signal G9056: std_logic; attribute dont_touch of G9056: signal is true;
	signal G9057: std_logic; attribute dont_touch of G9057: signal is true;
	signal G9058: std_logic; attribute dont_touch of G9058: signal is true;
	signal G9061: std_logic; attribute dont_touch of G9061: signal is true;
	signal G9062: std_logic; attribute dont_touch of G9062: signal is true;
	signal G9063: std_logic; attribute dont_touch of G9063: signal is true;
	signal G9064: std_logic; attribute dont_touch of G9064: signal is true;
	signal G9065: std_logic; attribute dont_touch of G9065: signal is true;
	signal G9066: std_logic; attribute dont_touch of G9066: signal is true;
	signal G9067: std_logic; attribute dont_touch of G9067: signal is true;
	signal G9073: std_logic; attribute dont_touch of G9073: signal is true;
	signal G9074: std_logic; attribute dont_touch of G9074: signal is true;
	signal G9075: std_logic; attribute dont_touch of G9075: signal is true;
	signal G9076: std_logic; attribute dont_touch of G9076: signal is true;
	signal G9077: std_logic; attribute dont_touch of G9077: signal is true;
	signal G9078: std_logic; attribute dont_touch of G9078: signal is true;
	signal G9079: std_logic; attribute dont_touch of G9079: signal is true;
	signal G9080: std_logic; attribute dont_touch of G9080: signal is true;
	signal G9081: std_logic; attribute dont_touch of G9081: signal is true;
	signal G9082: std_logic; attribute dont_touch of G9082: signal is true;
	signal G9083: std_logic; attribute dont_touch of G9083: signal is true;
	signal G9084: std_logic; attribute dont_touch of G9084: signal is true;
	signal G9090: std_logic; attribute dont_touch of G9090: signal is true;
	signal G9091: std_logic; attribute dont_touch of G9091: signal is true;
	signal G9092: std_logic; attribute dont_touch of G9092: signal is true;
	signal G9093: std_logic; attribute dont_touch of G9093: signal is true;
	signal G9094: std_logic; attribute dont_touch of G9094: signal is true;
	signal G9095: std_logic; attribute dont_touch of G9095: signal is true;
	signal G9096: std_logic; attribute dont_touch of G9096: signal is true;
	signal G9097: std_logic; attribute dont_touch of G9097: signal is true;
	signal G9098: std_logic; attribute dont_touch of G9098: signal is true;
	signal G9099: std_logic; attribute dont_touch of G9099: signal is true;
	signal G9100: std_logic; attribute dont_touch of G9100: signal is true;
	signal G9101: std_logic; attribute dont_touch of G9101: signal is true;
	signal G9102: std_logic; attribute dont_touch of G9102: signal is true;
	signal G9103: std_logic; attribute dont_touch of G9103: signal is true;
	signal G9104: std_logic; attribute dont_touch of G9104: signal is true;
	signal G9105: std_logic; attribute dont_touch of G9105: signal is true;
	signal G9106: std_logic; attribute dont_touch of G9106: signal is true;
	signal G9107: std_logic; attribute dont_touch of G9107: signal is true;
	signal G9108: std_logic; attribute dont_touch of G9108: signal is true;
	signal G9109: std_logic; attribute dont_touch of G9109: signal is true;
	signal G9110: std_logic; attribute dont_touch of G9110: signal is true;
	signal G9111: std_logic; attribute dont_touch of G9111: signal is true;
	signal G9112: std_logic; attribute dont_touch of G9112: signal is true;
	signal G9113: std_logic; attribute dont_touch of G9113: signal is true;
	signal G9114: std_logic; attribute dont_touch of G9114: signal is true;
	signal G9115: std_logic; attribute dont_touch of G9115: signal is true;
	signal G9116: std_logic; attribute dont_touch of G9116: signal is true;
	signal G9117: std_logic; attribute dont_touch of G9117: signal is true;
	signal G9118: std_logic; attribute dont_touch of G9118: signal is true;
	signal G9119: std_logic; attribute dont_touch of G9119: signal is true;
	signal G9120: std_logic; attribute dont_touch of G9120: signal is true;
	signal G9121: std_logic; attribute dont_touch of G9121: signal is true;
	signal G9122: std_logic; attribute dont_touch of G9122: signal is true;
	signal G9123: std_logic; attribute dont_touch of G9123: signal is true;
	signal G9124: std_logic; attribute dont_touch of G9124: signal is true;
	signal G9125: std_logic; attribute dont_touch of G9125: signal is true;
	signal G9126: std_logic; attribute dont_touch of G9126: signal is true;
	signal G9127: std_logic; attribute dont_touch of G9127: signal is true;
	signal G9128: std_logic; attribute dont_touch of G9128: signal is true;
	signal G9131: std_logic; attribute dont_touch of G9131: signal is true;
	signal G9132: std_logic; attribute dont_touch of G9132: signal is true;
	signal G9133: std_logic; attribute dont_touch of G9133: signal is true;
	signal G9134: std_logic; attribute dont_touch of G9134: signal is true;
	signal G9137: std_logic; attribute dont_touch of G9137: signal is true;
	signal G9138: std_logic; attribute dont_touch of G9138: signal is true;
	signal G9139: std_logic; attribute dont_touch of G9139: signal is true;
	signal G9140: std_logic; attribute dont_touch of G9140: signal is true;
	signal G9143: std_logic; attribute dont_touch of G9143: signal is true;
	signal G9144: std_logic; attribute dont_touch of G9144: signal is true;
	signal G9145: std_logic; attribute dont_touch of G9145: signal is true;
	signal G9146: std_logic; attribute dont_touch of G9146: signal is true;
	signal G9149: std_logic; attribute dont_touch of G9149: signal is true;
	signal G9150: std_logic; attribute dont_touch of G9150: signal is true;
	signal G9159: std_logic; attribute dont_touch of G9159: signal is true;
	signal G9160: std_logic; attribute dont_touch of G9160: signal is true;
	signal G9161: std_logic; attribute dont_touch of G9161: signal is true;
	signal G9170: std_logic; attribute dont_touch of G9170: signal is true;
	signal G9173: std_logic; attribute dont_touch of G9173: signal is true;
	signal G9174: std_logic; attribute dont_touch of G9174: signal is true;
	signal G9183: std_logic; attribute dont_touch of G9183: signal is true;
	signal G9184: std_logic; attribute dont_touch of G9184: signal is true;
	signal G9187: std_logic; attribute dont_touch of G9187: signal is true;
	signal G9196: std_logic; attribute dont_touch of G9196: signal is true;
	signal G9199: std_logic; attribute dont_touch of G9199: signal is true;
	signal G9202: std_logic; attribute dont_touch of G9202: signal is true;
	signal G9203: std_logic; attribute dont_touch of G9203: signal is true;
	signal G9212: std_logic; attribute dont_touch of G9212: signal is true;
	signal G9215: std_logic; attribute dont_touch of G9215: signal is true;
	signal G9216: std_logic; attribute dont_touch of G9216: signal is true;
	signal G9225: std_logic; attribute dont_touch of G9225: signal is true;
	signal G9226: std_logic; attribute dont_touch of G9226: signal is true;
	signal G9227: std_logic; attribute dont_touch of G9227: signal is true;
	signal G9228: std_logic; attribute dont_touch of G9228: signal is true;
	signal G9229: std_logic; attribute dont_touch of G9229: signal is true;
	signal G9232: std_logic; attribute dont_touch of G9232: signal is true;
	signal G9241: std_logic; attribute dont_touch of G9241: signal is true;
	signal G9242: std_logic; attribute dont_touch of G9242: signal is true;
	signal G9245: std_logic; attribute dont_touch of G9245: signal is true;
	signal G9248: std_logic; attribute dont_touch of G9248: signal is true;
	signal G9257: std_logic; attribute dont_touch of G9257: signal is true;
	signal G9260: std_logic; attribute dont_touch of G9260: signal is true;
	signal G9263: std_logic; attribute dont_touch of G9263: signal is true;
	signal G9264: std_logic; attribute dont_touch of G9264: signal is true;
	signal G9273: std_logic; attribute dont_touch of G9273: signal is true;
	signal G9276: std_logic; attribute dont_touch of G9276: signal is true;
	signal G9277: std_logic; attribute dont_touch of G9277: signal is true;
	signal G9286: std_logic; attribute dont_touch of G9286: signal is true;
	signal G9287: std_logic; attribute dont_touch of G9287: signal is true;
	signal G9288: std_logic; attribute dont_touch of G9288: signal is true;
	signal G9289: std_logic; attribute dont_touch of G9289: signal is true;
	signal G9290: std_logic; attribute dont_touch of G9290: signal is true;
	signal G9293: std_logic; attribute dont_touch of G9293: signal is true;
	signal G9301: std_logic; attribute dont_touch of G9301: signal is true;
	signal G9302: std_logic; attribute dont_touch of G9302: signal is true;
	signal G9303: std_logic; attribute dont_touch of G9303: signal is true;
	signal G9306: std_logic; attribute dont_touch of G9306: signal is true;
	signal G9309: std_logic; attribute dont_touch of G9309: signal is true;
	signal G9310: std_logic; attribute dont_touch of G9310: signal is true;
	signal G9319: std_logic; attribute dont_touch of G9319: signal is true;
	signal G9320: std_logic; attribute dont_touch of G9320: signal is true;
	signal G9323: std_logic; attribute dont_touch of G9323: signal is true;
	signal G9326: std_logic; attribute dont_touch of G9326: signal is true;
	signal G9335: std_logic; attribute dont_touch of G9335: signal is true;
	signal G9338: std_logic; attribute dont_touch of G9338: signal is true;
	signal G9341: std_logic; attribute dont_touch of G9341: signal is true;
	signal G9342: std_logic; attribute dont_touch of G9342: signal is true;
	signal G9351: std_logic; attribute dont_touch of G9351: signal is true;
	signal G9354: std_logic; attribute dont_touch of G9354: signal is true;
	signal G9355: std_logic; attribute dont_touch of G9355: signal is true;
	signal G9356: std_logic; attribute dont_touch of G9356: signal is true;
	signal G9364: std_logic; attribute dont_touch of G9364: signal is true;
	signal G9365: std_logic; attribute dont_touch of G9365: signal is true;
	signal G9366: std_logic; attribute dont_touch of G9366: signal is true;
	signal G9367: std_logic; attribute dont_touch of G9367: signal is true;
	signal G9368: std_logic; attribute dont_touch of G9368: signal is true;
	signal G9371: std_logic; attribute dont_touch of G9371: signal is true;
	signal G9374: std_logic; attribute dont_touch of G9374: signal is true;
	signal G9382: std_logic; attribute dont_touch of G9382: signal is true;
	signal G9383: std_logic; attribute dont_touch of G9383: signal is true;
	signal G9384: std_logic; attribute dont_touch of G9384: signal is true;
	signal G9387: std_logic; attribute dont_touch of G9387: signal is true;
	signal G9390: std_logic; attribute dont_touch of G9390: signal is true;
	signal G9391: std_logic; attribute dont_touch of G9391: signal is true;
	signal G9400: std_logic; attribute dont_touch of G9400: signal is true;
	signal G9401: std_logic; attribute dont_touch of G9401: signal is true;
	signal G9404: std_logic; attribute dont_touch of G9404: signal is true;
	signal G9407: std_logic; attribute dont_touch of G9407: signal is true;
	signal G9416: std_logic; attribute dont_touch of G9416: signal is true;
	signal G9419: std_logic; attribute dont_touch of G9419: signal is true;
	signal G9422: std_logic; attribute dont_touch of G9422: signal is true;
	signal G9423: std_logic; attribute dont_touch of G9423: signal is true;
	signal G9424: std_logic; attribute dont_touch of G9424: signal is true;
	signal G9425: std_logic; attribute dont_touch of G9425: signal is true;
	signal G9426: std_logic; attribute dont_touch of G9426: signal is true;
	signal G9427: std_logic; attribute dont_touch of G9427: signal is true;
	signal G9438: std_logic; attribute dont_touch of G9438: signal is true;
	signal G9439: std_logic; attribute dont_touch of G9439: signal is true;
	signal G9440: std_logic; attribute dont_touch of G9440: signal is true;
	signal G9441: std_logic; attribute dont_touch of G9441: signal is true;
	signal G9442: std_logic; attribute dont_touch of G9442: signal is true;
	signal G9443: std_logic; attribute dont_touch of G9443: signal is true;
	signal G9446: std_logic; attribute dont_touch of G9446: signal is true;
	signal G9449: std_logic; attribute dont_touch of G9449: signal is true;
	signal G9450: std_logic; attribute dont_touch of G9450: signal is true;
	signal G9453: std_logic; attribute dont_touch of G9453: signal is true;
	signal G9461: std_logic; attribute dont_touch of G9461: signal is true;
	signal G9462: std_logic; attribute dont_touch of G9462: signal is true;
	signal G9463: std_logic; attribute dont_touch of G9463: signal is true;
	signal G9464: std_logic; attribute dont_touch of G9464: signal is true;
	signal G9465: std_logic; attribute dont_touch of G9465: signal is true;
	signal G9468: std_logic; attribute dont_touch of G9468: signal is true;
	signal G9471: std_logic; attribute dont_touch of G9471: signal is true;
	signal G9479: std_logic; attribute dont_touch of G9479: signal is true;
	signal G9480: std_logic; attribute dont_touch of G9480: signal is true;
	signal G9481: std_logic; attribute dont_touch of G9481: signal is true;
	signal G9484: std_logic; attribute dont_touch of G9484: signal is true;
	signal G9487: std_logic; attribute dont_touch of G9487: signal is true;
	signal G9488: std_logic; attribute dont_touch of G9488: signal is true;
	signal G9497: std_logic; attribute dont_touch of G9497: signal is true;
	signal G9498: std_logic; attribute dont_touch of G9498: signal is true;
	signal G9501: std_logic; attribute dont_touch of G9501: signal is true;
	signal G9504: std_logic; attribute dont_touch of G9504: signal is true;
	signal G9505: std_logic; attribute dont_touch of G9505: signal is true;
	signal G9506: std_logic; attribute dont_touch of G9506: signal is true;
	signal G9507: std_logic; attribute dont_touch of G9507: signal is true;
	signal G9518: std_logic; attribute dont_touch of G9518: signal is true;
	signal G9519: std_logic; attribute dont_touch of G9519: signal is true;
	signal G9520: std_logic; attribute dont_touch of G9520: signal is true;
	signal G9521: std_logic; attribute dont_touch of G9521: signal is true;
	signal G9522: std_logic; attribute dont_touch of G9522: signal is true;
	signal G9523: std_logic; attribute dont_touch of G9523: signal is true;
	signal G9524: std_logic; attribute dont_touch of G9524: signal is true;
	signal G9527: std_logic; attribute dont_touch of G9527: signal is true;
	signal G9528: std_logic; attribute dont_touch of G9528: signal is true;
	signal G9531: std_logic; attribute dont_touch of G9531: signal is true;
	signal G9534: std_logic; attribute dont_touch of G9534: signal is true;
	signal G9569: std_logic; attribute dont_touch of G9569: signal is true;
	signal G9580: std_logic; attribute dont_touch of G9580: signal is true;
	signal G9581: std_logic; attribute dont_touch of G9581: signal is true;
	signal G9582: std_logic; attribute dont_touch of G9582: signal is true;
	signal G9583: std_logic; attribute dont_touch of G9583: signal is true;
	signal G9584: std_logic; attribute dont_touch of G9584: signal is true;
	signal G9585: std_logic; attribute dont_touch of G9585: signal is true;
	signal G9588: std_logic; attribute dont_touch of G9588: signal is true;
	signal G9591: std_logic; attribute dont_touch of G9591: signal is true;
	signal G9592: std_logic; attribute dont_touch of G9592: signal is true;
	signal G9595: std_logic; attribute dont_touch of G9595: signal is true;
	signal G9603: std_logic; attribute dont_touch of G9603: signal is true;
	signal G9604: std_logic; attribute dont_touch of G9604: signal is true;
	signal G9605: std_logic; attribute dont_touch of G9605: signal is true;
	signal G9606: std_logic; attribute dont_touch of G9606: signal is true;
	signal G9607: std_logic; attribute dont_touch of G9607: signal is true;
	signal G9610: std_logic; attribute dont_touch of G9610: signal is true;
	signal G9613: std_logic; attribute dont_touch of G9613: signal is true;
	signal G9621: std_logic; attribute dont_touch of G9621: signal is true;
	signal G9622: std_logic; attribute dont_touch of G9622: signal is true;
	signal G9623: std_logic; attribute dont_touch of G9623: signal is true;
	signal G9626: std_logic; attribute dont_touch of G9626: signal is true;
	signal G9629: std_logic; attribute dont_touch of G9629: signal is true;
	signal G9630: std_logic; attribute dont_touch of G9630: signal is true;
	signal G9631: std_logic; attribute dont_touch of G9631: signal is true;
	signal G9632: std_logic; attribute dont_touch of G9632: signal is true;
	signal G9633: std_logic; attribute dont_touch of G9633: signal is true;
	signal G9634: std_logic; attribute dont_touch of G9634: signal is true;
	signal G9635: std_logic; attribute dont_touch of G9635: signal is true;
	signal G9636: std_logic; attribute dont_touch of G9636: signal is true;
	signal G9639: std_logic; attribute dont_touch of G9639: signal is true;
	signal G9640: std_logic; attribute dont_touch of G9640: signal is true;
	signal G9641: std_logic; attribute dont_touch of G9641: signal is true;
	signal G9644: std_logic; attribute dont_touch of G9644: signal is true;
	signal G9647: std_logic; attribute dont_touch of G9647: signal is true;
	signal G9648: std_logic; attribute dont_touch of G9648: signal is true;
	signal G9649: std_logic; attribute dont_touch of G9649: signal is true;
	signal G9660: std_logic; attribute dont_touch of G9660: signal is true;
	signal G9661: std_logic; attribute dont_touch of G9661: signal is true;
	signal G9662: std_logic; attribute dont_touch of G9662: signal is true;
	signal G9663: std_logic; attribute dont_touch of G9663: signal is true;
	signal G9664: std_logic; attribute dont_touch of G9664: signal is true;
	signal G9665: std_logic; attribute dont_touch of G9665: signal is true;
	signal G9666: std_logic; attribute dont_touch of G9666: signal is true;
	signal G9669: std_logic; attribute dont_touch of G9669: signal is true;
	signal G9670: std_logic; attribute dont_touch of G9670: signal is true;
	signal G9673: std_logic; attribute dont_touch of G9673: signal is true;
	signal G9676: std_logic; attribute dont_touch of G9676: signal is true;
	signal G9711: std_logic; attribute dont_touch of G9711: signal is true;
	signal G9722: std_logic; attribute dont_touch of G9722: signal is true;
	signal G9723: std_logic; attribute dont_touch of G9723: signal is true;
	signal G9724: std_logic; attribute dont_touch of G9724: signal is true;
	signal G9725: std_logic; attribute dont_touch of G9725: signal is true;
	signal G9726: std_logic; attribute dont_touch of G9726: signal is true;
	signal G9727: std_logic; attribute dont_touch of G9727: signal is true;
	signal G9730: std_logic; attribute dont_touch of G9730: signal is true;
	signal G9733: std_logic; attribute dont_touch of G9733: signal is true;
	signal G9734: std_logic; attribute dont_touch of G9734: signal is true;
	signal G9737: std_logic; attribute dont_touch of G9737: signal is true;
	signal G9745: std_logic; attribute dont_touch of G9745: signal is true;
	signal G9746: std_logic; attribute dont_touch of G9746: signal is true;
	signal G9747: std_logic; attribute dont_touch of G9747: signal is true;
	signal G9748: std_logic; attribute dont_touch of G9748: signal is true;
	signal G9749: std_logic; attribute dont_touch of G9749: signal is true;
	signal G9752: std_logic; attribute dont_touch of G9752: signal is true;
	signal G9755: std_logic; attribute dont_touch of G9755: signal is true;
	signal G9756: std_logic; attribute dont_touch of G9756: signal is true;
	signal G9757: std_logic; attribute dont_touch of G9757: signal is true;
	signal G9758: std_logic; attribute dont_touch of G9758: signal is true;
	signal G9759: std_logic; attribute dont_touch of G9759: signal is true;
	signal G9760: std_logic; attribute dont_touch of G9760: signal is true;
	signal G9761: std_logic; attribute dont_touch of G9761: signal is true;
	signal G9762: std_logic; attribute dont_touch of G9762: signal is true;
	signal G9763: std_logic; attribute dont_touch of G9763: signal is true;
	signal G9764: std_logic; attribute dont_touch of G9764: signal is true;
	signal G9765: std_logic; attribute dont_touch of G9765: signal is true;
	signal G9766: std_logic; attribute dont_touch of G9766: signal is true;
	signal G9767: std_logic; attribute dont_touch of G9767: signal is true;
	signal G9770: std_logic; attribute dont_touch of G9770: signal is true;
	signal G9773: std_logic; attribute dont_touch of G9773: signal is true;
	signal G9774: std_logic; attribute dont_touch of G9774: signal is true;
	signal G9775: std_logic; attribute dont_touch of G9775: signal is true;
	signal G9776: std_logic; attribute dont_touch of G9776: signal is true;
	signal G9777: std_logic; attribute dont_touch of G9777: signal is true;
	signal G9778: std_logic; attribute dont_touch of G9778: signal is true;
	signal G9779: std_logic; attribute dont_touch of G9779: signal is true;
	signal G9780: std_logic; attribute dont_touch of G9780: signal is true;
	signal G9781: std_logic; attribute dont_touch of G9781: signal is true;
	signal G9782: std_logic; attribute dont_touch of G9782: signal is true;
	signal G9785: std_logic; attribute dont_touch of G9785: signal is true;
	signal G9786: std_logic; attribute dont_touch of G9786: signal is true;
	signal G9787: std_logic; attribute dont_touch of G9787: signal is true;
	signal G9790: std_logic; attribute dont_touch of G9790: signal is true;
	signal G9793: std_logic; attribute dont_touch of G9793: signal is true;
	signal G9794: std_logic; attribute dont_touch of G9794: signal is true;
	signal G9795: std_logic; attribute dont_touch of G9795: signal is true;
	signal G9806: std_logic; attribute dont_touch of G9806: signal is true;
	signal G9807: std_logic; attribute dont_touch of G9807: signal is true;
	signal G9808: std_logic; attribute dont_touch of G9808: signal is true;
	signal G9809: std_logic; attribute dont_touch of G9809: signal is true;
	signal G9810: std_logic; attribute dont_touch of G9810: signal is true;
	signal G9811: std_logic; attribute dont_touch of G9811: signal is true;
	signal G9812: std_logic; attribute dont_touch of G9812: signal is true;
	signal G9815: std_logic; attribute dont_touch of G9815: signal is true;
	signal G9816: std_logic; attribute dont_touch of G9816: signal is true;
	signal G9819: std_logic; attribute dont_touch of G9819: signal is true;
	signal G9822: std_logic; attribute dont_touch of G9822: signal is true;
	signal G9857: std_logic; attribute dont_touch of G9857: signal is true;
	signal G9868: std_logic; attribute dont_touch of G9868: signal is true;
	signal G9869: std_logic; attribute dont_touch of G9869: signal is true;
	signal G9870: std_logic; attribute dont_touch of G9870: signal is true;
	signal G9871: std_logic; attribute dont_touch of G9871: signal is true;
	signal G9872: std_logic; attribute dont_touch of G9872: signal is true;
	signal G9873: std_logic; attribute dont_touch of G9873: signal is true;
	signal G9876: std_logic; attribute dont_touch of G9876: signal is true;
	signal G9879: std_logic; attribute dont_touch of G9879: signal is true;
	signal G9880: std_logic; attribute dont_touch of G9880: signal is true;
	signal G9883: std_logic; attribute dont_touch of G9883: signal is true;
	signal G9884: std_logic; attribute dont_touch of G9884: signal is true;
	signal G9885: std_logic; attribute dont_touch of G9885: signal is true;
	signal G9886: std_logic; attribute dont_touch of G9886: signal is true;
	signal G9887: std_logic; attribute dont_touch of G9887: signal is true;
	signal G9888: std_logic; attribute dont_touch of G9888: signal is true;
	signal G9889: std_logic; attribute dont_touch of G9889: signal is true;
	signal G9890: std_logic; attribute dont_touch of G9890: signal is true;
	signal G9891: std_logic; attribute dont_touch of G9891: signal is true;
	signal G9892: std_logic; attribute dont_touch of G9892: signal is true;
	signal G9893: std_logic; attribute dont_touch of G9893: signal is true;
	signal G9894: std_logic; attribute dont_touch of G9894: signal is true;
	signal G9895: std_logic; attribute dont_touch of G9895: signal is true;
	signal G9898: std_logic; attribute dont_touch of G9898: signal is true;
	signal G9901: std_logic; attribute dont_touch of G9901: signal is true;
	signal G9902: std_logic; attribute dont_touch of G9902: signal is true;
	signal G9903: std_logic; attribute dont_touch of G9903: signal is true;
	signal G9904: std_logic; attribute dont_touch of G9904: signal is true;
	signal G9905: std_logic; attribute dont_touch of G9905: signal is true;
	signal G9906: std_logic; attribute dont_touch of G9906: signal is true;
	signal G9907: std_logic; attribute dont_touch of G9907: signal is true;
	signal G9908: std_logic; attribute dont_touch of G9908: signal is true;
	signal G9909: std_logic; attribute dont_touch of G9909: signal is true;
	signal G9910: std_logic; attribute dont_touch of G9910: signal is true;
	signal G9911: std_logic; attribute dont_touch of G9911: signal is true;
	signal G9912: std_logic; attribute dont_touch of G9912: signal is true;
	signal G9913: std_logic; attribute dont_touch of G9913: signal is true;
	signal G9916: std_logic; attribute dont_touch of G9916: signal is true;
	signal G9919: std_logic; attribute dont_touch of G9919: signal is true;
	signal G9920: std_logic; attribute dont_touch of G9920: signal is true;
	signal G9921: std_logic; attribute dont_touch of G9921: signal is true;
	signal G9922: std_logic; attribute dont_touch of G9922: signal is true;
	signal G9923: std_logic; attribute dont_touch of G9923: signal is true;
	signal G9924: std_logic; attribute dont_touch of G9924: signal is true;
	signal G9925: std_logic; attribute dont_touch of G9925: signal is true;
	signal G9926: std_logic; attribute dont_touch of G9926: signal is true;
	signal G9927: std_logic; attribute dont_touch of G9927: signal is true;
	signal G9928: std_logic; attribute dont_touch of G9928: signal is true;
	signal G9931: std_logic; attribute dont_touch of G9931: signal is true;
	signal G9932: std_logic; attribute dont_touch of G9932: signal is true;
	signal G9933: std_logic; attribute dont_touch of G9933: signal is true;
	signal G9936: std_logic; attribute dont_touch of G9936: signal is true;
	signal G9939: std_logic; attribute dont_touch of G9939: signal is true;
	signal G9940: std_logic; attribute dont_touch of G9940: signal is true;
	signal G9941: std_logic; attribute dont_touch of G9941: signal is true;
	signal G9952: std_logic; attribute dont_touch of G9952: signal is true;
	signal G9953: std_logic; attribute dont_touch of G9953: signal is true;
	signal G9954: std_logic; attribute dont_touch of G9954: signal is true;
	signal G9955: std_logic; attribute dont_touch of G9955: signal is true;
	signal G9956: std_logic; attribute dont_touch of G9956: signal is true;
	signal G9957: std_logic; attribute dont_touch of G9957: signal is true;
	signal G9958: std_logic; attribute dont_touch of G9958: signal is true;
	signal G9961: std_logic; attribute dont_touch of G9961: signal is true;
	signal G9962: std_logic; attribute dont_touch of G9962: signal is true;
	signal G9965: std_logic; attribute dont_touch of G9965: signal is true;
	signal G9968: std_logic; attribute dont_touch of G9968: signal is true;
	signal G10003: std_logic; attribute dont_touch of G10003: signal is true;
	signal G10004: std_logic; attribute dont_touch of G10004: signal is true;
	signal G10007: std_logic; attribute dont_touch of G10007: signal is true;
	signal G10008: std_logic; attribute dont_touch of G10008: signal is true;
	signal G10009: std_logic; attribute dont_touch of G10009: signal is true;
	signal G10010: std_logic; attribute dont_touch of G10010: signal is true;
	signal G10011: std_logic; attribute dont_touch of G10011: signal is true;
	signal G10012: std_logic; attribute dont_touch of G10012: signal is true;
	signal G10013: std_logic; attribute dont_touch of G10013: signal is true;
	signal G10014: std_logic; attribute dont_touch of G10014: signal is true;
	signal G10015: std_logic; attribute dont_touch of G10015: signal is true;
	signal G10016: std_logic; attribute dont_touch of G10016: signal is true;
	signal G10017: std_logic; attribute dont_touch of G10017: signal is true;
	signal G10018: std_logic; attribute dont_touch of G10018: signal is true;
	signal G10021: std_logic; attribute dont_touch of G10021: signal is true;
	signal G10024: std_logic; attribute dont_touch of G10024: signal is true;
	signal G10035: std_logic; attribute dont_touch of G10035: signal is true;
	signal G10036: std_logic; attribute dont_touch of G10036: signal is true;
	signal G10037: std_logic; attribute dont_touch of G10037: signal is true;
	signal G10038: std_logic; attribute dont_touch of G10038: signal is true;
	signal G10041: std_logic; attribute dont_touch of G10041: signal is true;
	signal G10042: std_logic; attribute dont_touch of G10042: signal is true;
	signal G10043: std_logic; attribute dont_touch of G10043: signal is true;
	signal G10044: std_logic; attribute dont_touch of G10044: signal is true;
	signal G10045: std_logic; attribute dont_touch of G10045: signal is true;
	signal G10046: std_logic; attribute dont_touch of G10046: signal is true;
	signal G10047: std_logic; attribute dont_touch of G10047: signal is true;
	signal G10048: std_logic; attribute dont_touch of G10048: signal is true;
	signal G10049: std_logic; attribute dont_touch of G10049: signal is true;
	signal G10052: std_logic; attribute dont_touch of G10052: signal is true;
	signal G10055: std_logic; attribute dont_touch of G10055: signal is true;
	signal G10056: std_logic; attribute dont_touch of G10056: signal is true;
	signal G10057: std_logic; attribute dont_touch of G10057: signal is true;
	signal G10058: std_logic; attribute dont_touch of G10058: signal is true;
	signal G10059: std_logic; attribute dont_touch of G10059: signal is true;
	signal G10060: std_logic; attribute dont_touch of G10060: signal is true;
	signal G10061: std_logic; attribute dont_touch of G10061: signal is true;
	signal G10062: std_logic; attribute dont_touch of G10062: signal is true;
	signal G10063: std_logic; attribute dont_touch of G10063: signal is true;
	signal G10064: std_logic; attribute dont_touch of G10064: signal is true;
	signal G10065: std_logic; attribute dont_touch of G10065: signal is true;
	signal G10066: std_logic; attribute dont_touch of G10066: signal is true;
	signal G10067: std_logic; attribute dont_touch of G10067: signal is true;
	signal G10070: std_logic; attribute dont_touch of G10070: signal is true;
	signal G10073: std_logic; attribute dont_touch of G10073: signal is true;
	signal G10074: std_logic; attribute dont_touch of G10074: signal is true;
	signal G10075: std_logic; attribute dont_touch of G10075: signal is true;
	signal G10076: std_logic; attribute dont_touch of G10076: signal is true;
	signal G10077: std_logic; attribute dont_touch of G10077: signal is true;
	signal G10078: std_logic; attribute dont_touch of G10078: signal is true;
	signal G10079: std_logic; attribute dont_touch of G10079: signal is true;
	signal G10080: std_logic; attribute dont_touch of G10080: signal is true;
	signal G10081: std_logic; attribute dont_touch of G10081: signal is true;
	signal G10082: std_logic; attribute dont_touch of G10082: signal is true;
	signal G10085: std_logic; attribute dont_touch of G10085: signal is true;
	signal G10086: std_logic; attribute dont_touch of G10086: signal is true;
	signal G10087: std_logic; attribute dont_touch of G10087: signal is true;
	signal G10090: std_logic; attribute dont_touch of G10090: signal is true;
	signal G10093: std_logic; attribute dont_touch of G10093: signal is true;
	signal G10094: std_logic; attribute dont_touch of G10094: signal is true;
	signal G10095: std_logic; attribute dont_touch of G10095: signal is true;
	signal G10096: std_logic; attribute dont_touch of G10096: signal is true;
	signal G10099: std_logic; attribute dont_touch of G10099: signal is true;
	signal G10100: std_logic; attribute dont_touch of G10100: signal is true;
	signal G10101: std_logic; attribute dont_touch of G10101: signal is true;
	signal G10102: std_logic; attribute dont_touch of G10102: signal is true;
	signal G10103: std_logic; attribute dont_touch of G10103: signal is true;
	signal G10104: std_logic; attribute dont_touch of G10104: signal is true;
	signal G10105: std_logic; attribute dont_touch of G10105: signal is true;
	signal G10106: std_logic; attribute dont_touch of G10106: signal is true;
	signal G10107: std_logic; attribute dont_touch of G10107: signal is true;
	signal G10108: std_logic; attribute dont_touch of G10108: signal is true;
	signal G10109: std_logic; attribute dont_touch of G10109: signal is true;
	signal G10112: std_logic; attribute dont_touch of G10112: signal is true;
	signal G10113: std_logic; attribute dont_touch of G10113: signal is true;
	signal G10114: std_logic; attribute dont_touch of G10114: signal is true;
	signal G10115: std_logic; attribute dont_touch of G10115: signal is true;
	signal G10116: std_logic; attribute dont_touch of G10116: signal is true;
	signal G10117: std_logic; attribute dont_touch of G10117: signal is true;
	signal G10118: std_logic; attribute dont_touch of G10118: signal is true;
	signal G10119: std_logic; attribute dont_touch of G10119: signal is true;
	signal G10120: std_logic; attribute dont_touch of G10120: signal is true;
	signal G10121: std_logic; attribute dont_touch of G10121: signal is true;
	signal G10122: std_logic; attribute dont_touch of G10122: signal is true;
	signal G10123: std_logic; attribute dont_touch of G10123: signal is true;
	signal G10124: std_logic; attribute dont_touch of G10124: signal is true;
	signal G10125: std_logic; attribute dont_touch of G10125: signal is true;
	signal G10126: std_logic; attribute dont_touch of G10126: signal is true;
	signal G10127: std_logic; attribute dont_touch of G10127: signal is true;
	signal G10130: std_logic; attribute dont_touch of G10130: signal is true;
	signal G10133: std_logic; attribute dont_touch of G10133: signal is true;
	signal G10144: std_logic; attribute dont_touch of G10144: signal is true;
	signal G10145: std_logic; attribute dont_touch of G10145: signal is true;
	signal G10146: std_logic; attribute dont_touch of G10146: signal is true;
	signal G10147: std_logic; attribute dont_touch of G10147: signal is true;
	signal G10150: std_logic; attribute dont_touch of G10150: signal is true;
	signal G10151: std_logic; attribute dont_touch of G10151: signal is true;
	signal G10152: std_logic; attribute dont_touch of G10152: signal is true;
	signal G10153: std_logic; attribute dont_touch of G10153: signal is true;
	signal G10154: std_logic; attribute dont_touch of G10154: signal is true;
	signal G10155: std_logic; attribute dont_touch of G10155: signal is true;
	signal G10156: std_logic; attribute dont_touch of G10156: signal is true;
	signal G10157: std_logic; attribute dont_touch of G10157: signal is true;
	signal G10158: std_logic; attribute dont_touch of G10158: signal is true;
	signal G10161: std_logic; attribute dont_touch of G10161: signal is true;
	signal G10164: std_logic; attribute dont_touch of G10164: signal is true;
	signal G10165: std_logic; attribute dont_touch of G10165: signal is true;
	signal G10166: std_logic; attribute dont_touch of G10166: signal is true;
	signal G10167: std_logic; attribute dont_touch of G10167: signal is true;
	signal G10168: std_logic; attribute dont_touch of G10168: signal is true;
	signal G10169: std_logic; attribute dont_touch of G10169: signal is true;
	signal G10170: std_logic; attribute dont_touch of G10170: signal is true;
	signal G10171: std_logic; attribute dont_touch of G10171: signal is true;
	signal G10172: std_logic; attribute dont_touch of G10172: signal is true;
	signal G10173: std_logic; attribute dont_touch of G10173: signal is true;
	signal G10174: std_logic; attribute dont_touch of G10174: signal is true;
	signal G10175: std_logic; attribute dont_touch of G10175: signal is true;
	signal G10176: std_logic; attribute dont_touch of G10176: signal is true;
	signal G10179: std_logic; attribute dont_touch of G10179: signal is true;
	signal G10182: std_logic; attribute dont_touch of G10182: signal is true;
	signal G10183: std_logic; attribute dont_touch of G10183: signal is true;
	signal G10184: std_logic; attribute dont_touch of G10184: signal is true;
	signal G10185: std_logic; attribute dont_touch of G10185: signal is true;
	signal G10186: std_logic; attribute dont_touch of G10186: signal is true;
	signal G10189: std_logic; attribute dont_touch of G10189: signal is true;
	signal G10192: std_logic; attribute dont_touch of G10192: signal is true;
	signal G10193: std_logic; attribute dont_touch of G10193: signal is true;
	signal G10194: std_logic; attribute dont_touch of G10194: signal is true;
	signal G10195: std_logic; attribute dont_touch of G10195: signal is true;
	signal G10196: std_logic; attribute dont_touch of G10196: signal is true;
	signal G10197: std_logic; attribute dont_touch of G10197: signal is true;
	signal G10198: std_logic; attribute dont_touch of G10198: signal is true;
	signal G10199: std_logic; attribute dont_touch of G10199: signal is true;
	signal G10200: std_logic; attribute dont_touch of G10200: signal is true;
	signal G10201: std_logic; attribute dont_touch of G10201: signal is true;
	signal G10202: std_logic; attribute dont_touch of G10202: signal is true;
	signal G10203: std_logic; attribute dont_touch of G10203: signal is true;
	signal G10204: std_logic; attribute dont_touch of G10204: signal is true;
	signal G10205: std_logic; attribute dont_touch of G10205: signal is true;
	signal G10206: std_logic; attribute dont_touch of G10206: signal is true;
	signal G10207: std_logic; attribute dont_touch of G10207: signal is true;
	signal G10208: std_logic; attribute dont_touch of G10208: signal is true;
	signal G10209: std_logic; attribute dont_touch of G10209: signal is true;
	signal G10210: std_logic; attribute dont_touch of G10210: signal is true;
	signal G10211: std_logic; attribute dont_touch of G10211: signal is true;
	signal G10212: std_logic; attribute dont_touch of G10212: signal is true;
	signal G10213: std_logic; attribute dont_touch of G10213: signal is true;
	signal G10214: std_logic; attribute dont_touch of G10214: signal is true;
	signal G10217: std_logic; attribute dont_touch of G10217: signal is true;
	signal G10218: std_logic; attribute dont_touch of G10218: signal is true;
	signal G10219: std_logic; attribute dont_touch of G10219: signal is true;
	signal G10220: std_logic; attribute dont_touch of G10220: signal is true;
	signal G10221: std_logic; attribute dont_touch of G10221: signal is true;
	signal G10222: std_logic; attribute dont_touch of G10222: signal is true;
	signal G10223: std_logic; attribute dont_touch of G10223: signal is true;
	signal G10224: std_logic; attribute dont_touch of G10224: signal is true;
	signal G10225: std_logic; attribute dont_touch of G10225: signal is true;
	signal G10226: std_logic; attribute dont_touch of G10226: signal is true;
	signal G10227: std_logic; attribute dont_touch of G10227: signal is true;
	signal G10228: std_logic; attribute dont_touch of G10228: signal is true;
	signal G10229: std_logic; attribute dont_touch of G10229: signal is true;
	signal G10230: std_logic; attribute dont_touch of G10230: signal is true;
	signal G10231: std_logic; attribute dont_touch of G10231: signal is true;
	signal G10232: std_logic; attribute dont_touch of G10232: signal is true;
	signal G10235: std_logic; attribute dont_touch of G10235: signal is true;
	signal G10238: std_logic; attribute dont_touch of G10238: signal is true;
	signal G10249: std_logic; attribute dont_touch of G10249: signal is true;
	signal G10250: std_logic; attribute dont_touch of G10250: signal is true;
	signal G10251: std_logic; attribute dont_touch of G10251: signal is true;
	signal G10252: std_logic; attribute dont_touch of G10252: signal is true;
	signal G10255: std_logic; attribute dont_touch of G10255: signal is true;
	signal G10256: std_logic; attribute dont_touch of G10256: signal is true;
	signal G10257: std_logic; attribute dont_touch of G10257: signal is true;
	signal G10258: std_logic; attribute dont_touch of G10258: signal is true;
	signal G10259: std_logic; attribute dont_touch of G10259: signal is true;
	signal G10260: std_logic; attribute dont_touch of G10260: signal is true;
	signal G10261: std_logic; attribute dont_touch of G10261: signal is true;
	signal G10262: std_logic; attribute dont_touch of G10262: signal is true;
	signal G10263: std_logic; attribute dont_touch of G10263: signal is true;
	signal G10266: std_logic; attribute dont_touch of G10266: signal is true;
	signal G10269: std_logic; attribute dont_touch of G10269: signal is true;
	signal G10270: std_logic; attribute dont_touch of G10270: signal is true;
	signal G10271: std_logic; attribute dont_touch of G10271: signal is true;
	signal G10272: std_logic; attribute dont_touch of G10272: signal is true;
	signal G10273: std_logic; attribute dont_touch of G10273: signal is true;
	signal G10276: std_logic; attribute dont_touch of G10276: signal is true;
	signal G10279: std_logic; attribute dont_touch of G10279: signal is true;
	signal G10280: std_logic; attribute dont_touch of G10280: signal is true;
	signal G10281: std_logic; attribute dont_touch of G10281: signal is true;
	signal G10282: std_logic; attribute dont_touch of G10282: signal is true;
	signal G10283: std_logic; attribute dont_touch of G10283: signal is true;
	signal G10284: std_logic; attribute dont_touch of G10284: signal is true;
	signal G10285: std_logic; attribute dont_touch of G10285: signal is true;
	signal G10286: std_logic; attribute dont_touch of G10286: signal is true;
	signal G10287: std_logic; attribute dont_touch of G10287: signal is true;
	signal G10288: std_logic; attribute dont_touch of G10288: signal is true;
	signal G10289: std_logic; attribute dont_touch of G10289: signal is true;
	signal G10290: std_logic; attribute dont_touch of G10290: signal is true;
	signal G10291: std_logic; attribute dont_touch of G10291: signal is true;
	signal G10292: std_logic; attribute dont_touch of G10292: signal is true;
	signal G10293: std_logic; attribute dont_touch of G10293: signal is true;
	signal G10294: std_logic; attribute dont_touch of G10294: signal is true;
	signal G10295: std_logic; attribute dont_touch of G10295: signal is true;
	signal G10296: std_logic; attribute dont_touch of G10296: signal is true;
	signal G10297: std_logic; attribute dont_touch of G10297: signal is true;
	signal G10298: std_logic; attribute dont_touch of G10298: signal is true;
	signal G10299: std_logic; attribute dont_touch of G10299: signal is true;
	signal G10300: std_logic; attribute dont_touch of G10300: signal is true;
	signal G10301: std_logic; attribute dont_touch of G10301: signal is true;
	signal G10302: std_logic; attribute dont_touch of G10302: signal is true;
	signal G10303: std_logic; attribute dont_touch of G10303: signal is true;
	signal G10304: std_logic; attribute dont_touch of G10304: signal is true;
	signal G10305: std_logic; attribute dont_touch of G10305: signal is true;
	signal G10306: std_logic; attribute dont_touch of G10306: signal is true;
	signal G10307: std_logic; attribute dont_touch of G10307: signal is true;
	signal G10308: std_logic; attribute dont_touch of G10308: signal is true;
	signal G10309: std_logic; attribute dont_touch of G10309: signal is true;
	signal G10310: std_logic; attribute dont_touch of G10310: signal is true;
	signal G10311: std_logic; attribute dont_touch of G10311: signal is true;
	signal G10312: std_logic; attribute dont_touch of G10312: signal is true;
	signal G10313: std_logic; attribute dont_touch of G10313: signal is true;
	signal G10314: std_logic; attribute dont_touch of G10314: signal is true;
	signal G10315: std_logic; attribute dont_touch of G10315: signal is true;
	signal G10316: std_logic; attribute dont_touch of G10316: signal is true;
	signal G10319: std_logic; attribute dont_touch of G10319: signal is true;
	signal G10320: std_logic; attribute dont_touch of G10320: signal is true;
	signal G10321: std_logic; attribute dont_touch of G10321: signal is true;
	signal G10322: std_logic; attribute dont_touch of G10322: signal is true;
	signal G10323: std_logic; attribute dont_touch of G10323: signal is true;
	signal G10324: std_logic; attribute dont_touch of G10324: signal is true;
	signal G10325: std_logic; attribute dont_touch of G10325: signal is true;
	signal G10326: std_logic; attribute dont_touch of G10326: signal is true;
	signal G10327: std_logic; attribute dont_touch of G10327: signal is true;
	signal G10328: std_logic; attribute dont_touch of G10328: signal is true;
	signal G10329: std_logic; attribute dont_touch of G10329: signal is true;
	signal G10330: std_logic; attribute dont_touch of G10330: signal is true;
	signal G10331: std_logic; attribute dont_touch of G10331: signal is true;
	signal G10332: std_logic; attribute dont_touch of G10332: signal is true;
	signal G10333: std_logic; attribute dont_touch of G10333: signal is true;
	signal G10334: std_logic; attribute dont_touch of G10334: signal is true;
	signal G10337: std_logic; attribute dont_touch of G10337: signal is true;
	signal G10340: std_logic; attribute dont_touch of G10340: signal is true;
	signal G10351: std_logic; attribute dont_touch of G10351: signal is true;
	signal G10352: std_logic; attribute dont_touch of G10352: signal is true;
	signal G10353: std_logic; attribute dont_touch of G10353: signal is true;
	signal G10354: std_logic; attribute dont_touch of G10354: signal is true;
	signal G10357: std_logic; attribute dont_touch of G10357: signal is true;
	signal G10360: std_logic; attribute dont_touch of G10360: signal is true;
	signal G10361: std_logic; attribute dont_touch of G10361: signal is true;
	signal G10362: std_logic; attribute dont_touch of G10362: signal is true;
	signal G10363: std_logic; attribute dont_touch of G10363: signal is true;
	signal G10364: std_logic; attribute dont_touch of G10364: signal is true;
	signal G10365: std_logic; attribute dont_touch of G10365: signal is true;
	signal G10366: std_logic; attribute dont_touch of G10366: signal is true;
	signal G10367: std_logic; attribute dont_touch of G10367: signal is true;
	signal G10368: std_logic; attribute dont_touch of G10368: signal is true;
	signal G10369: std_logic; attribute dont_touch of G10369: signal is true;
	signal G10370: std_logic; attribute dont_touch of G10370: signal is true;
	signal G10371: std_logic; attribute dont_touch of G10371: signal is true;
	signal G10372: std_logic; attribute dont_touch of G10372: signal is true;
	signal G10373: std_logic; attribute dont_touch of G10373: signal is true;
	signal G10374: std_logic; attribute dont_touch of G10374: signal is true;
	signal G10375: std_logic; attribute dont_touch of G10375: signal is true;
	signal G10376: std_logic; attribute dont_touch of G10376: signal is true;
	signal G10377: std_logic; attribute dont_touch of G10377: signal is true;
	signal G10378: std_logic; attribute dont_touch of G10378: signal is true;
	signal G10379: std_logic; attribute dont_touch of G10379: signal is true;
	signal G10380: std_logic; attribute dont_touch of G10380: signal is true;
	signal G10381: std_logic; attribute dont_touch of G10381: signal is true;
	signal G10382: std_logic; attribute dont_touch of G10382: signal is true;
	signal G10383: std_logic; attribute dont_touch of G10383: signal is true;
	signal G10384: std_logic; attribute dont_touch of G10384: signal is true;
	signal G10385: std_logic; attribute dont_touch of G10385: signal is true;
	signal G10386: std_logic; attribute dont_touch of G10386: signal is true;
	signal G10387: std_logic; attribute dont_touch of G10387: signal is true;
	signal G10388: std_logic; attribute dont_touch of G10388: signal is true;
	signal G10389: std_logic; attribute dont_touch of G10389: signal is true;
	signal G10390: std_logic; attribute dont_touch of G10390: signal is true;
	signal G10391: std_logic; attribute dont_touch of G10391: signal is true;
	signal G10392: std_logic; attribute dont_touch of G10392: signal is true;
	signal G10393: std_logic; attribute dont_touch of G10393: signal is true;
	signal G10394: std_logic; attribute dont_touch of G10394: signal is true;
	signal G10395: std_logic; attribute dont_touch of G10395: signal is true;
	signal G10396: std_logic; attribute dont_touch of G10396: signal is true;
	signal G10397: std_logic; attribute dont_touch of G10397: signal is true;
	signal G10398: std_logic; attribute dont_touch of G10398: signal is true;
	signal G10399: std_logic; attribute dont_touch of G10399: signal is true;
	signal G10400: std_logic; attribute dont_touch of G10400: signal is true;
	signal G10401: std_logic; attribute dont_touch of G10401: signal is true;
	signal G10402: std_logic; attribute dont_touch of G10402: signal is true;
	signal G10403: std_logic; attribute dont_touch of G10403: signal is true;
	signal G10404: std_logic; attribute dont_touch of G10404: signal is true;
	signal G10405: std_logic; attribute dont_touch of G10405: signal is true;
	signal G10406: std_logic; attribute dont_touch of G10406: signal is true;
	signal G10407: std_logic; attribute dont_touch of G10407: signal is true;
	signal G10408: std_logic; attribute dont_touch of G10408: signal is true;
	signal G10409: std_logic; attribute dont_touch of G10409: signal is true;
	signal G10412: std_logic; attribute dont_touch of G10412: signal is true;
	signal G10413: std_logic; attribute dont_touch of G10413: signal is true;
	signal G10414: std_logic; attribute dont_touch of G10414: signal is true;
	signal G10415: std_logic; attribute dont_touch of G10415: signal is true;
	signal G10416: std_logic; attribute dont_touch of G10416: signal is true;
	signal G10419: std_logic; attribute dont_touch of G10419: signal is true;
	signal G10422: std_logic; attribute dont_touch of G10422: signal is true;
	signal G10423: std_logic; attribute dont_touch of G10423: signal is true;
	signal G10424: std_logic; attribute dont_touch of G10424: signal is true;
	signal G10430: std_logic; attribute dont_touch of G10430: signal is true;
	signal G10431: std_logic; attribute dont_touch of G10431: signal is true;
	signal G10432: std_logic; attribute dont_touch of G10432: signal is true;
	signal G10433: std_logic; attribute dont_touch of G10433: signal is true;
	signal G10434: std_logic; attribute dont_touch of G10434: signal is true;
	signal G10435: std_logic; attribute dont_touch of G10435: signal is true;
	signal G10436: std_logic; attribute dont_touch of G10436: signal is true;
	signal G10437: std_logic; attribute dont_touch of G10437: signal is true;
	signal G10438: std_logic; attribute dont_touch of G10438: signal is true;
	signal G10439: std_logic; attribute dont_touch of G10439: signal is true;
	signal G10440: std_logic; attribute dont_touch of G10440: signal is true;
	signal G10441: std_logic; attribute dont_touch of G10441: signal is true;
	signal G10442: std_logic; attribute dont_touch of G10442: signal is true;
	signal G10443: std_logic; attribute dont_touch of G10443: signal is true;
	signal G10444: std_logic; attribute dont_touch of G10444: signal is true;
	signal G10445: std_logic; attribute dont_touch of G10445: signal is true;
	signal G10446: std_logic; attribute dont_touch of G10446: signal is true;
	signal G10447: std_logic; attribute dont_touch of G10447: signal is true;
	signal G10448: std_logic; attribute dont_touch of G10448: signal is true;
	signal G10449: std_logic; attribute dont_touch of G10449: signal is true;
	signal G10450: std_logic; attribute dont_touch of G10450: signal is true;
	signal G10451: std_logic; attribute dont_touch of G10451: signal is true;
	signal G10452: std_logic; attribute dont_touch of G10452: signal is true;
	signal G10453: std_logic; attribute dont_touch of G10453: signal is true;
	signal G10454: std_logic; attribute dont_touch of G10454: signal is true;
	signal G10455: std_logic; attribute dont_touch of G10455: signal is true;
	signal G10456: std_logic; attribute dont_touch of G10456: signal is true;
	signal G10457: std_logic; attribute dont_touch of G10457: signal is true;
	signal G10458: std_logic; attribute dont_touch of G10458: signal is true;
	signal G10459: std_logic; attribute dont_touch of G10459: signal is true;
	signal G10460: std_logic; attribute dont_touch of G10460: signal is true;
	signal G10461: std_logic; attribute dont_touch of G10461: signal is true;
	signal G10462: std_logic; attribute dont_touch of G10462: signal is true;
	signal G10463: std_logic; attribute dont_touch of G10463: signal is true;
	signal G10464: std_logic; attribute dont_touch of G10464: signal is true;
	signal G10465: std_logic; attribute dont_touch of G10465: signal is true;
	signal G10466: std_logic; attribute dont_touch of G10466: signal is true;
	signal G10467: std_logic; attribute dont_touch of G10467: signal is true;
	signal G10468: std_logic; attribute dont_touch of G10468: signal is true;
	signal G10469: std_logic; attribute dont_touch of G10469: signal is true;
	signal G10470: std_logic; attribute dont_touch of G10470: signal is true;
	signal G10471: std_logic; attribute dont_touch of G10471: signal is true;
	signal G10472: std_logic; attribute dont_touch of G10472: signal is true;
	signal G10473: std_logic; attribute dont_touch of G10473: signal is true;
	signal G10474: std_logic; attribute dont_touch of G10474: signal is true;
	signal G10475: std_logic; attribute dont_touch of G10475: signal is true;
	signal G10476: std_logic; attribute dont_touch of G10476: signal is true;
	signal G10477: std_logic; attribute dont_touch of G10477: signal is true;
	signal G10478: std_logic; attribute dont_touch of G10478: signal is true;
	signal G10479: std_logic; attribute dont_touch of G10479: signal is true;
	signal G10480: std_logic; attribute dont_touch of G10480: signal is true;
	signal G10481: std_logic; attribute dont_touch of G10481: signal is true;
	signal G10482: std_logic; attribute dont_touch of G10482: signal is true;
	signal G10485: std_logic; attribute dont_touch of G10485: signal is true;
	signal G10486: std_logic; attribute dont_touch of G10486: signal is true;
	signal G10492: std_logic; attribute dont_touch of G10492: signal is true;
	signal G10493: std_logic; attribute dont_touch of G10493: signal is true;
	signal G10494: std_logic; attribute dont_touch of G10494: signal is true;
	signal G10495: std_logic; attribute dont_touch of G10495: signal is true;
	signal G10496: std_logic; attribute dont_touch of G10496: signal is true;
	signal G10497: std_logic; attribute dont_touch of G10497: signal is true;
	signal G10498: std_logic; attribute dont_touch of G10498: signal is true;
	signal G10499: std_logic; attribute dont_touch of G10499: signal is true;
	signal G10500: std_logic; attribute dont_touch of G10500: signal is true;
	signal G10506: std_logic; attribute dont_touch of G10506: signal is true;
	signal G10507: std_logic; attribute dont_touch of G10507: signal is true;
	signal G10508: std_logic; attribute dont_touch of G10508: signal is true;
	signal G10509: std_logic; attribute dont_touch of G10509: signal is true;
	signal G10510: std_logic; attribute dont_touch of G10510: signal is true;
	signal G10511: std_logic; attribute dont_touch of G10511: signal is true;
	signal G10512: std_logic; attribute dont_touch of G10512: signal is true;
	signal G10513: std_logic; attribute dont_touch of G10513: signal is true;
	signal G10514: std_logic; attribute dont_touch of G10514: signal is true;
	signal G10515: std_logic; attribute dont_touch of G10515: signal is true;
	signal G10516: std_logic; attribute dont_touch of G10516: signal is true;
	signal G10517: std_logic; attribute dont_touch of G10517: signal is true;
	signal G10518: std_logic; attribute dont_touch of G10518: signal is true;
	signal G10519: std_logic; attribute dont_touch of G10519: signal is true;
	signal G10520: std_logic; attribute dont_touch of G10520: signal is true;
	signal G10521: std_logic; attribute dont_touch of G10521: signal is true;
	signal G10522: std_logic; attribute dont_touch of G10522: signal is true;
	signal G10523: std_logic; attribute dont_touch of G10523: signal is true;
	signal G10524: std_logic; attribute dont_touch of G10524: signal is true;
	signal G10525: std_logic; attribute dont_touch of G10525: signal is true;
	signal G10526: std_logic; attribute dont_touch of G10526: signal is true;
	signal G10527: std_logic; attribute dont_touch of G10527: signal is true;
	signal G10528: std_logic; attribute dont_touch of G10528: signal is true;
	signal G10529: std_logic; attribute dont_touch of G10529: signal is true;
	signal G10530: std_logic; attribute dont_touch of G10530: signal is true;
	signal G10531: std_logic; attribute dont_touch of G10531: signal is true;
	signal G10532: std_logic; attribute dont_touch of G10532: signal is true;
	signal G10533: std_logic; attribute dont_touch of G10533: signal is true;
	signal G10534: std_logic; attribute dont_touch of G10534: signal is true;
	signal G10535: std_logic; attribute dont_touch of G10535: signal is true;
	signal G10536: std_logic; attribute dont_touch of G10536: signal is true;
	signal G10537: std_logic; attribute dont_touch of G10537: signal is true;
	signal G10538: std_logic; attribute dont_touch of G10538: signal is true;
	signal G10539: std_logic; attribute dont_touch of G10539: signal is true;
	signal G10540: std_logic; attribute dont_touch of G10540: signal is true;
	signal G10541: std_logic; attribute dont_touch of G10541: signal is true;
	signal G10542: std_logic; attribute dont_touch of G10542: signal is true;
	signal G10545: std_logic; attribute dont_touch of G10545: signal is true;
	signal G10548: std_logic; attribute dont_touch of G10548: signal is true;
	signal G10549: std_logic; attribute dont_touch of G10549: signal is true;
	signal G10555: std_logic; attribute dont_touch of G10555: signal is true;
	signal G10556: std_logic; attribute dont_touch of G10556: signal is true;
	signal G10557: std_logic; attribute dont_touch of G10557: signal is true;
	signal G10558: std_logic; attribute dont_touch of G10558: signal is true;
	signal G10559: std_logic; attribute dont_touch of G10559: signal is true;
	signal G10560: std_logic; attribute dont_touch of G10560: signal is true;
	signal G10566: std_logic; attribute dont_touch of G10566: signal is true;
	signal G10567: std_logic; attribute dont_touch of G10567: signal is true;
	signal G10568: std_logic; attribute dont_touch of G10568: signal is true;
	signal G10569: std_logic; attribute dont_touch of G10569: signal is true;
	signal G10570: std_logic; attribute dont_touch of G10570: signal is true;
	signal G10571: std_logic; attribute dont_touch of G10571: signal is true;
	signal G10572: std_logic; attribute dont_touch of G10572: signal is true;
	signal G10573: std_logic; attribute dont_touch of G10573: signal is true;
	signal G10574: std_logic; attribute dont_touch of G10574: signal is true;
	signal G10580: std_logic; attribute dont_touch of G10580: signal is true;
	signal G10581: std_logic; attribute dont_touch of G10581: signal is true;
	signal G10582: std_logic; attribute dont_touch of G10582: signal is true;
	signal G10583: std_logic; attribute dont_touch of G10583: signal is true;
	signal G10584: std_logic; attribute dont_touch of G10584: signal is true;
	signal G10585: std_logic; attribute dont_touch of G10585: signal is true;
	signal G10586: std_logic; attribute dont_touch of G10586: signal is true;
	signal G10587: std_logic; attribute dont_touch of G10587: signal is true;
	signal G10588: std_logic; attribute dont_touch of G10588: signal is true;
	signal G10589: std_logic; attribute dont_touch of G10589: signal is true;
	signal G10590: std_logic; attribute dont_touch of G10590: signal is true;
	signal G10591: std_logic; attribute dont_touch of G10591: signal is true;
	signal G10592: std_logic; attribute dont_touch of G10592: signal is true;
	signal G10593: std_logic; attribute dont_touch of G10593: signal is true;
	signal G10594: std_logic; attribute dont_touch of G10594: signal is true;
	signal G10595: std_logic; attribute dont_touch of G10595: signal is true;
	signal G10596: std_logic; attribute dont_touch of G10596: signal is true;
	signal G10597: std_logic; attribute dont_touch of G10597: signal is true;
	signal G10598: std_logic; attribute dont_touch of G10598: signal is true;
	signal G10599: std_logic; attribute dont_touch of G10599: signal is true;
	signal G10600: std_logic; attribute dont_touch of G10600: signal is true;
	signal G10601: std_logic; attribute dont_touch of G10601: signal is true;
	signal G10604: std_logic; attribute dont_touch of G10604: signal is true;
	signal G10605: std_logic; attribute dont_touch of G10605: signal is true;
	signal G10606: std_logic; attribute dont_touch of G10606: signal is true;
	signal G10612: std_logic; attribute dont_touch of G10612: signal is true;
	signal G10613: std_logic; attribute dont_touch of G10613: signal is true;
	signal G10614: std_logic; attribute dont_touch of G10614: signal is true;
	signal G10615: std_logic; attribute dont_touch of G10615: signal is true;
	signal G10616: std_logic; attribute dont_touch of G10616: signal is true;
	signal G10617: std_logic; attribute dont_touch of G10617: signal is true;
	signal G10623: std_logic; attribute dont_touch of G10623: signal is true;
	signal G10624: std_logic; attribute dont_touch of G10624: signal is true;
	signal G10625: std_logic; attribute dont_touch of G10625: signal is true;
	signal G10626: std_logic; attribute dont_touch of G10626: signal is true;
	signal G10627: std_logic; attribute dont_touch of G10627: signal is true;
	signal G10628: std_logic; attribute dont_touch of G10628: signal is true;
	signal G10629: std_logic; attribute dont_touch of G10629: signal is true;
	signal G10630: std_logic; attribute dont_touch of G10630: signal is true;
	signal G10631: std_logic; attribute dont_touch of G10631: signal is true;
	signal G10637: std_logic; attribute dont_touch of G10637: signal is true;
	signal G10638: std_logic; attribute dont_touch of G10638: signal is true;
	signal G10639: std_logic; attribute dont_touch of G10639: signal is true;
	signal G10640: std_logic; attribute dont_touch of G10640: signal is true;
	signal G10641: std_logic; attribute dont_touch of G10641: signal is true;
	signal G10642: std_logic; attribute dont_touch of G10642: signal is true;
	signal G10643: std_logic; attribute dont_touch of G10643: signal is true;
	signal G10644: std_logic; attribute dont_touch of G10644: signal is true;
	signal G10645: std_logic; attribute dont_touch of G10645: signal is true;
	signal G10646: std_logic; attribute dont_touch of G10646: signal is true;
	signal G10649: std_logic; attribute dont_touch of G10649: signal is true;
	signal G10650: std_logic; attribute dont_touch of G10650: signal is true;
	signal G10651: std_logic; attribute dont_touch of G10651: signal is true;
	signal G10652: std_logic; attribute dont_touch of G10652: signal is true;
	signal G10653: std_logic; attribute dont_touch of G10653: signal is true;
	signal G10659: std_logic; attribute dont_touch of G10659: signal is true;
	signal G10660: std_logic; attribute dont_touch of G10660: signal is true;
	signal G10661: std_logic; attribute dont_touch of G10661: signal is true;
	signal G10662: std_logic; attribute dont_touch of G10662: signal is true;
	signal G10663: std_logic; attribute dont_touch of G10663: signal is true;
	signal G10664: std_logic; attribute dont_touch of G10664: signal is true;
	signal G10670: std_logic; attribute dont_touch of G10670: signal is true;
	signal G10671: std_logic; attribute dont_touch of G10671: signal is true;
	signal G10672: std_logic; attribute dont_touch of G10672: signal is true;
	signal G10673: std_logic; attribute dont_touch of G10673: signal is true;
	signal G10674: std_logic; attribute dont_touch of G10674: signal is true;
	signal G10675: std_logic; attribute dont_touch of G10675: signal is true;
	signal G10676: std_logic; attribute dont_touch of G10676: signal is true;
	signal G10677: std_logic; attribute dont_touch of G10677: signal is true;
	signal G10678: std_logic; attribute dont_touch of G10678: signal is true;
	signal G10679: std_logic; attribute dont_touch of G10679: signal is true;
	signal G10680: std_logic; attribute dont_touch of G10680: signal is true;
	signal G10681: std_logic; attribute dont_touch of G10681: signal is true;
	signal G10682: std_logic; attribute dont_touch of G10682: signal is true;
	signal G10683: std_logic; attribute dont_touch of G10683: signal is true;
	signal G10689: std_logic; attribute dont_touch of G10689: signal is true;
	signal G10690: std_logic; attribute dont_touch of G10690: signal is true;
	signal G10691: std_logic; attribute dont_touch of G10691: signal is true;
	signal G10692: std_logic; attribute dont_touch of G10692: signal is true;
	signal G10693: std_logic; attribute dont_touch of G10693: signal is true;
	signal G10694: std_logic; attribute dont_touch of G10694: signal is true;
	signal G10703: std_logic; attribute dont_touch of G10703: signal is true;
	signal G10704: std_logic; attribute dont_touch of G10704: signal is true;
	signal G10705: std_logic; attribute dont_touch of G10705: signal is true;
	signal G10706: std_logic; attribute dont_touch of G10706: signal is true;
	signal G10707: std_logic; attribute dont_touch of G10707: signal is true;
	signal G10708: std_logic; attribute dont_touch of G10708: signal is true;
	signal G10709: std_logic; attribute dont_touch of G10709: signal is true;
	signal G10710: std_logic; attribute dont_touch of G10710: signal is true;
	signal G10711: std_logic; attribute dont_touch of G10711: signal is true;
	signal G10714: std_logic; attribute dont_touch of G10714: signal is true;
	signal G10723: std_logic; attribute dont_touch of G10723: signal is true;
	signal G10724: std_logic; attribute dont_touch of G10724: signal is true;
	signal G10725: std_logic; attribute dont_touch of G10725: signal is true;
	signal G10726: std_logic; attribute dont_touch of G10726: signal is true;
	signal G10727: std_logic; attribute dont_touch of G10727: signal is true;
	signal G10728: std_logic; attribute dont_touch of G10728: signal is true;
	signal G10729: std_logic; attribute dont_touch of G10729: signal is true;
	signal G10730: std_logic; attribute dont_touch of G10730: signal is true;
	signal G10735: std_logic; attribute dont_touch of G10735: signal is true;
	signal G10744: std_logic; attribute dont_touch of G10744: signal is true;
	signal G10745: std_logic; attribute dont_touch of G10745: signal is true;
	signal G10746: std_logic; attribute dont_touch of G10746: signal is true;
	signal G10747: std_logic; attribute dont_touch of G10747: signal is true;
	signal G10748: std_logic; attribute dont_touch of G10748: signal is true;
	signal G10749: std_logic; attribute dont_touch of G10749: signal is true;
	signal G10754: std_logic; attribute dont_touch of G10754: signal is true;
	signal G10763: std_logic; attribute dont_touch of G10763: signal is true;
	signal G10764: std_logic; attribute dont_touch of G10764: signal is true;
	signal G10765: std_logic; attribute dont_touch of G10765: signal is true;
	signal G10766: std_logic; attribute dont_touch of G10766: signal is true;
	signal G10767: std_logic; attribute dont_touch of G10767: signal is true;
	signal G10772: std_logic; attribute dont_touch of G10772: signal is true;
	signal G10773: std_logic; attribute dont_touch of G10773: signal is true;
	signal G10778: std_logic; attribute dont_touch of G10778: signal is true;
	signal G10779: std_logic; attribute dont_touch of G10779: signal is true;
	signal G10783: std_logic; attribute dont_touch of G10783: signal is true;
	signal G10784: std_logic; attribute dont_touch of G10784: signal is true;
	signal G10787: std_logic; attribute dont_touch of G10787: signal is true;
	signal G10788: std_logic; attribute dont_touch of G10788: signal is true;
	signal G10789: std_logic; attribute dont_touch of G10789: signal is true;
	signal G10792: std_logic; attribute dont_touch of G10792: signal is true;
	signal G10793: std_logic; attribute dont_touch of G10793: signal is true;
	signal G10796: std_logic; attribute dont_touch of G10796: signal is true;
	signal G10797: std_logic; attribute dont_touch of G10797: signal is true;
	signal G10800: std_logic; attribute dont_touch of G10800: signal is true;
	signal G10801: std_logic; attribute dont_touch of G10801: signal is true;
	signal G10804: std_logic; attribute dont_touch of G10804: signal is true;
	signal G10805: std_logic; attribute dont_touch of G10805: signal is true;
	signal G10808: std_logic; attribute dont_touch of G10808: signal is true;
	signal G10809: std_logic; attribute dont_touch of G10809: signal is true;
	signal G10810: std_logic; attribute dont_touch of G10810: signal is true;
	signal G10813: std_logic; attribute dont_touch of G10813: signal is true;
	signal G10814: std_logic; attribute dont_touch of G10814: signal is true;
	signal G10817: std_logic; attribute dont_touch of G10817: signal is true;
	signal G10818: std_logic; attribute dont_touch of G10818: signal is true;
	signal G10821: std_logic; attribute dont_touch of G10821: signal is true;
	signal G10822: std_logic; attribute dont_touch of G10822: signal is true;
	signal G10825: std_logic; attribute dont_touch of G10825: signal is true;
	signal G10826: std_logic; attribute dont_touch of G10826: signal is true;
	signal G10829: std_logic; attribute dont_touch of G10829: signal is true;
	signal G10830: std_logic; attribute dont_touch of G10830: signal is true;
	signal G10831: std_logic; attribute dont_touch of G10831: signal is true;
	signal G10834: std_logic; attribute dont_touch of G10834: signal is true;
	signal G10835: std_logic; attribute dont_touch of G10835: signal is true;
	signal G10838: std_logic; attribute dont_touch of G10838: signal is true;
	signal G10839: std_logic; attribute dont_touch of G10839: signal is true;
	signal G10842: std_logic; attribute dont_touch of G10842: signal is true;
	signal G10843: std_logic; attribute dont_touch of G10843: signal is true;
	signal G10846: std_logic; attribute dont_touch of G10846: signal is true;
	signal G10847: std_logic; attribute dont_touch of G10847: signal is true;
	signal G10848: std_logic; attribute dont_touch of G10848: signal is true;
	signal G10849: std_logic; attribute dont_touch of G10849: signal is true;
	signal G10850: std_logic; attribute dont_touch of G10850: signal is true;
	signal G10851: std_logic; attribute dont_touch of G10851: signal is true;
	signal G10854: std_logic; attribute dont_touch of G10854: signal is true;
	signal G10855: std_logic; attribute dont_touch of G10855: signal is true;
	signal G10858: std_logic; attribute dont_touch of G10858: signal is true;
	signal G10859: std_logic; attribute dont_touch of G10859: signal is true;
	signal G10862: std_logic; attribute dont_touch of G10862: signal is true;
	signal G10865: std_logic; attribute dont_touch of G10865: signal is true;
	signal G10866: std_logic; attribute dont_touch of G10866: signal is true;
	signal G10867: std_logic; attribute dont_touch of G10867: signal is true;
	signal G10868: std_logic; attribute dont_touch of G10868: signal is true;
	signal G10869: std_logic; attribute dont_touch of G10869: signal is true;
	signal G10870: std_logic; attribute dont_touch of G10870: signal is true;
	signal G10871: std_logic; attribute dont_touch of G10871: signal is true;
	signal G10872: std_logic; attribute dont_touch of G10872: signal is true;
	signal G10875: std_logic; attribute dont_touch of G10875: signal is true;
	signal G10876: std_logic; attribute dont_touch of G10876: signal is true;
	signal G10877: std_logic; attribute dont_touch of G10877: signal is true;
	signal G10880: std_logic; attribute dont_touch of G10880: signal is true;
	signal G10883: std_logic; attribute dont_touch of G10883: signal is true;
	signal G10886: std_logic; attribute dont_touch of G10886: signal is true;
	signal G10887: std_logic; attribute dont_touch of G10887: signal is true;
	signal G10888: std_logic; attribute dont_touch of G10888: signal is true;
	signal G10889: std_logic; attribute dont_touch of G10889: signal is true;
	signal G10890: std_logic; attribute dont_touch of G10890: signal is true;
	signal G10891: std_logic; attribute dont_touch of G10891: signal is true;
	signal G10892: std_logic; attribute dont_touch of G10892: signal is true;
	signal G10895: std_logic; attribute dont_touch of G10895: signal is true;
	signal G10898: std_logic; attribute dont_touch of G10898: signal is true;
	signal G10901: std_logic; attribute dont_touch of G10901: signal is true;
	signal G10904: std_logic; attribute dont_touch of G10904: signal is true;
	signal G10905: std_logic; attribute dont_touch of G10905: signal is true;
	signal G10906: std_logic; attribute dont_touch of G10906: signal is true;
	signal G10907: std_logic; attribute dont_touch of G10907: signal is true;
	signal G10908: std_logic; attribute dont_touch of G10908: signal is true;
	signal G10909: std_logic; attribute dont_touch of G10909: signal is true;
	signal G10910: std_logic; attribute dont_touch of G10910: signal is true;
	signal G10911: std_logic; attribute dont_touch of G10911: signal is true;
	signal G10912: std_logic; attribute dont_touch of G10912: signal is true;
	signal G10915: std_logic; attribute dont_touch of G10915: signal is true;
	signal G10918: std_logic; attribute dont_touch of G10918: signal is true;
	signal G10921: std_logic; attribute dont_touch of G10921: signal is true;
	signal G10924: std_logic; attribute dont_touch of G10924: signal is true;
	signal G10927: std_logic; attribute dont_touch of G10927: signal is true;
	signal G10928: std_logic; attribute dont_touch of G10928: signal is true;
	signal G10929: std_logic; attribute dont_touch of G10929: signal is true;
	signal G10930: std_logic; attribute dont_touch of G10930: signal is true;
	signal G10931: std_logic; attribute dont_touch of G10931: signal is true;
	signal G10932: std_logic; attribute dont_touch of G10932: signal is true;
	signal G10933: std_logic; attribute dont_touch of G10933: signal is true;
	signal G10934: std_logic; attribute dont_touch of G10934: signal is true;
	signal G10935: std_logic; attribute dont_touch of G10935: signal is true;
	signal G10936: std_logic; attribute dont_touch of G10936: signal is true;
	signal G10937: std_logic; attribute dont_touch of G10937: signal is true;
	signal G10940: std_logic; attribute dont_touch of G10940: signal is true;
	signal G10943: std_logic; attribute dont_touch of G10943: signal is true;
	signal G10946: std_logic; attribute dont_touch of G10946: signal is true;
	signal G10949: std_logic; attribute dont_touch of G10949: signal is true;
	signal G10952: std_logic; attribute dont_touch of G10952: signal is true;
	signal G10961: std_logic; attribute dont_touch of G10961: signal is true;
	signal G10962: std_logic; attribute dont_touch of G10962: signal is true;
	signal G10963: std_logic; attribute dont_touch of G10963: signal is true;
	signal G10966: std_logic; attribute dont_touch of G10966: signal is true;
	signal G10967: std_logic; attribute dont_touch of G10967: signal is true;
	signal G10968: std_logic; attribute dont_touch of G10968: signal is true;
	signal G10969: std_logic; attribute dont_touch of G10969: signal is true;
	signal G10972: std_logic; attribute dont_touch of G10972: signal is true;
	signal G10973: std_logic; attribute dont_touch of G10973: signal is true;
	signal G10974: std_logic; attribute dont_touch of G10974: signal is true;
	signal G10977: std_logic; attribute dont_touch of G10977: signal is true;
	signal G10980: std_logic; attribute dont_touch of G10980: signal is true;
	signal G10983: std_logic; attribute dont_touch of G10983: signal is true;
	signal G10986: std_logic; attribute dont_touch of G10986: signal is true;
	signal G10987: std_logic; attribute dont_touch of G10987: signal is true;
	signal G10988: std_logic; attribute dont_touch of G10988: signal is true;
	signal G10991: std_logic; attribute dont_touch of G10991: signal is true;
	signal G10994: std_logic; attribute dont_touch of G10994: signal is true;
	signal G10995: std_logic; attribute dont_touch of G10995: signal is true;
	signal G10996: std_logic; attribute dont_touch of G10996: signal is true;
	signal G10999: std_logic; attribute dont_touch of G10999: signal is true;
	signal G11002: std_logic; attribute dont_touch of G11002: signal is true;
	signal G11003: std_logic; attribute dont_touch of G11003: signal is true;
	signal G11004: std_logic; attribute dont_touch of G11004: signal is true;
	signal G11007: std_logic; attribute dont_touch of G11007: signal is true;
	signal G11008: std_logic; attribute dont_touch of G11008: signal is true;
	signal G11011: std_logic; attribute dont_touch of G11011: signal is true;
	signal G11014: std_logic; attribute dont_touch of G11014: signal is true;
	signal G11017: std_logic; attribute dont_touch of G11017: signal is true;
	signal G11020: std_logic; attribute dont_touch of G11020: signal is true;
	signal G11021: std_logic; attribute dont_touch of G11021: signal is true;
	signal G11022: std_logic; attribute dont_touch of G11022: signal is true;
	signal G11025: std_logic; attribute dont_touch of G11025: signal is true;
	signal G11028: std_logic; attribute dont_touch of G11028: signal is true;
	signal G11031: std_logic; attribute dont_touch of G11031: signal is true;
	signal G11032: std_logic; attribute dont_touch of G11032: signal is true;
	signal G11035: std_logic; attribute dont_touch of G11035: signal is true;
	signal G11036: std_logic; attribute dont_touch of G11036: signal is true;
	signal G11039: std_logic; attribute dont_touch of G11039: signal is true;
	signal G11042: std_logic; attribute dont_touch of G11042: signal is true;
	signal G11045: std_logic; attribute dont_touch of G11045: signal is true;
	signal G11048: std_logic; attribute dont_touch of G11048: signal is true;
	signal G11051: std_logic; attribute dont_touch of G11051: signal is true;
	signal G11054: std_logic; attribute dont_touch of G11054: signal is true;
	signal G11055: std_logic; attribute dont_touch of G11055: signal is true;
	signal G11056: std_logic; attribute dont_touch of G11056: signal is true;
	signal G11059: std_logic; attribute dont_touch of G11059: signal is true;
	signal G11063: std_logic; attribute dont_touch of G11063: signal is true;
	signal G11066: std_logic; attribute dont_touch of G11066: signal is true;
	signal G11069: std_logic; attribute dont_touch of G11069: signal is true;
	signal G11078: std_logic; attribute dont_touch of G11078: signal is true;
	signal G11079: std_logic; attribute dont_touch of G11079: signal is true;
	signal G11082: std_logic; attribute dont_touch of G11082: signal is true;
	signal G11085: std_logic; attribute dont_touch of G11085: signal is true;
	signal G11088: std_logic; attribute dont_touch of G11088: signal is true;
	signal G11091: std_logic; attribute dont_touch of G11091: signal is true;
	signal G11092: std_logic; attribute dont_touch of G11092: signal is true;
	signal G11095: std_logic; attribute dont_touch of G11095: signal is true;
	signal G11098: std_logic; attribute dont_touch of G11098: signal is true;
	signal G11101: std_logic; attribute dont_touch of G11101: signal is true;
	signal G11102: std_logic; attribute dont_touch of G11102: signal is true;
	signal G11105: std_logic; attribute dont_touch of G11105: signal is true;
	signal G11108: std_logic; attribute dont_touch of G11108: signal is true;
	signal G11111: std_logic; attribute dont_touch of G11111: signal is true;
	signal G11114: std_logic; attribute dont_touch of G11114: signal is true;
	signal G11117: std_logic; attribute dont_touch of G11117: signal is true;
	signal G11120: std_logic; attribute dont_touch of G11120: signal is true;
	signal G11123: std_logic; attribute dont_touch of G11123: signal is true;
	signal G11126: std_logic; attribute dont_touch of G11126: signal is true;
	signal G11129: std_logic; attribute dont_touch of G11129: signal is true;
	signal G11132: std_logic; attribute dont_touch of G11132: signal is true;
	signal G11135: std_logic; attribute dont_touch of G11135: signal is true;
	signal G11138: std_logic; attribute dont_touch of G11138: signal is true;
	signal G11141: std_logic; attribute dont_touch of G11141: signal is true;
	signal G11144: std_logic; attribute dont_touch of G11144: signal is true;
	signal G11145: std_logic; attribute dont_touch of G11145: signal is true;
	signal G11148: std_logic; attribute dont_touch of G11148: signal is true;
	signal G11151: std_logic; attribute dont_touch of G11151: signal is true;
	signal G11154: std_logic; attribute dont_touch of G11154: signal is true;
	signal G11157: std_logic; attribute dont_touch of G11157: signal is true;
	signal G11160: std_logic; attribute dont_touch of G11160: signal is true;
	signal G11163: std_logic; attribute dont_touch of G11163: signal is true;
	signal G11166: std_logic; attribute dont_touch of G11166: signal is true;
	signal G11169: std_logic; attribute dont_touch of G11169: signal is true;
	signal G11170: std_logic; attribute dont_touch of G11170: signal is true;
	signal G11173: std_logic; attribute dont_touch of G11173: signal is true;
	signal G11176: std_logic; attribute dont_touch of G11176: signal is true;
	signal G11179: std_logic; attribute dont_touch of G11179: signal is true;
	signal G11182: std_logic; attribute dont_touch of G11182: signal is true;
	signal G11185: std_logic; attribute dont_touch of G11185: signal is true;
	signal G11188: std_logic; attribute dont_touch of G11188: signal is true;
	signal G11189: std_logic; attribute dont_touch of G11189: signal is true;
	signal G11190: std_logic; attribute dont_touch of G11190: signal is true;
	signal G11199: std_logic; attribute dont_touch of G11199: signal is true;
	signal G11202: std_logic; attribute dont_touch of G11202: signal is true;
	signal G11205: std_logic; attribute dont_touch of G11205: signal is true;
	signal G11208: std_logic; attribute dont_touch of G11208: signal is true;
	signal G11209: std_logic; attribute dont_touch of G11209: signal is true;
	signal G11210: std_logic; attribute dont_touch of G11210: signal is true;
	signal G11213: std_logic; attribute dont_touch of G11213: signal is true;
	signal G11216: std_logic; attribute dont_touch of G11216: signal is true;
	signal G11219: std_logic; attribute dont_touch of G11219: signal is true;
	signal G11222: std_logic; attribute dont_touch of G11222: signal is true;
	signal G11225: std_logic; attribute dont_touch of G11225: signal is true;
	signal G11228: std_logic; attribute dont_touch of G11228: signal is true;
	signal G11231: std_logic; attribute dont_touch of G11231: signal is true;
	signal G11234: std_logic; attribute dont_touch of G11234: signal is true;
	signal G11237: std_logic; attribute dont_touch of G11237: signal is true;
	signal G11240: std_logic; attribute dont_touch of G11240: signal is true;
	signal G11243: std_logic; attribute dont_touch of G11243: signal is true;
	signal G11246: std_logic; attribute dont_touch of G11246: signal is true;
	signal G11249: std_logic; attribute dont_touch of G11249: signal is true;
	signal G11252: std_logic; attribute dont_touch of G11252: signal is true;
	signal G11255: std_logic; attribute dont_touch of G11255: signal is true;
	signal G11256: std_logic; attribute dont_touch of G11256: signal is true;
	signal G11259: std_logic; attribute dont_touch of G11259: signal is true;
	signal G11262: std_logic; attribute dont_touch of G11262: signal is true;
	signal G11263: std_logic; attribute dont_touch of G11263: signal is true;
	signal G11264: std_logic; attribute dont_touch of G11264: signal is true;
	signal G11265: std_logic; attribute dont_touch of G11265: signal is true;
	signal G11268: std_logic; attribute dont_touch of G11268: signal is true;
	signal G11271: std_logic; attribute dont_touch of G11271: signal is true;
	signal G11274: std_logic; attribute dont_touch of G11274: signal is true;
	signal G11277: std_logic; attribute dont_touch of G11277: signal is true;
	signal G11278: std_logic; attribute dont_touch of G11278: signal is true;
	signal G11281: std_logic; attribute dont_touch of G11281: signal is true;
	signal G11284: std_logic; attribute dont_touch of G11284: signal is true;
	signal G11287: std_logic; attribute dont_touch of G11287: signal is true;
	signal G11290: std_logic; attribute dont_touch of G11290: signal is true;
	signal G11291: std_logic; attribute dont_touch of G11291: signal is true;
	signal G11294: std_logic; attribute dont_touch of G11294: signal is true;
	signal G11297: std_logic; attribute dont_touch of G11297: signal is true;
	signal G11300: std_logic; attribute dont_touch of G11300: signal is true;
	signal G11303: std_logic; attribute dont_touch of G11303: signal is true;
	signal G11306: std_logic; attribute dont_touch of G11306: signal is true;
	signal G11309: std_logic; attribute dont_touch of G11309: signal is true;
	signal G11312: std_logic; attribute dont_touch of G11312: signal is true;
	signal G11315: std_logic; attribute dont_touch of G11315: signal is true;
	signal G11318: std_logic; attribute dont_touch of G11318: signal is true;
	signal G11321: std_logic; attribute dont_touch of G11321: signal is true;
	signal G11324: std_logic; attribute dont_touch of G11324: signal is true;
	signal G11327: std_logic; attribute dont_touch of G11327: signal is true;
	signal G11330: std_logic; attribute dont_touch of G11330: signal is true;
	signal G11331: std_logic; attribute dont_touch of G11331: signal is true;
	signal G11332: std_logic; attribute dont_touch of G11332: signal is true;
	signal G11341: std_logic; attribute dont_touch of G11341: signal is true;
	signal G11344: std_logic; attribute dont_touch of G11344: signal is true;
	signal G11347: std_logic; attribute dont_touch of G11347: signal is true;
	signal G11348: std_logic; attribute dont_touch of G11348: signal is true;
	signal G11351: std_logic; attribute dont_touch of G11351: signal is true;
	signal G11354: std_logic; attribute dont_touch of G11354: signal is true;
	signal G11355: std_logic; attribute dont_touch of G11355: signal is true;
	signal G11358: std_logic; attribute dont_touch of G11358: signal is true;
	signal G11361: std_logic; attribute dont_touch of G11361: signal is true;
	signal G11364: std_logic; attribute dont_touch of G11364: signal is true;
	signal G11367: std_logic; attribute dont_touch of G11367: signal is true;
	signal G11370: std_logic; attribute dont_touch of G11370: signal is true;
	signal G11373: std_logic; attribute dont_touch of G11373: signal is true;
	signal G11376: std_logic; attribute dont_touch of G11376: signal is true;
	signal G11379: std_logic; attribute dont_touch of G11379: signal is true;
	signal G11382: std_logic; attribute dont_touch of G11382: signal is true;
	signal G11385: std_logic; attribute dont_touch of G11385: signal is true;
	signal G11386: std_logic; attribute dont_touch of G11386: signal is true;
	signal G11389: std_logic; attribute dont_touch of G11389: signal is true;
	signal G11392: std_logic; attribute dont_touch of G11392: signal is true;
	signal G11395: std_logic; attribute dont_touch of G11395: signal is true;
	signal G11398: std_logic; attribute dont_touch of G11398: signal is true;
	signal G11401: std_logic; attribute dont_touch of G11401: signal is true;
	signal G11404: std_logic; attribute dont_touch of G11404: signal is true;
	signal G11407: std_logic; attribute dont_touch of G11407: signal is true;
	signal G11410: std_logic; attribute dont_touch of G11410: signal is true;
	signal G11411: std_logic; attribute dont_touch of G11411: signal is true;
	signal G11414: std_logic; attribute dont_touch of G11414: signal is true;
	signal G11417: std_logic; attribute dont_touch of G11417: signal is true;
	signal G11420: std_logic; attribute dont_touch of G11420: signal is true;
	signal G11421: std_logic; attribute dont_touch of G11421: signal is true;
	signal G11422: std_logic; attribute dont_touch of G11422: signal is true;
	signal G11425: std_logic; attribute dont_touch of G11425: signal is true;
	signal G11428: std_logic; attribute dont_touch of G11428: signal is true;
	signal G11431: std_logic; attribute dont_touch of G11431: signal is true;
	signal G11432: std_logic; attribute dont_touch of G11432: signal is true;
	signal G11435: std_logic; attribute dont_touch of G11435: signal is true;
	signal G11438: std_logic; attribute dont_touch of G11438: signal is true;
	signal G11441: std_logic; attribute dont_touch of G11441: signal is true;
	signal G11444: std_logic; attribute dont_touch of G11444: signal is true;
	signal G11447: std_logic; attribute dont_touch of G11447: signal is true;
	signal G11450: std_logic; attribute dont_touch of G11450: signal is true;
	signal G11453: std_logic; attribute dont_touch of G11453: signal is true;
	signal G11456: std_logic; attribute dont_touch of G11456: signal is true;
	signal G11459: std_logic; attribute dont_touch of G11459: signal is true;
	signal G11462: std_logic; attribute dont_touch of G11462: signal is true;
	signal G11465: std_logic; attribute dont_touch of G11465: signal is true;
	signal G11468: std_logic; attribute dont_touch of G11468: signal is true;
	signal G11471: std_logic; attribute dont_touch of G11471: signal is true;
	signal G11472: std_logic; attribute dont_touch of G11472: signal is true;
	signal G11475: std_logic; attribute dont_touch of G11475: signal is true;
	signal G11478: std_logic; attribute dont_touch of G11478: signal is true;
	signal G11481: std_logic; attribute dont_touch of G11481: signal is true;
	signal G11490: std_logic; attribute dont_touch of G11490: signal is true;
	signal G11491: std_logic; attribute dont_touch of G11491: signal is true;
	signal G11492: std_logic; attribute dont_touch of G11492: signal is true;
	signal G11493: std_logic; attribute dont_touch of G11493: signal is true;
	signal G11494: std_logic; attribute dont_touch of G11494: signal is true;
	signal G11495: std_logic; attribute dont_touch of G11495: signal is true;
	signal G11496: std_logic; attribute dont_touch of G11496: signal is true;
	signal G11497: std_logic; attribute dont_touch of G11497: signal is true;
	signal G11498: std_logic; attribute dont_touch of G11498: signal is true;
	signal G11499: std_logic; attribute dont_touch of G11499: signal is true;
	signal G11500: std_logic; attribute dont_touch of G11500: signal is true;
	signal G11501: std_logic; attribute dont_touch of G11501: signal is true;
	signal G11502: std_logic; attribute dont_touch of G11502: signal is true;
	signal G11503: std_logic; attribute dont_touch of G11503: signal is true;
	signal G11504: std_logic; attribute dont_touch of G11504: signal is true;
	signal G11505: std_logic; attribute dont_touch of G11505: signal is true;
	signal G11506: std_logic; attribute dont_touch of G11506: signal is true;
	signal G11507: std_logic; attribute dont_touch of G11507: signal is true;
	signal G11508: std_logic; attribute dont_touch of G11508: signal is true;
	signal G11509: std_logic; attribute dont_touch of G11509: signal is true;
	signal G11510: std_logic; attribute dont_touch of G11510: signal is true;
	signal G11511: std_logic; attribute dont_touch of G11511: signal is true;
	signal G11512: std_logic; attribute dont_touch of G11512: signal is true;
	signal G11513: std_logic; attribute dont_touch of G11513: signal is true;
	signal G11514: std_logic; attribute dont_touch of G11514: signal is true;
	signal G11515: std_logic; attribute dont_touch of G11515: signal is true;
	signal G11516: std_logic; attribute dont_touch of G11516: signal is true;
	signal G11517: std_logic; attribute dont_touch of G11517: signal is true;
	signal G11518: std_logic; attribute dont_touch of G11518: signal is true;
	signal G11519: std_logic; attribute dont_touch of G11519: signal is true;
	signal G11520: std_logic; attribute dont_touch of G11520: signal is true;
	signal G11521: std_logic; attribute dont_touch of G11521: signal is true;
	signal G11522: std_logic; attribute dont_touch of G11522: signal is true;
	signal G11523: std_logic; attribute dont_touch of G11523: signal is true;
	signal G11524: std_logic; attribute dont_touch of G11524: signal is true;
	signal G11525: std_logic; attribute dont_touch of G11525: signal is true;
	signal G11526: std_logic; attribute dont_touch of G11526: signal is true;
	signal G11527: std_logic; attribute dont_touch of G11527: signal is true;
	signal G11528: std_logic; attribute dont_touch of G11528: signal is true;
	signal G11529: std_logic; attribute dont_touch of G11529: signal is true;
	signal G11530: std_logic; attribute dont_touch of G11530: signal is true;
	signal G11531: std_logic; attribute dont_touch of G11531: signal is true;
	signal G11532: std_logic; attribute dont_touch of G11532: signal is true;
	signal G11533: std_logic; attribute dont_touch of G11533: signal is true;
	signal G11534: std_logic; attribute dont_touch of G11534: signal is true;
	signal G11535: std_logic; attribute dont_touch of G11535: signal is true;
	signal G11536: std_logic; attribute dont_touch of G11536: signal is true;
	signal G11537: std_logic; attribute dont_touch of G11537: signal is true;
	signal G11538: std_logic; attribute dont_touch of G11538: signal is true;
	signal G11539: std_logic; attribute dont_touch of G11539: signal is true;
	signal G11540: std_logic; attribute dont_touch of G11540: signal is true;
	signal G11541: std_logic; attribute dont_touch of G11541: signal is true;
	signal G11542: std_logic; attribute dont_touch of G11542: signal is true;
	signal G11543: std_logic; attribute dont_touch of G11543: signal is true;
	signal G11544: std_logic; attribute dont_touch of G11544: signal is true;
	signal G11545: std_logic; attribute dont_touch of G11545: signal is true;
	signal G11546: std_logic; attribute dont_touch of G11546: signal is true;
	signal G11547: std_logic; attribute dont_touch of G11547: signal is true;
	signal G11548: std_logic; attribute dont_touch of G11548: signal is true;
	signal G11549: std_logic; attribute dont_touch of G11549: signal is true;
	signal G11550: std_logic; attribute dont_touch of G11550: signal is true;
	signal G11551: std_logic; attribute dont_touch of G11551: signal is true;
	signal G11552: std_logic; attribute dont_touch of G11552: signal is true;
	signal G11553: std_logic; attribute dont_touch of G11553: signal is true;
	signal G11554: std_logic; attribute dont_touch of G11554: signal is true;
	signal G11555: std_logic; attribute dont_touch of G11555: signal is true;
	signal G11556: std_logic; attribute dont_touch of G11556: signal is true;
	signal G11557: std_logic; attribute dont_touch of G11557: signal is true;
	signal G11558: std_logic; attribute dont_touch of G11558: signal is true;
	signal G11559: std_logic; attribute dont_touch of G11559: signal is true;
	signal G11560: std_logic; attribute dont_touch of G11560: signal is true;
	signal G11561: std_logic; attribute dont_touch of G11561: signal is true;
	signal G11562: std_logic; attribute dont_touch of G11562: signal is true;
	signal G11563: std_logic; attribute dont_touch of G11563: signal is true;
	signal G11564: std_logic; attribute dont_touch of G11564: signal is true;
	signal G11565: std_logic; attribute dont_touch of G11565: signal is true;
	signal G11566: std_logic; attribute dont_touch of G11566: signal is true;
	signal G11567: std_logic; attribute dont_touch of G11567: signal is true;
	signal G11568: std_logic; attribute dont_touch of G11568: signal is true;
	signal G11569: std_logic; attribute dont_touch of G11569: signal is true;
	signal G11570: std_logic; attribute dont_touch of G11570: signal is true;
	signal G11571: std_logic; attribute dont_touch of G11571: signal is true;
	signal G11572: std_logic; attribute dont_touch of G11572: signal is true;
	signal G11573: std_logic; attribute dont_touch of G11573: signal is true;
	signal G11574: std_logic; attribute dont_touch of G11574: signal is true;
	signal G11575: std_logic; attribute dont_touch of G11575: signal is true;
	signal G11576: std_logic; attribute dont_touch of G11576: signal is true;
	signal G11577: std_logic; attribute dont_touch of G11577: signal is true;
	signal G11578: std_logic; attribute dont_touch of G11578: signal is true;
	signal G11579: std_logic; attribute dont_touch of G11579: signal is true;
	signal G11580: std_logic; attribute dont_touch of G11580: signal is true;
	signal G11581: std_logic; attribute dont_touch of G11581: signal is true;
	signal G11582: std_logic; attribute dont_touch of G11582: signal is true;
	signal G11583: std_logic; attribute dont_touch of G11583: signal is true;
	signal G11584: std_logic; attribute dont_touch of G11584: signal is true;
	signal G11585: std_logic; attribute dont_touch of G11585: signal is true;
	signal G11586: std_logic; attribute dont_touch of G11586: signal is true;
	signal G11587: std_logic; attribute dont_touch of G11587: signal is true;
	signal G11588: std_logic; attribute dont_touch of G11588: signal is true;
	signal G11589: std_logic; attribute dont_touch of G11589: signal is true;
	signal G11590: std_logic; attribute dont_touch of G11590: signal is true;
	signal G11591: std_logic; attribute dont_touch of G11591: signal is true;
	signal G11592: std_logic; attribute dont_touch of G11592: signal is true;
	signal G11593: std_logic; attribute dont_touch of G11593: signal is true;
	signal G11594: std_logic; attribute dont_touch of G11594: signal is true;
	signal G11595: std_logic; attribute dont_touch of G11595: signal is true;
	signal G11596: std_logic; attribute dont_touch of G11596: signal is true;
	signal G11597: std_logic; attribute dont_touch of G11597: signal is true;
	signal G11598: std_logic; attribute dont_touch of G11598: signal is true;
	signal G11599: std_logic; attribute dont_touch of G11599: signal is true;
	signal G11600: std_logic; attribute dont_touch of G11600: signal is true;
	signal G11603: std_logic; attribute dont_touch of G11603: signal is true;
	signal G11606: std_logic; attribute dont_touch of G11606: signal is true;
	signal G11607: std_logic; attribute dont_touch of G11607: signal is true;
	signal G11608: std_logic; attribute dont_touch of G11608: signal is true;
	signal G11611: std_logic; attribute dont_touch of G11611: signal is true;
	signal G11612: std_logic; attribute dont_touch of G11612: signal is true;
	signal G11613: std_logic; attribute dont_touch of G11613: signal is true;
	signal G11616: std_logic; attribute dont_touch of G11616: signal is true;
	signal G11617: std_logic; attribute dont_touch of G11617: signal is true;
	signal G11620: std_logic; attribute dont_touch of G11620: signal is true;
	signal G11621: std_logic; attribute dont_touch of G11621: signal is true;
	signal G11622: std_logic; attribute dont_touch of G11622: signal is true;
	signal G11623: std_logic; attribute dont_touch of G11623: signal is true;
	signal G11624: std_logic; attribute dont_touch of G11624: signal is true;
	signal G11627: std_logic; attribute dont_touch of G11627: signal is true;
	signal G11628: std_logic; attribute dont_touch of G11628: signal is true;
	signal G11629: std_logic; attribute dont_touch of G11629: signal is true;
	signal G11630: std_logic; attribute dont_touch of G11630: signal is true;
	signal G11633: std_logic; attribute dont_touch of G11633: signal is true;
	signal G11636: std_logic; attribute dont_touch of G11636: signal is true;
	signal G11637: std_logic; attribute dont_touch of G11637: signal is true;
	signal G11638: std_logic; attribute dont_touch of G11638: signal is true;
	signal G11641: std_logic; attribute dont_touch of G11641: signal is true;
	signal G11642: std_logic; attribute dont_touch of G11642: signal is true;
	signal G11643: std_logic; attribute dont_touch of G11643: signal is true;
	signal G11644: std_logic; attribute dont_touch of G11644: signal is true;
	signal G11647: std_logic; attribute dont_touch of G11647: signal is true;
	signal G11650: std_logic; attribute dont_touch of G11650: signal is true;
	signal G11651: std_logic; attribute dont_touch of G11651: signal is true;
	signal G11652: std_logic; attribute dont_touch of G11652: signal is true;
	signal G11653: std_logic; attribute dont_touch of G11653: signal is true;
	signal G11656: std_logic; attribute dont_touch of G11656: signal is true;
	signal G11659: std_logic; attribute dont_touch of G11659: signal is true;
	signal G11660: std_logic; attribute dont_touch of G11660: signal is true;
	signal G11661: std_logic; attribute dont_touch of G11661: signal is true;
	signal G11662: std_logic; attribute dont_touch of G11662: signal is true;
	signal G11663: std_logic; attribute dont_touch of G11663: signal is true;
	signal G11666: std_logic; attribute dont_touch of G11666: signal is true;
	signal G11669: std_logic; attribute dont_touch of G11669: signal is true;
	signal G11670: std_logic; attribute dont_touch of G11670: signal is true;
	signal G11671: std_logic; attribute dont_touch of G11671: signal is true;
	signal G11672: std_logic; attribute dont_touch of G11672: signal is true;
	signal G11673: std_logic; attribute dont_touch of G11673: signal is true;
	signal G11674: std_logic; attribute dont_touch of G11674: signal is true;
	signal G11675: std_logic; attribute dont_touch of G11675: signal is true;
	signal G11678: std_logic; attribute dont_touch of G11678: signal is true;
	signal G11681: std_logic; attribute dont_touch of G11681: signal is true;
	signal G11682: std_logic; attribute dont_touch of G11682: signal is true;
	signal G11683: std_logic; attribute dont_touch of G11683: signal is true;
	signal G11684: std_logic; attribute dont_touch of G11684: signal is true;
	signal G11685: std_logic; attribute dont_touch of G11685: signal is true;
	signal G11686: std_logic; attribute dont_touch of G11686: signal is true;
	signal G11687: std_logic; attribute dont_touch of G11687: signal is true;
	signal G11690: std_logic; attribute dont_touch of G11690: signal is true;
	signal G11691: std_logic; attribute dont_touch of G11691: signal is true;
	signal G11692: std_logic; attribute dont_touch of G11692: signal is true;
	signal G11693: std_logic; attribute dont_touch of G11693: signal is true;
	signal G11694: std_logic; attribute dont_touch of G11694: signal is true;
	signal G11695: std_logic; attribute dont_touch of G11695: signal is true;
	signal G11696: std_logic; attribute dont_touch of G11696: signal is true;
	signal G11697: std_logic; attribute dont_touch of G11697: signal is true;
	signal G11698: std_logic; attribute dont_touch of G11698: signal is true;
	signal G11699: std_logic; attribute dont_touch of G11699: signal is true;
	signal G11700: std_logic; attribute dont_touch of G11700: signal is true;
	signal G11701: std_logic; attribute dont_touch of G11701: signal is true;
	signal G11702: std_logic; attribute dont_touch of G11702: signal is true;
	signal G11703: std_logic; attribute dont_touch of G11703: signal is true;
	signal G11704: std_logic; attribute dont_touch of G11704: signal is true;
	signal G11705: std_logic; attribute dont_touch of G11705: signal is true;
	signal G11706: std_logic; attribute dont_touch of G11706: signal is true;
	signal G11707: std_logic; attribute dont_touch of G11707: signal is true;
	signal G11708: std_logic; attribute dont_touch of G11708: signal is true;
	signal G11709: std_logic; attribute dont_touch of G11709: signal is true;
	signal G11710: std_logic; attribute dont_touch of G11710: signal is true;
	signal G11711: std_logic; attribute dont_touch of G11711: signal is true;
	signal G11712: std_logic; attribute dont_touch of G11712: signal is true;
	signal G11713: std_logic; attribute dont_touch of G11713: signal is true;
	signal G11716: std_logic; attribute dont_touch of G11716: signal is true;
	signal G11717: std_logic; attribute dont_touch of G11717: signal is true;
	signal G11718: std_logic; attribute dont_touch of G11718: signal is true;
	signal G11719: std_logic; attribute dont_touch of G11719: signal is true;
	signal G11720: std_logic; attribute dont_touch of G11720: signal is true;
	signal G11721: std_logic; attribute dont_touch of G11721: signal is true;
	signal G11722: std_logic; attribute dont_touch of G11722: signal is true;
	signal G11723: std_logic; attribute dont_touch of G11723: signal is true;
	signal G11724: std_logic; attribute dont_touch of G11724: signal is true;
	signal G11725: std_logic; attribute dont_touch of G11725: signal is true;
	signal G11726: std_logic; attribute dont_touch of G11726: signal is true;
	signal G11727: std_logic; attribute dont_touch of G11727: signal is true;
	signal G11728: std_logic; attribute dont_touch of G11728: signal is true;
	signal G11729: std_logic; attribute dont_touch of G11729: signal is true;
	signal G11730: std_logic; attribute dont_touch of G11730: signal is true;
	signal G11731: std_logic; attribute dont_touch of G11731: signal is true;
	signal G11732: std_logic; attribute dont_touch of G11732: signal is true;
	signal G11733: std_logic; attribute dont_touch of G11733: signal is true;
	signal G11734: std_logic; attribute dont_touch of G11734: signal is true;
	signal G11735: std_logic; attribute dont_touch of G11735: signal is true;
	signal G11736: std_logic; attribute dont_touch of G11736: signal is true;
	signal G11737: std_logic; attribute dont_touch of G11737: signal is true;
	signal G11740: std_logic; attribute dont_touch of G11740: signal is true;
	signal G11741: std_logic; attribute dont_touch of G11741: signal is true;
	signal G11742: std_logic; attribute dont_touch of G11742: signal is true;
	signal G11743: std_logic; attribute dont_touch of G11743: signal is true;
	signal G11744: std_logic; attribute dont_touch of G11744: signal is true;
	signal G11745: std_logic; attribute dont_touch of G11745: signal is true;
	signal G11746: std_logic; attribute dont_touch of G11746: signal is true;
	signal G11747: std_logic; attribute dont_touch of G11747: signal is true;
	signal G11748: std_logic; attribute dont_touch of G11748: signal is true;
	signal G11749: std_logic; attribute dont_touch of G11749: signal is true;
	signal G11758: std_logic; attribute dont_touch of G11758: signal is true;
	signal G11759: std_logic; attribute dont_touch of G11759: signal is true;
	signal G11760: std_logic; attribute dont_touch of G11760: signal is true;
	signal G11761: std_logic; attribute dont_touch of G11761: signal is true;
	signal G11762: std_logic; attribute dont_touch of G11762: signal is true;
	signal G11763: std_logic; attribute dont_touch of G11763: signal is true;
	signal G11764: std_logic; attribute dont_touch of G11764: signal is true;
	signal G11765: std_logic; attribute dont_touch of G11765: signal is true;
	signal G11766: std_logic; attribute dont_touch of G11766: signal is true;
	signal G11767: std_logic; attribute dont_touch of G11767: signal is true;
	signal G11768: std_logic; attribute dont_touch of G11768: signal is true;
	signal G11769: std_logic; attribute dont_touch of G11769: signal is true;
	signal G11770: std_logic; attribute dont_touch of G11770: signal is true;
	signal G11771: std_logic; attribute dont_touch of G11771: signal is true;
	signal G11772: std_logic; attribute dont_touch of G11772: signal is true;
	signal G11773: std_logic; attribute dont_touch of G11773: signal is true;
	signal G11774: std_logic; attribute dont_touch of G11774: signal is true;
	signal G11775: std_logic; attribute dont_touch of G11775: signal is true;
	signal G11776: std_logic; attribute dont_touch of G11776: signal is true;
	signal G11777: std_logic; attribute dont_touch of G11777: signal is true;
	signal G11778: std_logic; attribute dont_touch of G11778: signal is true;
	signal G11779: std_logic; attribute dont_touch of G11779: signal is true;
	signal G11780: std_logic; attribute dont_touch of G11780: signal is true;
	signal G11781: std_logic; attribute dont_touch of G11781: signal is true;
	signal G11782: std_logic; attribute dont_touch of G11782: signal is true;
	signal G11783: std_logic; attribute dont_touch of G11783: signal is true;
	signal G11784: std_logic; attribute dont_touch of G11784: signal is true;
	signal G11785: std_logic; attribute dont_touch of G11785: signal is true;
	signal G11786: std_logic; attribute dont_touch of G11786: signal is true;
	signal G11787: std_logic; attribute dont_touch of G11787: signal is true;
	signal G11788: std_logic; attribute dont_touch of G11788: signal is true;
	signal G11789: std_logic; attribute dont_touch of G11789: signal is true;
	signal G11790: std_logic; attribute dont_touch of G11790: signal is true;
	signal G11791: std_logic; attribute dont_touch of G11791: signal is true;
	signal G11794: std_logic; attribute dont_touch of G11794: signal is true;
	signal G11795: std_logic; attribute dont_touch of G11795: signal is true;
	signal G11796: std_logic; attribute dont_touch of G11796: signal is true;
	signal G11797: std_logic; attribute dont_touch of G11797: signal is true;
	signal G11798: std_logic; attribute dont_touch of G11798: signal is true;
	signal G11799: std_logic; attribute dont_touch of G11799: signal is true;
	signal G11800: std_logic; attribute dont_touch of G11800: signal is true;
	signal G11801: std_logic; attribute dont_touch of G11801: signal is true;
	signal G11802: std_logic; attribute dont_touch of G11802: signal is true;
	signal G11803: std_logic; attribute dont_touch of G11803: signal is true;
	signal G11804: std_logic; attribute dont_touch of G11804: signal is true;
	signal G11805: std_logic; attribute dont_touch of G11805: signal is true;
	signal G11806: std_logic; attribute dont_touch of G11806: signal is true;
	signal G11807: std_logic; attribute dont_touch of G11807: signal is true;
	signal G11808: std_logic; attribute dont_touch of G11808: signal is true;
	signal G11809: std_logic; attribute dont_touch of G11809: signal is true;
	signal G11810: std_logic; attribute dont_touch of G11810: signal is true;
	signal G11811: std_logic; attribute dont_touch of G11811: signal is true;
	signal G11812: std_logic; attribute dont_touch of G11812: signal is true;
	signal G11813: std_logic; attribute dont_touch of G11813: signal is true;
	signal G11814: std_logic; attribute dont_touch of G11814: signal is true;
	signal G11815: std_logic; attribute dont_touch of G11815: signal is true;
	signal G11816: std_logic; attribute dont_touch of G11816: signal is true;
	signal G11817: std_logic; attribute dont_touch of G11817: signal is true;
	signal G11818: std_logic; attribute dont_touch of G11818: signal is true;
	signal G11819: std_logic; attribute dont_touch of G11819: signal is true;
	signal G11820: std_logic; attribute dont_touch of G11820: signal is true;
	signal G11821: std_logic; attribute dont_touch of G11821: signal is true;
	signal G11822: std_logic; attribute dont_touch of G11822: signal is true;
	signal G11823: std_logic; attribute dont_touch of G11823: signal is true;
	signal G11824: std_logic; attribute dont_touch of G11824: signal is true;
	signal G11825: std_logic; attribute dont_touch of G11825: signal is true;
	signal G11826: std_logic; attribute dont_touch of G11826: signal is true;
	signal G11827: std_logic; attribute dont_touch of G11827: signal is true;
	signal G11828: std_logic; attribute dont_touch of G11828: signal is true;
	signal G11829: std_logic; attribute dont_touch of G11829: signal is true;
	signal G11830: std_logic; attribute dont_touch of G11830: signal is true;
	signal G11831: std_logic; attribute dont_touch of G11831: signal is true;
	signal G11832: std_logic; attribute dont_touch of G11832: signal is true;
	signal G11833: std_logic; attribute dont_touch of G11833: signal is true;
	signal G11834: std_logic; attribute dont_touch of G11834: signal is true;
	signal G11835: std_logic; attribute dont_touch of G11835: signal is true;
	signal G11836: std_logic; attribute dont_touch of G11836: signal is true;
	signal G11837: std_logic; attribute dont_touch of G11837: signal is true;
	signal G11838: std_logic; attribute dont_touch of G11838: signal is true;
	signal G11839: std_logic; attribute dont_touch of G11839: signal is true;
	signal G11840: std_logic; attribute dont_touch of G11840: signal is true;
	signal G11841: std_logic; attribute dont_touch of G11841: signal is true;
	signal G11842: std_logic; attribute dont_touch of G11842: signal is true;
	signal G11843: std_logic; attribute dont_touch of G11843: signal is true;
	signal G11844: std_logic; attribute dont_touch of G11844: signal is true;
	signal G11845: std_logic; attribute dont_touch of G11845: signal is true;
	signal G11846: std_logic; attribute dont_touch of G11846: signal is true;
	signal G11847: std_logic; attribute dont_touch of G11847: signal is true;
	signal G11848: std_logic; attribute dont_touch of G11848: signal is true;
	signal G11851: std_logic; attribute dont_touch of G11851: signal is true;
	signal G11852: std_logic; attribute dont_touch of G11852: signal is true;
	signal G11853: std_logic; attribute dont_touch of G11853: signal is true;
	signal G11854: std_logic; attribute dont_touch of G11854: signal is true;
	signal G11855: std_logic; attribute dont_touch of G11855: signal is true;
	signal G11856: std_logic; attribute dont_touch of G11856: signal is true;
	signal G11857: std_logic; attribute dont_touch of G11857: signal is true;
	signal G11858: std_logic; attribute dont_touch of G11858: signal is true;
	signal G11859: std_logic; attribute dont_touch of G11859: signal is true;
	signal G11860: std_logic; attribute dont_touch of G11860: signal is true;
	signal G11861: std_logic; attribute dont_touch of G11861: signal is true;
	signal G11862: std_logic; attribute dont_touch of G11862: signal is true;
	signal G11863: std_logic; attribute dont_touch of G11863: signal is true;
	signal G11864: std_logic; attribute dont_touch of G11864: signal is true;
	signal G11865: std_logic; attribute dont_touch of G11865: signal is true;
	signal G11866: std_logic; attribute dont_touch of G11866: signal is true;
	signal G11867: std_logic; attribute dont_touch of G11867: signal is true;
	signal G11868: std_logic; attribute dont_touch of G11868: signal is true;
	signal G11869: std_logic; attribute dont_touch of G11869: signal is true;
	signal G11870: std_logic; attribute dont_touch of G11870: signal is true;
	signal G11871: std_logic; attribute dont_touch of G11871: signal is true;
	signal G11872: std_logic; attribute dont_touch of G11872: signal is true;
	signal G11873: std_logic; attribute dont_touch of G11873: signal is true;
	signal G11874: std_logic; attribute dont_touch of G11874: signal is true;
	signal G11875: std_logic; attribute dont_touch of G11875: signal is true;
	signal G11876: std_logic; attribute dont_touch of G11876: signal is true;
	signal G11877: std_logic; attribute dont_touch of G11877: signal is true;
	signal G11878: std_logic; attribute dont_touch of G11878: signal is true;
	signal G11879: std_logic; attribute dont_touch of G11879: signal is true;
	signal G11880: std_logic; attribute dont_touch of G11880: signal is true;
	signal G11881: std_logic; attribute dont_touch of G11881: signal is true;
	signal G11882: std_logic; attribute dont_touch of G11882: signal is true;
	signal G11883: std_logic; attribute dont_touch of G11883: signal is true;
	signal G11884: std_logic; attribute dont_touch of G11884: signal is true;
	signal G11885: std_logic; attribute dont_touch of G11885: signal is true;
	signal G11886: std_logic; attribute dont_touch of G11886: signal is true;
	signal G11887: std_logic; attribute dont_touch of G11887: signal is true;
	signal G11888: std_logic; attribute dont_touch of G11888: signal is true;
	signal G11889: std_logic; attribute dont_touch of G11889: signal is true;
	signal G11890: std_logic; attribute dont_touch of G11890: signal is true;
	signal G11891: std_logic; attribute dont_touch of G11891: signal is true;
	signal G11892: std_logic; attribute dont_touch of G11892: signal is true;
	signal G11893: std_logic; attribute dont_touch of G11893: signal is true;
	signal G11894: std_logic; attribute dont_touch of G11894: signal is true;
	signal G11895: std_logic; attribute dont_touch of G11895: signal is true;
	signal G11896: std_logic; attribute dont_touch of G11896: signal is true;
	signal G11897: std_logic; attribute dont_touch of G11897: signal is true;
	signal G11898: std_logic; attribute dont_touch of G11898: signal is true;
	signal G11899: std_logic; attribute dont_touch of G11899: signal is true;
	signal G11900: std_logic; attribute dont_touch of G11900: signal is true;
	signal G11901: std_logic; attribute dont_touch of G11901: signal is true;
	signal G11902: std_logic; attribute dont_touch of G11902: signal is true;
	signal G11903: std_logic; attribute dont_touch of G11903: signal is true;
	signal G11904: std_logic; attribute dont_touch of G11904: signal is true;
	signal G11905: std_logic; attribute dont_touch of G11905: signal is true;
	signal G11906: std_logic; attribute dont_touch of G11906: signal is true;
	signal G11907: std_logic; attribute dont_touch of G11907: signal is true;
	signal G11908: std_logic; attribute dont_touch of G11908: signal is true;
	signal G11909: std_logic; attribute dont_touch of G11909: signal is true;
	signal G11910: std_logic; attribute dont_touch of G11910: signal is true;
	signal G11911: std_logic; attribute dont_touch of G11911: signal is true;
	signal G11912: std_logic; attribute dont_touch of G11912: signal is true;
	signal G11913: std_logic; attribute dont_touch of G11913: signal is true;
	signal G11914: std_logic; attribute dont_touch of G11914: signal is true;
	signal G11915: std_logic; attribute dont_touch of G11915: signal is true;
	signal G11916: std_logic; attribute dont_touch of G11916: signal is true;
	signal G11917: std_logic; attribute dont_touch of G11917: signal is true;
	signal G11918: std_logic; attribute dont_touch of G11918: signal is true;
	signal G11919: std_logic; attribute dont_touch of G11919: signal is true;
	signal G11920: std_logic; attribute dont_touch of G11920: signal is true;
	signal G11921: std_logic; attribute dont_touch of G11921: signal is true;
	signal G11922: std_logic; attribute dont_touch of G11922: signal is true;
	signal G11923: std_logic; attribute dont_touch of G11923: signal is true;
	signal G11926: std_logic; attribute dont_touch of G11926: signal is true;
	signal G11927: std_logic; attribute dont_touch of G11927: signal is true;
	signal G11928: std_logic; attribute dont_touch of G11928: signal is true;
	signal G11929: std_logic; attribute dont_touch of G11929: signal is true;
	signal G11930: std_logic; attribute dont_touch of G11930: signal is true;
	signal G11931: std_logic; attribute dont_touch of G11931: signal is true;
	signal G11932: std_logic; attribute dont_touch of G11932: signal is true;
	signal G11933: std_logic; attribute dont_touch of G11933: signal is true;
	signal G11934: std_logic; attribute dont_touch of G11934: signal is true;
	signal G11935: std_logic; attribute dont_touch of G11935: signal is true;
	signal G11936: std_logic; attribute dont_touch of G11936: signal is true;
	signal G11937: std_logic; attribute dont_touch of G11937: signal is true;
	signal G11938: std_logic; attribute dont_touch of G11938: signal is true;
	signal G11939: std_logic; attribute dont_touch of G11939: signal is true;
	signal G11940: std_logic; attribute dont_touch of G11940: signal is true;
	signal G11941: std_logic; attribute dont_touch of G11941: signal is true;
	signal G11942: std_logic; attribute dont_touch of G11942: signal is true;
	signal G11943: std_logic; attribute dont_touch of G11943: signal is true;
	signal G11944: std_logic; attribute dont_touch of G11944: signal is true;
	signal G11945: std_logic; attribute dont_touch of G11945: signal is true;
	signal G11946: std_logic; attribute dont_touch of G11946: signal is true;
	signal G11947: std_logic; attribute dont_touch of G11947: signal is true;
	signal G11948: std_logic; attribute dont_touch of G11948: signal is true;
	signal G11949: std_logic; attribute dont_touch of G11949: signal is true;
	signal G11950: std_logic; attribute dont_touch of G11950: signal is true;
	signal G11951: std_logic; attribute dont_touch of G11951: signal is true;
	signal G11952: std_logic; attribute dont_touch of G11952: signal is true;
	signal G11953: std_logic; attribute dont_touch of G11953: signal is true;
	signal G11954: std_logic; attribute dont_touch of G11954: signal is true;
	signal G11955: std_logic; attribute dont_touch of G11955: signal is true;
	signal G11956: std_logic; attribute dont_touch of G11956: signal is true;
	signal G11957: std_logic; attribute dont_touch of G11957: signal is true;
	signal G11958: std_logic; attribute dont_touch of G11958: signal is true;
	signal G11959: std_logic; attribute dont_touch of G11959: signal is true;
	signal G11960: std_logic; attribute dont_touch of G11960: signal is true;
	signal G11961: std_logic; attribute dont_touch of G11961: signal is true;
	signal G11962: std_logic; attribute dont_touch of G11962: signal is true;
	signal G11963: std_logic; attribute dont_touch of G11963: signal is true;
	signal G11964: std_logic; attribute dont_touch of G11964: signal is true;
	signal G11965: std_logic; attribute dont_touch of G11965: signal is true;
	signal G11966: std_logic; attribute dont_touch of G11966: signal is true;
	signal G11967: std_logic; attribute dont_touch of G11967: signal is true;
	signal G11968: std_logic; attribute dont_touch of G11968: signal is true;
	signal G11969: std_logic; attribute dont_touch of G11969: signal is true;
	signal G11970: std_logic; attribute dont_touch of G11970: signal is true;
	signal G11971: std_logic; attribute dont_touch of G11971: signal is true;
	signal G11972: std_logic; attribute dont_touch of G11972: signal is true;
	signal G11973: std_logic; attribute dont_touch of G11973: signal is true;
	signal G11974: std_logic; attribute dont_touch of G11974: signal is true;
	signal G11975: std_logic; attribute dont_touch of G11975: signal is true;
	signal G11976: std_logic; attribute dont_touch of G11976: signal is true;
	signal G11979: std_logic; attribute dont_touch of G11979: signal is true;
	signal G11980: std_logic; attribute dont_touch of G11980: signal is true;
	signal G11981: std_logic; attribute dont_touch of G11981: signal is true;
	signal G11982: std_logic; attribute dont_touch of G11982: signal is true;
	signal G11983: std_logic; attribute dont_touch of G11983: signal is true;
	signal G11984: std_logic; attribute dont_touch of G11984: signal is true;
	signal G11985: std_logic; attribute dont_touch of G11985: signal is true;
	signal G11986: std_logic; attribute dont_touch of G11986: signal is true;
	signal G11987: std_logic; attribute dont_touch of G11987: signal is true;
	signal G11988: std_logic; attribute dont_touch of G11988: signal is true;
	signal G11989: std_logic; attribute dont_touch of G11989: signal is true;
	signal G11990: std_logic; attribute dont_touch of G11990: signal is true;
	signal G11991: std_logic; attribute dont_touch of G11991: signal is true;
	signal G11992: std_logic; attribute dont_touch of G11992: signal is true;
	signal G11993: std_logic; attribute dont_touch of G11993: signal is true;
	signal G11994: std_logic; attribute dont_touch of G11994: signal is true;
	signal G11995: std_logic; attribute dont_touch of G11995: signal is true;
	signal G11996: std_logic; attribute dont_touch of G11996: signal is true;
	signal G11997: std_logic; attribute dont_touch of G11997: signal is true;
	signal G11998: std_logic; attribute dont_touch of G11998: signal is true;
	signal G11999: std_logic; attribute dont_touch of G11999: signal is true;
	signal G12000: std_logic; attribute dont_touch of G12000: signal is true;
	signal G12001: std_logic; attribute dont_touch of G12001: signal is true;
	signal G12002: std_logic; attribute dont_touch of G12002: signal is true;
	signal G12003: std_logic; attribute dont_touch of G12003: signal is true;
	signal G12004: std_logic; attribute dont_touch of G12004: signal is true;
	signal G12005: std_logic; attribute dont_touch of G12005: signal is true;
	signal G12006: std_logic; attribute dont_touch of G12006: signal is true;
	signal G12007: std_logic; attribute dont_touch of G12007: signal is true;
	signal G12008: std_logic; attribute dont_touch of G12008: signal is true;
	signal G12009: std_logic; attribute dont_touch of G12009: signal is true;
	signal G12012: std_logic; attribute dont_touch of G12012: signal is true;
	signal G12013: std_logic; attribute dont_touch of G12013: signal is true;
	signal G12017: std_logic; attribute dont_touch of G12017: signal is true;
	signal G12020: std_logic; attribute dont_touch of G12020: signal is true;
	signal G12021: std_logic; attribute dont_touch of G12021: signal is true;
	signal G12022: std_logic; attribute dont_touch of G12022: signal is true;
	signal G12023: std_logic; attribute dont_touch of G12023: signal is true;
	signal G12024: std_logic; attribute dont_touch of G12024: signal is true;
	signal G12025: std_logic; attribute dont_touch of G12025: signal is true;
	signal G12026: std_logic; attribute dont_touch of G12026: signal is true;
	signal G12027: std_logic; attribute dont_touch of G12027: signal is true;
	signal G12030: std_logic; attribute dont_touch of G12030: signal is true;
	signal G12033: std_logic; attribute dont_touch of G12033: signal is true;
	signal G12034: std_logic; attribute dont_touch of G12034: signal is true;
	signal G12035: std_logic; attribute dont_touch of G12035: signal is true;
	signal G12036: std_logic; attribute dont_touch of G12036: signal is true;
	signal G12037: std_logic; attribute dont_touch of G12037: signal is true;
	signal G12038: std_logic; attribute dont_touch of G12038: signal is true;
	signal G12039: std_logic; attribute dont_touch of G12039: signal is true;
	signal G12040: std_logic; attribute dont_touch of G12040: signal is true;
	signal G12041: std_logic; attribute dont_touch of G12041: signal is true;
	signal G12042: std_logic; attribute dont_touch of G12042: signal is true;
	signal G12043: std_logic; attribute dont_touch of G12043: signal is true;
	signal G12044: std_logic; attribute dont_touch of G12044: signal is true;
	signal G12045: std_logic; attribute dont_touch of G12045: signal is true;
	signal G12048: std_logic; attribute dont_touch of G12048: signal is true;
	signal G12049: std_logic; attribute dont_touch of G12049: signal is true;
	signal G12050: std_logic; attribute dont_touch of G12050: signal is true;
	signal G12051: std_logic; attribute dont_touch of G12051: signal is true;
	signal G12052: std_logic; attribute dont_touch of G12052: signal is true;
	signal G12053: std_logic; attribute dont_touch of G12053: signal is true;
	signal G12054: std_logic; attribute dont_touch of G12054: signal is true;
	signal G12055: std_logic; attribute dont_touch of G12055: signal is true;
	signal G12056: std_logic; attribute dont_touch of G12056: signal is true;
	signal G12057: std_logic; attribute dont_touch of G12057: signal is true;
	signal G12058: std_logic; attribute dont_touch of G12058: signal is true;
	signal G12059: std_logic; attribute dont_touch of G12059: signal is true;
	signal G12060: std_logic; attribute dont_touch of G12060: signal is true;
	signal G12061: std_logic; attribute dont_touch of G12061: signal is true;
	signal G12062: std_logic; attribute dont_touch of G12062: signal is true;
	signal G12063: std_logic; attribute dont_touch of G12063: signal is true;
	signal G12064: std_logic; attribute dont_touch of G12064: signal is true;
	signal G12065: std_logic; attribute dont_touch of G12065: signal is true;
	signal G12066: std_logic; attribute dont_touch of G12066: signal is true;
	signal G12067: std_logic; attribute dont_touch of G12067: signal is true;
	signal G12068: std_logic; attribute dont_touch of G12068: signal is true;
	signal G12069: std_logic; attribute dont_touch of G12069: signal is true;
	signal G12070: std_logic; attribute dont_touch of G12070: signal is true;
	signal G12071: std_logic; attribute dont_touch of G12071: signal is true;
	signal G12075: std_logic; attribute dont_touch of G12075: signal is true;
	signal G12076: std_logic; attribute dont_touch of G12076: signal is true;
	signal G12077: std_logic; attribute dont_touch of G12077: signal is true;
	signal G12078: std_logic; attribute dont_touch of G12078: signal is true;
	signal G12079: std_logic; attribute dont_touch of G12079: signal is true;
	signal G12080: std_logic; attribute dont_touch of G12080: signal is true;
	signal G12081: std_logic; attribute dont_touch of G12081: signal is true;
	signal G12082: std_logic; attribute dont_touch of G12082: signal is true;
	signal G12083: std_logic; attribute dont_touch of G12083: signal is true;
	signal G12084: std_logic; attribute dont_touch of G12084: signal is true;
	signal G12085: std_logic; attribute dont_touch of G12085: signal is true;
	signal G12086: std_logic; attribute dont_touch of G12086: signal is true;
	signal G12087: std_logic; attribute dont_touch of G12087: signal is true;
	signal G12088: std_logic; attribute dont_touch of G12088: signal is true;
	signal G12089: std_logic; attribute dont_touch of G12089: signal is true;
	signal G12090: std_logic; attribute dont_touch of G12090: signal is true;
	signal G12091: std_logic; attribute dont_touch of G12091: signal is true;
	signal G12094: std_logic; attribute dont_touch of G12094: signal is true;
	signal G12097: std_logic; attribute dont_touch of G12097: signal is true;
	signal G12098: std_logic; attribute dont_touch of G12098: signal is true;
	signal G12099: std_logic; attribute dont_touch of G12099: signal is true;
	signal G12100: std_logic; attribute dont_touch of G12100: signal is true;
	signal G12101: std_logic; attribute dont_touch of G12101: signal is true;
	signal G12102: std_logic; attribute dont_touch of G12102: signal is true;
	signal G12103: std_logic; attribute dont_touch of G12103: signal is true;
	signal G12104: std_logic; attribute dont_touch of G12104: signal is true;
	signal G12105: std_logic; attribute dont_touch of G12105: signal is true;
	signal G12106: std_logic; attribute dont_touch of G12106: signal is true;
	signal G12107: std_logic; attribute dont_touch of G12107: signal is true;
	signal G12108: std_logic; attribute dont_touch of G12108: signal is true;
	signal G12109: std_logic; attribute dont_touch of G12109: signal is true;
	signal G12112: std_logic; attribute dont_touch of G12112: signal is true;
	signal G12113: std_logic; attribute dont_touch of G12113: signal is true;
	signal G12114: std_logic; attribute dont_touch of G12114: signal is true;
	signal G12115: std_logic; attribute dont_touch of G12115: signal is true;
	signal G12116: std_logic; attribute dont_touch of G12116: signal is true;
	signal G12117: std_logic; attribute dont_touch of G12117: signal is true;
	signal G12118: std_logic; attribute dont_touch of G12118: signal is true;
	signal G12119: std_logic; attribute dont_touch of G12119: signal is true;
	signal G12120: std_logic; attribute dont_touch of G12120: signal is true;
	signal G12121: std_logic; attribute dont_touch of G12121: signal is true;
	signal G12122: std_logic; attribute dont_touch of G12122: signal is true;
	signal G12123: std_logic; attribute dont_touch of G12123: signal is true;
	signal G12124: std_logic; attribute dont_touch of G12124: signal is true;
	signal G12125: std_logic; attribute dont_touch of G12125: signal is true;
	signal G12128: std_logic; attribute dont_touch of G12128: signal is true;
	signal G12129: std_logic; attribute dont_touch of G12129: signal is true;
	signal G12130: std_logic; attribute dont_touch of G12130: signal is true;
	signal G12134: std_logic; attribute dont_touch of G12134: signal is true;
	signal G12135: std_logic; attribute dont_touch of G12135: signal is true;
	signal G12136: std_logic; attribute dont_touch of G12136: signal is true;
	signal G12139: std_logic; attribute dont_touch of G12139: signal is true;
	signal G12142: std_logic; attribute dont_touch of G12142: signal is true;
	signal G12145: std_logic; attribute dont_touch of G12145: signal is true;
	signal G12146: std_logic; attribute dont_touch of G12146: signal is true;
	signal G12147: std_logic; attribute dont_touch of G12147: signal is true;
	signal G12148: std_logic; attribute dont_touch of G12148: signal is true;
	signal G12149: std_logic; attribute dont_touch of G12149: signal is true;
	signal G12150: std_logic; attribute dont_touch of G12150: signal is true;
	signal G12151: std_logic; attribute dont_touch of G12151: signal is true;
	signal G12152: std_logic; attribute dont_touch of G12152: signal is true;
	signal G12153: std_logic; attribute dont_touch of G12153: signal is true;
	signal G12154: std_logic; attribute dont_touch of G12154: signal is true;
	signal G12155: std_logic; attribute dont_touch of G12155: signal is true;
	signal G12156: std_logic; attribute dont_touch of G12156: signal is true;
	signal G12157: std_logic; attribute dont_touch of G12157: signal is true;
	signal G12158: std_logic; attribute dont_touch of G12158: signal is true;
	signal G12159: std_logic; attribute dont_touch of G12159: signal is true;
	signal G12160: std_logic; attribute dont_touch of G12160: signal is true;
	signal G12161: std_logic; attribute dont_touch of G12161: signal is true;
	signal G12162: std_logic; attribute dont_touch of G12162: signal is true;
	signal G12163: std_logic; attribute dont_touch of G12163: signal is true;
	signal G12166: std_logic; attribute dont_touch of G12166: signal is true;
	signal G12169: std_logic; attribute dont_touch of G12169: signal is true;
	signal G12170: std_logic; attribute dont_touch of G12170: signal is true;
	signal G12171: std_logic; attribute dont_touch of G12171: signal is true;
	signal G12172: std_logic; attribute dont_touch of G12172: signal is true;
	signal G12173: std_logic; attribute dont_touch of G12173: signal is true;
	signal G12174: std_logic; attribute dont_touch of G12174: signal is true;
	signal G12175: std_logic; attribute dont_touch of G12175: signal is true;
	signal G12176: std_logic; attribute dont_touch of G12176: signal is true;
	signal G12177: std_logic; attribute dont_touch of G12177: signal is true;
	signal G12178: std_logic; attribute dont_touch of G12178: signal is true;
	signal G12179: std_logic; attribute dont_touch of G12179: signal is true;
	signal G12180: std_logic; attribute dont_touch of G12180: signal is true;
	signal G12181: std_logic; attribute dont_touch of G12181: signal is true;
	signal G12184: std_logic; attribute dont_touch of G12184: signal is true;
	signal G12185: std_logic; attribute dont_touch of G12185: signal is true;
	signal G12186: std_logic; attribute dont_touch of G12186: signal is true;
	signal G12187: std_logic; attribute dont_touch of G12187: signal is true;
	signal G12191: std_logic; attribute dont_touch of G12191: signal is true;
	signal G12192: std_logic; attribute dont_touch of G12192: signal is true;
	signal G12193: std_logic; attribute dont_touch of G12193: signal is true;
	signal G12194: std_logic; attribute dont_touch of G12194: signal is true;
	signal G12195: std_logic; attribute dont_touch of G12195: signal is true;
	signal G12196: std_logic; attribute dont_touch of G12196: signal is true;
	signal G12197: std_logic; attribute dont_touch of G12197: signal is true;
	signal G12198: std_logic; attribute dont_touch of G12198: signal is true;
	signal G12201: std_logic; attribute dont_touch of G12201: signal is true;
	signal G12204: std_logic; attribute dont_touch of G12204: signal is true;
	signal G12207: std_logic; attribute dont_touch of G12207: signal is true;
	signal G12208: std_logic; attribute dont_touch of G12208: signal is true;
	signal G12209: std_logic; attribute dont_touch of G12209: signal is true;
	signal G12210: std_logic; attribute dont_touch of G12210: signal is true;
	signal G12211: std_logic; attribute dont_touch of G12211: signal is true;
	signal G12212: std_logic; attribute dont_touch of G12212: signal is true;
	signal G12213: std_logic; attribute dont_touch of G12213: signal is true;
	signal G12214: std_logic; attribute dont_touch of G12214: signal is true;
	signal G12215: std_logic; attribute dont_touch of G12215: signal is true;
	signal G12216: std_logic; attribute dont_touch of G12216: signal is true;
	signal G12217: std_logic; attribute dont_touch of G12217: signal is true;
	signal G12218: std_logic; attribute dont_touch of G12218: signal is true;
	signal G12219: std_logic; attribute dont_touch of G12219: signal is true;
	signal G12220: std_logic; attribute dont_touch of G12220: signal is true;
	signal G12221: std_logic; attribute dont_touch of G12221: signal is true;
	signal G12222: std_logic; attribute dont_touch of G12222: signal is true;
	signal G12223: std_logic; attribute dont_touch of G12223: signal is true;
	signal G12224: std_logic; attribute dont_touch of G12224: signal is true;
	signal G12225: std_logic; attribute dont_touch of G12225: signal is true;
	signal G12228: std_logic; attribute dont_touch of G12228: signal is true;
	signal G12231: std_logic; attribute dont_touch of G12231: signal is true;
	signal G12232: std_logic; attribute dont_touch of G12232: signal is true;
	signal G12233: std_logic; attribute dont_touch of G12233: signal is true;
	signal G12234: std_logic; attribute dont_touch of G12234: signal is true;
	signal G12235: std_logic; attribute dont_touch of G12235: signal is true;
	signal G12239: std_logic; attribute dont_touch of G12239: signal is true;
	signal G12242: std_logic; attribute dont_touch of G12242: signal is true;
	signal G12245: std_logic; attribute dont_touch of G12245: signal is true;
	signal G12246: std_logic; attribute dont_touch of G12246: signal is true;
	signal G12247: std_logic; attribute dont_touch of G12247: signal is true;
	signal G12248: std_logic; attribute dont_touch of G12248: signal is true;
	signal G12249: std_logic; attribute dont_touch of G12249: signal is true;
	signal G12250: std_logic; attribute dont_touch of G12250: signal is true;
	signal G12251: std_logic; attribute dont_touch of G12251: signal is true;
	signal G12252: std_logic; attribute dont_touch of G12252: signal is true;
	signal G12253: std_logic; attribute dont_touch of G12253: signal is true;
	signal G12256: std_logic; attribute dont_touch of G12256: signal is true;
	signal G12259: std_logic; attribute dont_touch of G12259: signal is true;
	signal G12262: std_logic; attribute dont_touch of G12262: signal is true;
	signal G12263: std_logic; attribute dont_touch of G12263: signal is true;
	signal G12264: std_logic; attribute dont_touch of G12264: signal is true;
	signal G12265: std_logic; attribute dont_touch of G12265: signal is true;
	signal G12266: std_logic; attribute dont_touch of G12266: signal is true;
	signal G12267: std_logic; attribute dont_touch of G12267: signal is true;
	signal G12268: std_logic; attribute dont_touch of G12268: signal is true;
	signal G12269: std_logic; attribute dont_touch of G12269: signal is true;
	signal G12270: std_logic; attribute dont_touch of G12270: signal is true;
	signal G12271: std_logic; attribute dont_touch of G12271: signal is true;
	signal G12272: std_logic; attribute dont_touch of G12272: signal is true;
	signal G12273: std_logic; attribute dont_touch of G12273: signal is true;
	signal G12274: std_logic; attribute dont_touch of G12274: signal is true;
	signal G12275: std_logic; attribute dont_touch of G12275: signal is true;
	signal G12279: std_logic; attribute dont_touch of G12279: signal is true;
	signal G12282: std_logic; attribute dont_touch of G12282: signal is true;
	signal G12285: std_logic; attribute dont_touch of G12285: signal is true;
	signal G12288: std_logic; attribute dont_touch of G12288: signal is true;
	signal G12289: std_logic; attribute dont_touch of G12289: signal is true;
	signal G12290: std_logic; attribute dont_touch of G12290: signal is true;
	signal G12291: std_logic; attribute dont_touch of G12291: signal is true;
	signal G12292: std_logic; attribute dont_touch of G12292: signal is true;
	signal G12293: std_logic; attribute dont_touch of G12293: signal is true;
	signal G12294: std_logic; attribute dont_touch of G12294: signal is true;
	signal G12295: std_logic; attribute dont_touch of G12295: signal is true;
	signal G12296: std_logic; attribute dont_touch of G12296: signal is true;
	signal G12299: std_logic; attribute dont_touch of G12299: signal is true;
	signal G12302: std_logic; attribute dont_touch of G12302: signal is true;
	signal G12305: std_logic; attribute dont_touch of G12305: signal is true;
	signal G12306: std_logic; attribute dont_touch of G12306: signal is true;
	signal G12307: std_logic; attribute dont_touch of G12307: signal is true;
	signal G12308: std_logic; attribute dont_touch of G12308: signal is true;
	signal G12312: std_logic; attribute dont_touch of G12312: signal is true;
	signal G12315: std_logic; attribute dont_touch of G12315: signal is true;
	signal G12318: std_logic; attribute dont_touch of G12318: signal is true;
	signal G12321: std_logic; attribute dont_touch of G12321: signal is true;
	signal G12324: std_logic; attribute dont_touch of G12324: signal is true;
	signal G12325: std_logic; attribute dont_touch of G12325: signal is true;
	signal G12326: std_logic; attribute dont_touch of G12326: signal is true;
	signal G12327: std_logic; attribute dont_touch of G12327: signal is true;
	signal G12328: std_logic; attribute dont_touch of G12328: signal is true;
	signal G12329: std_logic; attribute dont_touch of G12329: signal is true;
	signal G12330: std_logic; attribute dont_touch of G12330: signal is true;
	signal G12331: std_logic; attribute dont_touch of G12331: signal is true;
	signal G12332: std_logic; attribute dont_touch of G12332: signal is true;
	signal G12333: std_logic; attribute dont_touch of G12333: signal is true;
	signal G12336: std_logic; attribute dont_touch of G12336: signal is true;
	signal G12339: std_logic; attribute dont_touch of G12339: signal is true;
	signal G12340: std_logic; attribute dont_touch of G12340: signal is true;
	signal G12343: std_logic; attribute dont_touch of G12343: signal is true;
	signal G12346: std_logic; attribute dont_touch of G12346: signal is true;
	signal G12349: std_logic; attribute dont_touch of G12349: signal is true;
	signal G12352: std_logic; attribute dont_touch of G12352: signal is true;
	signal G12353: std_logic; attribute dont_touch of G12353: signal is true;
	signal G12354: std_logic; attribute dont_touch of G12354: signal is true;
	signal G12362: std_logic; attribute dont_touch of G12362: signal is true;
	signal G12363: std_logic; attribute dont_touch of G12363: signal is true;
	signal G12366: std_logic; attribute dont_touch of G12366: signal is true;
	signal G12369: std_logic; attribute dont_touch of G12369: signal is true;
	signal G12370: std_logic; attribute dont_touch of G12370: signal is true;
	signal G12373: std_logic; attribute dont_touch of G12373: signal is true;
	signal G12376: std_logic; attribute dont_touch of G12376: signal is true;
	signal G12377: std_logic; attribute dont_touch of G12377: signal is true;
	signal G12378: std_logic; attribute dont_touch of G12378: signal is true;
	signal G12379: std_logic; attribute dont_touch of G12379: signal is true;
	signal G12382: std_logic; attribute dont_touch of G12382: signal is true;
	signal G12385: std_logic; attribute dont_touch of G12385: signal is true;
	signal G12388: std_logic; attribute dont_touch of G12388: signal is true;
	signal G12389: std_logic; attribute dont_touch of G12389: signal is true;
	signal G12392: std_logic; attribute dont_touch of G12392: signal is true;
	signal G12407: std_logic; attribute dont_touch of G12407: signal is true;
	signal G12408: std_logic; attribute dont_touch of G12408: signal is true;
	signal G12409: std_logic; attribute dont_touch of G12409: signal is true;
	signal G12412: std_logic; attribute dont_touch of G12412: signal is true;
	signal G12415: std_logic; attribute dont_touch of G12415: signal is true;
	signal G12418: std_logic; attribute dont_touch of G12418: signal is true;
	signal G12419: std_logic; attribute dont_touch of G12419: signal is true;
	signal G12420: std_logic; attribute dont_touch of G12420: signal is true;
	signal G12421: std_logic; attribute dont_touch of G12421: signal is true;
	signal G12424: std_logic; attribute dont_touch of G12424: signal is true;
	signal G12425: std_logic; attribute dont_touch of G12425: signal is true;
	signal G12426: std_logic; attribute dont_touch of G12426: signal is true;
	signal G12429: std_logic; attribute dont_touch of G12429: signal is true;
	signal G12430: std_logic; attribute dont_touch of G12430: signal is true;
	signal G12431: std_logic; attribute dont_touch of G12431: signal is true;
	signal G12432: std_logic; attribute dont_touch of G12432: signal is true;
	signal G12433: std_logic; attribute dont_touch of G12433: signal is true;
	signal G12434: std_logic; attribute dont_touch of G12434: signal is true;
	signal G12435: std_logic; attribute dont_touch of G12435: signal is true;
	signal G12436: std_logic; attribute dont_touch of G12436: signal is true;
	signal G12437: std_logic; attribute dont_touch of G12437: signal is true;
	signal G12438: std_logic; attribute dont_touch of G12438: signal is true;
	signal G12439: std_logic; attribute dont_touch of G12439: signal is true;
	signal G12440: std_logic; attribute dont_touch of G12440: signal is true;
	signal G12441: std_logic; attribute dont_touch of G12441: signal is true;
	signal G12442: std_logic; attribute dont_touch of G12442: signal is true;
	signal G12443: std_logic; attribute dont_touch of G12443: signal is true;
	signal G12444: std_logic; attribute dont_touch of G12444: signal is true;
	signal G12445: std_logic; attribute dont_touch of G12445: signal is true;
	signal G12446: std_logic; attribute dont_touch of G12446: signal is true;
	signal G12447: std_logic; attribute dont_touch of G12447: signal is true;
	signal G12448: std_logic; attribute dont_touch of G12448: signal is true;
	signal G12449: std_logic; attribute dont_touch of G12449: signal is true;
	signal G12450: std_logic; attribute dont_touch of G12450: signal is true;
	signal G12451: std_logic; attribute dont_touch of G12451: signal is true;
	signal G12452: std_logic; attribute dont_touch of G12452: signal is true;
	signal G12453: std_logic; attribute dont_touch of G12453: signal is true;
	signal G12454: std_logic; attribute dont_touch of G12454: signal is true;
	signal G12455: std_logic; attribute dont_touch of G12455: signal is true;
	signal G12456: std_logic; attribute dont_touch of G12456: signal is true;
	signal G12457: std_logic; attribute dont_touch of G12457: signal is true;
	signal G12460: std_logic; attribute dont_touch of G12460: signal is true;
	signal G12461: std_logic; attribute dont_touch of G12461: signal is true;
	signal G12462: std_logic; attribute dont_touch of G12462: signal is true;
	signal G12463: std_logic; attribute dont_touch of G12463: signal is true;
	signal G12466: std_logic; attribute dont_touch of G12466: signal is true;
	signal G12467: std_logic; attribute dont_touch of G12467: signal is true;
	signal G12470: std_logic; attribute dont_touch of G12470: signal is true;
	signal G12471: std_logic; attribute dont_touch of G12471: signal is true;
	signal G12472: std_logic; attribute dont_touch of G12472: signal is true;
	signal G12473: std_logic; attribute dont_touch of G12473: signal is true;
	signal G12476: std_logic; attribute dont_touch of G12476: signal is true;
	signal G12477: std_logic; attribute dont_touch of G12477: signal is true;
	signal G12478: std_logic; attribute dont_touch of G12478: signal is true;
	signal G12481: std_logic; attribute dont_touch of G12481: signal is true;
	signal G12482: std_logic; attribute dont_touch of G12482: signal is true;
	signal G12485: std_logic; attribute dont_touch of G12485: signal is true;
	signal G12486: std_logic; attribute dont_touch of G12486: signal is true;
	signal G12487: std_logic; attribute dont_touch of G12487: signal is true;
	signal G12490: std_logic; attribute dont_touch of G12490: signal is true;
	signal G12493: std_logic; attribute dont_touch of G12493: signal is true;
	signal G12494: std_logic; attribute dont_touch of G12494: signal is true;
	signal G12495: std_logic; attribute dont_touch of G12495: signal is true;
	signal G12498: std_logic; attribute dont_touch of G12498: signal is true;
	signal G12499: std_logic; attribute dont_touch of G12499: signal is true;
	signal G12502: std_logic; attribute dont_touch of G12502: signal is true;
	signal G12503: std_logic; attribute dont_touch of G12503: signal is true;
	signal G12504: std_logic; attribute dont_touch of G12504: signal is true;
	signal G12505: std_logic; attribute dont_touch of G12505: signal is true;
	signal G12506: std_logic; attribute dont_touch of G12506: signal is true;
	signal G12507: std_logic; attribute dont_touch of G12507: signal is true;
	signal G12510: std_logic; attribute dont_touch of G12510: signal is true;
	signal G12513: std_logic; attribute dont_touch of G12513: signal is true;
	signal G12514: std_logic; attribute dont_touch of G12514: signal is true;
	signal G12515: std_logic; attribute dont_touch of G12515: signal is true;
	signal G12518: std_logic; attribute dont_touch of G12518: signal is true;
	signal G12519: std_logic; attribute dont_touch of G12519: signal is true;
	signal G12520: std_logic; attribute dont_touch of G12520: signal is true;
	signal G12521: std_logic; attribute dont_touch of G12521: signal is true;
	signal G12522: std_logic; attribute dont_touch of G12522: signal is true;
	signal G12523: std_logic; attribute dont_touch of G12523: signal is true;
	signal G12524: std_logic; attribute dont_touch of G12524: signal is true;
	signal G12527: std_logic; attribute dont_touch of G12527: signal is true;
	signal G12530: std_logic; attribute dont_touch of G12530: signal is true;
	signal G12531: std_logic; attribute dont_touch of G12531: signal is true;
	signal G12532: std_logic; attribute dont_touch of G12532: signal is true;
	signal G12533: std_logic; attribute dont_touch of G12533: signal is true;
	signal G12534: std_logic; attribute dont_touch of G12534: signal is true;
	signal G12535: std_logic; attribute dont_touch of G12535: signal is true;
	signal G12536: std_logic; attribute dont_touch of G12536: signal is true;
	signal G12537: std_logic; attribute dont_touch of G12537: signal is true;
	signal G12538: std_logic; attribute dont_touch of G12538: signal is true;
	signal G12539: std_logic; attribute dont_touch of G12539: signal is true;
	signal G12542: std_logic; attribute dont_touch of G12542: signal is true;
	signal G12543: std_logic; attribute dont_touch of G12543: signal is true;
	signal G12544: std_logic; attribute dont_touch of G12544: signal is true;
	signal G12545: std_logic; attribute dont_touch of G12545: signal is true;
	signal G12546: std_logic; attribute dont_touch of G12546: signal is true;
	signal G12547: std_logic; attribute dont_touch of G12547: signal is true;
	signal G12548: std_logic; attribute dont_touch of G12548: signal is true;
	signal G12551: std_logic; attribute dont_touch of G12551: signal is true;
	signal G12552: std_logic; attribute dont_touch of G12552: signal is true;
	signal G12553: std_logic; attribute dont_touch of G12553: signal is true;
	signal G12554: std_logic; attribute dont_touch of G12554: signal is true;
	signal G12555: std_logic; attribute dont_touch of G12555: signal is true;
	signal G12558: std_logic; attribute dont_touch of G12558: signal is true;
	signal G12559: std_logic; attribute dont_touch of G12559: signal is true;
	signal G12560: std_logic; attribute dont_touch of G12560: signal is true;
	signal G12561: std_logic; attribute dont_touch of G12561: signal is true;
	signal G12564: std_logic; attribute dont_touch of G12564: signal is true;
	signal G12565: std_logic; attribute dont_touch of G12565: signal is true;
	signal G12596: std_logic; attribute dont_touch of G12596: signal is true;
	signal G12597: std_logic; attribute dont_touch of G12597: signal is true;
	signal G12598: std_logic; attribute dont_touch of G12598: signal is true;
	signal G12599: std_logic; attribute dont_touch of G12599: signal is true;
	signal G12600: std_logic; attribute dont_touch of G12600: signal is true;
	signal G12601: std_logic; attribute dont_touch of G12601: signal is true;
	signal G12604: std_logic; attribute dont_touch of G12604: signal is true;
	signal G12607: std_logic; attribute dont_touch of G12607: signal is true;
	signal G12608: std_logic; attribute dont_touch of G12608: signal is true;
	signal G12611: std_logic; attribute dont_touch of G12611: signal is true;
	signal G12642: std_logic; attribute dont_touch of G12642: signal is true;
	signal G12643: std_logic; attribute dont_touch of G12643: signal is true;
	signal G12644: std_logic; attribute dont_touch of G12644: signal is true;
	signal G12645: std_logic; attribute dont_touch of G12645: signal is true;
	signal G12646: std_logic; attribute dont_touch of G12646: signal is true;
	signal G12647: std_logic; attribute dont_touch of G12647: signal is true;
	signal G12650: std_logic; attribute dont_touch of G12650: signal is true;
	signal G12651: std_logic; attribute dont_touch of G12651: signal is true;
	signal G12654: std_logic; attribute dont_touch of G12654: signal is true;
	signal G12657: std_logic; attribute dont_touch of G12657: signal is true;
	signal G12688: std_logic; attribute dont_touch of G12688: signal is true;
	signal G12689: std_logic; attribute dont_touch of G12689: signal is true;
	signal G12690: std_logic; attribute dont_touch of G12690: signal is true;
	signal G12691: std_logic; attribute dont_touch of G12691: signal is true;
	signal G12692: std_logic; attribute dont_touch of G12692: signal is true;
	signal G12695: std_logic; attribute dont_touch of G12695: signal is true;
	signal G12698: std_logic; attribute dont_touch of G12698: signal is true;
	signal G12699: std_logic; attribute dont_touch of G12699: signal is true;
	signal G12702: std_logic; attribute dont_touch of G12702: signal is true;
	signal G12705: std_logic; attribute dont_touch of G12705: signal is true;
	signal G12708: std_logic; attribute dont_touch of G12708: signal is true;
	signal G12711: std_logic; attribute dont_touch of G12711: signal is true;
	signal G12742: std_logic; attribute dont_touch of G12742: signal is true;
	signal G12743: std_logic; attribute dont_touch of G12743: signal is true;
	signal G12744: std_logic; attribute dont_touch of G12744: signal is true;
	signal G12747: std_logic; attribute dont_touch of G12747: signal is true;
	signal G12748: std_logic; attribute dont_touch of G12748: signal is true;
	signal G12749: std_logic; attribute dont_touch of G12749: signal is true;
	signal G12752: std_logic; attribute dont_touch of G12752: signal is true;
	signal G12755: std_logic; attribute dont_touch of G12755: signal is true;
	signal G12756: std_logic; attribute dont_touch of G12756: signal is true;
	signal G12759: std_logic; attribute dont_touch of G12759: signal is true;
	signal G12762: std_logic; attribute dont_touch of G12762: signal is true;
	signal G12765: std_logic; attribute dont_touch of G12765: signal is true;
	signal G12768: std_logic; attribute dont_touch of G12768: signal is true;
	signal G12769: std_logic; attribute dont_touch of G12769: signal is true;
	signal G12772: std_logic; attribute dont_touch of G12772: signal is true;
	signal G12775: std_logic; attribute dont_touch of G12775: signal is true;
	signal G12776: std_logic; attribute dont_touch of G12776: signal is true;
	signal G12780: std_logic; attribute dont_touch of G12780: signal is true;
	signal G12781: std_logic; attribute dont_touch of G12781: signal is true;
	signal G12782: std_logic; attribute dont_touch of G12782: signal is true;
	signal G12783: std_logic; attribute dont_touch of G12783: signal is true;
	signal G12786: std_logic; attribute dont_touch of G12786: signal is true;
	signal G12789: std_logic; attribute dont_touch of G12789: signal is true;
	signal G12790: std_logic; attribute dont_touch of G12790: signal is true;
	signal G12791: std_logic; attribute dont_touch of G12791: signal is true;
	signal G12794: std_logic; attribute dont_touch of G12794: signal is true;
	signal G12797: std_logic; attribute dont_touch of G12797: signal is true;
	signal G12798: std_logic; attribute dont_touch of G12798: signal is true;
	signal G12801: std_logic; attribute dont_touch of G12801: signal is true;
	signal G12804: std_logic; attribute dont_touch of G12804: signal is true;
	signal G12807: std_logic; attribute dont_touch of G12807: signal is true;
	signal G12808: std_logic; attribute dont_touch of G12808: signal is true;
	signal G12811: std_logic; attribute dont_touch of G12811: signal is true;
	signal G12814: std_logic; attribute dont_touch of G12814: signal is true;
	signal G12815: std_logic; attribute dont_touch of G12815: signal is true;
	signal G12816: std_logic; attribute dont_touch of G12816: signal is true;
	signal G12819: std_logic; attribute dont_touch of G12819: signal is true;
	signal G12820: std_logic; attribute dont_touch of G12820: signal is true;
	signal G12821: std_logic; attribute dont_touch of G12821: signal is true;
	signal G12822: std_logic; attribute dont_touch of G12822: signal is true;
	signal G12825: std_logic; attribute dont_touch of G12825: signal is true;
	signal G12828: std_logic; attribute dont_touch of G12828: signal is true;
	signal G12829: std_logic; attribute dont_touch of G12829: signal is true;
	signal G12830: std_logic; attribute dont_touch of G12830: signal is true;
	signal G12833: std_logic; attribute dont_touch of G12833: signal is true;
	signal G12836: std_logic; attribute dont_touch of G12836: signal is true;
	signal G12837: std_logic; attribute dont_touch of G12837: signal is true;
	signal G12840: std_logic; attribute dont_touch of G12840: signal is true;
	signal G12843: std_logic; attribute dont_touch of G12843: signal is true;
	signal G12844: std_logic; attribute dont_touch of G12844: signal is true;
	signal G12847: std_logic; attribute dont_touch of G12847: signal is true;
	signal G12848: std_logic; attribute dont_touch of G12848: signal is true;
	signal G12849: std_logic; attribute dont_touch of G12849: signal is true;
	signal G12850: std_logic; attribute dont_touch of G12850: signal is true;
	signal G12851: std_logic; attribute dont_touch of G12851: signal is true;
	signal G12852: std_logic; attribute dont_touch of G12852: signal is true;
	signal G12853: std_logic; attribute dont_touch of G12853: signal is true;
	signal G12854: std_logic; attribute dont_touch of G12854: signal is true;
	signal G12857: std_logic; attribute dont_touch of G12857: signal is true;
	signal G12858: std_logic; attribute dont_touch of G12858: signal is true;
	signal G12859: std_logic; attribute dont_touch of G12859: signal is true;
	signal G12860: std_logic; attribute dont_touch of G12860: signal is true;
	signal G12863: std_logic; attribute dont_touch of G12863: signal is true;
	signal G12866: std_logic; attribute dont_touch of G12866: signal is true;
	signal G12867: std_logic; attribute dont_touch of G12867: signal is true;
	signal G12868: std_logic; attribute dont_touch of G12868: signal is true;
	signal G12871: std_logic; attribute dont_touch of G12871: signal is true;
	signal G12874: std_logic; attribute dont_touch of G12874: signal is true;
	signal G12875: std_logic; attribute dont_touch of G12875: signal is true;
	signal G12876: std_logic; attribute dont_touch of G12876: signal is true;
	signal G12880: std_logic; attribute dont_touch of G12880: signal is true;
	signal G12881: std_logic; attribute dont_touch of G12881: signal is true;
	signal G12882: std_logic; attribute dont_touch of G12882: signal is true;
	signal G12883: std_logic; attribute dont_touch of G12883: signal is true;
	signal G12886: std_logic; attribute dont_touch of G12886: signal is true;
	signal G12890: std_logic; attribute dont_touch of G12890: signal is true;
	signal G12891: std_logic; attribute dont_touch of G12891: signal is true;
	signal G12892: std_logic; attribute dont_touch of G12892: signal is true;
	signal G12893: std_logic; attribute dont_touch of G12893: signal is true;
	signal G12894: std_logic; attribute dont_touch of G12894: signal is true;
	signal G12895: std_logic; attribute dont_touch of G12895: signal is true;
	signal G12898: std_logic; attribute dont_touch of G12898: signal is true;
	signal G12899: std_logic; attribute dont_touch of G12899: signal is true;
	signal G12900: std_logic; attribute dont_touch of G12900: signal is true;
	signal G12901: std_logic; attribute dont_touch of G12901: signal is true;
	signal G12904: std_logic; attribute dont_touch of G12904: signal is true;
	signal G12907: std_logic; attribute dont_touch of G12907: signal is true;
	signal G12908: std_logic; attribute dont_touch of G12908: signal is true;
	signal G12909: std_logic; attribute dont_touch of G12909: signal is true;
	signal G12912: std_logic; attribute dont_touch of G12912: signal is true;
	signal G12913: std_logic; attribute dont_touch of G12913: signal is true;
	signal G12914: std_logic; attribute dont_touch of G12914: signal is true;
	signal G12915: std_logic; attribute dont_touch of G12915: signal is true;
	signal G12916: std_logic; attribute dont_touch of G12916: signal is true;
	signal G12920: std_logic; attribute dont_touch of G12920: signal is true;
	signal G12921: std_logic; attribute dont_touch of G12921: signal is true;
	signal G12922: std_logic; attribute dont_touch of G12922: signal is true;
	signal G12923: std_logic; attribute dont_touch of G12923: signal is true;
	signal G12926: std_logic; attribute dont_touch of G12926: signal is true;
	signal G12930: std_logic; attribute dont_touch of G12930: signal is true;
	signal G12931: std_logic; attribute dont_touch of G12931: signal is true;
	signal G12932: std_logic; attribute dont_touch of G12932: signal is true;
	signal G12933: std_logic; attribute dont_touch of G12933: signal is true;
	signal G12934: std_logic; attribute dont_touch of G12934: signal is true;
	signal G12935: std_logic; attribute dont_touch of G12935: signal is true;
	signal G12938: std_logic; attribute dont_touch of G12938: signal is true;
	signal G12939: std_logic; attribute dont_touch of G12939: signal is true;
	signal G12940: std_logic; attribute dont_touch of G12940: signal is true;
	signal G12941: std_logic; attribute dont_touch of G12941: signal is true;
	signal G12942: std_logic; attribute dont_touch of G12942: signal is true;
	signal G12943: std_logic; attribute dont_touch of G12943: signal is true;
	signal G12944: std_logic; attribute dont_touch of G12944: signal is true;
	signal G12945: std_logic; attribute dont_touch of G12945: signal is true;
	signal G12949: std_logic; attribute dont_touch of G12949: signal is true;
	signal G12950: std_logic; attribute dont_touch of G12950: signal is true;
	signal G12951: std_logic; attribute dont_touch of G12951: signal is true;
	signal G12952: std_logic; attribute dont_touch of G12952: signal is true;
	signal G12955: std_logic; attribute dont_touch of G12955: signal is true;
	signal G12959: std_logic; attribute dont_touch of G12959: signal is true;
	signal G12960: std_logic; attribute dont_touch of G12960: signal is true;
	signal G12961: std_logic; attribute dont_touch of G12961: signal is true;
	signal G12962: std_logic; attribute dont_touch of G12962: signal is true;
	signal G12965: std_logic; attribute dont_touch of G12965: signal is true;
	signal G12966: std_logic; attribute dont_touch of G12966: signal is true;
	signal G12967: std_logic; attribute dont_touch of G12967: signal is true;
	signal G12968: std_logic; attribute dont_touch of G12968: signal is true;
	signal G12969: std_logic; attribute dont_touch of G12969: signal is true;
	signal G12970: std_logic; attribute dont_touch of G12970: signal is true;
	signal G12971: std_logic; attribute dont_touch of G12971: signal is true;
	signal G12972: std_logic; attribute dont_touch of G12972: signal is true;
	signal G12973: std_logic; attribute dont_touch of G12973: signal is true;
	signal G12974: std_logic; attribute dont_touch of G12974: signal is true;
	signal G12978: std_logic; attribute dont_touch of G12978: signal is true;
	signal G12979: std_logic; attribute dont_touch of G12979: signal is true;
	signal G12980: std_logic; attribute dont_touch of G12980: signal is true;
	signal G12981: std_logic; attribute dont_touch of G12981: signal is true;
	signal G12984: std_logic; attribute dont_touch of G12984: signal is true;
	signal G12988: std_logic; attribute dont_touch of G12988: signal is true;
	signal G12989: std_logic; attribute dont_touch of G12989: signal is true;
	signal G12990: std_logic; attribute dont_touch of G12990: signal is true;
	signal G12991: std_logic; attribute dont_touch of G12991: signal is true;
	signal G12992: std_logic; attribute dont_touch of G12992: signal is true;
	signal G12993: std_logic; attribute dont_touch of G12993: signal is true;
	signal G12994: std_logic; attribute dont_touch of G12994: signal is true;
	signal G12995: std_logic; attribute dont_touch of G12995: signal is true;
	signal G12996: std_logic; attribute dont_touch of G12996: signal is true;
	signal G12997: std_logic; attribute dont_touch of G12997: signal is true;
	signal G12998: std_logic; attribute dont_touch of G12998: signal is true;
	signal G12999: std_logic; attribute dont_touch of G12999: signal is true;
	signal G13000: std_logic; attribute dont_touch of G13000: signal is true;
	signal G13001: std_logic; attribute dont_touch of G13001: signal is true;
	signal G13002: std_logic; attribute dont_touch of G13002: signal is true;
	signal G13003: std_logic; attribute dont_touch of G13003: signal is true;
	signal G13004: std_logic; attribute dont_touch of G13004: signal is true;
	signal G13009: std_logic; attribute dont_touch of G13009: signal is true;
	signal G13010: std_logic; attribute dont_touch of G13010: signal is true;
	signal G13011: std_logic; attribute dont_touch of G13011: signal is true;
	signal G13020: std_logic; attribute dont_touch of G13020: signal is true;
	signal G13021: std_logic; attribute dont_touch of G13021: signal is true;
	signal G13022: std_logic; attribute dont_touch of G13022: signal is true;
	signal G13023: std_logic; attribute dont_touch of G13023: signal is true;
	signal G13024: std_logic; attribute dont_touch of G13024: signal is true;
	signal G13025: std_logic; attribute dont_touch of G13025: signal is true;
	signal G13026: std_logic; attribute dont_touch of G13026: signal is true;
	signal G13027: std_logic; attribute dont_touch of G13027: signal is true;
	signal G13028: std_logic; attribute dont_touch of G13028: signal is true;
	signal G13029: std_logic; attribute dont_touch of G13029: signal is true;
	signal G13030: std_logic; attribute dont_touch of G13030: signal is true;
	signal G13031: std_logic; attribute dont_touch of G13031: signal is true;
	signal G13032: std_logic; attribute dont_touch of G13032: signal is true;
	signal G13033: std_logic; attribute dont_touch of G13033: signal is true;
	signal G13034: std_logic; attribute dont_touch of G13034: signal is true;
	signal G13035: std_logic; attribute dont_touch of G13035: signal is true;
	signal G13036: std_logic; attribute dont_touch of G13036: signal is true;
	signal G13037: std_logic; attribute dont_touch of G13037: signal is true;
	signal G13038: std_logic; attribute dont_touch of G13038: signal is true;
	signal G13039: std_logic; attribute dont_touch of G13039: signal is true;
	signal G13040: std_logic; attribute dont_touch of G13040: signal is true;
	signal G13041: std_logic; attribute dont_touch of G13041: signal is true;
	signal G13042: std_logic; attribute dont_touch of G13042: signal is true;
	signal G13043: std_logic; attribute dont_touch of G13043: signal is true;
	signal G13044: std_logic; attribute dont_touch of G13044: signal is true;
	signal G13045: std_logic; attribute dont_touch of G13045: signal is true;
	signal G13046: std_logic; attribute dont_touch of G13046: signal is true;
	signal G13047: std_logic; attribute dont_touch of G13047: signal is true;
	signal G13048: std_logic; attribute dont_touch of G13048: signal is true;
	signal G13049: std_logic; attribute dont_touch of G13049: signal is true;
	signal G13050: std_logic; attribute dont_touch of G13050: signal is true;
	signal G13051: std_logic; attribute dont_touch of G13051: signal is true;
	signal G13052: std_logic; attribute dont_touch of G13052: signal is true;
	signal G13053: std_logic; attribute dont_touch of G13053: signal is true;
	signal G13054: std_logic; attribute dont_touch of G13054: signal is true;
	signal G13055: std_logic; attribute dont_touch of G13055: signal is true;
	signal G13056: std_logic; attribute dont_touch of G13056: signal is true;
	signal G13057: std_logic; attribute dont_touch of G13057: signal is true;
	signal G13058: std_logic; attribute dont_touch of G13058: signal is true;
	signal G13059: std_logic; attribute dont_touch of G13059: signal is true;
	signal G13060: std_logic; attribute dont_touch of G13060: signal is true;
	signal G13061: std_logic; attribute dont_touch of G13061: signal is true;
	signal G13062: std_logic; attribute dont_touch of G13062: signal is true;
	signal G13063: std_logic; attribute dont_touch of G13063: signal is true;
	signal G13064: std_logic; attribute dont_touch of G13064: signal is true;
	signal G13065: std_logic; attribute dont_touch of G13065: signal is true;
	signal G13066: std_logic; attribute dont_touch of G13066: signal is true;
	signal G13067: std_logic; attribute dont_touch of G13067: signal is true;
	signal G13068: std_logic; attribute dont_touch of G13068: signal is true;
	signal G13069: std_logic; attribute dont_touch of G13069: signal is true;
	signal G13070: std_logic; attribute dont_touch of G13070: signal is true;
	signal G13071: std_logic; attribute dont_touch of G13071: signal is true;
	signal G13072: std_logic; attribute dont_touch of G13072: signal is true;
	signal G13073: std_logic; attribute dont_touch of G13073: signal is true;
	signal G13074: std_logic; attribute dont_touch of G13074: signal is true;
	signal G13075: std_logic; attribute dont_touch of G13075: signal is true;
	signal G13076: std_logic; attribute dont_touch of G13076: signal is true;
	signal G13077: std_logic; attribute dont_touch of G13077: signal is true;
	signal G13078: std_logic; attribute dont_touch of G13078: signal is true;
	signal G13079: std_logic; attribute dont_touch of G13079: signal is true;
	signal G13080: std_logic; attribute dont_touch of G13080: signal is true;
	signal G13081: std_logic; attribute dont_touch of G13081: signal is true;
	signal G13082: std_logic; attribute dont_touch of G13082: signal is true;
	signal G13087: std_logic; attribute dont_touch of G13087: signal is true;
	signal G13088: std_logic; attribute dont_touch of G13088: signal is true;
	signal G13089: std_logic; attribute dont_touch of G13089: signal is true;
	signal G13090: std_logic; attribute dont_touch of G13090: signal is true;
	signal G13091: std_logic; attribute dont_touch of G13091: signal is true;
	signal G13092: std_logic; attribute dont_touch of G13092: signal is true;
	signal G13093: std_logic; attribute dont_touch of G13093: signal is true;
	signal G13094: std_logic; attribute dont_touch of G13094: signal is true;
	signal G13095: std_logic; attribute dont_touch of G13095: signal is true;
	signal G13096: std_logic; attribute dont_touch of G13096: signal is true;
	signal G13097: std_logic; attribute dont_touch of G13097: signal is true;
	signal G13098: std_logic; attribute dont_touch of G13098: signal is true;
	signal G13099: std_logic; attribute dont_touch of G13099: signal is true;
	signal G13100: std_logic; attribute dont_touch of G13100: signal is true;
	signal G13101: std_logic; attribute dont_touch of G13101: signal is true;
	signal G13102: std_logic; attribute dont_touch of G13102: signal is true;
	signal G13103: std_logic; attribute dont_touch of G13103: signal is true;
	signal G13104: std_logic; attribute dont_touch of G13104: signal is true;
	signal G13105: std_logic; attribute dont_touch of G13105: signal is true;
	signal G13106: std_logic; attribute dont_touch of G13106: signal is true;
	signal G13107: std_logic; attribute dont_touch of G13107: signal is true;
	signal G13108: std_logic; attribute dont_touch of G13108: signal is true;
	signal G13109: std_logic; attribute dont_touch of G13109: signal is true;
	signal G13110: std_logic; attribute dont_touch of G13110: signal is true;
	signal G13111: std_logic; attribute dont_touch of G13111: signal is true;
	signal G13112: std_logic; attribute dont_touch of G13112: signal is true;
	signal G13113: std_logic; attribute dont_touch of G13113: signal is true;
	signal G13114: std_logic; attribute dont_touch of G13114: signal is true;
	signal G13115: std_logic; attribute dont_touch of G13115: signal is true;
	signal G13116: std_logic; attribute dont_touch of G13116: signal is true;
	signal G13117: std_logic; attribute dont_touch of G13117: signal is true;
	signal G13118: std_logic; attribute dont_touch of G13118: signal is true;
	signal G13119: std_logic; attribute dont_touch of G13119: signal is true;
	signal G13120: std_logic; attribute dont_touch of G13120: signal is true;
	signal G13121: std_logic; attribute dont_touch of G13121: signal is true;
	signal G13122: std_logic; attribute dont_touch of G13122: signal is true;
	signal G13123: std_logic; attribute dont_touch of G13123: signal is true;
	signal G13124: std_logic; attribute dont_touch of G13124: signal is true;
	signal G13125: std_logic; attribute dont_touch of G13125: signal is true;
	signal G13126: std_logic; attribute dont_touch of G13126: signal is true;
	signal G13127: std_logic; attribute dont_touch of G13127: signal is true;
	signal G13128: std_logic; attribute dont_touch of G13128: signal is true;
	signal G13129: std_logic; attribute dont_touch of G13129: signal is true;
	signal G13130: std_logic; attribute dont_touch of G13130: signal is true;
	signal G13131: std_logic; attribute dont_touch of G13131: signal is true;
	signal G13132: std_logic; attribute dont_touch of G13132: signal is true;
	signal G13133: std_logic; attribute dont_touch of G13133: signal is true;
	signal G13134: std_logic; attribute dont_touch of G13134: signal is true;
	signal G13135: std_logic; attribute dont_touch of G13135: signal is true;
	signal G13136: std_logic; attribute dont_touch of G13136: signal is true;
	signal G13137: std_logic; attribute dont_touch of G13137: signal is true;
	signal G13138: std_logic; attribute dont_touch of G13138: signal is true;
	signal G13139: std_logic; attribute dont_touch of G13139: signal is true;
	signal G13140: std_logic; attribute dont_touch of G13140: signal is true;
	signal G13141: std_logic; attribute dont_touch of G13141: signal is true;
	signal G13142: std_logic; attribute dont_touch of G13142: signal is true;
	signal G13143: std_logic; attribute dont_touch of G13143: signal is true;
	signal G13144: std_logic; attribute dont_touch of G13144: signal is true;
	signal G13145: std_logic; attribute dont_touch of G13145: signal is true;
	signal G13146: std_logic; attribute dont_touch of G13146: signal is true;
	signal G13147: std_logic; attribute dont_touch of G13147: signal is true;
	signal G13148: std_logic; attribute dont_touch of G13148: signal is true;
	signal G13149: std_logic; attribute dont_touch of G13149: signal is true;
	signal G13150: std_logic; attribute dont_touch of G13150: signal is true;
	signal G13151: std_logic; attribute dont_touch of G13151: signal is true;
	signal G13152: std_logic; attribute dont_touch of G13152: signal is true;
	signal G13153: std_logic; attribute dont_touch of G13153: signal is true;
	signal G13154: std_logic; attribute dont_touch of G13154: signal is true;
	signal G13155: std_logic; attribute dont_touch of G13155: signal is true;
	signal G13156: std_logic; attribute dont_touch of G13156: signal is true;
	signal G13157: std_logic; attribute dont_touch of G13157: signal is true;
	signal G13158: std_logic; attribute dont_touch of G13158: signal is true;
	signal G13159: std_logic; attribute dont_touch of G13159: signal is true;
	signal G13160: std_logic; attribute dont_touch of G13160: signal is true;
	signal G13161: std_logic; attribute dont_touch of G13161: signal is true;
	signal G13162: std_logic; attribute dont_touch of G13162: signal is true;
	signal G13163: std_logic; attribute dont_touch of G13163: signal is true;
	signal G13164: std_logic; attribute dont_touch of G13164: signal is true;
	signal G13165: std_logic; attribute dont_touch of G13165: signal is true;
	signal G13166: std_logic; attribute dont_touch of G13166: signal is true;
	signal G13167: std_logic; attribute dont_touch of G13167: signal is true;
	signal G13168: std_logic; attribute dont_touch of G13168: signal is true;
	signal G13169: std_logic; attribute dont_touch of G13169: signal is true;
	signal G13170: std_logic; attribute dont_touch of G13170: signal is true;
	signal G13171: std_logic; attribute dont_touch of G13171: signal is true;
	signal G13172: std_logic; attribute dont_touch of G13172: signal is true;
	signal G13173: std_logic; attribute dont_touch of G13173: signal is true;
	signal G13174: std_logic; attribute dont_touch of G13174: signal is true;
	signal G13175: std_logic; attribute dont_touch of G13175: signal is true;
	signal G13176: std_logic; attribute dont_touch of G13176: signal is true;
	signal G13177: std_logic; attribute dont_touch of G13177: signal is true;
	signal G13178: std_logic; attribute dont_touch of G13178: signal is true;
	signal G13179: std_logic; attribute dont_touch of G13179: signal is true;
	signal G13180: std_logic; attribute dont_touch of G13180: signal is true;
	signal G13181: std_logic; attribute dont_touch of G13181: signal is true;
	signal G13182: std_logic; attribute dont_touch of G13182: signal is true;
	signal G13183: std_logic; attribute dont_touch of G13183: signal is true;
	signal G13184: std_logic; attribute dont_touch of G13184: signal is true;
	signal G13185: std_logic; attribute dont_touch of G13185: signal is true;
	signal G13186: std_logic; attribute dont_touch of G13186: signal is true;
	signal G13187: std_logic; attribute dont_touch of G13187: signal is true;
	signal G13188: std_logic; attribute dont_touch of G13188: signal is true;
	signal G13189: std_logic; attribute dont_touch of G13189: signal is true;
	signal G13190: std_logic; attribute dont_touch of G13190: signal is true;
	signal G13191: std_logic; attribute dont_touch of G13191: signal is true;
	signal G13192: std_logic; attribute dont_touch of G13192: signal is true;
	signal G13193: std_logic; attribute dont_touch of G13193: signal is true;
	signal G13194: std_logic; attribute dont_touch of G13194: signal is true;
	signal G13195: std_logic; attribute dont_touch of G13195: signal is true;
	signal G13196: std_logic; attribute dont_touch of G13196: signal is true;
	signal G13197: std_logic; attribute dont_touch of G13197: signal is true;
	signal G13198: std_logic; attribute dont_touch of G13198: signal is true;
	signal G13199: std_logic; attribute dont_touch of G13199: signal is true;
	signal G13200: std_logic; attribute dont_touch of G13200: signal is true;
	signal G13201: std_logic; attribute dont_touch of G13201: signal is true;
	signal G13202: std_logic; attribute dont_touch of G13202: signal is true;
	signal G13203: std_logic; attribute dont_touch of G13203: signal is true;
	signal G13204: std_logic; attribute dont_touch of G13204: signal is true;
	signal G13205: std_logic; attribute dont_touch of G13205: signal is true;
	signal G13206: std_logic; attribute dont_touch of G13206: signal is true;
	signal G13207: std_logic; attribute dont_touch of G13207: signal is true;
	signal G13208: std_logic; attribute dont_touch of G13208: signal is true;
	signal G13209: std_logic; attribute dont_touch of G13209: signal is true;
	signal G13210: std_logic; attribute dont_touch of G13210: signal is true;
	signal G13211: std_logic; attribute dont_touch of G13211: signal is true;
	signal G13212: std_logic; attribute dont_touch of G13212: signal is true;
	signal G13213: std_logic; attribute dont_touch of G13213: signal is true;
	signal G13214: std_logic; attribute dont_touch of G13214: signal is true;
	signal G13215: std_logic; attribute dont_touch of G13215: signal is true;
	signal G13218: std_logic; attribute dont_touch of G13218: signal is true;
	signal G13219: std_logic; attribute dont_touch of G13219: signal is true;
	signal G13220: std_logic; attribute dont_touch of G13220: signal is true;
	signal G13221: std_logic; attribute dont_touch of G13221: signal is true;
	signal G13222: std_logic; attribute dont_touch of G13222: signal is true;
	signal G13223: std_logic; attribute dont_touch of G13223: signal is true;
	signal G13224: std_logic; attribute dont_touch of G13224: signal is true;
	signal G13225: std_logic; attribute dont_touch of G13225: signal is true;
	signal G13226: std_logic; attribute dont_touch of G13226: signal is true;
	signal G13227: std_logic; attribute dont_touch of G13227: signal is true;
	signal G13228: std_logic; attribute dont_touch of G13228: signal is true;
	signal G13229: std_logic; attribute dont_touch of G13229: signal is true;
	signal G13232: std_logic; attribute dont_touch of G13232: signal is true;
	signal G13233: std_logic; attribute dont_touch of G13233: signal is true;
	signal G13234: std_logic; attribute dont_touch of G13234: signal is true;
	signal G13237: std_logic; attribute dont_touch of G13237: signal is true;
	signal G13238: std_logic; attribute dont_touch of G13238: signal is true;
	signal G13239: std_logic; attribute dont_touch of G13239: signal is true;
	signal G13240: std_logic; attribute dont_touch of G13240: signal is true;
	signal G13241: std_logic; attribute dont_touch of G13241: signal is true;
	signal G13242: std_logic; attribute dont_touch of G13242: signal is true;
	signal G13243: std_logic; attribute dont_touch of G13243: signal is true;
	signal G13244: std_logic; attribute dont_touch of G13244: signal is true;
	signal G13245: std_logic; attribute dont_touch of G13245: signal is true;
	signal G13246: std_logic; attribute dont_touch of G13246: signal is true;
	signal G13247: std_logic; attribute dont_touch of G13247: signal is true;
	signal G13248: std_logic; attribute dont_touch of G13248: signal is true;
	signal G13249: std_logic; attribute dont_touch of G13249: signal is true;
	signal G13250: std_logic; attribute dont_touch of G13250: signal is true;
	signal G13251: std_logic; attribute dont_touch of G13251: signal is true;
	signal G13252: std_logic; attribute dont_touch of G13252: signal is true;
	signal G13255: std_logic; attribute dont_touch of G13255: signal is true;
	signal G13256: std_logic; attribute dont_touch of G13256: signal is true;
	signal G13257: std_logic; attribute dont_touch of G13257: signal is true;
	signal G13260: std_logic; attribute dont_touch of G13260: signal is true;
	signal G13261: std_logic; attribute dont_touch of G13261: signal is true;
	signal G13262: std_logic; attribute dont_touch of G13262: signal is true;
	signal G13263: std_logic; attribute dont_touch of G13263: signal is true;
	signal G13264: std_logic; attribute dont_touch of G13264: signal is true;
	signal G13265: std_logic; attribute dont_touch of G13265: signal is true;
	signal G13266: std_logic; attribute dont_touch of G13266: signal is true;
	signal G13267: std_logic; attribute dont_touch of G13267: signal is true;
	signal G13268: std_logic; attribute dont_touch of G13268: signal is true;
	signal G13269: std_logic; attribute dont_touch of G13269: signal is true;
	signal G13270: std_logic; attribute dont_touch of G13270: signal is true;
	signal G13271: std_logic; attribute dont_touch of G13271: signal is true;
	signal G13272: std_logic; attribute dont_touch of G13272: signal is true;
	signal G13273: std_logic; attribute dont_touch of G13273: signal is true;
	signal G13274: std_logic; attribute dont_touch of G13274: signal is true;
	signal G13275: std_logic; attribute dont_touch of G13275: signal is true;
	signal G13278: std_logic; attribute dont_touch of G13278: signal is true;
	signal G13279: std_logic; attribute dont_touch of G13279: signal is true;
	signal G13280: std_logic; attribute dont_touch of G13280: signal is true;
	signal G13283: std_logic; attribute dont_touch of G13283: signal is true;
	signal G13284: std_logic; attribute dont_touch of G13284: signal is true;
	signal G13285: std_logic; attribute dont_touch of G13285: signal is true;
	signal G13286: std_logic; attribute dont_touch of G13286: signal is true;
	signal G13289: std_logic; attribute dont_touch of G13289: signal is true;
	signal G13290: std_logic; attribute dont_touch of G13290: signal is true;
	signal G13291: std_logic; attribute dont_touch of G13291: signal is true;
	signal G13292: std_logic; attribute dont_touch of G13292: signal is true;
	signal G13293: std_logic; attribute dont_touch of G13293: signal is true;
	signal G13294: std_logic; attribute dont_touch of G13294: signal is true;
	signal G13295: std_logic; attribute dont_touch of G13295: signal is true;
	signal G13296: std_logic; attribute dont_touch of G13296: signal is true;
	signal G13297: std_logic; attribute dont_touch of G13297: signal is true;
	signal G13298: std_logic; attribute dont_touch of G13298: signal is true;
	signal G13299: std_logic; attribute dont_touch of G13299: signal is true;
	signal G13300: std_logic; attribute dont_touch of G13300: signal is true;
	signal G13303: std_logic; attribute dont_touch of G13303: signal is true;
	signal G13304: std_logic; attribute dont_touch of G13304: signal is true;
	signal G13305: std_logic; attribute dont_touch of G13305: signal is true;
	signal G13308: std_logic; attribute dont_touch of G13308: signal is true;
	signal G13309: std_logic; attribute dont_touch of G13309: signal is true;
	signal G13310: std_logic; attribute dont_touch of G13310: signal is true;
	signal G13313: std_logic; attribute dont_touch of G13313: signal is true;
	signal G13316: std_logic; attribute dont_touch of G13316: signal is true;
	signal G13317: std_logic; attribute dont_touch of G13317: signal is true;
	signal G13318: std_logic; attribute dont_touch of G13318: signal is true;
	signal G13319: std_logic; attribute dont_touch of G13319: signal is true;
	signal G13320: std_logic; attribute dont_touch of G13320: signal is true;
	signal G13321: std_logic; attribute dont_touch of G13321: signal is true;
	signal G13322: std_logic; attribute dont_touch of G13322: signal is true;
	signal G13323: std_logic; attribute dont_touch of G13323: signal is true;
	signal G13324: std_logic; attribute dont_touch of G13324: signal is true;
	signal G13325: std_logic; attribute dont_touch of G13325: signal is true;
	signal G13326: std_logic; attribute dont_touch of G13326: signal is true;
	signal G13327: std_logic; attribute dont_touch of G13327: signal is true;
	signal G13328: std_logic; attribute dont_touch of G13328: signal is true;
	signal G13329: std_logic; attribute dont_touch of G13329: signal is true;
	signal G13330: std_logic; attribute dont_touch of G13330: signal is true;
	signal G13331: std_logic; attribute dont_touch of G13331: signal is true;
	signal G13332: std_logic; attribute dont_touch of G13332: signal is true;
	signal G13335: std_logic; attribute dont_touch of G13335: signal is true;
	signal G13336: std_logic; attribute dont_touch of G13336: signal is true;
	signal G13339: std_logic; attribute dont_touch of G13339: signal is true;
	signal G13340: std_logic; attribute dont_touch of G13340: signal is true;
	signal G13341: std_logic; attribute dont_touch of G13341: signal is true;
	signal G13342: std_logic; attribute dont_touch of G13342: signal is true;
	signal G13343: std_logic; attribute dont_touch of G13343: signal is true;
	signal G13344: std_logic; attribute dont_touch of G13344: signal is true;
	signal G13345: std_logic; attribute dont_touch of G13345: signal is true;
	signal G13346: std_logic; attribute dont_touch of G13346: signal is true;
	signal G13347: std_logic; attribute dont_touch of G13347: signal is true;
	signal G13348: std_logic; attribute dont_touch of G13348: signal is true;
	signal G13351: std_logic; attribute dont_touch of G13351: signal is true;
	signal G13352: std_logic; attribute dont_touch of G13352: signal is true;
	signal G13353: std_logic; attribute dont_touch of G13353: signal is true;
	signal G13354: std_logic; attribute dont_touch of G13354: signal is true;
	signal G13355: std_logic; attribute dont_touch of G13355: signal is true;
	signal G13356: std_logic; attribute dont_touch of G13356: signal is true;
	signal G13359: std_logic; attribute dont_touch of G13359: signal is true;
	signal G13360: std_logic; attribute dont_touch of G13360: signal is true;
	signal G13361: std_logic; attribute dont_touch of G13361: signal is true;
	signal G13364: std_logic; attribute dont_touch of G13364: signal is true;
	signal G13365: std_logic; attribute dont_touch of G13365: signal is true;
	signal G13366: std_logic; attribute dont_touch of G13366: signal is true;
	signal G13367: std_logic; attribute dont_touch of G13367: signal is true;
	signal G13368: std_logic; attribute dont_touch of G13368: signal is true;
	signal G13369: std_logic; attribute dont_touch of G13369: signal is true;
	signal G13370: std_logic; attribute dont_touch of G13370: signal is true;
	signal G13373: std_logic; attribute dont_touch of G13373: signal is true;
	signal G13374: std_logic; attribute dont_touch of G13374: signal is true;
	signal G13375: std_logic; attribute dont_touch of G13375: signal is true;
	signal G13378: std_logic; attribute dont_touch of G13378: signal is true;
	signal G13381: std_logic; attribute dont_touch of G13381: signal is true;
	signal G13384: std_logic; attribute dont_touch of G13384: signal is true;
	signal G13385: std_logic; attribute dont_touch of G13385: signal is true;
	signal G13386: std_logic; attribute dont_touch of G13386: signal is true;
	signal G13389: std_logic; attribute dont_touch of G13389: signal is true;
	signal G13390: std_logic; attribute dont_touch of G13390: signal is true;
	signal G13391: std_logic; attribute dont_touch of G13391: signal is true;
	signal G13394: std_logic; attribute dont_touch of G13394: signal is true;
	signal G13395: std_logic; attribute dont_touch of G13395: signal is true;
	signal G13396: std_logic; attribute dont_touch of G13396: signal is true;
	signal G13397: std_logic; attribute dont_touch of G13397: signal is true;
	signal G13398: std_logic; attribute dont_touch of G13398: signal is true;
	signal G13399: std_logic; attribute dont_touch of G13399: signal is true;
	signal G13400: std_logic; attribute dont_touch of G13400: signal is true;
	signal G13401: std_logic; attribute dont_touch of G13401: signal is true;
	signal G13404: std_logic; attribute dont_touch of G13404: signal is true;
	signal G13405: std_logic; attribute dont_touch of G13405: signal is true;
	signal G13406: std_logic; attribute dont_touch of G13406: signal is true;
	signal G13407: std_logic; attribute dont_touch of G13407: signal is true;
	signal G13408: std_logic; attribute dont_touch of G13408: signal is true;
	signal G13409: std_logic; attribute dont_touch of G13409: signal is true;
	signal G13410: std_logic; attribute dont_touch of G13410: signal is true;
	signal G13411: std_logic; attribute dont_touch of G13411: signal is true;
	signal G13412: std_logic; attribute dont_touch of G13412: signal is true;
	signal G13413: std_logic; attribute dont_touch of G13413: signal is true;
	signal G13414: std_logic; attribute dont_touch of G13414: signal is true;
	signal G13415: std_logic; attribute dont_touch of G13415: signal is true;
	signal G13416: std_logic; attribute dont_touch of G13416: signal is true;
	signal G13417: std_logic; attribute dont_touch of G13417: signal is true;
	signal G13418: std_logic; attribute dont_touch of G13418: signal is true;
	signal G13419: std_logic; attribute dont_touch of G13419: signal is true;
	signal G13420: std_logic; attribute dont_touch of G13420: signal is true;
	signal G13421: std_logic; attribute dont_touch of G13421: signal is true;
	signal G13422: std_logic; attribute dont_touch of G13422: signal is true;
	signal G13423: std_logic; attribute dont_touch of G13423: signal is true;
	signal G13424: std_logic; attribute dont_touch of G13424: signal is true;
	signal G13425: std_logic; attribute dont_touch of G13425: signal is true;
	signal G13426: std_logic; attribute dont_touch of G13426: signal is true;
	signal G13427: std_logic; attribute dont_touch of G13427: signal is true;
	signal G13428: std_logic; attribute dont_touch of G13428: signal is true;
	signal G13429: std_logic; attribute dont_touch of G13429: signal is true;
	signal G13430: std_logic; attribute dont_touch of G13430: signal is true;
	signal G13431: std_logic; attribute dont_touch of G13431: signal is true;
	signal G13432: std_logic; attribute dont_touch of G13432: signal is true;
	signal G13433: std_logic; attribute dont_touch of G13433: signal is true;
	signal G13434: std_logic; attribute dont_touch of G13434: signal is true;
	signal G13435: std_logic; attribute dont_touch of G13435: signal is true;
	signal G13436: std_logic; attribute dont_touch of G13436: signal is true;
	signal G13437: std_logic; attribute dont_touch of G13437: signal is true;
	signal G13438: std_logic; attribute dont_touch of G13438: signal is true;
	signal G13439: std_logic; attribute dont_touch of G13439: signal is true;
	signal G13440: std_logic; attribute dont_touch of G13440: signal is true;
	signal G13441: std_logic; attribute dont_touch of G13441: signal is true;
	signal G13442: std_logic; attribute dont_touch of G13442: signal is true;
	signal G13443: std_logic; attribute dont_touch of G13443: signal is true;
	signal G13444: std_logic; attribute dont_touch of G13444: signal is true;
	signal G13445: std_logic; attribute dont_touch of G13445: signal is true;
	signal G13446: std_logic; attribute dont_touch of G13446: signal is true;
	signal G13447: std_logic; attribute dont_touch of G13447: signal is true;
	signal G13448: std_logic; attribute dont_touch of G13448: signal is true;
	signal G13449: std_logic; attribute dont_touch of G13449: signal is true;
	signal G13450: std_logic; attribute dont_touch of G13450: signal is true;
	signal G13451: std_logic; attribute dont_touch of G13451: signal is true;
	signal G13452: std_logic; attribute dont_touch of G13452: signal is true;
	signal G13453: std_logic; attribute dont_touch of G13453: signal is true;
	signal G13454: std_logic; attribute dont_touch of G13454: signal is true;
	signal G13455: std_logic; attribute dont_touch of G13455: signal is true;
	signal G13456: std_logic; attribute dont_touch of G13456: signal is true;
	signal G13457: std_logic; attribute dont_touch of G13457: signal is true;
	signal G13458: std_logic; attribute dont_touch of G13458: signal is true;
	signal G13459: std_logic; attribute dont_touch of G13459: signal is true;
	signal G13460: std_logic; attribute dont_touch of G13460: signal is true;
	signal G13461: std_logic; attribute dont_touch of G13461: signal is true;
	signal G13462: std_logic; attribute dont_touch of G13462: signal is true;
	signal G13463: std_logic; attribute dont_touch of G13463: signal is true;
	signal G13464: std_logic; attribute dont_touch of G13464: signal is true;
	signal G13465: std_logic; attribute dont_touch of G13465: signal is true;
	signal G13466: std_logic; attribute dont_touch of G13466: signal is true;
	signal G13467: std_logic; attribute dont_touch of G13467: signal is true;
	signal G13468: std_logic; attribute dont_touch of G13468: signal is true;
	signal G13469: std_logic; attribute dont_touch of G13469: signal is true;
	signal G13475: std_logic; attribute dont_touch of G13475: signal is true;
	signal G13476: std_logic; attribute dont_touch of G13476: signal is true;
	signal G13477: std_logic; attribute dont_touch of G13477: signal is true;
	signal G13478: std_logic; attribute dont_touch of G13478: signal is true;
	signal G13479: std_logic; attribute dont_touch of G13479: signal is true;
	signal G13480: std_logic; attribute dont_touch of G13480: signal is true;
	signal G13481: std_logic; attribute dont_touch of G13481: signal is true;
	signal G13482: std_logic; attribute dont_touch of G13482: signal is true;
	signal G13483: std_logic; attribute dont_touch of G13483: signal is true;
	signal G13484: std_logic; attribute dont_touch of G13484: signal is true;
	signal G13485: std_logic; attribute dont_touch of G13485: signal is true;
	signal G13486: std_logic; attribute dont_touch of G13486: signal is true;
	signal G13487: std_logic; attribute dont_touch of G13487: signal is true;
	signal G13488: std_logic; attribute dont_touch of G13488: signal is true;
	signal G13489: std_logic; attribute dont_touch of G13489: signal is true;
	signal G13490: std_logic; attribute dont_touch of G13490: signal is true;
	signal G13491: std_logic; attribute dont_touch of G13491: signal is true;
	signal G13492: std_logic; attribute dont_touch of G13492: signal is true;
	signal G13493: std_logic; attribute dont_touch of G13493: signal is true;
	signal G13494: std_logic; attribute dont_touch of G13494: signal is true;
	signal G13495: std_logic; attribute dont_touch of G13495: signal is true;
	signal G13496: std_logic; attribute dont_touch of G13496: signal is true;
	signal G13497: std_logic; attribute dont_touch of G13497: signal is true;
	signal G13498: std_logic; attribute dont_touch of G13498: signal is true;
	signal G13499: std_logic; attribute dont_touch of G13499: signal is true;
	signal G13500: std_logic; attribute dont_touch of G13500: signal is true;
	signal G13501: std_logic; attribute dont_touch of G13501: signal is true;
	signal G13502: std_logic; attribute dont_touch of G13502: signal is true;
	signal G13503: std_logic; attribute dont_touch of G13503: signal is true;
	signal G13504: std_logic; attribute dont_touch of G13504: signal is true;
	signal G13505: std_logic; attribute dont_touch of G13505: signal is true;
	signal G13506: std_logic; attribute dont_touch of G13506: signal is true;
	signal G13507: std_logic; attribute dont_touch of G13507: signal is true;
	signal G13510: std_logic; attribute dont_touch of G13510: signal is true;
	signal G13511: std_logic; attribute dont_touch of G13511: signal is true;
	signal G13512: std_logic; attribute dont_touch of G13512: signal is true;
	signal G13513: std_logic; attribute dont_touch of G13513: signal is true;
	signal G13514: std_logic; attribute dont_touch of G13514: signal is true;
	signal G13515: std_logic; attribute dont_touch of G13515: signal is true;
	signal G13516: std_logic; attribute dont_touch of G13516: signal is true;
	signal G13517: std_logic; attribute dont_touch of G13517: signal is true;
	signal G13518: std_logic; attribute dont_touch of G13518: signal is true;
	signal G13519: std_logic; attribute dont_touch of G13519: signal is true;
	signal G13524: std_logic; attribute dont_touch of G13524: signal is true;
	signal G13525: std_logic; attribute dont_touch of G13525: signal is true;
	signal G13526: std_logic; attribute dont_touch of G13526: signal is true;
	signal G13527: std_logic; attribute dont_touch of G13527: signal is true;
	signal G13528: std_logic; attribute dont_touch of G13528: signal is true;
	signal G13529: std_logic; attribute dont_touch of G13529: signal is true;
	signal G13530: std_logic; attribute dont_touch of G13530: signal is true;
	signal G13535: std_logic; attribute dont_touch of G13535: signal is true;
	signal G13536: std_logic; attribute dont_touch of G13536: signal is true;
	signal G13537: std_logic; attribute dont_touch of G13537: signal is true;
	signal G13538: std_logic; attribute dont_touch of G13538: signal is true;
	signal G13539: std_logic; attribute dont_touch of G13539: signal is true;
	signal G13540: std_logic; attribute dont_touch of G13540: signal is true;
	signal G13541: std_logic; attribute dont_touch of G13541: signal is true;
	signal G13546: std_logic; attribute dont_touch of G13546: signal is true;
	signal G13547: std_logic; attribute dont_touch of G13547: signal is true;
	signal G13548: std_logic; attribute dont_touch of G13548: signal is true;
	signal G13549: std_logic; attribute dont_touch of G13549: signal is true;
	signal G13550: std_logic; attribute dont_touch of G13550: signal is true;
	signal G13551: std_logic; attribute dont_touch of G13551: signal is true;
	signal G13552: std_logic; attribute dont_touch of G13552: signal is true;
	signal G13557: std_logic; attribute dont_touch of G13557: signal is true;
	signal G13558: std_logic; attribute dont_touch of G13558: signal is true;
	signal G13559: std_logic; attribute dont_touch of G13559: signal is true;
	signal G13560: std_logic; attribute dont_touch of G13560: signal is true;
	signal G13561: std_logic; attribute dont_touch of G13561: signal is true;
	signal G13562: std_logic; attribute dont_touch of G13562: signal is true;
	signal G13563: std_logic; attribute dont_touch of G13563: signal is true;
	signal G13564: std_logic; attribute dont_touch of G13564: signal is true;
	signal G13565: std_logic; attribute dont_touch of G13565: signal is true;
	signal G13568: std_logic; attribute dont_touch of G13568: signal is true;
	signal G13571: std_logic; attribute dont_touch of G13571: signal is true;
	signal G13572: std_logic; attribute dont_touch of G13572: signal is true;
	signal G13573: std_logic; attribute dont_touch of G13573: signal is true;
	signal G13576: std_logic; attribute dont_touch of G13576: signal is true;
	signal G13579: std_logic; attribute dont_touch of G13579: signal is true;
	signal G13580: std_logic; attribute dont_touch of G13580: signal is true;
	signal G13581: std_logic; attribute dont_touch of G13581: signal is true;
	signal G13582: std_logic; attribute dont_touch of G13582: signal is true;
	signal G13585: std_logic; attribute dont_touch of G13585: signal is true;
	signal G13588: std_logic; attribute dont_touch of G13588: signal is true;
	signal G13589: std_logic; attribute dont_touch of G13589: signal is true;
	signal G13598: std_logic; attribute dont_touch of G13598: signal is true;
	signal G13599: std_logic; attribute dont_touch of G13599: signal is true;
	signal G13600: std_logic; attribute dont_touch of G13600: signal is true;
	signal G13601: std_logic; attribute dont_touch of G13601: signal is true;
	signal G13602: std_logic; attribute dont_touch of G13602: signal is true;
	signal G13605: std_logic; attribute dont_touch of G13605: signal is true;
	signal G13608: std_logic; attribute dont_touch of G13608: signal is true;
	signal G13609: std_logic; attribute dont_touch of G13609: signal is true;
	signal G13610: std_logic; attribute dont_touch of G13610: signal is true;
	signal G13611: std_logic; attribute dont_touch of G13611: signal is true;
	signal G13612: std_logic; attribute dont_touch of G13612: signal is true;
	signal G13613: std_logic; attribute dont_touch of G13613: signal is true;
	signal G13614: std_logic; attribute dont_touch of G13614: signal is true;
	signal G13619: std_logic; attribute dont_touch of G13619: signal is true;
	signal G13620: std_logic; attribute dont_touch of G13620: signal is true;
	signal G13621: std_logic; attribute dont_touch of G13621: signal is true;
	signal G13622: std_logic; attribute dont_touch of G13622: signal is true;
	signal G13623: std_logic; attribute dont_touch of G13623: signal is true;
	signal G13624: std_logic; attribute dont_touch of G13624: signal is true;
	signal G13625: std_logic; attribute dont_touch of G13625: signal is true;
	signal G13626: std_logic; attribute dont_touch of G13626: signal is true;
	signal G13631: std_logic; attribute dont_touch of G13631: signal is true;
	signal G13632: std_logic; attribute dont_touch of G13632: signal is true;
	signal G13633: std_logic; attribute dont_touch of G13633: signal is true;
	signal G13634: std_logic; attribute dont_touch of G13634: signal is true;
	signal G13635: std_logic; attribute dont_touch of G13635: signal is true;
	signal G13636: std_logic; attribute dont_touch of G13636: signal is true;
	signal G13637: std_logic; attribute dont_touch of G13637: signal is true;
	signal G13642: std_logic; attribute dont_touch of G13642: signal is true;
	signal G13643: std_logic; attribute dont_touch of G13643: signal is true;
	signal G13644: std_logic; attribute dont_touch of G13644: signal is true;
	signal G13645: std_logic; attribute dont_touch of G13645: signal is true;
	signal G13646: std_logic; attribute dont_touch of G13646: signal is true;
	signal G13647: std_logic; attribute dont_touch of G13647: signal is true;
	signal G13648: std_logic; attribute dont_touch of G13648: signal is true;
	signal G13649: std_logic; attribute dont_touch of G13649: signal is true;
	signal G13654: std_logic; attribute dont_touch of G13654: signal is true;
	signal G13655: std_logic; attribute dont_touch of G13655: signal is true;
	signal G13656: std_logic; attribute dont_touch of G13656: signal is true;
	signal G13657: std_logic; attribute dont_touch of G13657: signal is true;
	signal G13669: std_logic; attribute dont_touch of G13669: signal is true;
	signal G13670: std_logic; attribute dont_touch of G13670: signal is true;
	signal G13671: std_logic; attribute dont_touch of G13671: signal is true;
	signal G13672: std_logic; attribute dont_touch of G13672: signal is true;
	signal G13673: std_logic; attribute dont_touch of G13673: signal is true;
	signal G13674: std_logic; attribute dont_touch of G13674: signal is true;
	signal G13675: std_logic; attribute dont_touch of G13675: signal is true;
	signal G13676: std_logic; attribute dont_touch of G13676: signal is true;
	signal G13677: std_logic; attribute dont_touch of G13677: signal is true;
	signal G13687: std_logic; attribute dont_touch of G13687: signal is true;
	signal G13699: std_logic; attribute dont_touch of G13699: signal is true;
	signal G13700: std_logic; attribute dont_touch of G13700: signal is true;
	signal G13701: std_logic; attribute dont_touch of G13701: signal is true;
	signal G13702: std_logic; attribute dont_touch of G13702: signal is true;
	signal G13703: std_logic; attribute dont_touch of G13703: signal is true;
	signal G13704: std_logic; attribute dont_touch of G13704: signal is true;
	signal G13705: std_logic; attribute dont_touch of G13705: signal is true;
	signal G13706: std_logic; attribute dont_touch of G13706: signal is true;
	signal G13714: std_logic; attribute dont_touch of G13714: signal is true;
	signal G13724: std_logic; attribute dont_touch of G13724: signal is true;
	signal G13736: std_logic; attribute dont_touch of G13736: signal is true;
	signal G13737: std_logic; attribute dont_touch of G13737: signal is true;
	signal G13738: std_logic; attribute dont_touch of G13738: signal is true;
	signal G13739: std_logic; attribute dont_touch of G13739: signal is true;
	signal G13740: std_logic; attribute dont_touch of G13740: signal is true;
	signal G13741: std_logic; attribute dont_touch of G13741: signal is true;
	signal G13750: std_logic; attribute dont_touch of G13750: signal is true;
	signal G13755: std_logic; attribute dont_touch of G13755: signal is true;
	signal G13756: std_logic; attribute dont_touch of G13756: signal is true;
	signal G13764: std_logic; attribute dont_touch of G13764: signal is true;
	signal G13774: std_logic; attribute dont_touch of G13774: signal is true;
	signal G13786: std_logic; attribute dont_touch of G13786: signal is true;
	signal G13787: std_logic; attribute dont_touch of G13787: signal is true;
	signal G13788: std_logic; attribute dont_touch of G13788: signal is true;
	signal G13789: std_logic; attribute dont_touch of G13789: signal is true;
	signal G13790: std_logic; attribute dont_touch of G13790: signal is true;
	signal G13791: std_logic; attribute dont_touch of G13791: signal is true;
	signal G13796: std_logic; attribute dont_touch of G13796: signal is true;
	signal G13797: std_logic; attribute dont_touch of G13797: signal is true;
	signal G13805: std_logic; attribute dont_touch of G13805: signal is true;
	signal G13815: std_logic; attribute dont_touch of G13815: signal is true;
	signal G13816: std_logic; attribute dont_touch of G13816: signal is true;
	signal G13817: std_logic; attribute dont_touch of G13817: signal is true;
	signal G13818: std_logic; attribute dont_touch of G13818: signal is true;
	signal G13819: std_logic; attribute dont_touch of G13819: signal is true;
	signal G13824: std_logic; attribute dont_touch of G13824: signal is true;
	signal G13825: std_logic; attribute dont_touch of G13825: signal is true;
	signal G13833: std_logic; attribute dont_touch of G13833: signal is true;
	signal G13834: std_logic; attribute dont_touch of G13834: signal is true;
	signal G13835: std_logic; attribute dont_touch of G13835: signal is true;
	signal G13836: std_logic; attribute dont_touch of G13836: signal is true;
	signal G13837: std_logic; attribute dont_touch of G13837: signal is true;
	signal G13838: std_logic; attribute dont_touch of G13838: signal is true;
	signal G13839: std_logic; attribute dont_touch of G13839: signal is true;
	signal G13840: std_logic; attribute dont_touch of G13840: signal is true;
	signal G13845: std_logic; attribute dont_touch of G13845: signal is true;
	signal G13846: std_logic; attribute dont_touch of G13846: signal is true;
	signal G13847: std_logic; attribute dont_touch of G13847: signal is true;
	signal G13848: std_logic; attribute dont_touch of G13848: signal is true;
	signal G13849: std_logic; attribute dont_touch of G13849: signal is true;
	signal G13850: std_logic; attribute dont_touch of G13850: signal is true;
	signal G13851: std_logic; attribute dont_touch of G13851: signal is true;
	signal G13852: std_logic; attribute dont_touch of G13852: signal is true;
	signal G13853: std_logic; attribute dont_touch of G13853: signal is true;
	signal G13854: std_logic; attribute dont_touch of G13854: signal is true;
	signal G13855: std_logic; attribute dont_touch of G13855: signal is true;
	signal G13856: std_logic; attribute dont_touch of G13856: signal is true;
	signal G13857: std_logic; attribute dont_touch of G13857: signal is true;
	signal G13858: std_logic; attribute dont_touch of G13858: signal is true;
	signal G13859: std_logic; attribute dont_touch of G13859: signal is true;
	signal G13860: std_logic; attribute dont_touch of G13860: signal is true;
	signal G13861: std_logic; attribute dont_touch of G13861: signal is true;
	signal G13862: std_logic; attribute dont_touch of G13862: signal is true;
	signal G13863: std_logic; attribute dont_touch of G13863: signal is true;
	signal G13864: std_logic; attribute dont_touch of G13864: signal is true;
	signal G13865: std_logic; attribute dont_touch of G13865: signal is true;
	signal G13866: std_logic; attribute dont_touch of G13866: signal is true;
	signal G13867: std_logic; attribute dont_touch of G13867: signal is true;
	signal G13868: std_logic; attribute dont_touch of G13868: signal is true;
	signal G13869: std_logic; attribute dont_touch of G13869: signal is true;
	signal G13870: std_logic; attribute dont_touch of G13870: signal is true;
	signal G13871: std_logic; attribute dont_touch of G13871: signal is true;
	signal G13872: std_logic; attribute dont_touch of G13872: signal is true;
	signal G13873: std_logic; attribute dont_touch of G13873: signal is true;
	signal G13878: std_logic; attribute dont_touch of G13878: signal is true;
	signal G13879: std_logic; attribute dont_touch of G13879: signal is true;
	signal G13880: std_logic; attribute dont_touch of G13880: signal is true;
	signal G13881: std_logic; attribute dont_touch of G13881: signal is true;
	signal G13882: std_logic; attribute dont_touch of G13882: signal is true;
	signal G13883: std_logic; attribute dont_touch of G13883: signal is true;
	signal G13884: std_logic; attribute dont_touch of G13884: signal is true;
	signal G13885: std_logic; attribute dont_touch of G13885: signal is true;
	signal G13886: std_logic; attribute dont_touch of G13886: signal is true;
	signal G13892: std_logic; attribute dont_touch of G13892: signal is true;
	signal G13893: std_logic; attribute dont_touch of G13893: signal is true;
	signal G13894: std_logic; attribute dont_touch of G13894: signal is true;
	signal G13895: std_logic; attribute dont_touch of G13895: signal is true;
	signal G13900: std_logic; attribute dont_touch of G13900: signal is true;
	signal G13901: std_logic; attribute dont_touch of G13901: signal is true;
	signal G13902: std_logic; attribute dont_touch of G13902: signal is true;
	signal G13903: std_logic; attribute dont_touch of G13903: signal is true;
	signal G13904: std_logic; attribute dont_touch of G13904: signal is true;
	signal G13905: std_logic; attribute dont_touch of G13905: signal is true;
	signal G13906: std_logic; attribute dont_touch of G13906: signal is true;
	signal G13907: std_logic; attribute dont_touch of G13907: signal is true;
	signal G13913: std_logic; attribute dont_touch of G13913: signal is true;
	signal G13914: std_logic; attribute dont_touch of G13914: signal is true;
	signal G13915: std_logic; attribute dont_touch of G13915: signal is true;
	signal G13918: std_logic; attribute dont_touch of G13918: signal is true;
	signal G13922: std_logic; attribute dont_touch of G13922: signal is true;
	signal G13926: std_logic; attribute dont_touch of G13926: signal is true;
	signal G13927: std_logic; attribute dont_touch of G13927: signal is true;
	signal G13933: std_logic; attribute dont_touch of G13933: signal is true;
	signal G13934: std_logic; attribute dont_touch of G13934: signal is true;
	signal G13935: std_logic; attribute dont_touch of G13935: signal is true;
	signal G13936: std_logic; attribute dont_touch of G13936: signal is true;
	signal G13941: std_logic; attribute dont_touch of G13941: signal is true;
	signal G13942: std_logic; attribute dont_touch of G13942: signal is true;
	signal G13943: std_logic; attribute dont_touch of G13943: signal is true;
	signal G13944: std_logic; attribute dont_touch of G13944: signal is true;
	signal G13945: std_logic; attribute dont_touch of G13945: signal is true;
	signal G13946: std_logic; attribute dont_touch of G13946: signal is true;
	signal G13952: std_logic; attribute dont_touch of G13952: signal is true;
	signal G13953: std_logic; attribute dont_touch of G13953: signal is true;
	signal G13954: std_logic; attribute dont_touch of G13954: signal is true;
	signal G13957: std_logic; attribute dont_touch of G13957: signal is true;
	signal G13958: std_logic; attribute dont_touch of G13958: signal is true;
	signal G13962: std_logic; attribute dont_touch of G13962: signal is true;
	signal G13963: std_logic; attribute dont_touch of G13963: signal is true;
	signal G13969: std_logic; attribute dont_touch of G13969: signal is true;
	signal G13970: std_logic; attribute dont_touch of G13970: signal is true;
	signal G13971: std_logic; attribute dont_touch of G13971: signal is true;
	signal G13974: std_logic; attribute dont_touch of G13974: signal is true;
	signal G13978: std_logic; attribute dont_touch of G13978: signal is true;
	signal G13982: std_logic; attribute dont_touch of G13982: signal is true;
	signal G13983: std_logic; attribute dont_touch of G13983: signal is true;
	signal G13989: std_logic; attribute dont_touch of G13989: signal is true;
	signal G13990: std_logic; attribute dont_touch of G13990: signal is true;
	signal G13991: std_logic; attribute dont_touch of G13991: signal is true;
	signal G13992: std_logic; attribute dont_touch of G13992: signal is true;
	signal G13997: std_logic; attribute dont_touch of G13997: signal is true;
	signal G13998: std_logic; attribute dont_touch of G13998: signal is true;
	signal G13999: std_logic; attribute dont_touch of G13999: signal is true;
	signal G14000: std_logic; attribute dont_touch of G14000: signal is true;
	signal G14001: std_logic; attribute dont_touch of G14001: signal is true;
	signal G14006: std_logic; attribute dont_touch of G14006: signal is true;
	signal G14007: std_logic; attribute dont_touch of G14007: signal is true;
	signal G14008: std_logic; attribute dont_touch of G14008: signal is true;
	signal G14011: std_logic; attribute dont_touch of G14011: signal is true;
	signal G14015: std_logic; attribute dont_touch of G14015: signal is true;
	signal G14016: std_logic; attribute dont_touch of G14016: signal is true;
	signal G14022: std_logic; attribute dont_touch of G14022: signal is true;
	signal G14023: std_logic; attribute dont_touch of G14023: signal is true;
	signal G14024: std_logic; attribute dont_touch of G14024: signal is true;
	signal G14027: std_logic; attribute dont_touch of G14027: signal is true;
	signal G14028: std_logic; attribute dont_touch of G14028: signal is true;
	signal G14032: std_logic; attribute dont_touch of G14032: signal is true;
	signal G14033: std_logic; attribute dont_touch of G14033: signal is true;
	signal G14039: std_logic; attribute dont_touch of G14039: signal is true;
	signal G14040: std_logic; attribute dont_touch of G14040: signal is true;
	signal G14041: std_logic; attribute dont_touch of G14041: signal is true;
	signal G14044: std_logic; attribute dont_touch of G14044: signal is true;
	signal G14048: std_logic; attribute dont_touch of G14048: signal is true;
	signal G14052: std_logic; attribute dont_touch of G14052: signal is true;
	signal G14053: std_logic; attribute dont_touch of G14053: signal is true;
	signal G14059: std_logic; attribute dont_touch of G14059: signal is true;
	signal G14060: std_logic; attribute dont_touch of G14060: signal is true;
	signal G14061: std_logic; attribute dont_touch of G14061: signal is true;
	signal G14062: std_logic; attribute dont_touch of G14062: signal is true;
	signal G14067: std_logic; attribute dont_touch of G14067: signal is true;
	signal G14068: std_logic; attribute dont_touch of G14068: signal is true;
	signal G14071: std_logic; attribute dont_touch of G14071: signal is true;
	signal G14079: std_logic; attribute dont_touch of G14079: signal is true;
	signal G14086: std_logic; attribute dont_touch of G14086: signal is true;
	signal G14090: std_logic; attribute dont_touch of G14090: signal is true;
	signal G14091: std_logic; attribute dont_touch of G14091: signal is true;
	signal G14092: std_logic; attribute dont_touch of G14092: signal is true;
	signal G14097: std_logic; attribute dont_touch of G14097: signal is true;
	signal G14098: std_logic; attribute dont_touch of G14098: signal is true;
	signal G14099: std_logic; attribute dont_touch of G14099: signal is true;
	signal G14102: std_logic; attribute dont_touch of G14102: signal is true;
	signal G14106: std_logic; attribute dont_touch of G14106: signal is true;
	signal G14107: std_logic; attribute dont_touch of G14107: signal is true;
	signal G14113: std_logic; attribute dont_touch of G14113: signal is true;
	signal G14114: std_logic; attribute dont_touch of G14114: signal is true;
	signal G14115: std_logic; attribute dont_touch of G14115: signal is true;
	signal G14118: std_logic; attribute dont_touch of G14118: signal is true;
	signal G14119: std_logic; attribute dont_touch of G14119: signal is true;
	signal G14123: std_logic; attribute dont_touch of G14123: signal is true;
	signal G14124: std_logic; attribute dont_touch of G14124: signal is true;
	signal G14130: std_logic; attribute dont_touch of G14130: signal is true;
	signal G14131: std_logic; attribute dont_touch of G14131: signal is true;
	signal G14132: std_logic; attribute dont_touch of G14132: signal is true;
	signal G14135: std_logic; attribute dont_touch of G14135: signal is true;
	signal G14139: std_logic; attribute dont_touch of G14139: signal is true;
	signal G14143: std_logic; attribute dont_touch of G14143: signal is true;
	signal G14144: std_logic; attribute dont_touch of G14144: signal is true;
	signal G14148: std_logic; attribute dont_touch of G14148: signal is true;
	signal G14153: std_logic; attribute dont_touch of G14153: signal is true;
	signal G14158: std_logic; attribute dont_touch of G14158: signal is true;
	signal G14165: std_logic; attribute dont_touch of G14165: signal is true;
	signal G14171: std_logic; attribute dont_touch of G14171: signal is true;
	signal G14175: std_logic; attribute dont_touch of G14175: signal is true;
	signal G14176: std_logic; attribute dont_touch of G14176: signal is true;
	signal G14177: std_logic; attribute dont_touch of G14177: signal is true;
	signal G14182: std_logic; attribute dont_touch of G14182: signal is true;
	signal G14183: std_logic; attribute dont_touch of G14183: signal is true;
	signal G14186: std_logic; attribute dont_touch of G14186: signal is true;
	signal G14194: std_logic; attribute dont_touch of G14194: signal is true;
	signal G14201: std_logic; attribute dont_touch of G14201: signal is true;
	signal G14205: std_logic; attribute dont_touch of G14205: signal is true;
	signal G14206: std_logic; attribute dont_touch of G14206: signal is true;
	signal G14207: std_logic; attribute dont_touch of G14207: signal is true;
	signal G14212: std_logic; attribute dont_touch of G14212: signal is true;
	signal G14213: std_logic; attribute dont_touch of G14213: signal is true;
	signal G14214: std_logic; attribute dont_touch of G14214: signal is true;
	signal G14217: std_logic; attribute dont_touch of G14217: signal is true;
	signal G14221: std_logic; attribute dont_touch of G14221: signal is true;
	signal G14222: std_logic; attribute dont_touch of G14222: signal is true;
	signal G14228: std_logic; attribute dont_touch of G14228: signal is true;
	signal G14229: std_logic; attribute dont_touch of G14229: signal is true;
	signal G14230: std_logic; attribute dont_touch of G14230: signal is true;
	signal G14233: std_logic; attribute dont_touch of G14233: signal is true;
	signal G14234: std_logic; attribute dont_touch of G14234: signal is true;
	signal G14238: std_logic; attribute dont_touch of G14238: signal is true;
	signal G14244: std_logic; attribute dont_touch of G14244: signal is true;
	signal G14249: std_logic; attribute dont_touch of G14249: signal is true;
	signal G14252: std_logic; attribute dont_touch of G14252: signal is true;
	signal G14256: std_logic; attribute dont_touch of G14256: signal is true;
	signal G14259: std_logic; attribute dont_touch of G14259: signal is true;
	signal G14263: std_logic; attribute dont_touch of G14263: signal is true;
	signal G14268: std_logic; attribute dont_touch of G14268: signal is true;
	signal G14273: std_logic; attribute dont_touch of G14273: signal is true;
	signal G14280: std_logic; attribute dont_touch of G14280: signal is true;
	signal G14286: std_logic; attribute dont_touch of G14286: signal is true;
	signal G14290: std_logic; attribute dont_touch of G14290: signal is true;
	signal G14291: std_logic; attribute dont_touch of G14291: signal is true;
	signal G14292: std_logic; attribute dont_touch of G14292: signal is true;
	signal G14297: std_logic; attribute dont_touch of G14297: signal is true;
	signal G14298: std_logic; attribute dont_touch of G14298: signal is true;
	signal G14301: std_logic; attribute dont_touch of G14301: signal is true;
	signal G14309: std_logic; attribute dont_touch of G14309: signal is true;
	signal G14316: std_logic; attribute dont_touch of G14316: signal is true;
	signal G14320: std_logic; attribute dont_touch of G14320: signal is true;
	signal G14321: std_logic; attribute dont_touch of G14321: signal is true;
	signal G14322: std_logic; attribute dont_touch of G14322: signal is true;
	signal G14327: std_logic; attribute dont_touch of G14327: signal is true;
	signal G14328: std_logic; attribute dont_touch of G14328: signal is true;
	signal G14329: std_logic; attribute dont_touch of G14329: signal is true;
	signal G14332: std_logic; attribute dont_touch of G14332: signal is true;
	signal G14336: std_logic; attribute dont_touch of G14336: signal is true;
	signal G14337: std_logic; attribute dont_touch of G14337: signal is true;
	signal G14342: std_logic; attribute dont_touch of G14342: signal is true;
	signal G14347: std_logic; attribute dont_touch of G14347: signal is true;
	signal G14352: std_logic; attribute dont_touch of G14352: signal is true;
	signal G14355: std_logic; attribute dont_touch of G14355: signal is true;
	signal G14359: std_logic; attribute dont_touch of G14359: signal is true;
	signal G14360: std_logic; attribute dont_touch of G14360: signal is true;
	signal G14366: std_logic; attribute dont_touch of G14366: signal is true;
	signal G14371: std_logic; attribute dont_touch of G14371: signal is true;
	signal G14374: std_logic; attribute dont_touch of G14374: signal is true;
	signal G14378: std_logic; attribute dont_touch of G14378: signal is true;
	signal G14381: std_logic; attribute dont_touch of G14381: signal is true;
	signal G14385: std_logic; attribute dont_touch of G14385: signal is true;
	signal G14390: std_logic; attribute dont_touch of G14390: signal is true;
	signal G14395: std_logic; attribute dont_touch of G14395: signal is true;
	signal G14402: std_logic; attribute dont_touch of G14402: signal is true;
	signal G14408: std_logic; attribute dont_touch of G14408: signal is true;
	signal G14412: std_logic; attribute dont_touch of G14412: signal is true;
	signal G14413: std_logic; attribute dont_touch of G14413: signal is true;
	signal G14414: std_logic; attribute dont_touch of G14414: signal is true;
	signal G14419: std_logic; attribute dont_touch of G14419: signal is true;
	signal G14420: std_logic; attribute dont_touch of G14420: signal is true;
	signal G14423: std_logic; attribute dont_touch of G14423: signal is true;
	signal G14431: std_logic; attribute dont_touch of G14431: signal is true;
	signal G14438: std_logic; attribute dont_touch of G14438: signal is true;
	signal G14442: std_logic; attribute dont_touch of G14442: signal is true;
	signal G14450: std_logic; attribute dont_touch of G14450: signal is true;
	signal G14454: std_logic; attribute dont_touch of G14454: signal is true;
	signal G14459: std_logic; attribute dont_touch of G14459: signal is true;
	signal G14464: std_logic; attribute dont_touch of G14464: signal is true;
	signal G14467: std_logic; attribute dont_touch of G14467: signal is true;
	signal G14471: std_logic; attribute dont_touch of G14471: signal is true;
	signal G14472: std_logic; attribute dont_touch of G14472: signal is true;
	signal G14478: std_logic; attribute dont_touch of G14478: signal is true;
	signal G14483: std_logic; attribute dont_touch of G14483: signal is true;
	signal G14486: std_logic; attribute dont_touch of G14486: signal is true;
	signal G14490: std_logic; attribute dont_touch of G14490: signal is true;
	signal G14493: std_logic; attribute dont_touch of G14493: signal is true;
	signal G14497: std_logic; attribute dont_touch of G14497: signal is true;
	signal G14502: std_logic; attribute dont_touch of G14502: signal is true;
	signal G14507: std_logic; attribute dont_touch of G14507: signal is true;
	signal G14514: std_logic; attribute dont_touch of G14514: signal is true;
	signal G14520: std_logic; attribute dont_touch of G14520: signal is true;
	signal G14524: std_logic; attribute dont_touch of G14524: signal is true;
	signal G14525: std_logic; attribute dont_touch of G14525: signal is true;
	signal G14529: std_logic; attribute dont_touch of G14529: signal is true;
	signal G14537: std_logic; attribute dont_touch of G14537: signal is true;
	signal G14541: std_logic; attribute dont_touch of G14541: signal is true;
	signal G14546: std_logic; attribute dont_touch of G14546: signal is true;
	signal G14551: std_logic; attribute dont_touch of G14551: signal is true;
	signal G14554: std_logic; attribute dont_touch of G14554: signal is true;
	signal G14558: std_logic; attribute dont_touch of G14558: signal is true;
	signal G14559: std_logic; attribute dont_touch of G14559: signal is true;
	signal G14565: std_logic; attribute dont_touch of G14565: signal is true;
	signal G14570: std_logic; attribute dont_touch of G14570: signal is true;
	signal G14573: std_logic; attribute dont_touch of G14573: signal is true;
	signal G14577: std_logic; attribute dont_touch of G14577: signal is true;
	signal G14580: std_logic; attribute dont_touch of G14580: signal is true;
	signal G14584: std_logic; attribute dont_touch of G14584: signal is true;
	signal G14592: std_logic; attribute dont_touch of G14592: signal is true;
	signal G14596: std_logic; attribute dont_touch of G14596: signal is true;
	signal G14601: std_logic; attribute dont_touch of G14601: signal is true;
	signal G14606: std_logic; attribute dont_touch of G14606: signal is true;
	signal G14609: std_logic; attribute dont_touch of G14609: signal is true;
	signal G14613: std_logic; attribute dont_touch of G14613: signal is true;
	signal G14614: std_logic; attribute dont_touch of G14614: signal is true;
	signal G14618: std_logic; attribute dont_touch of G14618: signal is true;
	signal G14626: std_logic; attribute dont_touch of G14626: signal is true;
	signal G14630: std_logic; attribute dont_touch of G14630: signal is true;
	signal G14637: std_logic; attribute dont_touch of G14637: signal is true;
	signal G14641: std_logic; attribute dont_touch of G14641: signal is true;
	signal G14642: std_logic; attribute dont_touch of G14642: signal is true;
	signal G14650: std_logic; attribute dont_touch of G14650: signal is true;
	signal G14657: std_logic; attribute dont_touch of G14657: signal is true;
	signal G14668: std_logic; attribute dont_touch of G14668: signal is true;
	signal G14669: std_logic; attribute dont_touch of G14669: signal is true;
	signal G14677: std_logic; attribute dont_touch of G14677: signal is true;
	signal G14684: std_logic; attribute dont_touch of G14684: signal is true;
	signal G14685: std_logic; attribute dont_touch of G14685: signal is true;
	signal G14690: std_logic; attribute dont_touch of G14690: signal is true;
	signal G14691: std_logic; attribute dont_touch of G14691: signal is true;
	signal G14702: std_logic; attribute dont_touch of G14702: signal is true;
	signal G14703: std_logic; attribute dont_touch of G14703: signal is true;
	signal G14711: std_logic; attribute dont_touch of G14711: signal is true;
	signal G14718: std_logic; attribute dont_touch of G14718: signal is true;
	signal G14719: std_logic; attribute dont_touch of G14719: signal is true;
	signal G14724: std_logic; attribute dont_touch of G14724: signal is true;
	signal G14725: std_logic; attribute dont_touch of G14725: signal is true;
	signal G14736: std_logic; attribute dont_touch of G14736: signal is true;
	signal G14737: std_logic; attribute dont_touch of G14737: signal is true;
	signal G14745: std_logic; attribute dont_touch of G14745: signal is true;
	signal G14746: std_logic; attribute dont_touch of G14746: signal is true;
	signal G14747: std_logic; attribute dont_touch of G14747: signal is true;
	signal G14752: std_logic; attribute dont_touch of G14752: signal is true;
	signal G14753: std_logic; attribute dont_touch of G14753: signal is true;
	signal G14764: std_logic; attribute dont_touch of G14764: signal is true;
	signal G14765: std_logic; attribute dont_touch of G14765: signal is true;
	signal G14766: std_logic; attribute dont_touch of G14766: signal is true;
	signal G14767: std_logic; attribute dont_touch of G14767: signal is true;
	signal G14768: std_logic; attribute dont_touch of G14768: signal is true;
	signal G14773: std_logic; attribute dont_touch of G14773: signal is true;
	signal G14774: std_logic; attribute dont_touch of G14774: signal is true;
	signal G14775: std_logic; attribute dont_touch of G14775: signal is true;
	signal G14776: std_logic; attribute dont_touch of G14776: signal is true;
	signal G14794: std_logic; attribute dont_touch of G14794: signal is true;
	signal G14795: std_logic; attribute dont_touch of G14795: signal is true;
	signal G14796: std_logic; attribute dont_touch of G14796: signal is true;
	signal G14797: std_logic; attribute dont_touch of G14797: signal is true;
	signal G14811: std_logic; attribute dont_touch of G14811: signal is true;
	signal G14829: std_logic; attribute dont_touch of G14829: signal is true;
	signal G14830: std_logic; attribute dont_touch of G14830: signal is true;
	signal G14831: std_logic; attribute dont_touch of G14831: signal is true;
	signal G14837: std_logic; attribute dont_touch of G14837: signal is true;
	signal G14849: std_logic; attribute dont_touch of G14849: signal is true;
	signal G14863: std_logic; attribute dont_touch of G14863: signal is true;
	signal G14881: std_logic; attribute dont_touch of G14881: signal is true;
	signal G14882: std_logic; attribute dont_touch of G14882: signal is true;
	signal G14883: std_logic; attribute dont_touch of G14883: signal is true;
	signal G14884: std_logic; attribute dont_touch of G14884: signal is true;
	signal G14885: std_logic; attribute dont_touch of G14885: signal is true;
	signal G14894: std_logic; attribute dont_touch of G14894: signal is true;
	signal G14895: std_logic; attribute dont_touch of G14895: signal is true;
	signal G14904: std_logic; attribute dont_touch of G14904: signal is true;
	signal G14910: std_logic; attribute dont_touch of G14910: signal is true;
	signal G14922: std_logic; attribute dont_touch of G14922: signal is true;
	signal G14936: std_logic; attribute dont_touch of G14936: signal is true;
	signal G14954: std_logic; attribute dont_touch of G14954: signal is true;
	signal G14955: std_logic; attribute dont_touch of G14955: signal is true;
	signal G14956: std_logic; attribute dont_touch of G14956: signal is true;
	signal G14957: std_logic; attribute dont_touch of G14957: signal is true;
	signal G14958: std_logic; attribute dont_touch of G14958: signal is true;
	signal G14959: std_logic; attribute dont_touch of G14959: signal is true;
	signal G14960: std_logic; attribute dont_touch of G14960: signal is true;
	signal G14963: std_logic; attribute dont_touch of G14963: signal is true;
	signal G14966: std_logic; attribute dont_touch of G14966: signal is true;
	signal G14975: std_logic; attribute dont_touch of G14975: signal is true;
	signal G14976: std_logic; attribute dont_touch of G14976: signal is true;
	signal G14985: std_logic; attribute dont_touch of G14985: signal is true;
	signal G14991: std_logic; attribute dont_touch of G14991: signal is true;
	signal G15003: std_logic; attribute dont_touch of G15003: signal is true;
	signal G15017: std_logic; attribute dont_touch of G15017: signal is true;
	signal G15018: std_logic; attribute dont_touch of G15018: signal is true;
	signal G15019: std_logic; attribute dont_touch of G15019: signal is true;
	signal G15020: std_logic; attribute dont_touch of G15020: signal is true;
	signal G15021: std_logic; attribute dont_touch of G15021: signal is true;
	signal G15022: std_logic; attribute dont_touch of G15022: signal is true;
	signal G15030: std_logic; attribute dont_touch of G15030: signal is true;
	signal G15031: std_logic; attribute dont_touch of G15031: signal is true;
	signal G15032: std_logic; attribute dont_touch of G15032: signal is true;
	signal G15033: std_logic; attribute dont_touch of G15033: signal is true;
	signal G15034: std_logic; attribute dont_touch of G15034: signal is true;
	signal G15037: std_logic; attribute dont_touch of G15037: signal is true;
	signal G15040: std_logic; attribute dont_touch of G15040: signal is true;
	signal G15043: std_logic; attribute dont_touch of G15043: signal is true;
	signal G15046: std_logic; attribute dont_touch of G15046: signal is true;
	signal G15047: std_logic; attribute dont_touch of G15047: signal is true;
	signal G15048: std_logic; attribute dont_touch of G15048: signal is true;
	signal G15049: std_logic; attribute dont_touch of G15049: signal is true;
	signal G15052: std_logic; attribute dont_touch of G15052: signal is true;
	signal G15055: std_logic; attribute dont_touch of G15055: signal is true;
	signal G15064: std_logic; attribute dont_touch of G15064: signal is true;
	signal G15065: std_logic; attribute dont_touch of G15065: signal is true;
	signal G15074: std_logic; attribute dont_touch of G15074: signal is true;
	signal G15080: std_logic; attribute dont_touch of G15080: signal is true;
	signal G15092: std_logic; attribute dont_touch of G15092: signal is true;
	signal G15093: std_logic; attribute dont_touch of G15093: signal is true;
	signal G15094: std_logic; attribute dont_touch of G15094: signal is true;
	signal G15095: std_logic; attribute dont_touch of G15095: signal is true;
	signal G15096: std_logic; attribute dont_touch of G15096: signal is true;
	signal G15104: std_logic; attribute dont_touch of G15104: signal is true;
	signal G15105: std_logic; attribute dont_touch of G15105: signal is true;
	signal G15106: std_logic; attribute dont_touch of G15106: signal is true;
	signal G15109: std_logic; attribute dont_touch of G15109: signal is true;
	signal G15112: std_logic; attribute dont_touch of G15112: signal is true;
	signal G15115: std_logic; attribute dont_touch of G15115: signal is true;
	signal G15118: std_logic; attribute dont_touch of G15118: signal is true;
	signal G15126: std_logic; attribute dont_touch of G15126: signal is true;
	signal G15127: std_logic; attribute dont_touch of G15127: signal is true;
	signal G15128: std_logic; attribute dont_touch of G15128: signal is true;
	signal G15129: std_logic; attribute dont_touch of G15129: signal is true;
	signal G15130: std_logic; attribute dont_touch of G15130: signal is true;
	signal G15133: std_logic; attribute dont_touch of G15133: signal is true;
	signal G15136: std_logic; attribute dont_touch of G15136: signal is true;
	signal G15139: std_logic; attribute dont_touch of G15139: signal is true;
	signal G15142: std_logic; attribute dont_touch of G15142: signal is true;
	signal G15143: std_logic; attribute dont_touch of G15143: signal is true;
	signal G15144: std_logic; attribute dont_touch of G15144: signal is true;
	signal G15145: std_logic; attribute dont_touch of G15145: signal is true;
	signal G15148: std_logic; attribute dont_touch of G15148: signal is true;
	signal G15151: std_logic; attribute dont_touch of G15151: signal is true;
	signal G15160: std_logic; attribute dont_touch of G15160: signal is true;
	signal G15161: std_logic; attribute dont_touch of G15161: signal is true;
	signal G15170: std_logic; attribute dont_touch of G15170: signal is true;
	signal G15171: std_logic; attribute dont_touch of G15171: signal is true;
	signal G15172: std_logic; attribute dont_touch of G15172: signal is true;
	signal G15173: std_logic; attribute dont_touch of G15173: signal is true;
	signal G15174: std_logic; attribute dont_touch of G15174: signal is true;
	signal G15175: std_logic; attribute dont_touch of G15175: signal is true;
	signal G15176: std_logic; attribute dont_touch of G15176: signal is true;
	signal G15177: std_logic; attribute dont_touch of G15177: signal is true;
	signal G15178: std_logic; attribute dont_touch of G15178: signal is true;
	signal G15179: std_logic; attribute dont_touch of G15179: signal is true;
	signal G15182: std_logic; attribute dont_touch of G15182: signal is true;
	signal G15185: std_logic; attribute dont_touch of G15185: signal is true;
	signal G15188: std_logic; attribute dont_touch of G15188: signal is true;
	signal G15196: std_logic; attribute dont_touch of G15196: signal is true;
	signal G15197: std_logic; attribute dont_touch of G15197: signal is true;
	signal G15198: std_logic; attribute dont_touch of G15198: signal is true;
	signal G15201: std_logic; attribute dont_touch of G15201: signal is true;
	signal G15204: std_logic; attribute dont_touch of G15204: signal is true;
	signal G15207: std_logic; attribute dont_touch of G15207: signal is true;
	signal G15210: std_logic; attribute dont_touch of G15210: signal is true;
	signal G15218: std_logic; attribute dont_touch of G15218: signal is true;
	signal G15219: std_logic; attribute dont_touch of G15219: signal is true;
	signal G15220: std_logic; attribute dont_touch of G15220: signal is true;
	signal G15221: std_logic; attribute dont_touch of G15221: signal is true;
	signal G15222: std_logic; attribute dont_touch of G15222: signal is true;
	signal G15225: std_logic; attribute dont_touch of G15225: signal is true;
	signal G15228: std_logic; attribute dont_touch of G15228: signal is true;
	signal G15231: std_logic; attribute dont_touch of G15231: signal is true;
	signal G15234: std_logic; attribute dont_touch of G15234: signal is true;
	signal G15235: std_logic; attribute dont_touch of G15235: signal is true;
	signal G15236: std_logic; attribute dont_touch of G15236: signal is true;
	signal G15237: std_logic; attribute dont_touch of G15237: signal is true;
	signal G15240: std_logic; attribute dont_touch of G15240: signal is true;
	signal G15243: std_logic; attribute dont_touch of G15243: signal is true;
	signal G15244: std_logic; attribute dont_touch of G15244: signal is true;
	signal G15245: std_logic; attribute dont_touch of G15245: signal is true;
	signal G15246: std_logic; attribute dont_touch of G15246: signal is true;
	signal G15247: std_logic; attribute dont_touch of G15247: signal is true;
	signal G15248: std_logic; attribute dont_touch of G15248: signal is true;
	signal G15251: std_logic; attribute dont_touch of G15251: signal is true;
	signal G15254: std_logic; attribute dont_touch of G15254: signal is true;
	signal G15257: std_logic; attribute dont_touch of G15257: signal is true;
	signal G15258: std_logic; attribute dont_touch of G15258: signal is true;
	signal G15259: std_logic; attribute dont_touch of G15259: signal is true;
	signal G15260: std_logic; attribute dont_touch of G15260: signal is true;
	signal G15261: std_logic; attribute dont_touch of G15261: signal is true;
	signal G15262: std_logic; attribute dont_touch of G15262: signal is true;
	signal G15263: std_logic; attribute dont_touch of G15263: signal is true;
	signal G15264: std_logic; attribute dont_touch of G15264: signal is true;
	signal G15265: std_logic; attribute dont_touch of G15265: signal is true;
	signal G15268: std_logic; attribute dont_touch of G15268: signal is true;
	signal G15271: std_logic; attribute dont_touch of G15271: signal is true;
	signal G15274: std_logic; attribute dont_touch of G15274: signal is true;
	signal G15282: std_logic; attribute dont_touch of G15282: signal is true;
	signal G15283: std_logic; attribute dont_touch of G15283: signal is true;
	signal G15284: std_logic; attribute dont_touch of G15284: signal is true;
	signal G15287: std_logic; attribute dont_touch of G15287: signal is true;
	signal G15290: std_logic; attribute dont_touch of G15290: signal is true;
	signal G15293: std_logic; attribute dont_touch of G15293: signal is true;
	signal G15296: std_logic; attribute dont_touch of G15296: signal is true;
	signal G15304: std_logic; attribute dont_touch of G15304: signal is true;
	signal G15305: std_logic; attribute dont_touch of G15305: signal is true;
	signal G15306: std_logic; attribute dont_touch of G15306: signal is true;
	signal G15307: std_logic; attribute dont_touch of G15307: signal is true;
	signal G15308: std_logic; attribute dont_touch of G15308: signal is true;
	signal G15311: std_logic; attribute dont_touch of G15311: signal is true;
	signal G15314: std_logic; attribute dont_touch of G15314: signal is true;
	signal G15317: std_logic; attribute dont_touch of G15317: signal is true;
	signal G15320: std_logic; attribute dont_touch of G15320: signal is true;
	signal G15321: std_logic; attribute dont_touch of G15321: signal is true;
	signal G15322: std_logic; attribute dont_touch of G15322: signal is true;
	signal G15323: std_logic; attribute dont_touch of G15323: signal is true;
	signal G15324: std_logic; attribute dont_touch of G15324: signal is true;
	signal G15325: std_logic; attribute dont_touch of G15325: signal is true;
	signal G15326: std_logic; attribute dont_touch of G15326: signal is true;
	signal G15329: std_logic; attribute dont_touch of G15329: signal is true;
	signal G15332: std_logic; attribute dont_touch of G15332: signal is true;
	signal G15335: std_logic; attribute dont_touch of G15335: signal is true;
	signal G15336: std_logic; attribute dont_touch of G15336: signal is true;
	signal G15337: std_logic; attribute dont_touch of G15337: signal is true;
	signal G15338: std_logic; attribute dont_touch of G15338: signal is true;
	signal G15339: std_logic; attribute dont_touch of G15339: signal is true;
	signal G15340: std_logic; attribute dont_touch of G15340: signal is true;
	signal G15343: std_logic; attribute dont_touch of G15343: signal is true;
	signal G15346: std_logic; attribute dont_touch of G15346: signal is true;
	signal G15349: std_logic; attribute dont_touch of G15349: signal is true;
	signal G15350: std_logic; attribute dont_touch of G15350: signal is true;
	signal G15351: std_logic; attribute dont_touch of G15351: signal is true;
	signal G15352: std_logic; attribute dont_touch of G15352: signal is true;
	signal G15353: std_logic; attribute dont_touch of G15353: signal is true;
	signal G15354: std_logic; attribute dont_touch of G15354: signal is true;
	signal G15355: std_logic; attribute dont_touch of G15355: signal is true;
	signal G15356: std_logic; attribute dont_touch of G15356: signal is true;
	signal G15357: std_logic; attribute dont_touch of G15357: signal is true;
	signal G15360: std_logic; attribute dont_touch of G15360: signal is true;
	signal G15363: std_logic; attribute dont_touch of G15363: signal is true;
	signal G15366: std_logic; attribute dont_touch of G15366: signal is true;
	signal G15374: std_logic; attribute dont_touch of G15374: signal is true;
	signal G15375: std_logic; attribute dont_touch of G15375: signal is true;
	signal G15376: std_logic; attribute dont_touch of G15376: signal is true;
	signal G15379: std_logic; attribute dont_touch of G15379: signal is true;
	signal G15382: std_logic; attribute dont_touch of G15382: signal is true;
	signal G15385: std_logic; attribute dont_touch of G15385: signal is true;
	signal G15388: std_logic; attribute dont_touch of G15388: signal is true;
	signal G15389: std_logic; attribute dont_touch of G15389: signal is true;
	signal G15390: std_logic; attribute dont_touch of G15390: signal is true;
	signal G15391: std_logic; attribute dont_touch of G15391: signal is true;
	signal G15392: std_logic; attribute dont_touch of G15392: signal is true;
	signal G15393: std_logic; attribute dont_touch of G15393: signal is true;
	signal G15396: std_logic; attribute dont_touch of G15396: signal is true;
	signal G15399: std_logic; attribute dont_touch of G15399: signal is true;
	signal G15402: std_logic; attribute dont_touch of G15402: signal is true;
	signal G15403: std_logic; attribute dont_touch of G15403: signal is true;
	signal G15404: std_logic; attribute dont_touch of G15404: signal is true;
	signal G15407: std_logic; attribute dont_touch of G15407: signal is true;
	signal G15408: std_logic; attribute dont_touch of G15408: signal is true;
	signal G15409: std_logic; attribute dont_touch of G15409: signal is true;
	signal G15410: std_logic; attribute dont_touch of G15410: signal is true;
	signal G15411: std_logic; attribute dont_touch of G15411: signal is true;
	signal G15412: std_logic; attribute dont_touch of G15412: signal is true;
	signal G15415: std_logic; attribute dont_touch of G15415: signal is true;
	signal G15418: std_logic; attribute dont_touch of G15418: signal is true;
	signal G15421: std_logic; attribute dont_touch of G15421: signal is true;
	signal G15422: std_logic; attribute dont_touch of G15422: signal is true;
	signal G15423: std_logic; attribute dont_touch of G15423: signal is true;
	signal G15424: std_logic; attribute dont_touch of G15424: signal is true;
	signal G15425: std_logic; attribute dont_touch of G15425: signal is true;
	signal G15426: std_logic; attribute dont_touch of G15426: signal is true;
	signal G15429: std_logic; attribute dont_touch of G15429: signal is true;
	signal G15432: std_logic; attribute dont_touch of G15432: signal is true;
	signal G15435: std_logic; attribute dont_touch of G15435: signal is true;
	signal G15436: std_logic; attribute dont_touch of G15436: signal is true;
	signal G15437: std_logic; attribute dont_touch of G15437: signal is true;
	signal G15438: std_logic; attribute dont_touch of G15438: signal is true;
	signal G15439: std_logic; attribute dont_touch of G15439: signal is true;
	signal G15440: std_logic; attribute dont_touch of G15440: signal is true;
	signal G15441: std_logic; attribute dont_touch of G15441: signal is true;
	signal G15442: std_logic; attribute dont_touch of G15442: signal is true;
	signal G15443: std_logic; attribute dont_touch of G15443: signal is true;
	signal G15446: std_logic; attribute dont_touch of G15446: signal is true;
	signal G15449: std_logic; attribute dont_touch of G15449: signal is true;
	signal G15452: std_logic; attribute dont_touch of G15452: signal is true;
	signal G15453: std_logic; attribute dont_touch of G15453: signal is true;
	signal G15454: std_logic; attribute dont_touch of G15454: signal is true;
	signal G15458: std_logic; attribute dont_touch of G15458: signal is true;
	signal G15459: std_logic; attribute dont_touch of G15459: signal is true;
	signal G15460: std_logic; attribute dont_touch of G15460: signal is true;
	signal G15461: std_logic; attribute dont_touch of G15461: signal is true;
	signal G15464: std_logic; attribute dont_touch of G15464: signal is true;
	signal G15467: std_logic; attribute dont_touch of G15467: signal is true;
	signal G15470: std_logic; attribute dont_touch of G15470: signal is true;
	signal G15471: std_logic; attribute dont_touch of G15471: signal is true;
	signal G15474: std_logic; attribute dont_touch of G15474: signal is true;
	signal G15475: std_logic; attribute dont_touch of G15475: signal is true;
	signal G15476: std_logic; attribute dont_touch of G15476: signal is true;
	signal G15477: std_logic; attribute dont_touch of G15477: signal is true;
	signal G15480: std_logic; attribute dont_touch of G15480: signal is true;
	signal G15483: std_logic; attribute dont_touch of G15483: signal is true;
	signal G15486: std_logic; attribute dont_touch of G15486: signal is true;
	signal G15487: std_logic; attribute dont_touch of G15487: signal is true;
	signal G15488: std_logic; attribute dont_touch of G15488: signal is true;
	signal G15491: std_logic; attribute dont_touch of G15491: signal is true;
	signal G15492: std_logic; attribute dont_touch of G15492: signal is true;
	signal G15493: std_logic; attribute dont_touch of G15493: signal is true;
	signal G15494: std_logic; attribute dont_touch of G15494: signal is true;
	signal G15495: std_logic; attribute dont_touch of G15495: signal is true;
	signal G15496: std_logic; attribute dont_touch of G15496: signal is true;
	signal G15499: std_logic; attribute dont_touch of G15499: signal is true;
	signal G15502: std_logic; attribute dont_touch of G15502: signal is true;
	signal G15505: std_logic; attribute dont_touch of G15505: signal is true;
	signal G15506: std_logic; attribute dont_touch of G15506: signal is true;
	signal G15507: std_logic; attribute dont_touch of G15507: signal is true;
	signal G15508: std_logic; attribute dont_touch of G15508: signal is true;
	signal G15509: std_logic; attribute dont_touch of G15509: signal is true;
	signal G15510: std_logic; attribute dont_touch of G15510: signal is true;
	signal G15513: std_logic; attribute dont_touch of G15513: signal is true;
	signal G15516: std_logic; attribute dont_touch of G15516: signal is true;
	signal G15519: std_logic; attribute dont_touch of G15519: signal is true;
	signal G15520: std_logic; attribute dont_touch of G15520: signal is true;
	signal G15521: std_logic; attribute dont_touch of G15521: signal is true;
	signal G15524: std_logic; attribute dont_touch of G15524: signal is true;
	signal G15525: std_logic; attribute dont_touch of G15525: signal is true;
	signal G15526: std_logic; attribute dont_touch of G15526: signal is true;
	signal G15527: std_logic; attribute dont_touch of G15527: signal is true;
	signal G15528: std_logic; attribute dont_touch of G15528: signal is true;
	signal G15531: std_logic; attribute dont_touch of G15531: signal is true;
	signal G15534: std_logic; attribute dont_touch of G15534: signal is true;
	signal G15537: std_logic; attribute dont_touch of G15537: signal is true;
	signal G15540: std_logic; attribute dont_touch of G15540: signal is true;
	signal G15544: std_logic; attribute dont_touch of G15544: signal is true;
	signal G15545: std_logic; attribute dont_touch of G15545: signal is true;
	signal G15546: std_logic; attribute dont_touch of G15546: signal is true;
	signal G15547: std_logic; attribute dont_touch of G15547: signal is true;
	signal G15550: std_logic; attribute dont_touch of G15550: signal is true;
	signal G15553: std_logic; attribute dont_touch of G15553: signal is true;
	signal G15556: std_logic; attribute dont_touch of G15556: signal is true;
	signal G15557: std_logic; attribute dont_touch of G15557: signal is true;
	signal G15560: std_logic; attribute dont_touch of G15560: signal is true;
	signal G15561: std_logic; attribute dont_touch of G15561: signal is true;
	signal G15562: std_logic; attribute dont_touch of G15562: signal is true;
	signal G15563: std_logic; attribute dont_touch of G15563: signal is true;
	signal G15566: std_logic; attribute dont_touch of G15566: signal is true;
	signal G15569: std_logic; attribute dont_touch of G15569: signal is true;
	signal G15572: std_logic; attribute dont_touch of G15572: signal is true;
	signal G15573: std_logic; attribute dont_touch of G15573: signal is true;
	signal G15574: std_logic; attribute dont_touch of G15574: signal is true;
	signal G15577: std_logic; attribute dont_touch of G15577: signal is true;
	signal G15578: std_logic; attribute dont_touch of G15578: signal is true;
	signal G15579: std_logic; attribute dont_touch of G15579: signal is true;
	signal G15580: std_logic; attribute dont_touch of G15580: signal is true;
	signal G15581: std_logic; attribute dont_touch of G15581: signal is true;
	signal G15582: std_logic; attribute dont_touch of G15582: signal is true;
	signal G15585: std_logic; attribute dont_touch of G15585: signal is true;
	signal G15588: std_logic; attribute dont_touch of G15588: signal is true;
	signal G15591: std_logic; attribute dont_touch of G15591: signal is true;
	signal G15592: std_logic; attribute dont_touch of G15592: signal is true;
	signal G15593: std_logic; attribute dont_touch of G15593: signal is true;
	signal G15594: std_logic; attribute dont_touch of G15594: signal is true;
	signal G15595: std_logic; attribute dont_touch of G15595: signal is true;
	signal G15596: std_logic; attribute dont_touch of G15596: signal is true;
	signal G15599: std_logic; attribute dont_touch of G15599: signal is true;
	signal G15602: std_logic; attribute dont_touch of G15602: signal is true;
	signal G15603: std_logic; attribute dont_touch of G15603: signal is true;
	signal G15604: std_logic; attribute dont_touch of G15604: signal is true;
	signal G15605: std_logic; attribute dont_touch of G15605: signal is true;
	signal G15606: std_logic; attribute dont_touch of G15606: signal is true;
	signal G15609: std_logic; attribute dont_touch of G15609: signal is true;
	signal G15612: std_logic; attribute dont_touch of G15612: signal is true;
	signal G15615: std_logic; attribute dont_touch of G15615: signal is true;
	signal G15618: std_logic; attribute dont_touch of G15618: signal is true;
	signal G15622: std_logic; attribute dont_touch of G15622: signal is true;
	signal G15623: std_logic; attribute dont_touch of G15623: signal is true;
	signal G15624: std_logic; attribute dont_touch of G15624: signal is true;
	signal G15625: std_logic; attribute dont_touch of G15625: signal is true;
	signal G15628: std_logic; attribute dont_touch of G15628: signal is true;
	signal G15631: std_logic; attribute dont_touch of G15631: signal is true;
	signal G15634: std_logic; attribute dont_touch of G15634: signal is true;
	signal G15635: std_logic; attribute dont_touch of G15635: signal is true;
	signal G15638: std_logic; attribute dont_touch of G15638: signal is true;
	signal G15639: std_logic; attribute dont_touch of G15639: signal is true;
	signal G15640: std_logic; attribute dont_touch of G15640: signal is true;
	signal G15641: std_logic; attribute dont_touch of G15641: signal is true;
	signal G15644: std_logic; attribute dont_touch of G15644: signal is true;
	signal G15647: std_logic; attribute dont_touch of G15647: signal is true;
	signal G15650: std_logic; attribute dont_touch of G15650: signal is true;
	signal G15651: std_logic; attribute dont_touch of G15651: signal is true;
	signal G15652: std_logic; attribute dont_touch of G15652: signal is true;
	signal G15655: std_logic; attribute dont_touch of G15655: signal is true;
	signal G15658: std_logic; attribute dont_touch of G15658: signal is true;
	signal G15659: std_logic; attribute dont_touch of G15659: signal is true;
	signal G15660: std_logic; attribute dont_touch of G15660: signal is true;
	signal G15661: std_logic; attribute dont_touch of G15661: signal is true;
	signal G15664: std_logic; attribute dont_touch of G15664: signal is true;
	signal G15665: std_logic; attribute dont_touch of G15665: signal is true;
	signal G15666: std_logic; attribute dont_touch of G15666: signal is true;
	signal G15667: std_logic; attribute dont_touch of G15667: signal is true;
	signal G15670: std_logic; attribute dont_touch of G15670: signal is true;
	signal G15671: std_logic; attribute dont_touch of G15671: signal is true;
	signal G15672: std_logic; attribute dont_touch of G15672: signal is true;
	signal G15675: std_logic; attribute dont_touch of G15675: signal is true;
	signal G15678: std_logic; attribute dont_touch of G15678: signal is true;
	signal G15679: std_logic; attribute dont_touch of G15679: signal is true;
	signal G15680: std_logic; attribute dont_touch of G15680: signal is true;
	signal G15681: std_logic; attribute dont_touch of G15681: signal is true;
	signal G15682: std_logic; attribute dont_touch of G15682: signal is true;
	signal G15685: std_logic; attribute dont_touch of G15685: signal is true;
	signal G15688: std_logic; attribute dont_touch of G15688: signal is true;
	signal G15691: std_logic; attribute dont_touch of G15691: signal is true;
	signal G15694: std_logic; attribute dont_touch of G15694: signal is true;
	signal G15698: std_logic; attribute dont_touch of G15698: signal is true;
	signal G15699: std_logic; attribute dont_touch of G15699: signal is true;
	signal G15700: std_logic; attribute dont_touch of G15700: signal is true;
	signal G15701: std_logic; attribute dont_touch of G15701: signal is true;
	signal G15704: std_logic; attribute dont_touch of G15704: signal is true;
	signal G15707: std_logic; attribute dont_touch of G15707: signal is true;
	signal G15710: std_logic; attribute dont_touch of G15710: signal is true;
	signal G15711: std_logic; attribute dont_touch of G15711: signal is true;
	signal G15714: std_logic; attribute dont_touch of G15714: signal is true;
	signal G15717: std_logic; attribute dont_touch of G15717: signal is true;
	signal G15718: std_logic; attribute dont_touch of G15718: signal is true;
	signal G15719: std_logic; attribute dont_touch of G15719: signal is true;
	signal G15720: std_logic; attribute dont_touch of G15720: signal is true;
	signal G15721: std_logic; attribute dont_touch of G15721: signal is true;
	signal G15722: std_logic; attribute dont_touch of G15722: signal is true;
	signal G15723: std_logic; attribute dont_touch of G15723: signal is true;
	signal G15724: std_logic; attribute dont_touch of G15724: signal is true;
	signal G15725: std_logic; attribute dont_touch of G15725: signal is true;
	signal G15726: std_logic; attribute dont_touch of G15726: signal is true;
	signal G15729: std_logic; attribute dont_touch of G15729: signal is true;
	signal G15730: std_logic; attribute dont_touch of G15730: signal is true;
	signal G15731: std_logic; attribute dont_touch of G15731: signal is true;
	signal G15734: std_logic; attribute dont_touch of G15734: signal is true;
	signal G15737: std_logic; attribute dont_touch of G15737: signal is true;
	signal G15738: std_logic; attribute dont_touch of G15738: signal is true;
	signal G15739: std_logic; attribute dont_touch of G15739: signal is true;
	signal G15740: std_logic; attribute dont_touch of G15740: signal is true;
	signal G15741: std_logic; attribute dont_touch of G15741: signal is true;
	signal G15744: std_logic; attribute dont_touch of G15744: signal is true;
	signal G15747: std_logic; attribute dont_touch of G15747: signal is true;
	signal G15750: std_logic; attribute dont_touch of G15750: signal is true;
	signal G15753: std_logic; attribute dont_touch of G15753: signal is true;
	signal G15754: std_logic; attribute dont_touch of G15754: signal is true;
	signal G15755: std_logic; attribute dont_touch of G15755: signal is true;
	signal G15756: std_logic; attribute dont_touch of G15756: signal is true;
	signal G15757: std_logic; attribute dont_touch of G15757: signal is true;
	signal G15758: std_logic; attribute dont_touch of G15758: signal is true;
	signal G15759: std_logic; attribute dont_touch of G15759: signal is true;
	signal G15760: std_logic; attribute dont_touch of G15760: signal is true;
	signal G15761: std_logic; attribute dont_touch of G15761: signal is true;
	signal G15762: std_logic; attribute dont_touch of G15762: signal is true;
	signal G15763: std_logic; attribute dont_touch of G15763: signal is true;
	signal G15764: std_logic; attribute dont_touch of G15764: signal is true;
	signal G15765: std_logic; attribute dont_touch of G15765: signal is true;
	signal G15766: std_logic; attribute dont_touch of G15766: signal is true;
	signal G15769: std_logic; attribute dont_touch of G15769: signal is true;
	signal G15770: std_logic; attribute dont_touch of G15770: signal is true;
	signal G15771: std_logic; attribute dont_touch of G15771: signal is true;
	signal G15774: std_logic; attribute dont_touch of G15774: signal is true;
	signal G15777: std_logic; attribute dont_touch of G15777: signal is true;
	signal G15780: std_logic; attribute dont_touch of G15780: signal is true;
	signal G15781: std_logic; attribute dont_touch of G15781: signal is true;
	signal G15782: std_logic; attribute dont_touch of G15782: signal is true;
	signal G15783: std_logic; attribute dont_touch of G15783: signal is true;
	signal G15784: std_logic; attribute dont_touch of G15784: signal is true;
	signal G15785: std_logic; attribute dont_touch of G15785: signal is true;
	signal G15786: std_logic; attribute dont_touch of G15786: signal is true;
	signal G15787: std_logic; attribute dont_touch of G15787: signal is true;
	signal G15788: std_logic; attribute dont_touch of G15788: signal is true;
	signal G15789: std_logic; attribute dont_touch of G15789: signal is true;
	signal G15790: std_logic; attribute dont_touch of G15790: signal is true;
	signal G15791: std_logic; attribute dont_touch of G15791: signal is true;
	signal G15792: std_logic; attribute dont_touch of G15792: signal is true;
	signal G15793: std_logic; attribute dont_touch of G15793: signal is true;
	signal G15794: std_logic; attribute dont_touch of G15794: signal is true;
	signal G15797: std_logic; attribute dont_touch of G15797: signal is true;
	signal G15800: std_logic; attribute dont_touch of G15800: signal is true;
	signal G15801: std_logic; attribute dont_touch of G15801: signal is true;
	signal G15802: std_logic; attribute dont_touch of G15802: signal is true;
	signal G15803: std_logic; attribute dont_touch of G15803: signal is true;
	signal G15804: std_logic; attribute dont_touch of G15804: signal is true;
	signal G15805: std_logic; attribute dont_touch of G15805: signal is true;
	signal G15806: std_logic; attribute dont_touch of G15806: signal is true;
	signal G15807: std_logic; attribute dont_touch of G15807: signal is true;
	signal G15808: std_logic; attribute dont_touch of G15808: signal is true;
	signal G15809: std_logic; attribute dont_touch of G15809: signal is true;
	signal G15810: std_logic; attribute dont_touch of G15810: signal is true;
	signal G15811: std_logic; attribute dont_touch of G15811: signal is true;
	signal G15812: std_logic; attribute dont_touch of G15812: signal is true;
	signal G15813: std_logic; attribute dont_touch of G15813: signal is true;
	signal G15814: std_logic; attribute dont_touch of G15814: signal is true;
	signal G15817: std_logic; attribute dont_touch of G15817: signal is true;
	signal G15818: std_logic; attribute dont_touch of G15818: signal is true;
	signal G15819: std_logic; attribute dont_touch of G15819: signal is true;
	signal G15820: std_logic; attribute dont_touch of G15820: signal is true;
	signal G15821: std_logic; attribute dont_touch of G15821: signal is true;
	signal G15822: std_logic; attribute dont_touch of G15822: signal is true;
	signal G15823: std_logic; attribute dont_touch of G15823: signal is true;
	signal G15824: std_logic; attribute dont_touch of G15824: signal is true;
	signal G15825: std_logic; attribute dont_touch of G15825: signal is true;
	signal G15826: std_logic; attribute dont_touch of G15826: signal is true;
	signal G15827: std_logic; attribute dont_touch of G15827: signal is true;
	signal G15828: std_logic; attribute dont_touch of G15828: signal is true;
	signal G15829: std_logic; attribute dont_touch of G15829: signal is true;
	signal G15830: std_logic; attribute dont_touch of G15830: signal is true;
	signal G15831: std_logic; attribute dont_touch of G15831: signal is true;
	signal G15832: std_logic; attribute dont_touch of G15832: signal is true;
	signal G15833: std_logic; attribute dont_touch of G15833: signal is true;
	signal G15834: std_logic; attribute dont_touch of G15834: signal is true;
	signal G15835: std_logic; attribute dont_touch of G15835: signal is true;
	signal G15836: std_logic; attribute dont_touch of G15836: signal is true;
	signal G15837: std_logic; attribute dont_touch of G15837: signal is true;
	signal G15838: std_logic; attribute dont_touch of G15838: signal is true;
	signal G15839: std_logic; attribute dont_touch of G15839: signal is true;
	signal G15840: std_logic; attribute dont_touch of G15840: signal is true;
	signal G15841: std_logic; attribute dont_touch of G15841: signal is true;
	signal G15842: std_logic; attribute dont_touch of G15842: signal is true;
	signal G15843: std_logic; attribute dont_touch of G15843: signal is true;
	signal G15844: std_logic; attribute dont_touch of G15844: signal is true;
	signal G15845: std_logic; attribute dont_touch of G15845: signal is true;
	signal G15846: std_logic; attribute dont_touch of G15846: signal is true;
	signal G15847: std_logic; attribute dont_touch of G15847: signal is true;
	signal G15848: std_logic; attribute dont_touch of G15848: signal is true;
	signal G15849: std_logic; attribute dont_touch of G15849: signal is true;
	signal G15850: std_logic; attribute dont_touch of G15850: signal is true;
	signal G15851: std_logic; attribute dont_touch of G15851: signal is true;
	signal G15852: std_logic; attribute dont_touch of G15852: signal is true;
	signal G15853: std_logic; attribute dont_touch of G15853: signal is true;
	signal G15854: std_logic; attribute dont_touch of G15854: signal is true;
	signal G15855: std_logic; attribute dont_touch of G15855: signal is true;
	signal G15856: std_logic; attribute dont_touch of G15856: signal is true;
	signal G15857: std_logic; attribute dont_touch of G15857: signal is true;
	signal G15858: std_logic; attribute dont_touch of G15858: signal is true;
	signal G15859: std_logic; attribute dont_touch of G15859: signal is true;
	signal G15866: std_logic; attribute dont_touch of G15866: signal is true;
	signal G15867: std_logic; attribute dont_touch of G15867: signal is true;
	signal G15868: std_logic; attribute dont_touch of G15868: signal is true;
	signal G15869: std_logic; attribute dont_touch of G15869: signal is true;
	signal G15870: std_logic; attribute dont_touch of G15870: signal is true;
	signal G15871: std_logic; attribute dont_touch of G15871: signal is true;
	signal G15872: std_logic; attribute dont_touch of G15872: signal is true;
	signal G15873: std_logic; attribute dont_touch of G15873: signal is true;
	signal G15876: std_logic; attribute dont_touch of G15876: signal is true;
	signal G15877: std_logic; attribute dont_touch of G15877: signal is true;
	signal G15878: std_logic; attribute dont_touch of G15878: signal is true;
	signal G15879: std_logic; attribute dont_touch of G15879: signal is true;
	signal G15880: std_logic; attribute dont_touch of G15880: signal is true;
	signal G15887: std_logic; attribute dont_touch of G15887: signal is true;
	signal G15888: std_logic; attribute dont_touch of G15888: signal is true;
	signal G15889: std_logic; attribute dont_touch of G15889: signal is true;
	signal G15890: std_logic; attribute dont_touch of G15890: signal is true;
	signal G15897: std_logic; attribute dont_touch of G15897: signal is true;
	signal G15898: std_logic; attribute dont_touch of G15898: signal is true;
	signal G15899: std_logic; attribute dont_touch of G15899: signal is true;
	signal G15900: std_logic; attribute dont_touch of G15900: signal is true;
	signal G15901: std_logic; attribute dont_touch of G15901: signal is true;
	signal G15902: std_logic; attribute dont_touch of G15902: signal is true;
	signal G15903: std_logic; attribute dont_touch of G15903: signal is true;
	signal G15904: std_logic; attribute dont_touch of G15904: signal is true;
	signal G15912: std_logic; attribute dont_touch of G15912: signal is true;
	signal G15913: std_logic; attribute dont_touch of G15913: signal is true;
	signal G15920: std_logic; attribute dont_touch of G15920: signal is true;
	signal G15921: std_logic; attribute dont_touch of G15921: signal is true;
	signal G15922: std_logic; attribute dont_touch of G15922: signal is true;
	signal G15923: std_logic; attribute dont_touch of G15923: signal is true;
	signal G15930: std_logic; attribute dont_touch of G15930: signal is true;
	signal G15931: std_logic; attribute dont_touch of G15931: signal is true;
	signal G15932: std_logic; attribute dont_touch of G15932: signal is true;
	signal G15933: std_logic; attribute dont_touch of G15933: signal is true;
	signal G15941: std_logic; attribute dont_touch of G15941: signal is true;
	signal G15942: std_logic; attribute dont_touch of G15942: signal is true;
	signal G15949: std_logic; attribute dont_touch of G15949: signal is true;
	signal G15950: std_logic; attribute dont_touch of G15950: signal is true;
	signal G15951: std_logic; attribute dont_touch of G15951: signal is true;
	signal G15952: std_logic; attribute dont_touch of G15952: signal is true;
	signal G15959: std_logic; attribute dont_touch of G15959: signal is true;
	signal G15962: std_logic; attribute dont_touch of G15962: signal is true;
	signal G15970: std_logic; attribute dont_touch of G15970: signal is true;
	signal G15971: std_logic; attribute dont_touch of G15971: signal is true;
	signal G15978: std_logic; attribute dont_touch of G15978: signal is true;
	signal G15981: std_logic; attribute dont_touch of G15981: signal is true;
	signal G15989: std_logic; attribute dont_touch of G15989: signal is true;
	signal G15990: std_logic; attribute dont_touch of G15990: signal is true;
	signal G15991: std_logic; attribute dont_touch of G15991: signal is true;
	signal G15992: std_logic; attribute dont_touch of G15992: signal is true;
	signal G15993: std_logic; attribute dont_touch of G15993: signal is true;
	signal G15994: std_logic; attribute dont_touch of G15994: signal is true;
	signal G15995: std_logic; attribute dont_touch of G15995: signal is true;
	signal G15996: std_logic; attribute dont_touch of G15996: signal is true;
	signal G15997: std_logic; attribute dont_touch of G15997: signal is true;
	signal G15998: std_logic; attribute dont_touch of G15998: signal is true;
	signal G15999: std_logic; attribute dont_touch of G15999: signal is true;
	signal G16000: std_logic; attribute dont_touch of G16000: signal is true;
	signal G16001: std_logic; attribute dont_touch of G16001: signal is true;
	signal G16002: std_logic; attribute dont_touch of G16002: signal is true;
	signal G16003: std_logic; attribute dont_touch of G16003: signal is true;
	signal G16004: std_logic; attribute dont_touch of G16004: signal is true;
	signal G16005: std_logic; attribute dont_touch of G16005: signal is true;
	signal G16006: std_logic; attribute dont_touch of G16006: signal is true;
	signal G16007: std_logic; attribute dont_touch of G16007: signal is true;
	signal G16008: std_logic; attribute dont_touch of G16008: signal is true;
	signal G16009: std_logic; attribute dont_touch of G16009: signal is true;
	signal G16010: std_logic; attribute dont_touch of G16010: signal is true;
	signal G16011: std_logic; attribute dont_touch of G16011: signal is true;
	signal G16012: std_logic; attribute dont_touch of G16012: signal is true;
	signal G16013: std_logic; attribute dont_touch of G16013: signal is true;
	signal G16014: std_logic; attribute dont_touch of G16014: signal is true;
	signal G16015: std_logic; attribute dont_touch of G16015: signal is true;
	signal G16016: std_logic; attribute dont_touch of G16016: signal is true;
	signal G16017: std_logic; attribute dont_touch of G16017: signal is true;
	signal G16018: std_logic; attribute dont_touch of G16018: signal is true;
	signal G16019: std_logic; attribute dont_touch of G16019: signal is true;
	signal G16020: std_logic; attribute dont_touch of G16020: signal is true;
	signal G16023: std_logic; attribute dont_touch of G16023: signal is true;
	signal G16024: std_logic; attribute dont_touch of G16024: signal is true;
	signal G16025: std_logic; attribute dont_touch of G16025: signal is true;
	signal G16026: std_logic; attribute dont_touch of G16026: signal is true;
	signal G16027: std_logic; attribute dont_touch of G16027: signal is true;
	signal G16028: std_logic; attribute dont_touch of G16028: signal is true;
	signal G16029: std_logic; attribute dont_touch of G16029: signal is true;
	signal G16030: std_logic; attribute dont_touch of G16030: signal is true;
	signal G16031: std_logic; attribute dont_touch of G16031: signal is true;
	signal G16032: std_logic; attribute dont_touch of G16032: signal is true;
	signal G16033: std_logic; attribute dont_touch of G16033: signal is true;
	signal G16034: std_logic; attribute dont_touch of G16034: signal is true;
	signal G16035: std_logic; attribute dont_touch of G16035: signal is true;
	signal G16036: std_logic; attribute dont_touch of G16036: signal is true;
	signal G16039: std_logic; attribute dont_touch of G16039: signal is true;
	signal G16040: std_logic; attribute dont_touch of G16040: signal is true;
	signal G16041: std_logic; attribute dont_touch of G16041: signal is true;
	signal G16042: std_logic; attribute dont_touch of G16042: signal is true;
	signal G16043: std_logic; attribute dont_touch of G16043: signal is true;
	signal G16044: std_logic; attribute dont_touch of G16044: signal is true;
	signal G16045: std_logic; attribute dont_touch of G16045: signal is true;
	signal G16046: std_logic; attribute dont_touch of G16046: signal is true;
	signal G16047: std_logic; attribute dont_touch of G16047: signal is true;
	signal G16048: std_logic; attribute dont_touch of G16048: signal is true;
	signal G16049: std_logic; attribute dont_touch of G16049: signal is true;
	signal G16050: std_logic; attribute dont_touch of G16050: signal is true;
	signal G16051: std_logic; attribute dont_touch of G16051: signal is true;
	signal G16052: std_logic; attribute dont_touch of G16052: signal is true;
	signal G16053: std_logic; attribute dont_touch of G16053: signal is true;
	signal G16054: std_logic; attribute dont_touch of G16054: signal is true;
	signal G16055: std_logic; attribute dont_touch of G16055: signal is true;
	signal G16056: std_logic; attribute dont_touch of G16056: signal is true;
	signal G16057: std_logic; attribute dont_touch of G16057: signal is true;
	signal G16058: std_logic; attribute dont_touch of G16058: signal is true;
	signal G16061: std_logic; attribute dont_touch of G16061: signal is true;
	signal G16062: std_logic; attribute dont_touch of G16062: signal is true;
	signal G16063: std_logic; attribute dont_touch of G16063: signal is true;
	signal G16064: std_logic; attribute dont_touch of G16064: signal is true;
	signal G16065: std_logic; attribute dont_touch of G16065: signal is true;
	signal G16066: std_logic; attribute dont_touch of G16066: signal is true;
	signal G16067: std_logic; attribute dont_touch of G16067: signal is true;
	signal G16068: std_logic; attribute dont_touch of G16068: signal is true;
	signal G16069: std_logic; attribute dont_touch of G16069: signal is true;
	signal G16070: std_logic; attribute dont_touch of G16070: signal is true;
	signal G16071: std_logic; attribute dont_touch of G16071: signal is true;
	signal G16072: std_logic; attribute dont_touch of G16072: signal is true;
	signal G16073: std_logic; attribute dont_touch of G16073: signal is true;
	signal G16074: std_logic; attribute dont_touch of G16074: signal is true;
	signal G16075: std_logic; attribute dont_touch of G16075: signal is true;
	signal G16081: std_logic; attribute dont_touch of G16081: signal is true;
	signal G16082: std_logic; attribute dont_touch of G16082: signal is true;
	signal G16085: std_logic; attribute dont_touch of G16085: signal is true;
	signal G16088: std_logic; attribute dont_touch of G16088: signal is true;
	signal G16089: std_logic; attribute dont_touch of G16089: signal is true;
	signal G16090: std_logic; attribute dont_touch of G16090: signal is true;
	signal G16091: std_logic; attribute dont_touch of G16091: signal is true;
	signal G16092: std_logic; attribute dont_touch of G16092: signal is true;
	signal G16093: std_logic; attribute dont_touch of G16093: signal is true;
	signal G16094: std_logic; attribute dont_touch of G16094: signal is true;
	signal G16097: std_logic; attribute dont_touch of G16097: signal is true;
	signal G16098: std_logic; attribute dont_touch of G16098: signal is true;
	signal G16099: std_logic; attribute dont_touch of G16099: signal is true;
	signal G16100: std_logic; attribute dont_touch of G16100: signal is true;
	signal G16101: std_logic; attribute dont_touch of G16101: signal is true;
	signal G16102: std_logic; attribute dont_touch of G16102: signal is true;
	signal G16103: std_logic; attribute dont_touch of G16103: signal is true;
	signal G16104: std_logic; attribute dont_touch of G16104: signal is true;
	signal G16105: std_logic; attribute dont_touch of G16105: signal is true;
	signal G16106: std_logic; attribute dont_touch of G16106: signal is true;
	signal G16107: std_logic; attribute dont_touch of G16107: signal is true;
	signal G16108: std_logic; attribute dont_touch of G16108: signal is true;
	signal G16109: std_logic; attribute dont_touch of G16109: signal is true;
	signal G16110: std_logic; attribute dont_touch of G16110: signal is true;
	signal G16111: std_logic; attribute dont_touch of G16111: signal is true;
	signal G16112: std_logic; attribute dont_touch of G16112: signal is true;
	signal G16113: std_logic; attribute dont_touch of G16113: signal is true;
	signal G16119: std_logic; attribute dont_touch of G16119: signal is true;
	signal G16120: std_logic; attribute dont_touch of G16120: signal is true;
	signal G16123: std_logic; attribute dont_touch of G16123: signal is true;
	signal G16126: std_logic; attribute dont_touch of G16126: signal is true;
	signal G16127: std_logic; attribute dont_touch of G16127: signal is true;
	signal G16128: std_logic; attribute dont_touch of G16128: signal is true;
	signal G16129: std_logic; attribute dont_touch of G16129: signal is true;
	signal G16130: std_logic; attribute dont_touch of G16130: signal is true;
	signal G16131: std_logic; attribute dont_touch of G16131: signal is true;
	signal G16132: std_logic; attribute dont_touch of G16132: signal is true;
	signal G16133: std_logic; attribute dont_touch of G16133: signal is true;
	signal G16134: std_logic; attribute dont_touch of G16134: signal is true;
	signal G16135: std_logic; attribute dont_touch of G16135: signal is true;
	signal G16136: std_logic; attribute dont_touch of G16136: signal is true;
	signal G16137: std_logic; attribute dont_touch of G16137: signal is true;
	signal G16138: std_logic; attribute dont_touch of G16138: signal is true;
	signal G16139: std_logic; attribute dont_touch of G16139: signal is true;
	signal G16140: std_logic; attribute dont_touch of G16140: signal is true;
	signal G16141: std_logic; attribute dont_touch of G16141: signal is true;
	signal G16142: std_logic; attribute dont_touch of G16142: signal is true;
	signal G16152: std_logic; attribute dont_touch of G16152: signal is true;
	signal G16153: std_logic; attribute dont_touch of G16153: signal is true;
	signal G16154: std_logic; attribute dont_touch of G16154: signal is true;
	signal G16158: std_logic; attribute dont_touch of G16158: signal is true;
	signal G16159: std_logic; attribute dont_touch of G16159: signal is true;
	signal G16160: std_logic; attribute dont_touch of G16160: signal is true;
	signal G16161: std_logic; attribute dont_touch of G16161: signal is true;
	signal G16162: std_logic; attribute dont_touch of G16162: signal is true;
	signal G16163: std_logic; attribute dont_touch of G16163: signal is true;
	signal G16164: std_logic; attribute dont_touch of G16164: signal is true;
	signal G16170: std_logic; attribute dont_touch of G16170: signal is true;
	signal G16171: std_logic; attribute dont_touch of G16171: signal is true;
	signal G16174: std_logic; attribute dont_touch of G16174: signal is true;
	signal G16177: std_logic; attribute dont_touch of G16177: signal is true;
	signal G16178: std_logic; attribute dont_touch of G16178: signal is true;
	signal G16179: std_logic; attribute dont_touch of G16179: signal is true;
	signal G16180: std_logic; attribute dont_touch of G16180: signal is true;
	signal G16181: std_logic; attribute dont_touch of G16181: signal is true;
	signal G16182: std_logic; attribute dont_touch of G16182: signal is true;
	signal G16183: std_logic; attribute dont_touch of G16183: signal is true;
	signal G16184: std_logic; attribute dont_touch of G16184: signal is true;
	signal G16185: std_logic; attribute dont_touch of G16185: signal is true;
	signal G16186: std_logic; attribute dont_touch of G16186: signal is true;
	signal G16187: std_logic; attribute dont_touch of G16187: signal is true;
	signal G16188: std_logic; attribute dont_touch of G16188: signal is true;
	signal G16189: std_logic; attribute dont_touch of G16189: signal is true;
	signal G16197: std_logic; attribute dont_touch of G16197: signal is true;
	signal G16198: std_logic; attribute dont_touch of G16198: signal is true;
	signal G16199: std_logic; attribute dont_touch of G16199: signal is true;
	signal G16200: std_logic; attribute dont_touch of G16200: signal is true;
	signal G16201: std_logic; attribute dont_touch of G16201: signal is true;
	signal G16211: std_logic; attribute dont_touch of G16211: signal is true;
	signal G16212: std_logic; attribute dont_touch of G16212: signal is true;
	signal G16213: std_logic; attribute dont_touch of G16213: signal is true;
	signal G16217: std_logic; attribute dont_touch of G16217: signal is true;
	signal G16218: std_logic; attribute dont_touch of G16218: signal is true;
	signal G16219: std_logic; attribute dont_touch of G16219: signal is true;
	signal G16220: std_logic; attribute dont_touch of G16220: signal is true;
	signal G16221: std_logic; attribute dont_touch of G16221: signal is true;
	signal G16222: std_logic; attribute dont_touch of G16222: signal is true;
	signal G16223: std_logic; attribute dont_touch of G16223: signal is true;
	signal G16229: std_logic; attribute dont_touch of G16229: signal is true;
	signal G16230: std_logic; attribute dont_touch of G16230: signal is true;
	signal G16233: std_logic; attribute dont_touch of G16233: signal is true;
	signal G16236: std_logic; attribute dont_touch of G16236: signal is true;
	signal G16237: std_logic; attribute dont_touch of G16237: signal is true;
	signal G16238: std_logic; attribute dont_touch of G16238: signal is true;
	signal G16239: std_logic; attribute dont_touch of G16239: signal is true;
	signal G16240: std_logic; attribute dont_touch of G16240: signal is true;
	signal G16241: std_logic; attribute dont_touch of G16241: signal is true;
	signal G16242: std_logic; attribute dont_touch of G16242: signal is true;
	signal G16243: std_logic; attribute dont_touch of G16243: signal is true;
	signal G16250: std_logic; attribute dont_touch of G16250: signal is true;
	signal G16251: std_logic; attribute dont_touch of G16251: signal is true;
	signal G16252: std_logic; attribute dont_touch of G16252: signal is true;
	signal G16253: std_logic; attribute dont_touch of G16253: signal is true;
	signal G16254: std_logic; attribute dont_touch of G16254: signal is true;
	signal G16262: std_logic; attribute dont_touch of G16262: signal is true;
	signal G16263: std_logic; attribute dont_touch of G16263: signal is true;
	signal G16264: std_logic; attribute dont_touch of G16264: signal is true;
	signal G16265: std_logic; attribute dont_touch of G16265: signal is true;
	signal G16266: std_logic; attribute dont_touch of G16266: signal is true;
	signal G16276: std_logic; attribute dont_touch of G16276: signal is true;
	signal G16277: std_logic; attribute dont_touch of G16277: signal is true;
	signal G16278: std_logic; attribute dont_touch of G16278: signal is true;
	signal G16282: std_logic; attribute dont_touch of G16282: signal is true;
	signal G16283: std_logic; attribute dont_touch of G16283: signal is true;
	signal G16284: std_logic; attribute dont_touch of G16284: signal is true;
	signal G16285: std_logic; attribute dont_touch of G16285: signal is true;
	signal G16286: std_logic; attribute dont_touch of G16286: signal is true;
	signal G16287: std_logic; attribute dont_touch of G16287: signal is true;
	signal G16288: std_logic; attribute dont_touch of G16288: signal is true;
	signal G16289: std_logic; attribute dont_touch of G16289: signal is true;
	signal G16290: std_logic; attribute dont_touch of G16290: signal is true;
	signal G16291: std_logic; attribute dont_touch of G16291: signal is true;
	signal G16292: std_logic; attribute dont_touch of G16292: signal is true;
	signal G16293: std_logic; attribute dont_touch of G16293: signal is true;
	signal G16298: std_logic; attribute dont_touch of G16298: signal is true;
	signal G16299: std_logic; attribute dont_touch of G16299: signal is true;
	signal G16300: std_logic; attribute dont_touch of G16300: signal is true;
	signal G16301: std_logic; attribute dont_touch of G16301: signal is true;
	signal G16302: std_logic; attribute dont_touch of G16302: signal is true;
	signal G16309: std_logic; attribute dont_touch of G16309: signal is true;
	signal G16310: std_logic; attribute dont_touch of G16310: signal is true;
	signal G16311: std_logic; attribute dont_touch of G16311: signal is true;
	signal G16312: std_logic; attribute dont_touch of G16312: signal is true;
	signal G16313: std_logic; attribute dont_touch of G16313: signal is true;
	signal G16321: std_logic; attribute dont_touch of G16321: signal is true;
	signal G16322: std_logic; attribute dont_touch of G16322: signal is true;
	signal G16323: std_logic; attribute dont_touch of G16323: signal is true;
	signal G16324: std_logic; attribute dont_touch of G16324: signal is true;
	signal G16325: std_logic; attribute dont_touch of G16325: signal is true;
	signal G16335: std_logic; attribute dont_touch of G16335: signal is true;
	signal G16336: std_logic; attribute dont_touch of G16336: signal is true;
	signal G16337: std_logic; attribute dont_touch of G16337: signal is true;
	signal G16341: std_logic; attribute dont_touch of G16341: signal is true;
	signal G16342: std_logic; attribute dont_touch of G16342: signal is true;
	signal G16343: std_logic; attribute dont_touch of G16343: signal is true;
	signal G16344: std_logic; attribute dont_touch of G16344: signal is true;
	signal G16345: std_logic; attribute dont_touch of G16345: signal is true;
	signal G16346: std_logic; attribute dont_touch of G16346: signal is true;
	signal G16347: std_logic; attribute dont_touch of G16347: signal is true;
	signal G16348: std_logic; attribute dont_touch of G16348: signal is true;
	signal G16349: std_logic; attribute dont_touch of G16349: signal is true;
	signal G16350: std_logic; attribute dont_touch of G16350: signal is true;
	signal G16351: std_logic; attribute dont_touch of G16351: signal is true;
	signal G16356: std_logic; attribute dont_touch of G16356: signal is true;
	signal G16357: std_logic; attribute dont_touch of G16357: signal is true;
	signal G16358: std_logic; attribute dont_touch of G16358: signal is true;
	signal G16359: std_logic; attribute dont_touch of G16359: signal is true;
	signal G16360: std_logic; attribute dont_touch of G16360: signal is true;
	signal G16367: std_logic; attribute dont_touch of G16367: signal is true;
	signal G16368: std_logic; attribute dont_touch of G16368: signal is true;
	signal G16369: std_logic; attribute dont_touch of G16369: signal is true;
	signal G16370: std_logic; attribute dont_touch of G16370: signal is true;
	signal G16371: std_logic; attribute dont_touch of G16371: signal is true;
	signal G16379: std_logic; attribute dont_touch of G16379: signal is true;
	signal G16380: std_logic; attribute dont_touch of G16380: signal is true;
	signal G16381: std_logic; attribute dont_touch of G16381: signal is true;
	signal G16382: std_logic; attribute dont_touch of G16382: signal is true;
	signal G16383: std_logic; attribute dont_touch of G16383: signal is true;
	signal G16384: std_logic; attribute dont_touch of G16384: signal is true;
	signal G16385: std_logic; attribute dont_touch of G16385: signal is true;
	signal G16386: std_logic; attribute dont_touch of G16386: signal is true;
	signal G16387: std_logic; attribute dont_touch of G16387: signal is true;
	signal G16388: std_logic; attribute dont_touch of G16388: signal is true;
	signal G16389: std_logic; attribute dont_touch of G16389: signal is true;
	signal G16390: std_logic; attribute dont_touch of G16390: signal is true;
	signal G16391: std_logic; attribute dont_touch of G16391: signal is true;
	signal G16392: std_logic; attribute dont_touch of G16392: signal is true;
	signal G16393: std_logic; attribute dont_touch of G16393: signal is true;
	signal G16394: std_logic; attribute dont_touch of G16394: signal is true;
	signal G16395: std_logic; attribute dont_touch of G16395: signal is true;
	signal G16400: std_logic; attribute dont_touch of G16400: signal is true;
	signal G16401: std_logic; attribute dont_touch of G16401: signal is true;
	signal G16402: std_logic; attribute dont_touch of G16402: signal is true;
	signal G16403: std_logic; attribute dont_touch of G16403: signal is true;
	signal G16404: std_logic; attribute dont_touch of G16404: signal is true;
	signal G16411: std_logic; attribute dont_touch of G16411: signal is true;
	signal G16412: std_logic; attribute dont_touch of G16412: signal is true;
	signal G16413: std_logic; attribute dont_touch of G16413: signal is true;
	signal G16414: std_logic; attribute dont_touch of G16414: signal is true;
	signal G16415: std_logic; attribute dont_touch of G16415: signal is true;
	signal G16416: std_logic; attribute dont_touch of G16416: signal is true;
	signal G16417: std_logic; attribute dont_touch of G16417: signal is true;
	signal G16418: std_logic; attribute dont_touch of G16418: signal is true;
	signal G16419: std_logic; attribute dont_touch of G16419: signal is true;
	signal G16420: std_logic; attribute dont_touch of G16420: signal is true;
	signal G16421: std_logic; attribute dont_touch of G16421: signal is true;
	signal G16422: std_logic; attribute dont_touch of G16422: signal is true;
	signal G16423: std_logic; attribute dont_touch of G16423: signal is true;
	signal G16424: std_logic; attribute dont_touch of G16424: signal is true;
	signal G16425: std_logic; attribute dont_touch of G16425: signal is true;
	signal G16426: std_logic; attribute dont_touch of G16426: signal is true;
	signal G16427: std_logic; attribute dont_touch of G16427: signal is true;
	signal G16428: std_logic; attribute dont_touch of G16428: signal is true;
	signal G16429: std_logic; attribute dont_touch of G16429: signal is true;
	signal G16430: std_logic; attribute dont_touch of G16430: signal is true;
	signal G16431: std_logic; attribute dont_touch of G16431: signal is true;
	signal G16432: std_logic; attribute dont_touch of G16432: signal is true;
	signal G16433: std_logic; attribute dont_touch of G16433: signal is true;
	signal G16438: std_logic; attribute dont_touch of G16438: signal is true;
	signal G16439: std_logic; attribute dont_touch of G16439: signal is true;
	signal G16442: std_logic; attribute dont_touch of G16442: signal is true;
	signal G16443: std_logic; attribute dont_touch of G16443: signal is true;
	signal G16444: std_logic; attribute dont_touch of G16444: signal is true;
	signal G16445: std_logic; attribute dont_touch of G16445: signal is true;
	signal G16446: std_logic; attribute dont_touch of G16446: signal is true;
	signal G16447: std_logic; attribute dont_touch of G16447: signal is true;
	signal G16448: std_logic; attribute dont_touch of G16448: signal is true;
	signal G16449: std_logic; attribute dont_touch of G16449: signal is true;
	signal G16450: std_logic; attribute dont_touch of G16450: signal is true;
	signal G16451: std_logic; attribute dont_touch of G16451: signal is true;
	signal G16452: std_logic; attribute dont_touch of G16452: signal is true;
	signal G16453: std_logic; attribute dont_touch of G16453: signal is true;
	signal G16454: std_logic; attribute dont_touch of G16454: signal is true;
	signal G16455: std_logic; attribute dont_touch of G16455: signal is true;
	signal G16456: std_logic; attribute dont_touch of G16456: signal is true;
	signal G16457: std_logic; attribute dont_touch of G16457: signal is true;
	signal G16458: std_logic; attribute dont_touch of G16458: signal is true;
	signal G16459: std_logic; attribute dont_touch of G16459: signal is true;
	signal G16460: std_logic; attribute dont_touch of G16460: signal is true;
	signal G16461: std_logic; attribute dont_touch of G16461: signal is true;
	signal G16462: std_logic; attribute dont_touch of G16462: signal is true;
	signal G16463: std_logic; attribute dont_touch of G16463: signal is true;
	signal G16466: std_logic; attribute dont_touch of G16466: signal is true;
	signal G16467: std_logic; attribute dont_touch of G16467: signal is true;
	signal G16468: std_logic; attribute dont_touch of G16468: signal is true;
	signal G16469: std_logic; attribute dont_touch of G16469: signal is true;
	signal G16470: std_logic; attribute dont_touch of G16470: signal is true;
	signal G16471: std_logic; attribute dont_touch of G16471: signal is true;
	signal G16472: std_logic; attribute dont_touch of G16472: signal is true;
	signal G16473: std_logic; attribute dont_touch of G16473: signal is true;
	signal G16474: std_logic; attribute dont_touch of G16474: signal is true;
	signal G16475: std_logic; attribute dont_touch of G16475: signal is true;
	signal G16476: std_logic; attribute dont_touch of G16476: signal is true;
	signal G16477: std_logic; attribute dont_touch of G16477: signal is true;
	signal G16478: std_logic; attribute dont_touch of G16478: signal is true;
	signal G16479: std_logic; attribute dont_touch of G16479: signal is true;
	signal G16480: std_logic; attribute dont_touch of G16480: signal is true;
	signal G16481: std_logic; attribute dont_touch of G16481: signal is true;
	signal G16482: std_logic; attribute dont_touch of G16482: signal is true;
	signal G16483: std_logic; attribute dont_touch of G16483: signal is true;
	signal G16484: std_logic; attribute dont_touch of G16484: signal is true;
	signal G16485: std_logic; attribute dont_touch of G16485: signal is true;
	signal G16486: std_logic; attribute dont_touch of G16486: signal is true;
	signal G16487: std_logic; attribute dont_touch of G16487: signal is true;
	signal G16488: std_logic; attribute dont_touch of G16488: signal is true;
	signal G16489: std_logic; attribute dont_touch of G16489: signal is true;
	signal G16490: std_logic; attribute dont_touch of G16490: signal is true;
	signal G16491: std_logic; attribute dont_touch of G16491: signal is true;
	signal G16492: std_logic; attribute dont_touch of G16492: signal is true;
	signal G16493: std_logic; attribute dont_touch of G16493: signal is true;
	signal G16494: std_logic; attribute dont_touch of G16494: signal is true;
	signal G16495: std_logic; attribute dont_touch of G16495: signal is true;
	signal G16497: std_logic; attribute dont_touch of G16497: signal is true;
	signal G16498: std_logic; attribute dont_touch of G16498: signal is true;
	signal G16501: std_logic; attribute dont_touch of G16501: signal is true;
	signal G16505: std_logic; attribute dont_touch of G16505: signal is true;
	signal G16506: std_logic; attribute dont_touch of G16506: signal is true;
	signal G16507: std_logic; attribute dont_touch of G16507: signal is true;
	signal G16513: std_logic; attribute dont_touch of G16513: signal is true;
	signal G16514: std_logic; attribute dont_touch of G16514: signal is true;
	signal G16515: std_logic; attribute dont_touch of G16515: signal is true;
	signal G16520: std_logic; attribute dont_touch of G16520: signal is true;
	signal G16523: std_logic; attribute dont_touch of G16523: signal is true;
	signal G16527: std_logic; attribute dont_touch of G16527: signal is true;
	signal G16528: std_logic; attribute dont_touch of G16528: signal is true;
	signal G16529: std_logic; attribute dont_touch of G16529: signal is true;
	signal G16535: std_logic; attribute dont_touch of G16535: signal is true;
	signal G16536: std_logic; attribute dont_touch of G16536: signal is true;
	signal G16539: std_logic; attribute dont_touch of G16539: signal is true;
	signal G16540: std_logic; attribute dont_touch of G16540: signal is true;
	signal G16543: std_logic; attribute dont_touch of G16543: signal is true;
	signal G16546: std_logic; attribute dont_touch of G16546: signal is true;
	signal G16551: std_logic; attribute dont_touch of G16551: signal is true;
	signal G16554: std_logic; attribute dont_touch of G16554: signal is true;
	signal G16558: std_logic; attribute dont_touch of G16558: signal is true;
	signal G16559: std_logic; attribute dont_touch of G16559: signal is true;
	signal G16560: std_logic; attribute dont_touch of G16560: signal is true;
	signal G16566: std_logic; attribute dont_touch of G16566: signal is true;
	signal G16567: std_logic; attribute dont_touch of G16567: signal is true;
	signal G16570: std_logic; attribute dont_touch of G16570: signal is true;
	signal G16571: std_logic; attribute dont_touch of G16571: signal is true;
	signal G16572: std_logic; attribute dont_touch of G16572: signal is true;
	signal G16575: std_logic; attribute dont_touch of G16575: signal is true;
	signal G16578: std_logic; attribute dont_touch of G16578: signal is true;
	signal G16583: std_logic; attribute dont_touch of G16583: signal is true;
	signal G16586: std_logic; attribute dont_touch of G16586: signal is true;
	signal G16590: std_logic; attribute dont_touch of G16590: signal is true;
	signal G16591: std_logic; attribute dont_touch of G16591: signal is true;
	signal G16594: std_logic; attribute dont_touch of G16594: signal is true;
	signal G16595: std_logic; attribute dont_touch of G16595: signal is true;
	signal G16596: std_logic; attribute dont_touch of G16596: signal is true;
	signal G16599: std_logic; attribute dont_touch of G16599: signal is true;
	signal G16602: std_logic; attribute dont_touch of G16602: signal is true;
	signal G16607: std_logic; attribute dont_touch of G16607: signal is true;
	signal G16608: std_logic; attribute dont_touch of G16608: signal is true;
	signal G16611: std_logic; attribute dont_touch of G16611: signal is true;
	signal G16614: std_logic; attribute dont_touch of G16614: signal is true;
	signal G16615: std_logic; attribute dont_touch of G16615: signal is true;
	signal G16616: std_logic; attribute dont_touch of G16616: signal is true;
	signal G16619: std_logic; attribute dont_touch of G16619: signal is true;
	signal G16622: std_logic; attribute dont_touch of G16622: signal is true;
	signal G16625: std_logic; attribute dont_touch of G16625: signal is true;
	signal G16626: std_logic; attribute dont_touch of G16626: signal is true;
	signal G16629: std_logic; attribute dont_touch of G16629: signal is true;
	signal G16632: std_logic; attribute dont_touch of G16632: signal is true;
	signal G16633: std_logic; attribute dont_touch of G16633: signal is true;
	signal G16636: std_logic; attribute dont_touch of G16636: signal is true;
	signal G16639: std_logic; attribute dont_touch of G16639: signal is true;
	signal G16640: std_logic; attribute dont_touch of G16640: signal is true;
	signal G16643: std_logic; attribute dont_touch of G16643: signal is true;
	signal G16644: std_logic; attribute dont_touch of G16644: signal is true;
	signal G16647: std_logic; attribute dont_touch of G16647: signal is true;
	signal G16650: std_logic; attribute dont_touch of G16650: signal is true;
	signal G16651: std_logic; attribute dont_touch of G16651: signal is true;
	signal G16654: std_logic; attribute dont_touch of G16654: signal is true;
	signal G16655: std_logic; attribute dont_touch of G16655: signal is true;
	signal G16656: std_logic; attribute dont_touch of G16656: signal is true;
	signal G16659: std_logic; attribute dont_touch of G16659: signal is true;
	signal G16662: std_logic; attribute dont_touch of G16662: signal is true;
	signal G16665: std_logic; attribute dont_touch of G16665: signal is true;
	signal G16671: std_logic; attribute dont_touch of G16671: signal is true;
	signal G16672: std_logic; attribute dont_touch of G16672: signal is true;
	signal G16673: std_logic; attribute dont_touch of G16673: signal is true;
	signal G16676: std_logic; attribute dont_touch of G16676: signal is true;
	signal G16679: std_logic; attribute dont_touch of G16679: signal is true;
	signal G16682: std_logic; attribute dont_touch of G16682: signal is true;
	signal G16686: std_logic; attribute dont_touch of G16686: signal is true;
	signal G16692: std_logic; attribute dont_touch of G16692: signal is true;
	signal G16693: std_logic; attribute dont_touch of G16693: signal is true;
	signal G16694: std_logic; attribute dont_touch of G16694: signal is true;
	signal G16697: std_logic; attribute dont_touch of G16697: signal is true;
	signal G16702: std_logic; attribute dont_touch of G16702: signal is true;
	signal G16705: std_logic; attribute dont_touch of G16705: signal is true;
	signal G16708: std_logic; attribute dont_touch of G16708: signal is true;
	signal G16712: std_logic; attribute dont_touch of G16712: signal is true;
	signal G16718: std_logic; attribute dont_touch of G16718: signal is true;
	signal G16719: std_logic; attribute dont_touch of G16719: signal is true;
	signal G16722: std_logic; attribute dont_touch of G16722: signal is true;
	signal G16725: std_logic; attribute dont_touch of G16725: signal is true;
	signal G16728: std_logic; attribute dont_touch of G16728: signal is true;
	signal G16733: std_logic; attribute dont_touch of G16733: signal is true;
	signal G16736: std_logic; attribute dont_touch of G16736: signal is true;
	signal G16739: std_logic; attribute dont_touch of G16739: signal is true;
	signal G16743: std_logic; attribute dont_touch of G16743: signal is true;
	signal G16749: std_logic; attribute dont_touch of G16749: signal is true;
	signal G16758: std_logic; attribute dont_touch of G16758: signal is true;
	signal G16761: std_logic; attribute dont_touch of G16761: signal is true;
	signal G16764: std_logic; attribute dont_touch of G16764: signal is true;
	signal G16767: std_logic; attribute dont_touch of G16767: signal is true;
	signal G16770: std_logic; attribute dont_touch of G16770: signal is true;
	signal G16775: std_logic; attribute dont_touch of G16775: signal is true;
	signal G16778: std_logic; attribute dont_touch of G16778: signal is true;
	signal G16781: std_logic; attribute dont_touch of G16781: signal is true;
	signal G16785: std_logic; attribute dont_touch of G16785: signal is true;
	signal G16788: std_logic; attribute dont_touch of G16788: signal is true;
	signal G16791: std_logic; attribute dont_touch of G16791: signal is true;
	signal G16794: std_logic; attribute dont_touch of G16794: signal is true;
	signal G16797: std_logic; attribute dont_touch of G16797: signal is true;
	signal G16802: std_logic; attribute dont_touch of G16802: signal is true;
	signal G16803: std_logic; attribute dont_touch of G16803: signal is true;
	signal G16804: std_logic; attribute dont_touch of G16804: signal is true;
	signal G16809: std_logic; attribute dont_touch of G16809: signal is true;
	signal G16813: std_logic; attribute dont_touch of G16813: signal is true;
	signal G16814: std_logic; attribute dont_touch of G16814: signal is true;
	signal G16817: std_logic; attribute dont_touch of G16817: signal is true;
	signal G16820: std_logic; attribute dont_touch of G16820: signal is true;
	signal G16823: std_logic; attribute dont_touch of G16823: signal is true;
	signal G16824: std_logic; attribute dont_touch of G16824: signal is true;
	signal G16825: std_logic; attribute dont_touch of G16825: signal is true;
	signal G16829: std_logic; attribute dont_touch of G16829: signal is true;
	signal G16830: std_logic; attribute dont_touch of G16830: signal is true;
	signal G16831: std_logic; attribute dont_touch of G16831: signal is true;
	signal G16832: std_logic; attribute dont_touch of G16832: signal is true;
	signal G16835: std_logic; attribute dont_touch of G16835: signal is true;
	signal G16836: std_logic; attribute dont_touch of G16836: signal is true;
	signal G16840: std_logic; attribute dont_touch of G16840: signal is true;
	signal G16841: std_logic; attribute dont_touch of G16841: signal is true;
	signal G16842: std_logic; attribute dont_touch of G16842: signal is true;
	signal G16843: std_logic; attribute dont_touch of G16843: signal is true;
	signal G16844: std_logic; attribute dont_touch of G16844: signal is true;
	signal G16845: std_logic; attribute dont_touch of G16845: signal is true;
	signal G16846: std_logic; attribute dont_touch of G16846: signal is true;
	signal G16847: std_logic; attribute dont_touch of G16847: signal is true;
	signal G16848: std_logic; attribute dont_touch of G16848: signal is true;
	signal G16849: std_logic; attribute dont_touch of G16849: signal is true;
	signal G16850: std_logic; attribute dont_touch of G16850: signal is true;
	signal G16851: std_logic; attribute dont_touch of G16851: signal is true;
	signal G16852: std_logic; attribute dont_touch of G16852: signal is true;
	signal G16853: std_logic; attribute dont_touch of G16853: signal is true;
	signal G16854: std_logic; attribute dont_touch of G16854: signal is true;
	signal G16855: std_logic; attribute dont_touch of G16855: signal is true;
	signal G16856: std_logic; attribute dont_touch of G16856: signal is true;
	signal G16857: std_logic; attribute dont_touch of G16857: signal is true;
	signal G16858: std_logic; attribute dont_touch of G16858: signal is true;
	signal G16859: std_logic; attribute dont_touch of G16859: signal is true;
	signal G16860: std_logic; attribute dont_touch of G16860: signal is true;
	signal G16861: std_logic; attribute dont_touch of G16861: signal is true;
	signal G16862: std_logic; attribute dont_touch of G16862: signal is true;
	signal G16863: std_logic; attribute dont_touch of G16863: signal is true;
	signal G16864: std_logic; attribute dont_touch of G16864: signal is true;
	signal G16865: std_logic; attribute dont_touch of G16865: signal is true;
	signal G16866: std_logic; attribute dont_touch of G16866: signal is true;
	signal G16867: std_logic; attribute dont_touch of G16867: signal is true;
	signal G16877: std_logic; attribute dont_touch of G16877: signal is true;
	signal G16878: std_logic; attribute dont_touch of G16878: signal is true;
	signal G16879: std_logic; attribute dont_touch of G16879: signal is true;
	signal G16880: std_logic; attribute dont_touch of G16880: signal is true;
	signal G16881: std_logic; attribute dont_touch of G16881: signal is true;
	signal G16884: std_logic; attribute dont_touch of G16884: signal is true;
	signal G16894: std_logic; attribute dont_touch of G16894: signal is true;
	signal G16895: std_logic; attribute dont_touch of G16895: signal is true;
	signal G16905: std_logic; attribute dont_touch of G16905: signal is true;
	signal G16906: std_logic; attribute dont_touch of G16906: signal is true;
	signal G16907: std_logic; attribute dont_touch of G16907: signal is true;
	signal G16908: std_logic; attribute dont_touch of G16908: signal is true;
	signal G16909: std_logic; attribute dont_touch of G16909: signal is true;
	signal G16910: std_logic; attribute dont_touch of G16910: signal is true;
	signal G16913: std_logic; attribute dont_touch of G16913: signal is true;
	signal G16923: std_logic; attribute dont_touch of G16923: signal is true;
	signal G16924: std_logic; attribute dont_touch of G16924: signal is true;
	signal G16934: std_logic; attribute dont_touch of G16934: signal is true;
	signal G16935: std_logic; attribute dont_touch of G16935: signal is true;
	signal G16938: std_logic; attribute dont_touch of G16938: signal is true;
	signal G16939: std_logic; attribute dont_touch of G16939: signal is true;
	signal G16940: std_logic; attribute dont_touch of G16940: signal is true;
	signal G16943: std_logic; attribute dont_touch of G16943: signal is true;
	signal G16953: std_logic; attribute dont_touch of G16953: signal is true;
	signal G16954: std_logic; attribute dont_touch of G16954: signal is true;
	signal G16964: std_logic; attribute dont_touch of G16964: signal is true;
	signal G16965: std_logic; attribute dont_touch of G16965: signal is true;
	signal G16966: std_logic; attribute dont_touch of G16966: signal is true;
	signal G16967: std_logic; attribute dont_touch of G16967: signal is true;
	signal G16968: std_logic; attribute dont_touch of G16968: signal is true;
	signal G16969: std_logic; attribute dont_touch of G16969: signal is true;
	signal G16970: std_logic; attribute dont_touch of G16970: signal is true;
	signal G16971: std_logic; attribute dont_touch of G16971: signal is true;
	signal G16974: std_logic; attribute dont_touch of G16974: signal is true;
	signal G16984: std_logic; attribute dont_touch of G16984: signal is true;
	signal G16985: std_logic; attribute dont_touch of G16985: signal is true;
	signal G16986: std_logic; attribute dont_touch of G16986: signal is true;
	signal G16987: std_logic; attribute dont_touch of G16987: signal is true;
	signal G16988: std_logic; attribute dont_touch of G16988: signal is true;
	signal G16989: std_logic; attribute dont_touch of G16989: signal is true;
	signal G16990: std_logic; attribute dont_touch of G16990: signal is true;
	signal G16991: std_logic; attribute dont_touch of G16991: signal is true;
	signal G16992: std_logic; attribute dont_touch of G16992: signal is true;
	signal G16993: std_logic; attribute dont_touch of G16993: signal is true;
	signal G16994: std_logic; attribute dont_touch of G16994: signal is true;
	signal G16995: std_logic; attribute dont_touch of G16995: signal is true;
	signal G16996: std_logic; attribute dont_touch of G16996: signal is true;
	signal G16997: std_logic; attribute dont_touch of G16997: signal is true;
	signal G16998: std_logic; attribute dont_touch of G16998: signal is true;
	signal G16999: std_logic; attribute dont_touch of G16999: signal is true;
	signal G17000: std_logic; attribute dont_touch of G17000: signal is true;
	signal G17001: std_logic; attribute dont_touch of G17001: signal is true;
	signal G17012: std_logic; attribute dont_touch of G17012: signal is true;
	signal G17015: std_logic; attribute dont_touch of G17015: signal is true;
	signal G17016: std_logic; attribute dont_touch of G17016: signal is true;
	signal G17017: std_logic; attribute dont_touch of G17017: signal is true;
	signal G17018: std_logic; attribute dont_touch of G17018: signal is true;
	signal G17019: std_logic; attribute dont_touch of G17019: signal is true;
	signal G17020: std_logic; attribute dont_touch of G17020: signal is true;
	signal G17021: std_logic; attribute dont_touch of G17021: signal is true;
	signal G17022: std_logic; attribute dont_touch of G17022: signal is true;
	signal G17023: std_logic; attribute dont_touch of G17023: signal is true;
	signal G17024: std_logic; attribute dont_touch of G17024: signal is true;
	signal G17025: std_logic; attribute dont_touch of G17025: signal is true;
	signal G17028: std_logic; attribute dont_touch of G17028: signal is true;
	signal G17029: std_logic; attribute dont_touch of G17029: signal is true;
	signal G17030: std_logic; attribute dont_touch of G17030: signal is true;
	signal G17031: std_logic; attribute dont_touch of G17031: signal is true;
	signal G17042: std_logic; attribute dont_touch of G17042: signal is true;
	signal G17045: std_logic; attribute dont_touch of G17045: signal is true;
	signal G17046: std_logic; attribute dont_touch of G17046: signal is true;
	signal G17047: std_logic; attribute dont_touch of G17047: signal is true;
	signal G17048: std_logic; attribute dont_touch of G17048: signal is true;
	signal G17049: std_logic; attribute dont_touch of G17049: signal is true;
	signal G17050: std_logic; attribute dont_touch of G17050: signal is true;
	signal G17051: std_logic; attribute dont_touch of G17051: signal is true;
	signal G17055: std_logic; attribute dont_touch of G17055: signal is true;
	signal G17056: std_logic; attribute dont_touch of G17056: signal is true;
	signal G17057: std_logic; attribute dont_touch of G17057: signal is true;
	signal G17058: std_logic; attribute dont_touch of G17058: signal is true;
	signal G17059: std_logic; attribute dont_touch of G17059: signal is true;
	signal G17062: std_logic; attribute dont_touch of G17062: signal is true;
	signal G17063: std_logic; attribute dont_touch of G17063: signal is true;
	signal G17064: std_logic; attribute dont_touch of G17064: signal is true;
	signal G17065: std_logic; attribute dont_touch of G17065: signal is true;
	signal G17076: std_logic; attribute dont_touch of G17076: signal is true;
	signal G17079: std_logic; attribute dont_touch of G17079: signal is true;
	signal G17080: std_logic; attribute dont_touch of G17080: signal is true;
	signal G17081: std_logic; attribute dont_touch of G17081: signal is true;
	signal G17082: std_logic; attribute dont_touch of G17082: signal is true;
	signal G17083: std_logic; attribute dont_touch of G17083: signal is true;
	signal G17084: std_logic; attribute dont_touch of G17084: signal is true;
	signal G17085: std_logic; attribute dont_touch of G17085: signal is true;
	signal G17086: std_logic; attribute dont_touch of G17086: signal is true;
	signal G17090: std_logic; attribute dont_touch of G17090: signal is true;
	signal G17091: std_logic; attribute dont_touch of G17091: signal is true;
	signal G17092: std_logic; attribute dont_touch of G17092: signal is true;
	signal G17093: std_logic; attribute dont_touch of G17093: signal is true;
	signal G17094: std_logic; attribute dont_touch of G17094: signal is true;
	signal G17097: std_logic; attribute dont_touch of G17097: signal is true;
	signal G17098: std_logic; attribute dont_touch of G17098: signal is true;
	signal G17099: std_logic; attribute dont_touch of G17099: signal is true;
	signal G17100: std_logic; attribute dont_touch of G17100: signal is true;
	signal G17111: std_logic; attribute dont_touch of G17111: signal is true;
	signal G17114: std_logic; attribute dont_touch of G17114: signal is true;
	signal G17115: std_logic; attribute dont_touch of G17115: signal is true;
	signal G17116: std_logic; attribute dont_touch of G17116: signal is true;
	signal G17117: std_logic; attribute dont_touch of G17117: signal is true;
	signal G17118: std_logic; attribute dont_touch of G17118: signal is true;
	signal G17121: std_logic; attribute dont_touch of G17121: signal is true;
	signal G17122: std_logic; attribute dont_touch of G17122: signal is true;
	signal G17123: std_logic; attribute dont_touch of G17123: signal is true;
	signal G17124: std_logic; attribute dont_touch of G17124: signal is true;
	signal G17128: std_logic; attribute dont_touch of G17128: signal is true;
	signal G17129: std_logic; attribute dont_touch of G17129: signal is true;
	signal G17130: std_logic; attribute dont_touch of G17130: signal is true;
	signal G17131: std_logic; attribute dont_touch of G17131: signal is true;
	signal G17132: std_logic; attribute dont_touch of G17132: signal is true;
	signal G17135: std_logic; attribute dont_touch of G17135: signal is true;
	signal G17136: std_logic; attribute dont_touch of G17136: signal is true;
	signal G17137: std_logic; attribute dont_touch of G17137: signal is true;
	signal G17138: std_logic; attribute dont_touch of G17138: signal is true;
	signal G17139: std_logic; attribute dont_touch of G17139: signal is true;
	signal G17142: std_logic; attribute dont_touch of G17142: signal is true;
	signal G17143: std_logic; attribute dont_touch of G17143: signal is true;
	signal G17144: std_logic; attribute dont_touch of G17144: signal is true;
	signal G17145: std_logic; attribute dont_touch of G17145: signal is true;
	signal G17148: std_logic; attribute dont_touch of G17148: signal is true;
	signal G17149: std_logic; attribute dont_touch of G17149: signal is true;
	signal G17150: std_logic; attribute dont_touch of G17150: signal is true;
	signal G17151: std_logic; attribute dont_touch of G17151: signal is true;
	signal G17155: std_logic; attribute dont_touch of G17155: signal is true;
	signal G17156: std_logic; attribute dont_touch of G17156: signal is true;
	signal G17157: std_logic; attribute dont_touch of G17157: signal is true;
	signal G17158: std_logic; attribute dont_touch of G17158: signal is true;
	signal G17159: std_logic; attribute dont_touch of G17159: signal is true;
	signal G17160: std_logic; attribute dont_touch of G17160: signal is true;
	signal G17161: std_logic; attribute dont_touch of G17161: signal is true;
	signal G17162: std_logic; attribute dont_touch of G17162: signal is true;
	signal G17165: std_logic; attribute dont_touch of G17165: signal is true;
	signal G17166: std_logic; attribute dont_touch of G17166: signal is true;
	signal G17167: std_logic; attribute dont_touch of G17167: signal is true;
	signal G17168: std_logic; attribute dont_touch of G17168: signal is true;
	signal G17171: std_logic; attribute dont_touch of G17171: signal is true;
	signal G17172: std_logic; attribute dont_touch of G17172: signal is true;
	signal G17173: std_logic; attribute dont_touch of G17173: signal is true;
	signal G17174: std_logic; attribute dont_touch of G17174: signal is true;
	signal G17175: std_logic; attribute dont_touch of G17175: signal is true;
	signal G17176: std_logic; attribute dont_touch of G17176: signal is true;
	signal G17177: std_logic; attribute dont_touch of G17177: signal is true;
	signal G17180: std_logic; attribute dont_touch of G17180: signal is true;
	signal G17181: std_logic; attribute dont_touch of G17181: signal is true;
	signal G17182: std_logic; attribute dont_touch of G17182: signal is true;
	signal G17183: std_logic; attribute dont_touch of G17183: signal is true;
	signal G17186: std_logic; attribute dont_touch of G17186: signal is true;
	signal G17189: std_logic; attribute dont_touch of G17189: signal is true;
	signal G17190: std_logic; attribute dont_touch of G17190: signal is true;
	signal G17191: std_logic; attribute dont_touch of G17191: signal is true;
	signal G17192: std_logic; attribute dont_touch of G17192: signal is true;
	signal G17193: std_logic; attribute dont_touch of G17193: signal is true;
	signal G17194: std_logic; attribute dont_touch of G17194: signal is true;
	signal G17197: std_logic; attribute dont_touch of G17197: signal is true;
	signal G17200: std_logic; attribute dont_touch of G17200: signal is true;
	signal G17201: std_logic; attribute dont_touch of G17201: signal is true;
	signal G17202: std_logic; attribute dont_touch of G17202: signal is true;
	signal G17203: std_logic; attribute dont_touch of G17203: signal is true;
	signal G17204: std_logic; attribute dont_touch of G17204: signal is true;
	signal G17207: std_logic; attribute dont_touch of G17207: signal is true;
	signal G17208: std_logic; attribute dont_touch of G17208: signal is true;
	signal G17209: std_logic; attribute dont_touch of G17209: signal is true;
	signal G17212: std_logic; attribute dont_touch of G17212: signal is true;
	signal G17213: std_logic; attribute dont_touch of G17213: signal is true;
	signal G17214: std_logic; attribute dont_touch of G17214: signal is true;
	signal G17215: std_logic; attribute dont_touch of G17215: signal is true;
	signal G17216: std_logic; attribute dont_touch of G17216: signal is true;
	signal G17217: std_logic; attribute dont_touch of G17217: signal is true;
	signal G17218: std_logic; attribute dont_touch of G17218: signal is true;
	signal G17219: std_logic; attribute dont_touch of G17219: signal is true;
	signal G17220: std_logic; attribute dont_touch of G17220: signal is true;
	signal G17221: std_logic; attribute dont_touch of G17221: signal is true;
	signal G17222: std_logic; attribute dont_touch of G17222: signal is true;
	signal G17223: std_logic; attribute dont_touch of G17223: signal is true;
	signal G17224: std_logic; attribute dont_touch of G17224: signal is true;
	signal G17225: std_logic; attribute dont_touch of G17225: signal is true;
	signal G17226: std_logic; attribute dont_touch of G17226: signal is true;
	signal G17227: std_logic; attribute dont_touch of G17227: signal is true;
	signal G17228: std_logic; attribute dont_touch of G17228: signal is true;
	signal G17229: std_logic; attribute dont_touch of G17229: signal is true;
	signal G17230: std_logic; attribute dont_touch of G17230: signal is true;
	signal G17233: std_logic; attribute dont_touch of G17233: signal is true;
	signal G17234: std_logic; attribute dont_touch of G17234: signal is true;
	signal G17235: std_logic; attribute dont_touch of G17235: signal is true;
	signal G17236: std_logic; attribute dont_touch of G17236: signal is true;
	signal G17237: std_logic; attribute dont_touch of G17237: signal is true;
	signal G17240: std_logic; attribute dont_touch of G17240: signal is true;
	signal G17243: std_logic; attribute dont_touch of G17243: signal is true;
	signal G17246: std_logic; attribute dont_touch of G17246: signal is true;
	signal G17247: std_logic; attribute dont_touch of G17247: signal is true;
	signal G17248: std_logic; attribute dont_touch of G17248: signal is true;
	signal G17249: std_logic; attribute dont_touch of G17249: signal is true;
	signal G17252: std_logic; attribute dont_touch of G17252: signal is true;
	signal G17255: std_logic; attribute dont_touch of G17255: signal is true;
	signal G17258: std_logic; attribute dont_touch of G17258: signal is true;
	signal G17259: std_logic; attribute dont_touch of G17259: signal is true;
	signal G17262: std_logic; attribute dont_touch of G17262: signal is true;
	signal G17265: std_logic; attribute dont_touch of G17265: signal is true;
	signal G17268: std_logic; attribute dont_touch of G17268: signal is true;
	signal G17269: std_logic; attribute dont_touch of G17269: signal is true;
	signal G17270: std_logic; attribute dont_touch of G17270: signal is true;
	signal G17271: std_logic; attribute dont_touch of G17271: signal is true;
	signal G17272: std_logic; attribute dont_touch of G17272: signal is true;
	signal G17275: std_logic; attribute dont_touch of G17275: signal is true;
	signal G17278: std_logic; attribute dont_touch of G17278: signal is true;
	signal G17281: std_logic; attribute dont_touch of G17281: signal is true;
	signal G17282: std_logic; attribute dont_touch of G17282: signal is true;
	signal G17285: std_logic; attribute dont_touch of G17285: signal is true;
	signal G17288: std_logic; attribute dont_touch of G17288: signal is true;
	signal G17291: std_logic; attribute dont_touch of G17291: signal is true;
	signal G17294: std_logic; attribute dont_touch of G17294: signal is true;
	signal G17297: std_logic; attribute dont_touch of G17297: signal is true;
	signal G17300: std_logic; attribute dont_touch of G17300: signal is true;
	signal G17301: std_logic; attribute dont_touch of G17301: signal is true;
	signal G17302: std_logic; attribute dont_touch of G17302: signal is true;
	signal G17303: std_logic; attribute dont_touch of G17303: signal is true;
	signal G17304: std_logic; attribute dont_touch of G17304: signal is true;
	signal G17307: std_logic; attribute dont_touch of G17307: signal is true;
	signal G17310: std_logic; attribute dont_touch of G17310: signal is true;
	signal G17313: std_logic; attribute dont_touch of G17313: signal is true;
	signal G17314: std_logic; attribute dont_touch of G17314: signal is true;
	signal G17315: std_logic; attribute dont_touch of G17315: signal is true;
	signal G17318: std_logic; attribute dont_touch of G17318: signal is true;
	signal G17321: std_logic; attribute dont_touch of G17321: signal is true;
	signal G17324: std_logic; attribute dont_touch of G17324: signal is true;
	signal G17327: std_logic; attribute dont_touch of G17327: signal is true;
	signal G17330: std_logic; attribute dont_touch of G17330: signal is true;
	signal G17333: std_logic; attribute dont_touch of G17333: signal is true;
	signal G17336: std_logic; attribute dont_touch of G17336: signal is true;
	signal G17339: std_logic; attribute dont_touch of G17339: signal is true;
	signal G17340: std_logic; attribute dont_touch of G17340: signal is true;
	signal G17341: std_logic; attribute dont_touch of G17341: signal is true;
	signal G17342: std_logic; attribute dont_touch of G17342: signal is true;
	signal G17345: std_logic; attribute dont_touch of G17345: signal is true;
	signal G17348: std_logic; attribute dont_touch of G17348: signal is true;
	signal G17351: std_logic; attribute dont_touch of G17351: signal is true;
	signal G17352: std_logic; attribute dont_touch of G17352: signal is true;
	signal G17353: std_logic; attribute dont_touch of G17353: signal is true;
	signal G17354: std_logic; attribute dont_touch of G17354: signal is true;
	signal G17357: std_logic; attribute dont_touch of G17357: signal is true;
	signal G17360: std_logic; attribute dont_touch of G17360: signal is true;
	signal G17363: std_logic; attribute dont_touch of G17363: signal is true;
	signal G17366: std_logic; attribute dont_touch of G17366: signal is true;
	signal G17369: std_logic; attribute dont_touch of G17369: signal is true;
	signal G17372: std_logic; attribute dont_touch of G17372: signal is true;
	signal G17375: std_logic; attribute dont_touch of G17375: signal is true;
	signal G17378: std_logic; attribute dont_touch of G17378: signal is true;
	signal G17381: std_logic; attribute dont_touch of G17381: signal is true;
	signal G17382: std_logic; attribute dont_touch of G17382: signal is true;
	signal G17383: std_logic; attribute dont_touch of G17383: signal is true;
	signal G17384: std_logic; attribute dont_touch of G17384: signal is true;
	signal G17387: std_logic; attribute dont_touch of G17387: signal is true;
	signal G17390: std_logic; attribute dont_touch of G17390: signal is true;
	signal G17393: std_logic; attribute dont_touch of G17393: signal is true;
	signal G17394: std_logic; attribute dont_touch of G17394: signal is true;
	signal G17395: std_logic; attribute dont_touch of G17395: signal is true;
	signal G17396: std_logic; attribute dont_touch of G17396: signal is true;
	signal G17397: std_logic; attribute dont_touch of G17397: signal is true;
	signal G17398: std_logic; attribute dont_touch of G17398: signal is true;
	signal G17399: std_logic; attribute dont_touch of G17399: signal is true;
	signal G17402: std_logic; attribute dont_touch of G17402: signal is true;
	signal G17405: std_logic; attribute dont_touch of G17405: signal is true;
	signal G17408: std_logic; attribute dont_touch of G17408: signal is true;
	signal G17409: std_logic; attribute dont_touch of G17409: signal is true;
	signal G17410: std_logic; attribute dont_touch of G17410: signal is true;
	signal G17413: std_logic; attribute dont_touch of G17413: signal is true;
	signal G17416: std_logic; attribute dont_touch of G17416: signal is true;
	signal G17419: std_logic; attribute dont_touch of G17419: signal is true;
	signal G17422: std_logic; attribute dont_touch of G17422: signal is true;
	signal G17425: std_logic; attribute dont_touch of G17425: signal is true;
	signal G17428: std_logic; attribute dont_touch of G17428: signal is true;
	signal G17429: std_logic; attribute dont_touch of G17429: signal is true;
	signal G17430: std_logic; attribute dont_touch of G17430: signal is true;
	signal G17433: std_logic; attribute dont_touch of G17433: signal is true;
	signal G17436: std_logic; attribute dont_touch of G17436: signal is true;
	signal G17439: std_logic; attribute dont_touch of G17439: signal is true;
	signal G17442: std_logic; attribute dont_touch of G17442: signal is true;
	signal G17445: std_logic; attribute dont_touch of G17445: signal is true;
	signal G17446: std_logic; attribute dont_touch of G17446: signal is true;
	signal G17447: std_logic; attribute dont_touch of G17447: signal is true;
	signal G17448: std_logic; attribute dont_touch of G17448: signal is true;
	signal G17449: std_logic; attribute dont_touch of G17449: signal is true;
	signal G17450: std_logic; attribute dont_touch of G17450: signal is true;
	signal G17451: std_logic; attribute dont_touch of G17451: signal is true;
	signal G17454: std_logic; attribute dont_touch of G17454: signal is true;
	signal G17457: std_logic; attribute dont_touch of G17457: signal is true;
	signal G17460: std_logic; attribute dont_touch of G17460: signal is true;
	signal G17461: std_logic; attribute dont_touch of G17461: signal is true;
	signal G17462: std_logic; attribute dont_touch of G17462: signal is true;
	signal G17463: std_logic; attribute dont_touch of G17463: signal is true;
	signal G17464: std_logic; attribute dont_touch of G17464: signal is true;
	signal G17465: std_logic; attribute dont_touch of G17465: signal is true;
	signal G17468: std_logic; attribute dont_touch of G17468: signal is true;
	signal G17471: std_logic; attribute dont_touch of G17471: signal is true;
	signal G17474: std_logic; attribute dont_touch of G17474: signal is true;
	signal G17475: std_logic; attribute dont_touch of G17475: signal is true;
	signal G17476: std_logic; attribute dont_touch of G17476: signal is true;
	signal G17479: std_logic; attribute dont_touch of G17479: signal is true;
	signal G17482: std_logic; attribute dont_touch of G17482: signal is true;
	signal G17485: std_logic; attribute dont_touch of G17485: signal is true;
	signal G17486: std_logic; attribute dont_touch of G17486: signal is true;
	signal G17487: std_logic; attribute dont_touch of G17487: signal is true;
	signal G17490: std_logic; attribute dont_touch of G17490: signal is true;
	signal G17493: std_logic; attribute dont_touch of G17493: signal is true;
	signal G17496: std_logic; attribute dont_touch of G17496: signal is true;
	signal G17499: std_logic; attribute dont_touch of G17499: signal is true;
	signal G17500: std_logic; attribute dont_touch of G17500: signal is true;
	signal G17503: std_logic; attribute dont_touch of G17503: signal is true;
	signal G17506: std_logic; attribute dont_touch of G17506: signal is true;
	signal G17507: std_logic; attribute dont_touch of G17507: signal is true;
	signal G17508: std_logic; attribute dont_touch of G17508: signal is true;
	signal G17509: std_logic; attribute dont_touch of G17509: signal is true;
	signal G17510: std_logic; attribute dont_touch of G17510: signal is true;
	signal G17511: std_logic; attribute dont_touch of G17511: signal is true;
	signal G17514: std_logic; attribute dont_touch of G17514: signal is true;
	signal G17517: std_logic; attribute dont_touch of G17517: signal is true;
	signal G17520: std_logic; attribute dont_touch of G17520: signal is true;
	signal G17523: std_logic; attribute dont_touch of G17523: signal is true;
	signal G17526: std_logic; attribute dont_touch of G17526: signal is true;
	signal G17527: std_logic; attribute dont_touch of G17527: signal is true;
	signal G17528: std_logic; attribute dont_touch of G17528: signal is true;
	signal G17529: std_logic; attribute dont_touch of G17529: signal is true;
	signal G17530: std_logic; attribute dont_touch of G17530: signal is true;
	signal G17531: std_logic; attribute dont_touch of G17531: signal is true;
	signal G17534: std_logic; attribute dont_touch of G17534: signal is true;
	signal G17537: std_logic; attribute dont_touch of G17537: signal is true;
	signal G17540: std_logic; attribute dont_touch of G17540: signal is true;
	signal G17541: std_logic; attribute dont_touch of G17541: signal is true;
	signal G17542: std_logic; attribute dont_touch of G17542: signal is true;
	signal G17543: std_logic; attribute dont_touch of G17543: signal is true;
	signal G17544: std_logic; attribute dont_touch of G17544: signal is true;
	signal G17545: std_logic; attribute dont_touch of G17545: signal is true;
	signal G17548: std_logic; attribute dont_touch of G17548: signal is true;
	signal G17551: std_logic; attribute dont_touch of G17551: signal is true;
	signal G17554: std_logic; attribute dont_touch of G17554: signal is true;
	signal G17555: std_logic; attribute dont_touch of G17555: signal is true;
	signal G17556: std_logic; attribute dont_touch of G17556: signal is true;
	signal G17557: std_logic; attribute dont_touch of G17557: signal is true;
	signal G17560: std_logic; attribute dont_touch of G17560: signal is true;
	signal G17563: std_logic; attribute dont_touch of G17563: signal is true;
	signal G17566: std_logic; attribute dont_touch of G17566: signal is true;
	signal G17567: std_logic; attribute dont_touch of G17567: signal is true;
	signal G17570: std_logic; attribute dont_touch of G17570: signal is true;
	signal G17573: std_logic; attribute dont_touch of G17573: signal is true;
	signal G17576: std_logic; attribute dont_touch of G17576: signal is true;
	signal G17577: std_logic; attribute dont_touch of G17577: signal is true;
	signal G17578: std_logic; attribute dont_touch of G17578: signal is true;
	signal G17579: std_logic; attribute dont_touch of G17579: signal is true;
	signal G17582: std_logic; attribute dont_touch of G17582: signal is true;
	signal G17585: std_logic; attribute dont_touch of G17585: signal is true;
	signal G17588: std_logic; attribute dont_touch of G17588: signal is true;
	signal G17591: std_logic; attribute dont_touch of G17591: signal is true;
	signal G17594: std_logic; attribute dont_touch of G17594: signal is true;
	signal G17597: std_logic; attribute dont_touch of G17597: signal is true;
	signal G17598: std_logic; attribute dont_touch of G17598: signal is true;
	signal G17599: std_logic; attribute dont_touch of G17599: signal is true;
	signal G17600: std_logic; attribute dont_touch of G17600: signal is true;
	signal G17601: std_logic; attribute dont_touch of G17601: signal is true;
	signal G17604: std_logic; attribute dont_touch of G17604: signal is true;
	signal G17607: std_logic; attribute dont_touch of G17607: signal is true;
	signal G17610: std_logic; attribute dont_touch of G17610: signal is true;
	signal G17613: std_logic; attribute dont_touch of G17613: signal is true;
	signal G17616: std_logic; attribute dont_touch of G17616: signal is true;
	signal G17617: std_logic; attribute dont_touch of G17617: signal is true;
	signal G17618: std_logic; attribute dont_touch of G17618: signal is true;
	signal G17619: std_logic; attribute dont_touch of G17619: signal is true;
	signal G17620: std_logic; attribute dont_touch of G17620: signal is true;
	signal G17621: std_logic; attribute dont_touch of G17621: signal is true;
	signal G17624: std_logic; attribute dont_touch of G17624: signal is true;
	signal G17627: std_logic; attribute dont_touch of G17627: signal is true;
	signal G17630: std_logic; attribute dont_touch of G17630: signal is true;
	signal G17631: std_logic; attribute dont_touch of G17631: signal is true;
	signal G17632: std_logic; attribute dont_touch of G17632: signal is true;
	signal G17633: std_logic; attribute dont_touch of G17633: signal is true;
	signal G17634: std_logic; attribute dont_touch of G17634: signal is true;
	signal G17635: std_logic; attribute dont_touch of G17635: signal is true;
	signal G17636: std_logic; attribute dont_touch of G17636: signal is true;
	signal G17637: std_logic; attribute dont_touch of G17637: signal is true;
	signal G17640: std_logic; attribute dont_touch of G17640: signal is true;
	signal G17645: std_logic; attribute dont_touch of G17645: signal is true;
	signal G17648: std_logic; attribute dont_touch of G17648: signal is true;
	signal G17649: std_logic; attribute dont_touch of G17649: signal is true;
	signal G17652: std_logic; attribute dont_touch of G17652: signal is true;
	signal G17653: std_logic; attribute dont_touch of G17653: signal is true;
	signal G17654: std_logic; attribute dont_touch of G17654: signal is true;
	signal G17655: std_logic; attribute dont_touch of G17655: signal is true;
	signal G17658: std_logic; attribute dont_touch of G17658: signal is true;
	signal G17661: std_logic; attribute dont_touch of G17661: signal is true;
	signal G17664: std_logic; attribute dont_touch of G17664: signal is true;
	signal G17667: std_logic; attribute dont_touch of G17667: signal is true;
	signal G17670: std_logic; attribute dont_touch of G17670: signal is true;
	signal G17673: std_logic; attribute dont_touch of G17673: signal is true;
	signal G17674: std_logic; attribute dont_touch of G17674: signal is true;
	signal G17675: std_logic; attribute dont_touch of G17675: signal is true;
	signal G17676: std_logic; attribute dont_touch of G17676: signal is true;
	signal G17679: std_logic; attribute dont_touch of G17679: signal is true;
	signal G17682: std_logic; attribute dont_touch of G17682: signal is true;
	signal G17685: std_logic; attribute dont_touch of G17685: signal is true;
	signal G17688: std_logic; attribute dont_touch of G17688: signal is true;
	signal G17691: std_logic; attribute dont_touch of G17691: signal is true;
	signal G17694: std_logic; attribute dont_touch of G17694: signal is true;
	signal G17695: std_logic; attribute dont_touch of G17695: signal is true;
	signal G17696: std_logic; attribute dont_touch of G17696: signal is true;
	signal G17697: std_logic; attribute dont_touch of G17697: signal is true;
	signal G17698: std_logic; attribute dont_touch of G17698: signal is true;
	signal G17701: std_logic; attribute dont_touch of G17701: signal is true;
	signal G17704: std_logic; attribute dont_touch of G17704: signal is true;
	signal G17707: std_logic; attribute dont_touch of G17707: signal is true;
	signal G17710: std_logic; attribute dont_touch of G17710: signal is true;
	signal G17713: std_logic; attribute dont_touch of G17713: signal is true;
	signal G17714: std_logic; attribute dont_touch of G17714: signal is true;
	signal G17715: std_logic; attribute dont_touch of G17715: signal is true;
	signal G17716: std_logic; attribute dont_touch of G17716: signal is true;
	signal G17717: std_logic; attribute dont_touch of G17717: signal is true;
	signal G17718: std_logic; attribute dont_touch of G17718: signal is true;
	signal G17719: std_logic; attribute dont_touch of G17719: signal is true;
	signal G17720: std_logic; attribute dont_touch of G17720: signal is true;
	signal G17724: std_logic; attribute dont_touch of G17724: signal is true;
	signal G17729: std_logic; attribute dont_touch of G17729: signal is true;
	signal G17734: std_logic; attribute dont_touch of G17734: signal is true;
	signal G17735: std_logic; attribute dont_touch of G17735: signal is true;
	signal G17736: std_logic; attribute dont_touch of G17736: signal is true;
	signal G17737: std_logic; attribute dont_touch of G17737: signal is true;
	signal G17738: std_logic; attribute dont_touch of G17738: signal is true;
	signal G17741: std_logic; attribute dont_touch of G17741: signal is true;
	signal G17746: std_logic; attribute dont_touch of G17746: signal is true;
	signal G17749: std_logic; attribute dont_touch of G17749: signal is true;
	signal G17752: std_logic; attribute dont_touch of G17752: signal is true;
	signal G17753: std_logic; attribute dont_touch of G17753: signal is true;
	signal G17754: std_logic; attribute dont_touch of G17754: signal is true;
	signal G17755: std_logic; attribute dont_touch of G17755: signal is true;
	signal G17758: std_logic; attribute dont_touch of G17758: signal is true;
	signal G17761: std_logic; attribute dont_touch of G17761: signal is true;
	signal G17764: std_logic; attribute dont_touch of G17764: signal is true;
	signal G17767: std_logic; attribute dont_touch of G17767: signal is true;
	signal G17770: std_logic; attribute dont_touch of G17770: signal is true;
	signal G17773: std_logic; attribute dont_touch of G17773: signal is true;
	signal G17774: std_logic; attribute dont_touch of G17774: signal is true;
	signal G17775: std_logic; attribute dont_touch of G17775: signal is true;
	signal G17776: std_logic; attribute dont_touch of G17776: signal is true;
	signal G17779: std_logic; attribute dont_touch of G17779: signal is true;
	signal G17782: std_logic; attribute dont_touch of G17782: signal is true;
	signal G17785: std_logic; attribute dont_touch of G17785: signal is true;
	signal G17788: std_logic; attribute dont_touch of G17788: signal is true;
	signal G17791: std_logic; attribute dont_touch of G17791: signal is true;
	signal G17794: std_logic; attribute dont_touch of G17794: signal is true;
	signal G17795: std_logic; attribute dont_touch of G17795: signal is true;
	signal G17796: std_logic; attribute dont_touch of G17796: signal is true;
	signal G17797: std_logic; attribute dont_touch of G17797: signal is true;
	signal G17798: std_logic; attribute dont_touch of G17798: signal is true;
	signal G17799: std_logic; attribute dont_touch of G17799: signal is true;
	signal G17802: std_logic; attribute dont_touch of G17802: signal is true;
	signal G17807: std_logic; attribute dont_touch of G17807: signal is true;
	signal G17812: std_logic; attribute dont_touch of G17812: signal is true;
	signal G17813: std_logic; attribute dont_touch of G17813: signal is true;
	signal G17814: std_logic; attribute dont_touch of G17814: signal is true;
	signal G17815: std_logic; attribute dont_touch of G17815: signal is true;
	signal G17824: std_logic; attribute dont_touch of G17824: signal is true;
	signal G17825: std_logic; attribute dont_touch of G17825: signal is true;
	signal G17830: std_logic; attribute dont_touch of G17830: signal is true;
	signal G17835: std_logic; attribute dont_touch of G17835: signal is true;
	signal G17836: std_logic; attribute dont_touch of G17836: signal is true;
	signal G17837: std_logic; attribute dont_touch of G17837: signal is true;
	signal G17838: std_logic; attribute dont_touch of G17838: signal is true;
	signal G17839: std_logic; attribute dont_touch of G17839: signal is true;
	signal G17842: std_logic; attribute dont_touch of G17842: signal is true;
	signal G17847: std_logic; attribute dont_touch of G17847: signal is true;
	signal G17850: std_logic; attribute dont_touch of G17850: signal is true;
	signal G17853: std_logic; attribute dont_touch of G17853: signal is true;
	signal G17854: std_logic; attribute dont_touch of G17854: signal is true;
	signal G17855: std_logic; attribute dont_touch of G17855: signal is true;
	signal G17856: std_logic; attribute dont_touch of G17856: signal is true;
	signal G17859: std_logic; attribute dont_touch of G17859: signal is true;
	signal G17862: std_logic; attribute dont_touch of G17862: signal is true;
	signal G17865: std_logic; attribute dont_touch of G17865: signal is true;
	signal G17868: std_logic; attribute dont_touch of G17868: signal is true;
	signal G17871: std_logic; attribute dont_touch of G17871: signal is true;
	signal G17874: std_logic; attribute dont_touch of G17874: signal is true;
	signal G17875: std_logic; attribute dont_touch of G17875: signal is true;
	signal G17876: std_logic; attribute dont_touch of G17876: signal is true;
	signal G17877: std_logic; attribute dont_touch of G17877: signal is true;
	signal G17878: std_logic; attribute dont_touch of G17878: signal is true;
	signal G17882: std_logic; attribute dont_touch of G17882: signal is true;
	signal G17887: std_logic; attribute dont_touch of G17887: signal is true;
	signal G17892: std_logic; attribute dont_touch of G17892: signal is true;
	signal G17893: std_logic; attribute dont_touch of G17893: signal is true;
	signal G17896: std_logic; attribute dont_touch of G17896: signal is true;
	signal G17900: std_logic; attribute dont_touch of G17900: signal is true;
	signal G17901: std_logic; attribute dont_touch of G17901: signal is true;
	signal G17902: std_logic; attribute dont_touch of G17902: signal is true;
	signal G17903: std_logic; attribute dont_touch of G17903: signal is true;
	signal G17912: std_logic; attribute dont_touch of G17912: signal is true;
	signal G17913: std_logic; attribute dont_touch of G17913: signal is true;
	signal G17914: std_logic; attribute dont_touch of G17914: signal is true;
	signal G17919: std_logic; attribute dont_touch of G17919: signal is true;
	signal G17924: std_logic; attribute dont_touch of G17924: signal is true;
	signal G17925: std_logic; attribute dont_touch of G17925: signal is true;
	signal G17926: std_logic; attribute dont_touch of G17926: signal is true;
	signal G17927: std_logic; attribute dont_touch of G17927: signal is true;
	signal G17936: std_logic; attribute dont_touch of G17936: signal is true;
	signal G17937: std_logic; attribute dont_touch of G17937: signal is true;
	signal G17942: std_logic; attribute dont_touch of G17942: signal is true;
	signal G17947: std_logic; attribute dont_touch of G17947: signal is true;
	signal G17948: std_logic; attribute dont_touch of G17948: signal is true;
	signal G17949: std_logic; attribute dont_touch of G17949: signal is true;
	signal G17950: std_logic; attribute dont_touch of G17950: signal is true;
	signal G17951: std_logic; attribute dont_touch of G17951: signal is true;
	signal G17954: std_logic; attribute dont_touch of G17954: signal is true;
	signal G17959: std_logic; attribute dont_touch of G17959: signal is true;
	signal G17962: std_logic; attribute dont_touch of G17962: signal is true;
	signal G17965: std_logic; attribute dont_touch of G17965: signal is true;
	signal G17966: std_logic; attribute dont_touch of G17966: signal is true;
	signal G17967: std_logic; attribute dont_touch of G17967: signal is true;
	signal G17968: std_logic; attribute dont_touch of G17968: signal is true;
	signal G17969: std_logic; attribute dont_touch of G17969: signal is true;
	signal G17973: std_logic; attribute dont_touch of G17973: signal is true;
	signal G17974: std_logic; attribute dont_touch of G17974: signal is true;
	signal G17979: std_logic; attribute dont_touch of G17979: signal is true;
	signal G17984: std_logic; attribute dont_touch of G17984: signal is true;
	signal G17985: std_logic; attribute dont_touch of G17985: signal is true;
	signal G17988: std_logic; attribute dont_touch of G17988: signal is true;
	signal G17989: std_logic; attribute dont_touch of G17989: signal is true;
	signal G17990: std_logic; attribute dont_touch of G17990: signal is true;
	signal G17991: std_logic; attribute dont_touch of G17991: signal is true;
	signal G17992: std_logic; attribute dont_touch of G17992: signal is true;
	signal G17993: std_logic; attribute dont_touch of G17993: signal is true;
	signal G17998: std_logic; attribute dont_touch of G17998: signal is true;
	signal G18003: std_logic; attribute dont_touch of G18003: signal is true;
	signal G18004: std_logic; attribute dont_touch of G18004: signal is true;
	signal G18007: std_logic; attribute dont_touch of G18007: signal is true;
	signal G18011: std_logic; attribute dont_touch of G18011: signal is true;
	signal G18012: std_logic; attribute dont_touch of G18012: signal is true;
	signal G18013: std_logic; attribute dont_touch of G18013: signal is true;
	signal G18014: std_logic; attribute dont_touch of G18014: signal is true;
	signal G18023: std_logic; attribute dont_touch of G18023: signal is true;
	signal G18024: std_logic; attribute dont_touch of G18024: signal is true;
	signal G18025: std_logic; attribute dont_touch of G18025: signal is true;
	signal G18030: std_logic; attribute dont_touch of G18030: signal is true;
	signal G18035: std_logic; attribute dont_touch of G18035: signal is true;
	signal G18036: std_logic; attribute dont_touch of G18036: signal is true;
	signal G18037: std_logic; attribute dont_touch of G18037: signal is true;
	signal G18038: std_logic; attribute dont_touch of G18038: signal is true;
	signal G18047: std_logic; attribute dont_touch of G18047: signal is true;
	signal G18048: std_logic; attribute dont_touch of G18048: signal is true;
	signal G18053: std_logic; attribute dont_touch of G18053: signal is true;
	signal G18058: std_logic; attribute dont_touch of G18058: signal is true;
	signal G18059: std_logic; attribute dont_touch of G18059: signal is true;
	signal G18060: std_logic; attribute dont_touch of G18060: signal is true;
	signal G18061: std_logic; attribute dont_touch of G18061: signal is true;
	signal G18062: std_logic; attribute dont_touch of G18062: signal is true;
	signal G18063: std_logic; attribute dont_touch of G18063: signal is true;
	signal G18070: std_logic; attribute dont_touch of G18070: signal is true;
	signal G18074: std_logic; attribute dont_touch of G18074: signal is true;
	signal G18079: std_logic; attribute dont_touch of G18079: signal is true;
	signal G18084: std_logic; attribute dont_touch of G18084: signal is true;
	signal G18085: std_logic; attribute dont_touch of G18085: signal is true;
	signal G18088: std_logic; attribute dont_touch of G18088: signal is true;
	signal G18089: std_logic; attribute dont_touch of G18089: signal is true;
	signal G18090: std_logic; attribute dont_touch of G18090: signal is true;
	signal G18091: std_logic; attribute dont_touch of G18091: signal is true;
	signal G18096: std_logic; attribute dont_touch of G18096: signal is true;
	signal G18101: std_logic; attribute dont_touch of G18101: signal is true;
	signal G18102: std_logic; attribute dont_touch of G18102: signal is true;
	signal G18105: std_logic; attribute dont_touch of G18105: signal is true;
	signal G18106: std_logic; attribute dont_touch of G18106: signal is true;
	signal G18107: std_logic; attribute dont_touch of G18107: signal is true;
	signal G18108: std_logic; attribute dont_touch of G18108: signal is true;
	signal G18109: std_logic; attribute dont_touch of G18109: signal is true;
	signal G18110: std_logic; attribute dont_touch of G18110: signal is true;
	signal G18115: std_logic; attribute dont_touch of G18115: signal is true;
	signal G18120: std_logic; attribute dont_touch of G18120: signal is true;
	signal G18121: std_logic; attribute dont_touch of G18121: signal is true;
	signal G18124: std_logic; attribute dont_touch of G18124: signal is true;
	signal G18128: std_logic; attribute dont_touch of G18128: signal is true;
	signal G18129: std_logic; attribute dont_touch of G18129: signal is true;
	signal G18130: std_logic; attribute dont_touch of G18130: signal is true;
	signal G18131: std_logic; attribute dont_touch of G18131: signal is true;
	signal G18140: std_logic; attribute dont_touch of G18140: signal is true;
	signal G18141: std_logic; attribute dont_touch of G18141: signal is true;
	signal G18142: std_logic; attribute dont_touch of G18142: signal is true;
	signal G18147: std_logic; attribute dont_touch of G18147: signal is true;
	signal G18152: std_logic; attribute dont_touch of G18152: signal is true;
	signal G18153: std_logic; attribute dont_touch of G18153: signal is true;
	signal G18154: std_logic; attribute dont_touch of G18154: signal is true;
	signal G18155: std_logic; attribute dont_touch of G18155: signal is true;
	signal G18164: std_logic; attribute dont_touch of G18164: signal is true;
	signal G18165: std_logic; attribute dont_touch of G18165: signal is true;
	signal G18166: std_logic; attribute dont_touch of G18166: signal is true;
	signal G18169: std_logic; attribute dont_touch of G18169: signal is true;
	signal G18170: std_logic; attribute dont_touch of G18170: signal is true;
	signal G18174: std_logic; attribute dont_touch of G18174: signal is true;
	signal G18179: std_logic; attribute dont_touch of G18179: signal is true;
	signal G18183: std_logic; attribute dont_touch of G18183: signal is true;
	signal G18188: std_logic; attribute dont_touch of G18188: signal is true;
	signal G18189: std_logic; attribute dont_touch of G18189: signal is true;
	signal G18190: std_logic; attribute dont_touch of G18190: signal is true;
	signal G18195: std_logic; attribute dont_touch of G18195: signal is true;
	signal G18200: std_logic; attribute dont_touch of G18200: signal is true;
	signal G18201: std_logic; attribute dont_touch of G18201: signal is true;
	signal G18204: std_logic; attribute dont_touch of G18204: signal is true;
	signal G18205: std_logic; attribute dont_touch of G18205: signal is true;
	signal G18206: std_logic; attribute dont_touch of G18206: signal is true;
	signal G18207: std_logic; attribute dont_touch of G18207: signal is true;
	signal G18212: std_logic; attribute dont_touch of G18212: signal is true;
	signal G18217: std_logic; attribute dont_touch of G18217: signal is true;
	signal G18218: std_logic; attribute dont_touch of G18218: signal is true;
	signal G18221: std_logic; attribute dont_touch of G18221: signal is true;
	signal G18222: std_logic; attribute dont_touch of G18222: signal is true;
	signal G18223: std_logic; attribute dont_touch of G18223: signal is true;
	signal G18224: std_logic; attribute dont_touch of G18224: signal is true;
	signal G18225: std_logic; attribute dont_touch of G18225: signal is true;
	signal G18226: std_logic; attribute dont_touch of G18226: signal is true;
	signal G18231: std_logic; attribute dont_touch of G18231: signal is true;
	signal G18236: std_logic; attribute dont_touch of G18236: signal is true;
	signal G18237: std_logic; attribute dont_touch of G18237: signal is true;
	signal G18240: std_logic; attribute dont_touch of G18240: signal is true;
	signal G18244: std_logic; attribute dont_touch of G18244: signal is true;
	signal G18245: std_logic; attribute dont_touch of G18245: signal is true;
	signal G18246: std_logic; attribute dont_touch of G18246: signal is true;
	signal G18247: std_logic; attribute dont_touch of G18247: signal is true;
	signal G18256: std_logic; attribute dont_touch of G18256: signal is true;
	signal G18257: std_logic; attribute dont_touch of G18257: signal is true;
	signal G18258: std_logic; attribute dont_touch of G18258: signal is true;
	signal G18261: std_logic; attribute dont_touch of G18261: signal is true;
	signal G18265: std_logic; attribute dont_touch of G18265: signal is true;
	signal G18270: std_logic; attribute dont_touch of G18270: signal is true;
	signal G18275: std_logic; attribute dont_touch of G18275: signal is true;
	signal G18276: std_logic; attribute dont_touch of G18276: signal is true;
	signal G18277: std_logic; attribute dont_touch of G18277: signal is true;
	signal G18278: std_logic; attribute dont_touch of G18278: signal is true;
	signal G18281: std_logic; attribute dont_touch of G18281: signal is true;
	signal G18286: std_logic; attribute dont_touch of G18286: signal is true;
	signal G18290: std_logic; attribute dont_touch of G18290: signal is true;
	signal G18295: std_logic; attribute dont_touch of G18295: signal is true;
	signal G18296: std_logic; attribute dont_touch of G18296: signal is true;
	signal G18297: std_logic; attribute dont_touch of G18297: signal is true;
	signal G18302: std_logic; attribute dont_touch of G18302: signal is true;
	signal G18307: std_logic; attribute dont_touch of G18307: signal is true;
	signal G18308: std_logic; attribute dont_touch of G18308: signal is true;
	signal G18311: std_logic; attribute dont_touch of G18311: signal is true;
	signal G18312: std_logic; attribute dont_touch of G18312: signal is true;
	signal G18313: std_logic; attribute dont_touch of G18313: signal is true;
	signal G18314: std_logic; attribute dont_touch of G18314: signal is true;
	signal G18319: std_logic; attribute dont_touch of G18319: signal is true;
	signal G18324: std_logic; attribute dont_touch of G18324: signal is true;
	signal G18325: std_logic; attribute dont_touch of G18325: signal is true;
	signal G18328: std_logic; attribute dont_touch of G18328: signal is true;
	signal G18329: std_logic; attribute dont_touch of G18329: signal is true;
	signal G18330: std_logic; attribute dont_touch of G18330: signal is true;
	signal G18331: std_logic; attribute dont_touch of G18331: signal is true;
	signal G18332: std_logic; attribute dont_touch of G18332: signal is true;
	signal G18333: std_logic; attribute dont_touch of G18333: signal is true;
	signal G18334: std_logic; attribute dont_touch of G18334: signal is true;
	signal G18337: std_logic; attribute dont_touch of G18337: signal is true;
	signal G18341: std_logic; attribute dont_touch of G18341: signal is true;
	signal G18346: std_logic; attribute dont_touch of G18346: signal is true;
	signal G18351: std_logic; attribute dont_touch of G18351: signal is true;
	signal G18352: std_logic; attribute dont_touch of G18352: signal is true;
	signal G18353: std_logic; attribute dont_touch of G18353: signal is true;
	signal G18354: std_logic; attribute dont_touch of G18354: signal is true;
	signal G18355: std_logic; attribute dont_touch of G18355: signal is true;
	signal G18358: std_logic; attribute dont_touch of G18358: signal is true;
	signal G18363: std_logic; attribute dont_touch of G18363: signal is true;
	signal G18368: std_logic; attribute dont_touch of G18368: signal is true;
	signal G18369: std_logic; attribute dont_touch of G18369: signal is true;
	signal G18370: std_logic; attribute dont_touch of G18370: signal is true;
	signal G18371: std_logic; attribute dont_touch of G18371: signal is true;
	signal G18374: std_logic; attribute dont_touch of G18374: signal is true;
	signal G18379: std_logic; attribute dont_touch of G18379: signal is true;
	signal G18383: std_logic; attribute dont_touch of G18383: signal is true;
	signal G18388: std_logic; attribute dont_touch of G18388: signal is true;
	signal G18389: std_logic; attribute dont_touch of G18389: signal is true;
	signal G18390: std_logic; attribute dont_touch of G18390: signal is true;
	signal G18395: std_logic; attribute dont_touch of G18395: signal is true;
	signal G18400: std_logic; attribute dont_touch of G18400: signal is true;
	signal G18401: std_logic; attribute dont_touch of G18401: signal is true;
	signal G18404: std_logic; attribute dont_touch of G18404: signal is true;
	signal G18405: std_logic; attribute dont_touch of G18405: signal is true;
	signal G18406: std_logic; attribute dont_touch of G18406: signal is true;
	signal G18407: std_logic; attribute dont_touch of G18407: signal is true;
	signal G18414: std_logic; attribute dont_touch of G18414: signal is true;
	signal G18415: std_logic; attribute dont_touch of G18415: signal is true;
	signal G18419: std_logic; attribute dont_touch of G18419: signal is true;
	signal G18424: std_logic; attribute dont_touch of G18424: signal is true;
	signal G18429: std_logic; attribute dont_touch of G18429: signal is true;
	signal G18430: std_logic; attribute dont_touch of G18430: signal is true;
	signal G18431: std_logic; attribute dont_touch of G18431: signal is true;
	signal G18432: std_logic; attribute dont_touch of G18432: signal is true;
	signal G18435: std_logic; attribute dont_touch of G18435: signal is true;
	signal G18436: std_logic; attribute dont_touch of G18436: signal is true;
	signal G18441: std_logic; attribute dont_touch of G18441: signal is true;
	signal G18446: std_logic; attribute dont_touch of G18446: signal is true;
	signal G18447: std_logic; attribute dont_touch of G18447: signal is true;
	signal G18448: std_logic; attribute dont_touch of G18448: signal is true;
	signal G18449: std_logic; attribute dont_touch of G18449: signal is true;
	signal G18450: std_logic; attribute dont_touch of G18450: signal is true;
	signal G18453: std_logic; attribute dont_touch of G18453: signal is true;
	signal G18458: std_logic; attribute dont_touch of G18458: signal is true;
	signal G18463: std_logic; attribute dont_touch of G18463: signal is true;
	signal G18464: std_logic; attribute dont_touch of G18464: signal is true;
	signal G18465: std_logic; attribute dont_touch of G18465: signal is true;
	signal G18466: std_logic; attribute dont_touch of G18466: signal is true;
	signal G18469: std_logic; attribute dont_touch of G18469: signal is true;
	signal G18474: std_logic; attribute dont_touch of G18474: signal is true;
	signal G18478: std_logic; attribute dont_touch of G18478: signal is true;
	signal G18483: std_logic; attribute dont_touch of G18483: signal is true;
	signal G18484: std_logic; attribute dont_touch of G18484: signal is true;
	signal G18485: std_logic; attribute dont_touch of G18485: signal is true;
	signal G18486: std_logic; attribute dont_touch of G18486: signal is true;
	signal G18490: std_logic; attribute dont_touch of G18490: signal is true;
	signal G18491: std_logic; attribute dont_touch of G18491: signal is true;
	signal G18492: std_logic; attribute dont_touch of G18492: signal is true;
	signal G18497: std_logic; attribute dont_touch of G18497: signal is true;
	signal G18502: std_logic; attribute dont_touch of G18502: signal is true;
	signal G18503: std_logic; attribute dont_touch of G18503: signal is true;
	signal G18504: std_logic; attribute dont_touch of G18504: signal is true;
	signal G18505: std_logic; attribute dont_touch of G18505: signal is true;
	signal G18508: std_logic; attribute dont_touch of G18508: signal is true;
	signal G18509: std_logic; attribute dont_touch of G18509: signal is true;
	signal G18514: std_logic; attribute dont_touch of G18514: signal is true;
	signal G18519: std_logic; attribute dont_touch of G18519: signal is true;
	signal G18520: std_logic; attribute dont_touch of G18520: signal is true;
	signal G18521: std_logic; attribute dont_touch of G18521: signal is true;
	signal G18522: std_logic; attribute dont_touch of G18522: signal is true;
	signal G18523: std_logic; attribute dont_touch of G18523: signal is true;
	signal G18526: std_logic; attribute dont_touch of G18526: signal is true;
	signal G18531: std_logic; attribute dont_touch of G18531: signal is true;
	signal G18536: std_logic; attribute dont_touch of G18536: signal is true;
	signal G18537: std_logic; attribute dont_touch of G18537: signal is true;
	signal G18538: std_logic; attribute dont_touch of G18538: signal is true;
	signal G18539: std_logic; attribute dont_touch of G18539: signal is true;
	signal G18542: std_logic; attribute dont_touch of G18542: signal is true;
	signal G18543: std_logic; attribute dont_touch of G18543: signal is true;
	signal G18547: std_logic; attribute dont_touch of G18547: signal is true;
	signal G18548: std_logic; attribute dont_touch of G18548: signal is true;
	signal G18552: std_logic; attribute dont_touch of G18552: signal is true;
	signal G18553: std_logic; attribute dont_touch of G18553: signal is true;
	signal G18554: std_logic; attribute dont_touch of G18554: signal is true;
	signal G18555: std_logic; attribute dont_touch of G18555: signal is true;
	signal G18556: std_logic; attribute dont_touch of G18556: signal is true;
	signal G18561: std_logic; attribute dont_touch of G18561: signal is true;
	signal G18566: std_logic; attribute dont_touch of G18566: signal is true;
	signal G18567: std_logic; attribute dont_touch of G18567: signal is true;
	signal G18568: std_logic; attribute dont_touch of G18568: signal is true;
	signal G18569: std_logic; attribute dont_touch of G18569: signal is true;
	signal G18572: std_logic; attribute dont_touch of G18572: signal is true;
	signal G18573: std_logic; attribute dont_touch of G18573: signal is true;
	signal G18578: std_logic; attribute dont_touch of G18578: signal is true;
	signal G18583: std_logic; attribute dont_touch of G18583: signal is true;
	signal G18584: std_logic; attribute dont_touch of G18584: signal is true;
	signal G18585: std_logic; attribute dont_touch of G18585: signal is true;
	signal G18586: std_logic; attribute dont_touch of G18586: signal is true;
	signal G18587: std_logic; attribute dont_touch of G18587: signal is true;
	signal G18590: std_logic; attribute dont_touch of G18590: signal is true;
	signal G18593: std_logic; attribute dont_touch of G18593: signal is true;
	signal G18597: std_logic; attribute dont_touch of G18597: signal is true;
	signal G18598: std_logic; attribute dont_touch of G18598: signal is true;
	signal G18602: std_logic; attribute dont_touch of G18602: signal is true;
	signal G18603: std_logic; attribute dont_touch of G18603: signal is true;
	signal G18604: std_logic; attribute dont_touch of G18604: signal is true;
	signal G18605: std_logic; attribute dont_touch of G18605: signal is true;
	signal G18606: std_logic; attribute dont_touch of G18606: signal is true;
	signal G18611: std_logic; attribute dont_touch of G18611: signal is true;
	signal G18616: std_logic; attribute dont_touch of G18616: signal is true;
	signal G18617: std_logic; attribute dont_touch of G18617: signal is true;
	signal G18618: std_logic; attribute dont_touch of G18618: signal is true;
	signal G18619: std_logic; attribute dont_touch of G18619: signal is true;
	signal G18622: std_logic; attribute dont_touch of G18622: signal is true;
	signal G18623: std_logic; attribute dont_touch of G18623: signal is true;
	signal G18626: std_logic; attribute dont_touch of G18626: signal is true;
	signal G18629: std_logic; attribute dont_touch of G18629: signal is true;
	signal G18630: std_logic; attribute dont_touch of G18630: signal is true;
	signal G18634: std_logic; attribute dont_touch of G18634: signal is true;
	signal G18635: std_logic; attribute dont_touch of G18635: signal is true;
	signal G18636: std_logic; attribute dont_touch of G18636: signal is true;
	signal G18637: std_logic; attribute dont_touch of G18637: signal is true;
	signal G18638: std_logic; attribute dont_touch of G18638: signal is true;
	signal G18639: std_logic; attribute dont_touch of G18639: signal is true;
	signal G18643: std_logic; attribute dont_touch of G18643: signal is true;
	signal G18644: std_logic; attribute dont_touch of G18644: signal is true;
	signal G18645: std_logic; attribute dont_touch of G18645: signal is true;
	signal G18646: std_logic; attribute dont_touch of G18646: signal is true;
	signal G18647: std_logic; attribute dont_touch of G18647: signal is true;
	signal G18648: std_logic; attribute dont_touch of G18648: signal is true;
	signal G18649: std_logic; attribute dont_touch of G18649: signal is true;
	signal G18650: std_logic; attribute dont_touch of G18650: signal is true;
	signal G18651: std_logic; attribute dont_touch of G18651: signal is true;
	signal G18652: std_logic; attribute dont_touch of G18652: signal is true;
	signal G18653: std_logic; attribute dont_touch of G18653: signal is true;
	signal G18654: std_logic; attribute dont_touch of G18654: signal is true;
	signal G18655: std_logic; attribute dont_touch of G18655: signal is true;
	signal G18656: std_logic; attribute dont_touch of G18656: signal is true;
	signal G18665: std_logic; attribute dont_touch of G18665: signal is true;
	signal G18666: std_logic; attribute dont_touch of G18666: signal is true;
	signal G18667: std_logic; attribute dont_touch of G18667: signal is true;
	signal G18668: std_logic; attribute dont_touch of G18668: signal is true;
	signal G18669: std_logic; attribute dont_touch of G18669: signal is true;
	signal G18670: std_logic; attribute dont_touch of G18670: signal is true;
	signal G18678: std_logic; attribute dont_touch of G18678: signal is true;
	signal G18679: std_logic; attribute dont_touch of G18679: signal is true;
	signal G18688: std_logic; attribute dont_touch of G18688: signal is true;
	signal G18689: std_logic; attribute dont_touch of G18689: signal is true;
	signal G18690: std_logic; attribute dont_touch of G18690: signal is true;
	signal G18691: std_logic; attribute dont_touch of G18691: signal is true;
	signal G18692: std_logic; attribute dont_touch of G18692: signal is true;
	signal G18699: std_logic; attribute dont_touch of G18699: signal is true;
	signal G18707: std_logic; attribute dont_touch of G18707: signal is true;
	signal G18708: std_logic; attribute dont_touch of G18708: signal is true;
	signal G18717: std_logic; attribute dont_touch of G18717: signal is true;
	signal G18718: std_logic; attribute dont_touch of G18718: signal is true;
	signal G18719: std_logic; attribute dont_touch of G18719: signal is true;
	signal G18720: std_logic; attribute dont_touch of G18720: signal is true;
	signal G18725: std_logic; attribute dont_touch of G18725: signal is true;
	signal G18726: std_logic; attribute dont_touch of G18726: signal is true;
	signal G18727: std_logic; attribute dont_touch of G18727: signal is true;
	signal G18728: std_logic; attribute dont_touch of G18728: signal is true;
	signal G18735: std_logic; attribute dont_touch of G18735: signal is true;
	signal G18743: std_logic; attribute dont_touch of G18743: signal is true;
	signal G18744: std_logic; attribute dont_touch of G18744: signal is true;
	signal G18753: std_logic; attribute dont_touch of G18753: signal is true;
	signal G18754: std_logic; attribute dont_touch of G18754: signal is true;
	signal G18755: std_logic; attribute dont_touch of G18755: signal is true;
	signal G18756: std_logic; attribute dont_touch of G18756: signal is true;
	signal G18757: std_logic; attribute dont_touch of G18757: signal is true;
	signal G18758: std_logic; attribute dont_touch of G18758: signal is true;
	signal G18763: std_logic; attribute dont_touch of G18763: signal is true;
	signal G18764: std_logic; attribute dont_touch of G18764: signal is true;
	signal G18765: std_logic; attribute dont_touch of G18765: signal is true;
	signal G18772: std_logic; attribute dont_touch of G18772: signal is true;
	signal G18780: std_logic; attribute dont_touch of G18780: signal is true;
	signal G18781: std_logic; attribute dont_touch of G18781: signal is true;
	signal G18782: std_logic; attribute dont_touch of G18782: signal is true;
	signal G18783: std_logic; attribute dont_touch of G18783: signal is true;
	signal G18784: std_logic; attribute dont_touch of G18784: signal is true;
	signal G18785: std_logic; attribute dont_touch of G18785: signal is true;
	signal G18786: std_logic; attribute dont_touch of G18786: signal is true;
	signal G18787: std_logic; attribute dont_touch of G18787: signal is true;
	signal G18788: std_logic; attribute dont_touch of G18788: signal is true;
	signal G18789: std_logic; attribute dont_touch of G18789: signal is true;
	signal G18794: std_logic; attribute dont_touch of G18794: signal is true;
	signal G18795: std_logic; attribute dont_touch of G18795: signal is true;
	signal G18796: std_logic; attribute dont_touch of G18796: signal is true;
	signal G18803: std_logic; attribute dont_touch of G18803: signal is true;
	signal G18804: std_logic; attribute dont_touch of G18804: signal is true;
	signal G18805: std_logic; attribute dont_touch of G18805: signal is true;
	signal G18806: std_logic; attribute dont_touch of G18806: signal is true;
	signal G18807: std_logic; attribute dont_touch of G18807: signal is true;
	signal G18808: std_logic; attribute dont_touch of G18808: signal is true;
	signal G18809: std_logic; attribute dont_touch of G18809: signal is true;
	signal G18810: std_logic; attribute dont_touch of G18810: signal is true;
	signal G18811: std_logic; attribute dont_touch of G18811: signal is true;
	signal G18812: std_logic; attribute dont_touch of G18812: signal is true;
	signal G18813: std_logic; attribute dont_touch of G18813: signal is true;
	signal G18814: std_logic; attribute dont_touch of G18814: signal is true;
	signal G18815: std_logic; attribute dont_touch of G18815: signal is true;
	signal G18820: std_logic; attribute dont_touch of G18820: signal is true;
	signal G18821: std_logic; attribute dont_touch of G18821: signal is true;
	signal G18822: std_logic; attribute dont_touch of G18822: signal is true;
	signal G18823: std_logic; attribute dont_touch of G18823: signal is true;
	signal G18824: std_logic; attribute dont_touch of G18824: signal is true;
	signal G18825: std_logic; attribute dont_touch of G18825: signal is true;
	signal G18826: std_logic; attribute dont_touch of G18826: signal is true;
	signal G18827: std_logic; attribute dont_touch of G18827: signal is true;
	signal G18828: std_logic; attribute dont_touch of G18828: signal is true;
	signal G18829: std_logic; attribute dont_touch of G18829: signal is true;
	signal G18830: std_logic; attribute dont_touch of G18830: signal is true;
	signal G18831: std_logic; attribute dont_touch of G18831: signal is true;
	signal G18832: std_logic; attribute dont_touch of G18832: signal is true;
	signal G18833: std_logic; attribute dont_touch of G18833: signal is true;
	signal G18834: std_logic; attribute dont_touch of G18834: signal is true;
	signal G18835: std_logic; attribute dont_touch of G18835: signal is true;
	signal G18836: std_logic; attribute dont_touch of G18836: signal is true;
	signal G18837: std_logic; attribute dont_touch of G18837: signal is true;
	signal G18838: std_logic; attribute dont_touch of G18838: signal is true;
	signal G18839: std_logic; attribute dont_touch of G18839: signal is true;
	signal G18840: std_logic; attribute dont_touch of G18840: signal is true;
	signal G18841: std_logic; attribute dont_touch of G18841: signal is true;
	signal G18842: std_logic; attribute dont_touch of G18842: signal is true;
	signal G18843: std_logic; attribute dont_touch of G18843: signal is true;
	signal G18844: std_logic; attribute dont_touch of G18844: signal is true;
	signal G18845: std_logic; attribute dont_touch of G18845: signal is true;
	signal G18846: std_logic; attribute dont_touch of G18846: signal is true;
	signal G18847: std_logic; attribute dont_touch of G18847: signal is true;
	signal G18848: std_logic; attribute dont_touch of G18848: signal is true;
	signal G18849: std_logic; attribute dont_touch of G18849: signal is true;
	signal G18850: std_logic; attribute dont_touch of G18850: signal is true;
	signal G18851: std_logic; attribute dont_touch of G18851: signal is true;
	signal G18852: std_logic; attribute dont_touch of G18852: signal is true;
	signal G18853: std_logic; attribute dont_touch of G18853: signal is true;
	signal G18854: std_logic; attribute dont_touch of G18854: signal is true;
	signal G18855: std_logic; attribute dont_touch of G18855: signal is true;
	signal G18856: std_logic; attribute dont_touch of G18856: signal is true;
	signal G18857: std_logic; attribute dont_touch of G18857: signal is true;
	signal G18858: std_logic; attribute dont_touch of G18858: signal is true;
	signal G18859: std_logic; attribute dont_touch of G18859: signal is true;
	signal G18860: std_logic; attribute dont_touch of G18860: signal is true;
	signal G18861: std_logic; attribute dont_touch of G18861: signal is true;
	signal G18862: std_logic; attribute dont_touch of G18862: signal is true;
	signal G18863: std_logic; attribute dont_touch of G18863: signal is true;
	signal G18864: std_logic; attribute dont_touch of G18864: signal is true;
	signal G18865: std_logic; attribute dont_touch of G18865: signal is true;
	signal G18866: std_logic; attribute dont_touch of G18866: signal is true;
	signal G18867: std_logic; attribute dont_touch of G18867: signal is true;
	signal G18868: std_logic; attribute dont_touch of G18868: signal is true;
	signal G18869: std_logic; attribute dont_touch of G18869: signal is true;
	signal G18870: std_logic; attribute dont_touch of G18870: signal is true;
	signal G18871: std_logic; attribute dont_touch of G18871: signal is true;
	signal G18872: std_logic; attribute dont_touch of G18872: signal is true;
	signal G18873: std_logic; attribute dont_touch of G18873: signal is true;
	signal G18874: std_logic; attribute dont_touch of G18874: signal is true;
	signal G18875: std_logic; attribute dont_touch of G18875: signal is true;
	signal G18876: std_logic; attribute dont_touch of G18876: signal is true;
	signal G18877: std_logic; attribute dont_touch of G18877: signal is true;
	signal G18878: std_logic; attribute dont_touch of G18878: signal is true;
	signal G18879: std_logic; attribute dont_touch of G18879: signal is true;
	signal G18880: std_logic; attribute dont_touch of G18880: signal is true;
	signal G18881: std_logic; attribute dont_touch of G18881: signal is true;
	signal G18882: std_logic; attribute dont_touch of G18882: signal is true;
	signal G18883: std_logic; attribute dont_touch of G18883: signal is true;
	signal G18884: std_logic; attribute dont_touch of G18884: signal is true;
	signal G18885: std_logic; attribute dont_touch of G18885: signal is true;
	signal G18886: std_logic; attribute dont_touch of G18886: signal is true;
	signal G18890: std_logic; attribute dont_touch of G18890: signal is true;
	signal G18891: std_logic; attribute dont_touch of G18891: signal is true;
	signal G18892: std_logic; attribute dont_touch of G18892: signal is true;
	signal G18893: std_logic; attribute dont_touch of G18893: signal is true;
	signal G18894: std_logic; attribute dont_touch of G18894: signal is true;
	signal G18895: std_logic; attribute dont_touch of G18895: signal is true;
	signal G18896: std_logic; attribute dont_touch of G18896: signal is true;
	signal G18897: std_logic; attribute dont_touch of G18897: signal is true;
	signal G18898: std_logic; attribute dont_touch of G18898: signal is true;
	signal G18899: std_logic; attribute dont_touch of G18899: signal is true;
	signal G18900: std_logic; attribute dont_touch of G18900: signal is true;
	signal G18901: std_logic; attribute dont_touch of G18901: signal is true;
	signal G18902: std_logic; attribute dont_touch of G18902: signal is true;
	signal G18903: std_logic; attribute dont_touch of G18903: signal is true;
	signal G18904: std_logic; attribute dont_touch of G18904: signal is true;
	signal G18905: std_logic; attribute dont_touch of G18905: signal is true;
	signal G18906: std_logic; attribute dont_touch of G18906: signal is true;
	signal G18907: std_logic; attribute dont_touch of G18907: signal is true;
	signal G18908: std_logic; attribute dont_touch of G18908: signal is true;
	signal G18909: std_logic; attribute dont_touch of G18909: signal is true;
	signal G18910: std_logic; attribute dont_touch of G18910: signal is true;
	signal G18911: std_logic; attribute dont_touch of G18911: signal is true;
	signal G18912: std_logic; attribute dont_touch of G18912: signal is true;
	signal G18913: std_logic; attribute dont_touch of G18913: signal is true;
	signal G18914: std_logic; attribute dont_touch of G18914: signal is true;
	signal G18915: std_logic; attribute dont_touch of G18915: signal is true;
	signal G18916: std_logic; attribute dont_touch of G18916: signal is true;
	signal G18917: std_logic; attribute dont_touch of G18917: signal is true;
	signal G18918: std_logic; attribute dont_touch of G18918: signal is true;
	signal G18919: std_logic; attribute dont_touch of G18919: signal is true;
	signal G18920: std_logic; attribute dont_touch of G18920: signal is true;
	signal G18921: std_logic; attribute dont_touch of G18921: signal is true;
	signal G18922: std_logic; attribute dont_touch of G18922: signal is true;
	signal G18923: std_logic; attribute dont_touch of G18923: signal is true;
	signal G18924: std_logic; attribute dont_touch of G18924: signal is true;
	signal G18925: std_logic; attribute dont_touch of G18925: signal is true;
	signal G18926: std_logic; attribute dont_touch of G18926: signal is true;
	signal G18927: std_logic; attribute dont_touch of G18927: signal is true;
	signal G18928: std_logic; attribute dont_touch of G18928: signal is true;
	signal G18929: std_logic; attribute dont_touch of G18929: signal is true;
	signal G18930: std_logic; attribute dont_touch of G18930: signal is true;
	signal G18931: std_logic; attribute dont_touch of G18931: signal is true;
	signal G18932: std_logic; attribute dont_touch of G18932: signal is true;
	signal G18933: std_logic; attribute dont_touch of G18933: signal is true;
	signal G18934: std_logic; attribute dont_touch of G18934: signal is true;
	signal G18935: std_logic; attribute dont_touch of G18935: signal is true;
	signal G18936: std_logic; attribute dont_touch of G18936: signal is true;
	signal G18937: std_logic; attribute dont_touch of G18937: signal is true;
	signal G18938: std_logic; attribute dont_touch of G18938: signal is true;
	signal G18939: std_logic; attribute dont_touch of G18939: signal is true;
	signal G18940: std_logic; attribute dont_touch of G18940: signal is true;
	signal G18941: std_logic; attribute dont_touch of G18941: signal is true;
	signal G18942: std_logic; attribute dont_touch of G18942: signal is true;
	signal G18943: std_logic; attribute dont_touch of G18943: signal is true;
	signal G18944: std_logic; attribute dont_touch of G18944: signal is true;
	signal G18945: std_logic; attribute dont_touch of G18945: signal is true;
	signal G18946: std_logic; attribute dont_touch of G18946: signal is true;
	signal G18947: std_logic; attribute dont_touch of G18947: signal is true;
	signal G18948: std_logic; attribute dont_touch of G18948: signal is true;
	signal G18949: std_logic; attribute dont_touch of G18949: signal is true;
	signal G18950: std_logic; attribute dont_touch of G18950: signal is true;
	signal G18951: std_logic; attribute dont_touch of G18951: signal is true;
	signal G18952: std_logic; attribute dont_touch of G18952: signal is true;
	signal G18953: std_logic; attribute dont_touch of G18953: signal is true;
	signal G18954: std_logic; attribute dont_touch of G18954: signal is true;
	signal G18955: std_logic; attribute dont_touch of G18955: signal is true;
	signal G18956: std_logic; attribute dont_touch of G18956: signal is true;
	signal G18957: std_logic; attribute dont_touch of G18957: signal is true;
	signal G18958: std_logic; attribute dont_touch of G18958: signal is true;
	signal G18959: std_logic; attribute dont_touch of G18959: signal is true;
	signal G18960: std_logic; attribute dont_touch of G18960: signal is true;
	signal G18961: std_logic; attribute dont_touch of G18961: signal is true;
	signal G18962: std_logic; attribute dont_touch of G18962: signal is true;
	signal G18963: std_logic; attribute dont_touch of G18963: signal is true;
	signal G18964: std_logic; attribute dont_touch of G18964: signal is true;
	signal G18965: std_logic; attribute dont_touch of G18965: signal is true;
	signal G18966: std_logic; attribute dont_touch of G18966: signal is true;
	signal G18967: std_logic; attribute dont_touch of G18967: signal is true;
	signal G18968: std_logic; attribute dont_touch of G18968: signal is true;
	signal G18969: std_logic; attribute dont_touch of G18969: signal is true;
	signal G18970: std_logic; attribute dont_touch of G18970: signal is true;
	signal G18971: std_logic; attribute dont_touch of G18971: signal is true;
	signal G18972: std_logic; attribute dont_touch of G18972: signal is true;
	signal G18973: std_logic; attribute dont_touch of G18973: signal is true;
	signal G18974: std_logic; attribute dont_touch of G18974: signal is true;
	signal G18975: std_logic; attribute dont_touch of G18975: signal is true;
	signal G18976: std_logic; attribute dont_touch of G18976: signal is true;
	signal G18977: std_logic; attribute dont_touch of G18977: signal is true;
	signal G18980: std_logic; attribute dont_touch of G18980: signal is true;
	signal G18981: std_logic; attribute dont_touch of G18981: signal is true;
	signal G18982: std_logic; attribute dont_touch of G18982: signal is true;
	signal G18983: std_logic; attribute dont_touch of G18983: signal is true;
	signal G18984: std_logic; attribute dont_touch of G18984: signal is true;
	signal G18985: std_logic; attribute dont_touch of G18985: signal is true;
	signal G18986: std_logic; attribute dont_touch of G18986: signal is true;
	signal G18987: std_logic; attribute dont_touch of G18987: signal is true;
	signal G18988: std_logic; attribute dont_touch of G18988: signal is true;
	signal G18989: std_logic; attribute dont_touch of G18989: signal is true;
	signal G18990: std_logic; attribute dont_touch of G18990: signal is true;
	signal G18991: std_logic; attribute dont_touch of G18991: signal is true;
	signal G18992: std_logic; attribute dont_touch of G18992: signal is true;
	signal G18993: std_logic; attribute dont_touch of G18993: signal is true;
	signal G18994: std_logic; attribute dont_touch of G18994: signal is true;
	signal G18995: std_logic; attribute dont_touch of G18995: signal is true;
	signal G18996: std_logic; attribute dont_touch of G18996: signal is true;
	signal G18997: std_logic; attribute dont_touch of G18997: signal is true;
	signal G18998: std_logic; attribute dont_touch of G18998: signal is true;
	signal G18999: std_logic; attribute dont_touch of G18999: signal is true;
	signal G19000: std_logic; attribute dont_touch of G19000: signal is true;
	signal G19001: std_logic; attribute dont_touch of G19001: signal is true;
	signal G19007: std_logic; attribute dont_touch of G19007: signal is true;
	signal G19008: std_logic; attribute dont_touch of G19008: signal is true;
	signal G19009: std_logic; attribute dont_touch of G19009: signal is true;
	signal G19010: std_logic; attribute dont_touch of G19010: signal is true;
	signal G19011: std_logic; attribute dont_touch of G19011: signal is true;
	signal G19012: std_logic; attribute dont_touch of G19012: signal is true;
	signal G19013: std_logic; attribute dont_touch of G19013: signal is true;
	signal G19014: std_logic; attribute dont_touch of G19014: signal is true;
	signal G19015: std_logic; attribute dont_touch of G19015: signal is true;
	signal G19016: std_logic; attribute dont_touch of G19016: signal is true;
	signal G19017: std_logic; attribute dont_touch of G19017: signal is true;
	signal G19018: std_logic; attribute dont_touch of G19018: signal is true;
	signal G19019: std_logic; attribute dont_touch of G19019: signal is true;
	signal G19020: std_logic; attribute dont_touch of G19020: signal is true;
	signal G19021: std_logic; attribute dont_touch of G19021: signal is true;
	signal G19022: std_logic; attribute dont_touch of G19022: signal is true;
	signal G19023: std_logic; attribute dont_touch of G19023: signal is true;
	signal G19024: std_logic; attribute dont_touch of G19024: signal is true;
	signal G19025: std_logic; attribute dont_touch of G19025: signal is true;
	signal G19026: std_logic; attribute dont_touch of G19026: signal is true;
	signal G19027: std_logic; attribute dont_touch of G19027: signal is true;
	signal G19028: std_logic; attribute dont_touch of G19028: signal is true;
	signal G19029: std_logic; attribute dont_touch of G19029: signal is true;
	signal G19030: std_logic; attribute dont_touch of G19030: signal is true;
	signal G19031: std_logic; attribute dont_touch of G19031: signal is true;
	signal G19032: std_logic; attribute dont_touch of G19032: signal is true;
	signal G19033: std_logic; attribute dont_touch of G19033: signal is true;
	signal G19034: std_logic; attribute dont_touch of G19034: signal is true;
	signal G19035: std_logic; attribute dont_touch of G19035: signal is true;
	signal G19036: std_logic; attribute dont_touch of G19036: signal is true;
	signal G19037: std_logic; attribute dont_touch of G19037: signal is true;
	signal G19038: std_logic; attribute dont_touch of G19038: signal is true;
	signal G19039: std_logic; attribute dont_touch of G19039: signal is true;
	signal G19040: std_logic; attribute dont_touch of G19040: signal is true;
	signal G19041: std_logic; attribute dont_touch of G19041: signal is true;
	signal G19042: std_logic; attribute dont_touch of G19042: signal is true;
	signal G19043: std_logic; attribute dont_touch of G19043: signal is true;
	signal G19044: std_logic; attribute dont_touch of G19044: signal is true;
	signal G19045: std_logic; attribute dont_touch of G19045: signal is true;
	signal G19046: std_logic; attribute dont_touch of G19046: signal is true;
	signal G19047: std_logic; attribute dont_touch of G19047: signal is true;
	signal G19048: std_logic; attribute dont_touch of G19048: signal is true;
	signal G19049: std_logic; attribute dont_touch of G19049: signal is true;
	signal G19050: std_logic; attribute dont_touch of G19050: signal is true;
	signal G19051: std_logic; attribute dont_touch of G19051: signal is true;
	signal G19052: std_logic; attribute dont_touch of G19052: signal is true;
	signal G19053: std_logic; attribute dont_touch of G19053: signal is true;
	signal G19054: std_logic; attribute dont_touch of G19054: signal is true;
	signal G19055: std_logic; attribute dont_touch of G19055: signal is true;
	signal G19056: std_logic; attribute dont_touch of G19056: signal is true;
	signal G19057: std_logic; attribute dont_touch of G19057: signal is true;
	signal G19058: std_logic; attribute dont_touch of G19058: signal is true;
	signal G19059: std_logic; attribute dont_touch of G19059: signal is true;
	signal G19060: std_logic; attribute dont_touch of G19060: signal is true;
	signal G19061: std_logic; attribute dont_touch of G19061: signal is true;
	signal G19062: std_logic; attribute dont_touch of G19062: signal is true;
	signal G19063: std_logic; attribute dont_touch of G19063: signal is true;
	signal G19064: std_logic; attribute dont_touch of G19064: signal is true;
	signal G19067: std_logic; attribute dont_touch of G19067: signal is true;
	signal G19070: std_logic; attribute dont_touch of G19070: signal is true;
	signal G19075: std_logic; attribute dont_touch of G19075: signal is true;
	signal G19078: std_logic; attribute dont_touch of G19078: signal is true;
	signal G19079: std_logic; attribute dont_touch of G19079: signal is true;
	signal G19080: std_logic; attribute dont_touch of G19080: signal is true;
	signal G19081: std_logic; attribute dont_touch of G19081: signal is true;
	signal G19084: std_logic; attribute dont_touch of G19084: signal is true;
	signal G19087: std_logic; attribute dont_touch of G19087: signal is true;
	signal G19088: std_logic; attribute dont_touch of G19088: signal is true;
	signal G19089: std_logic; attribute dont_touch of G19089: signal is true;
	signal G19090: std_logic; attribute dont_touch of G19090: signal is true;
	signal G19091: std_logic; attribute dont_touch of G19091: signal is true;
	signal G19092: std_logic; attribute dont_touch of G19092: signal is true;
	signal G19093: std_logic; attribute dont_touch of G19093: signal is true;
	signal G19094: std_logic; attribute dont_touch of G19094: signal is true;
	signal G19095: std_logic; attribute dont_touch of G19095: signal is true;
	signal G19096: std_logic; attribute dont_touch of G19096: signal is true;
	signal G19097: std_logic; attribute dont_touch of G19097: signal is true;
	signal G19098: std_logic; attribute dont_touch of G19098: signal is true;
	signal G19099: std_logic; attribute dont_touch of G19099: signal is true;
	signal G19100: std_logic; attribute dont_touch of G19100: signal is true;
	signal G19101: std_logic; attribute dont_touch of G19101: signal is true;
	signal G19102: std_logic; attribute dont_touch of G19102: signal is true;
	signal G19103: std_logic; attribute dont_touch of G19103: signal is true;
	signal G19104: std_logic; attribute dont_touch of G19104: signal is true;
	signal G19105: std_logic; attribute dont_touch of G19105: signal is true;
	signal G19106: std_logic; attribute dont_touch of G19106: signal is true;
	signal G19107: std_logic; attribute dont_touch of G19107: signal is true;
	signal G19108: std_logic; attribute dont_touch of G19108: signal is true;
	signal G19109: std_logic; attribute dont_touch of G19109: signal is true;
	signal G19110: std_logic; attribute dont_touch of G19110: signal is true;
	signal G19111: std_logic; attribute dont_touch of G19111: signal is true;
	signal G19112: std_logic; attribute dont_touch of G19112: signal is true;
	signal G19113: std_logic; attribute dont_touch of G19113: signal is true;
	signal G19116: std_logic; attribute dont_touch of G19116: signal is true;
	signal G19117: std_logic; attribute dont_touch of G19117: signal is true;
	signal G19118: std_logic; attribute dont_touch of G19118: signal is true;
	signal G19121: std_logic; attribute dont_touch of G19121: signal is true;
	signal G19124: std_logic; attribute dont_touch of G19124: signal is true;
	signal G19125: std_logic; attribute dont_touch of G19125: signal is true;
	signal G19128: std_logic; attribute dont_touch of G19128: signal is true;
	signal G19131: std_logic; attribute dont_touch of G19131: signal is true;
	signal G19132: std_logic; attribute dont_touch of G19132: signal is true;
	signal G19135: std_logic; attribute dont_touch of G19135: signal is true;
	signal G19138: std_logic; attribute dont_touch of G19138: signal is true;
	signal G19141: std_logic; attribute dont_touch of G19141: signal is true;
	signal G19142: std_logic; attribute dont_touch of G19142: signal is true;
	signal G19143: std_logic; attribute dont_touch of G19143: signal is true;
	signal G19144: std_logic; attribute dont_touch of G19144: signal is true;
	signal G19145: std_logic; attribute dont_touch of G19145: signal is true;
	signal G19146: std_logic; attribute dont_touch of G19146: signal is true;
	signal G19147: std_logic; attribute dont_touch of G19147: signal is true;
	signal G19148: std_logic; attribute dont_touch of G19148: signal is true;
	signal G19149: std_logic; attribute dont_touch of G19149: signal is true;
	signal G19150: std_logic; attribute dont_touch of G19150: signal is true;
	signal G19151: std_logic; attribute dont_touch of G19151: signal is true;
	signal G19152: std_logic; attribute dont_touch of G19152: signal is true;
	signal G19153: std_logic; attribute dont_touch of G19153: signal is true;
	signal G19154: std_logic; attribute dont_touch of G19154: signal is true;
	signal G19155: std_logic; attribute dont_touch of G19155: signal is true;
	signal G19156: std_logic; attribute dont_touch of G19156: signal is true;
	signal G19157: std_logic; attribute dont_touch of G19157: signal is true;
	signal G19158: std_logic; attribute dont_touch of G19158: signal is true;
	signal G19159: std_logic; attribute dont_touch of G19159: signal is true;
	signal G19160: std_logic; attribute dont_touch of G19160: signal is true;
	signal G19161: std_logic; attribute dont_touch of G19161: signal is true;
	signal G19162: std_logic; attribute dont_touch of G19162: signal is true;
	signal G19163: std_logic; attribute dont_touch of G19163: signal is true;
	signal G19164: std_logic; attribute dont_touch of G19164: signal is true;
	signal G19165: std_logic; attribute dont_touch of G19165: signal is true;
	signal G19166: std_logic; attribute dont_touch of G19166: signal is true;
	signal G19167: std_logic; attribute dont_touch of G19167: signal is true;
	signal G19168: std_logic; attribute dont_touch of G19168: signal is true;
	signal G19169: std_logic; attribute dont_touch of G19169: signal is true;
	signal G19170: std_logic; attribute dont_touch of G19170: signal is true;
	signal G19171: std_logic; attribute dont_touch of G19171: signal is true;
	signal G19172: std_logic; attribute dont_touch of G19172: signal is true;
	signal G19173: std_logic; attribute dont_touch of G19173: signal is true;
	signal G19174: std_logic; attribute dont_touch of G19174: signal is true;
	signal G19175: std_logic; attribute dont_touch of G19175: signal is true;
	signal G19176: std_logic; attribute dont_touch of G19176: signal is true;
	signal G19177: std_logic; attribute dont_touch of G19177: signal is true;
	signal G19178: std_logic; attribute dont_touch of G19178: signal is true;
	signal G19179: std_logic; attribute dont_touch of G19179: signal is true;
	signal G19180: std_logic; attribute dont_touch of G19180: signal is true;
	signal G19181: std_logic; attribute dont_touch of G19181: signal is true;
	signal G19182: std_logic; attribute dont_touch of G19182: signal is true;
	signal G19183: std_logic; attribute dont_touch of G19183: signal is true;
	signal G19184: std_logic; attribute dont_touch of G19184: signal is true;
	signal G19185: std_logic; attribute dont_touch of G19185: signal is true;
	signal G19186: std_logic; attribute dont_touch of G19186: signal is true;
	signal G19187: std_logic; attribute dont_touch of G19187: signal is true;
	signal G19188: std_logic; attribute dont_touch of G19188: signal is true;
	signal G19189: std_logic; attribute dont_touch of G19189: signal is true;
	signal G19190: std_logic; attribute dont_touch of G19190: signal is true;
	signal G19191: std_logic; attribute dont_touch of G19191: signal is true;
	signal G19192: std_logic; attribute dont_touch of G19192: signal is true;
	signal G19193: std_logic; attribute dont_touch of G19193: signal is true;
	signal G19194: std_logic; attribute dont_touch of G19194: signal is true;
	signal G19195: std_logic; attribute dont_touch of G19195: signal is true;
	signal G19196: std_logic; attribute dont_touch of G19196: signal is true;
	signal G19197: std_logic; attribute dont_touch of G19197: signal is true;
	signal G19198: std_logic; attribute dont_touch of G19198: signal is true;
	signal G19199: std_logic; attribute dont_touch of G19199: signal is true;
	signal G19200: std_logic; attribute dont_touch of G19200: signal is true;
	signal G19201: std_logic; attribute dont_touch of G19201: signal is true;
	signal G19202: std_logic; attribute dont_touch of G19202: signal is true;
	signal G19203: std_logic; attribute dont_touch of G19203: signal is true;
	signal G19204: std_logic; attribute dont_touch of G19204: signal is true;
	signal G19205: std_logic; attribute dont_touch of G19205: signal is true;
	signal G19206: std_logic; attribute dont_touch of G19206: signal is true;
	signal G19207: std_logic; attribute dont_touch of G19207: signal is true;
	signal G19208: std_logic; attribute dont_touch of G19208: signal is true;
	signal G19209: std_logic; attribute dont_touch of G19209: signal is true;
	signal G19210: std_logic; attribute dont_touch of G19210: signal is true;
	signal G19211: std_logic; attribute dont_touch of G19211: signal is true;
	signal G19212: std_logic; attribute dont_touch of G19212: signal is true;
	signal G19213: std_logic; attribute dont_touch of G19213: signal is true;
	signal G19214: std_logic; attribute dont_touch of G19214: signal is true;
	signal G19215: std_logic; attribute dont_touch of G19215: signal is true;
	signal G19216: std_logic; attribute dont_touch of G19216: signal is true;
	signal G19217: std_logic; attribute dont_touch of G19217: signal is true;
	signal G19218: std_logic; attribute dont_touch of G19218: signal is true;
	signal G19219: std_logic; attribute dont_touch of G19219: signal is true;
	signal G19220: std_logic; attribute dont_touch of G19220: signal is true;
	signal G19221: std_logic; attribute dont_touch of G19221: signal is true;
	signal G19222: std_logic; attribute dont_touch of G19222: signal is true;
	signal G19223: std_logic; attribute dont_touch of G19223: signal is true;
	signal G19224: std_logic; attribute dont_touch of G19224: signal is true;
	signal G19225: std_logic; attribute dont_touch of G19225: signal is true;
	signal G19226: std_logic; attribute dont_touch of G19226: signal is true;
	signal G19227: std_logic; attribute dont_touch of G19227: signal is true;
	signal G19228: std_logic; attribute dont_touch of G19228: signal is true;
	signal G19229: std_logic; attribute dont_touch of G19229: signal is true;
	signal G19230: std_logic; attribute dont_touch of G19230: signal is true;
	signal G19231: std_logic; attribute dont_touch of G19231: signal is true;
	signal G19232: std_logic; attribute dont_touch of G19232: signal is true;
	signal G19233: std_logic; attribute dont_touch of G19233: signal is true;
	signal G19234: std_logic; attribute dont_touch of G19234: signal is true;
	signal G19235: std_logic; attribute dont_touch of G19235: signal is true;
	signal G19236: std_logic; attribute dont_touch of G19236: signal is true;
	signal G19237: std_logic; attribute dont_touch of G19237: signal is true;
	signal G19238: std_logic; attribute dont_touch of G19238: signal is true;
	signal G19239: std_logic; attribute dont_touch of G19239: signal is true;
	signal G19240: std_logic; attribute dont_touch of G19240: signal is true;
	signal G19241: std_logic; attribute dont_touch of G19241: signal is true;
	signal G19242: std_logic; attribute dont_touch of G19242: signal is true;
	signal G19243: std_logic; attribute dont_touch of G19243: signal is true;
	signal G19244: std_logic; attribute dont_touch of G19244: signal is true;
	signal G19245: std_logic; attribute dont_touch of G19245: signal is true;
	signal G19246: std_logic; attribute dont_touch of G19246: signal is true;
	signal G19247: std_logic; attribute dont_touch of G19247: signal is true;
	signal G19248: std_logic; attribute dont_touch of G19248: signal is true;
	signal G19249: std_logic; attribute dont_touch of G19249: signal is true;
	signal G19250: std_logic; attribute dont_touch of G19250: signal is true;
	signal G19251: std_logic; attribute dont_touch of G19251: signal is true;
	signal G19252: std_logic; attribute dont_touch of G19252: signal is true;
	signal G19253: std_logic; attribute dont_touch of G19253: signal is true;
	signal G19254: std_logic; attribute dont_touch of G19254: signal is true;
	signal G19255: std_logic; attribute dont_touch of G19255: signal is true;
	signal G19256: std_logic; attribute dont_touch of G19256: signal is true;
	signal G19257: std_logic; attribute dont_touch of G19257: signal is true;
	signal G19258: std_logic; attribute dont_touch of G19258: signal is true;
	signal G19259: std_logic; attribute dont_touch of G19259: signal is true;
	signal G19260: std_logic; attribute dont_touch of G19260: signal is true;
	signal G19261: std_logic; attribute dont_touch of G19261: signal is true;
	signal G19262: std_logic; attribute dont_touch of G19262: signal is true;
	signal G19263: std_logic; attribute dont_touch of G19263: signal is true;
	signal G19264: std_logic; attribute dont_touch of G19264: signal is true;
	signal G19265: std_logic; attribute dont_touch of G19265: signal is true;
	signal G19266: std_logic; attribute dont_touch of G19266: signal is true;
	signal G19267: std_logic; attribute dont_touch of G19267: signal is true;
	signal G19268: std_logic; attribute dont_touch of G19268: signal is true;
	signal G19269: std_logic; attribute dont_touch of G19269: signal is true;
	signal G19270: std_logic; attribute dont_touch of G19270: signal is true;
	signal G19271: std_logic; attribute dont_touch of G19271: signal is true;
	signal G19272: std_logic; attribute dont_touch of G19272: signal is true;
	signal G19275: std_logic; attribute dont_touch of G19275: signal is true;
	signal G19276: std_logic; attribute dont_touch of G19276: signal is true;
	signal G19277: std_logic; attribute dont_touch of G19277: signal is true;
	signal G19278: std_logic; attribute dont_touch of G19278: signal is true;
	signal G19279: std_logic; attribute dont_touch of G19279: signal is true;
	signal G19280: std_logic; attribute dont_touch of G19280: signal is true;
	signal G19281: std_logic; attribute dont_touch of G19281: signal is true;
	signal G19282: std_logic; attribute dont_touch of G19282: signal is true;
	signal G19283: std_logic; attribute dont_touch of G19283: signal is true;
	signal G19284: std_logic; attribute dont_touch of G19284: signal is true;
	signal G19285: std_logic; attribute dont_touch of G19285: signal is true;
	signal G19286: std_logic; attribute dont_touch of G19286: signal is true;
	signal G19287: std_logic; attribute dont_touch of G19287: signal is true;
	signal G19288: std_logic; attribute dont_touch of G19288: signal is true;
	signal G19289: std_logic; attribute dont_touch of G19289: signal is true;
	signal G19290: std_logic; attribute dont_touch of G19290: signal is true;
	signal G19291: std_logic; attribute dont_touch of G19291: signal is true;
	signal G19294: std_logic; attribute dont_touch of G19294: signal is true;
	signal G19295: std_logic; attribute dont_touch of G19295: signal is true;
	signal G19296: std_logic; attribute dont_touch of G19296: signal is true;
	signal G19297: std_logic; attribute dont_touch of G19297: signal is true;
	signal G19298: std_logic; attribute dont_touch of G19298: signal is true;
	signal G19299: std_logic; attribute dont_touch of G19299: signal is true;
	signal G19300: std_logic; attribute dont_touch of G19300: signal is true;
	signal G19301: std_logic; attribute dont_touch of G19301: signal is true;
	signal G19302: std_logic; attribute dont_touch of G19302: signal is true;
	signal G19303: std_logic; attribute dont_touch of G19303: signal is true;
	signal G19304: std_logic; attribute dont_touch of G19304: signal is true;
	signal G19305: std_logic; attribute dont_touch of G19305: signal is true;
	signal G19306: std_logic; attribute dont_touch of G19306: signal is true;
	signal G19307: std_logic; attribute dont_touch of G19307: signal is true;
	signal G19308: std_logic; attribute dont_touch of G19308: signal is true;
	signal G19309: std_logic; attribute dont_touch of G19309: signal is true;
	signal G19312: std_logic; attribute dont_touch of G19312: signal is true;
	signal G19313: std_logic; attribute dont_touch of G19313: signal is true;
	signal G19314: std_logic; attribute dont_touch of G19314: signal is true;
	signal G19315: std_logic; attribute dont_touch of G19315: signal is true;
	signal G19316: std_logic; attribute dont_touch of G19316: signal is true;
	signal G19317: std_logic; attribute dont_touch of G19317: signal is true;
	signal G19318: std_logic; attribute dont_touch of G19318: signal is true;
	signal G19319: std_logic; attribute dont_touch of G19319: signal is true;
	signal G19320: std_logic; attribute dont_touch of G19320: signal is true;
	signal G19321: std_logic; attribute dont_touch of G19321: signal is true;
	signal G19322: std_logic; attribute dont_touch of G19322: signal is true;
	signal G19323: std_logic; attribute dont_touch of G19323: signal is true;
	signal G19324: std_logic; attribute dont_touch of G19324: signal is true;
	signal G19325: std_logic; attribute dont_touch of G19325: signal is true;
	signal G19326: std_logic; attribute dont_touch of G19326: signal is true;
	signal G19327: std_logic; attribute dont_touch of G19327: signal is true;
	signal G19328: std_logic; attribute dont_touch of G19328: signal is true;
	signal G19329: std_logic; attribute dont_touch of G19329: signal is true;
	signal G19330: std_logic; attribute dont_touch of G19330: signal is true;
	signal G19333: std_logic; attribute dont_touch of G19333: signal is true;
	signal G19334: std_logic; attribute dont_touch of G19334: signal is true;
	signal G19335: std_logic; attribute dont_touch of G19335: signal is true;
	signal G19345: std_logic; attribute dont_touch of G19345: signal is true;
	signal G19346: std_logic; attribute dont_touch of G19346: signal is true;
	signal G19347: std_logic; attribute dont_touch of G19347: signal is true;
	signal G19348: std_logic; attribute dont_touch of G19348: signal is true;
	signal G19349: std_logic; attribute dont_touch of G19349: signal is true;
	signal G19350: std_logic; attribute dont_touch of G19350: signal is true;
	signal G19351: std_logic; attribute dont_touch of G19351: signal is true;
	signal G19352: std_logic; attribute dont_touch of G19352: signal is true;
	signal G19353: std_logic; attribute dont_touch of G19353: signal is true;
	signal G19354: std_logic; attribute dont_touch of G19354: signal is true;
	signal G19355: std_logic; attribute dont_touch of G19355: signal is true;
	signal G19356: std_logic; attribute dont_touch of G19356: signal is true;
	signal G19357: std_logic; attribute dont_touch of G19357: signal is true;
	signal G19358: std_logic; attribute dont_touch of G19358: signal is true;
	signal G19368: std_logic; attribute dont_touch of G19368: signal is true;
	signal G19369: std_logic; attribute dont_touch of G19369: signal is true;
	signal G19379: std_logic; attribute dont_touch of G19379: signal is true;
	signal G19380: std_logic; attribute dont_touch of G19380: signal is true;
	signal G19381: std_logic; attribute dont_touch of G19381: signal is true;
	signal G19382: std_logic; attribute dont_touch of G19382: signal is true;
	signal G19383: std_logic; attribute dont_touch of G19383: signal is true;
	signal G19384: std_logic; attribute dont_touch of G19384: signal is true;
	signal G19385: std_logic; attribute dont_touch of G19385: signal is true;
	signal G19386: std_logic; attribute dont_touch of G19386: signal is true;
	signal G19387: std_logic; attribute dont_touch of G19387: signal is true;
	signal G19388: std_logic; attribute dont_touch of G19388: signal is true;
	signal G19389: std_logic; attribute dont_touch of G19389: signal is true;
	signal G19390: std_logic; attribute dont_touch of G19390: signal is true;
	signal G19400: std_logic; attribute dont_touch of G19400: signal is true;
	signal G19401: std_logic; attribute dont_touch of G19401: signal is true;
	signal G19411: std_logic; attribute dont_touch of G19411: signal is true;
	signal G19412: std_logic; attribute dont_touch of G19412: signal is true;
	signal G19413: std_logic; attribute dont_touch of G19413: signal is true;
	signal G19414: std_logic; attribute dont_touch of G19414: signal is true;
	signal G19415: std_logic; attribute dont_touch of G19415: signal is true;
	signal G19416: std_logic; attribute dont_touch of G19416: signal is true;
	signal G19417: std_logic; attribute dont_touch of G19417: signal is true;
	signal G19418: std_logic; attribute dont_touch of G19418: signal is true;
	signal G19419: std_logic; attribute dont_touch of G19419: signal is true;
	signal G19420: std_logic; attribute dont_touch of G19420: signal is true;
	signal G19430: std_logic; attribute dont_touch of G19430: signal is true;
	signal G19431: std_logic; attribute dont_touch of G19431: signal is true;
	signal G19441: std_logic; attribute dont_touch of G19441: signal is true;
	signal G19444: std_logic; attribute dont_touch of G19444: signal is true;
	signal G19448: std_logic; attribute dont_touch of G19448: signal is true;
	signal G19449: std_logic; attribute dont_touch of G19449: signal is true;
	signal G19450: std_logic; attribute dont_touch of G19450: signal is true;
	signal G19451: std_logic; attribute dont_touch of G19451: signal is true;
	signal G19452: std_logic; attribute dont_touch of G19452: signal is true;
	signal G19453: std_logic; attribute dont_touch of G19453: signal is true;
	signal G19454: std_logic; attribute dont_touch of G19454: signal is true;
	signal G19455: std_logic; attribute dont_touch of G19455: signal is true;
	signal G19456: std_logic; attribute dont_touch of G19456: signal is true;
	signal G19457: std_logic; attribute dont_touch of G19457: signal is true;
	signal G19467: std_logic; attribute dont_touch of G19467: signal is true;
	signal G19468: std_logic; attribute dont_touch of G19468: signal is true;
	signal G19471: std_logic; attribute dont_touch of G19471: signal is true;
	signal G19475: std_logic; attribute dont_touch of G19475: signal is true;
	signal G19476: std_logic; attribute dont_touch of G19476: signal is true;
	signal G19477: std_logic; attribute dont_touch of G19477: signal is true;
	signal G19478: std_logic; attribute dont_touch of G19478: signal is true;
	signal G19479: std_logic; attribute dont_touch of G19479: signal is true;
	signal G19480: std_logic; attribute dont_touch of G19480: signal is true;
	signal G19481: std_logic; attribute dont_touch of G19481: signal is true;
	signal G19482: std_logic; attribute dont_touch of G19482: signal is true;
	signal G19483: std_logic; attribute dont_touch of G19483: signal is true;
	signal G19484: std_logic; attribute dont_touch of G19484: signal is true;
	signal G19490: std_logic; attribute dont_touch of G19490: signal is true;
	signal G19491: std_logic; attribute dont_touch of G19491: signal is true;
	signal G19494: std_logic; attribute dont_touch of G19494: signal is true;
	signal G19498: std_logic; attribute dont_touch of G19498: signal is true;
	signal G19499: std_logic; attribute dont_touch of G19499: signal is true;
	signal G19500: std_logic; attribute dont_touch of G19500: signal is true;
	signal G19501: std_logic; attribute dont_touch of G19501: signal is true;
	signal G19502: std_logic; attribute dont_touch of G19502: signal is true;
	signal G19503: std_logic; attribute dont_touch of G19503: signal is true;
	signal G19504: std_logic; attribute dont_touch of G19504: signal is true;
	signal G19505: std_logic; attribute dont_touch of G19505: signal is true;
	signal G19511: std_logic; attribute dont_touch of G19511: signal is true;
	signal G19512: std_logic; attribute dont_touch of G19512: signal is true;
	signal G19515: std_logic; attribute dont_touch of G19515: signal is true;
	signal G19519: std_logic; attribute dont_touch of G19519: signal is true;
	signal G19520: std_logic; attribute dont_touch of G19520: signal is true;
	signal G19521: std_logic; attribute dont_touch of G19521: signal is true;
	signal G19522: std_logic; attribute dont_touch of G19522: signal is true;
	signal G19523: std_logic; attribute dont_touch of G19523: signal is true;
	signal G19524: std_logic; attribute dont_touch of G19524: signal is true;
	signal G19530: std_logic; attribute dont_touch of G19530: signal is true;
	signal G19531: std_logic; attribute dont_touch of G19531: signal is true;
	signal G19532: std_logic; attribute dont_touch of G19532: signal is true;
	signal G19533: std_logic; attribute dont_touch of G19533: signal is true;
	signal G19534: std_logic; attribute dont_touch of G19534: signal is true;
	signal G19540: std_logic; attribute dont_touch of G19540: signal is true;
	signal G19541: std_logic; attribute dont_touch of G19541: signal is true;
	signal G19542: std_logic; attribute dont_touch of G19542: signal is true;
	signal G19543: std_logic; attribute dont_touch of G19543: signal is true;
	signal G19544: std_logic; attribute dont_touch of G19544: signal is true;
	signal G19545: std_logic; attribute dont_touch of G19545: signal is true;
	signal G19546: std_logic; attribute dont_touch of G19546: signal is true;
	signal G19547: std_logic; attribute dont_touch of G19547: signal is true;
	signal G19548: std_logic; attribute dont_touch of G19548: signal is true;
	signal G19549: std_logic; attribute dont_touch of G19549: signal is true;
	signal G19550: std_logic; attribute dont_touch of G19550: signal is true;
	signal G19551: std_logic; attribute dont_touch of G19551: signal is true;
	signal G19552: std_logic; attribute dont_touch of G19552: signal is true;
	signal G19553: std_logic; attribute dont_touch of G19553: signal is true;
	signal G19554: std_logic; attribute dont_touch of G19554: signal is true;
	signal G19555: std_logic; attribute dont_touch of G19555: signal is true;
	signal G19556: std_logic; attribute dont_touch of G19556: signal is true;
	signal G19557: std_logic; attribute dont_touch of G19557: signal is true;
	signal G19558: std_logic; attribute dont_touch of G19558: signal is true;
	signal G19559: std_logic; attribute dont_touch of G19559: signal is true;
	signal G19560: std_logic; attribute dont_touch of G19560: signal is true;
	signal G19561: std_logic; attribute dont_touch of G19561: signal is true;
	signal G19562: std_logic; attribute dont_touch of G19562: signal is true;
	signal G19563: std_logic; attribute dont_touch of G19563: signal is true;
	signal G19564: std_logic; attribute dont_touch of G19564: signal is true;
	signal G19565: std_logic; attribute dont_touch of G19565: signal is true;
	signal G19566: std_logic; attribute dont_touch of G19566: signal is true;
	signal G19567: std_logic; attribute dont_touch of G19567: signal is true;
	signal G19568: std_logic; attribute dont_touch of G19568: signal is true;
	signal G19569: std_logic; attribute dont_touch of G19569: signal is true;
	signal G19570: std_logic; attribute dont_touch of G19570: signal is true;
	signal G19571: std_logic; attribute dont_touch of G19571: signal is true;
	signal G19572: std_logic; attribute dont_touch of G19572: signal is true;
	signal G19573: std_logic; attribute dont_touch of G19573: signal is true;
	signal G19574: std_logic; attribute dont_touch of G19574: signal is true;
	signal G19575: std_logic; attribute dont_touch of G19575: signal is true;
	signal G19576: std_logic; attribute dont_touch of G19576: signal is true;
	signal G19577: std_logic; attribute dont_touch of G19577: signal is true;
	signal G19578: std_logic; attribute dont_touch of G19578: signal is true;
	signal G19584: std_logic; attribute dont_touch of G19584: signal is true;
	signal G19585: std_logic; attribute dont_touch of G19585: signal is true;
	signal G19586: std_logic; attribute dont_touch of G19586: signal is true;
	signal G19587: std_logic; attribute dont_touch of G19587: signal is true;
	signal G19588: std_logic; attribute dont_touch of G19588: signal is true;
	signal G19589: std_logic; attribute dont_touch of G19589: signal is true;
	signal G19590: std_logic; attribute dont_touch of G19590: signal is true;
	signal G19591: std_logic; attribute dont_touch of G19591: signal is true;
	signal G19592: std_logic; attribute dont_touch of G19592: signal is true;
	signal G19593: std_logic; attribute dont_touch of G19593: signal is true;
	signal G19594: std_logic; attribute dont_touch of G19594: signal is true;
	signal G19595: std_logic; attribute dont_touch of G19595: signal is true;
	signal G19596: std_logic; attribute dont_touch of G19596: signal is true;
	signal G19597: std_logic; attribute dont_touch of G19597: signal is true;
	signal G19598: std_logic; attribute dont_touch of G19598: signal is true;
	signal G19599: std_logic; attribute dont_touch of G19599: signal is true;
	signal G19600: std_logic; attribute dont_touch of G19600: signal is true;
	signal G19601: std_logic; attribute dont_touch of G19601: signal is true;
	signal G19602: std_logic; attribute dont_touch of G19602: signal is true;
	signal G19603: std_logic; attribute dont_touch of G19603: signal is true;
	signal G19604: std_logic; attribute dont_touch of G19604: signal is true;
	signal G19605: std_logic; attribute dont_touch of G19605: signal is true;
	signal G19606: std_logic; attribute dont_touch of G19606: signal is true;
	signal G19607: std_logic; attribute dont_touch of G19607: signal is true;
	signal G19608: std_logic; attribute dont_touch of G19608: signal is true;
	signal G19614: std_logic; attribute dont_touch of G19614: signal is true;
	signal G19615: std_logic; attribute dont_touch of G19615: signal is true;
	signal G19616: std_logic; attribute dont_touch of G19616: signal is true;
	signal G19617: std_logic; attribute dont_touch of G19617: signal is true;
	signal G19618: std_logic; attribute dont_touch of G19618: signal is true;
	signal G19619: std_logic; attribute dont_touch of G19619: signal is true;
	signal G19620: std_logic; attribute dont_touch of G19620: signal is true;
	signal G19621: std_logic; attribute dont_touch of G19621: signal is true;
	signal G19622: std_logic; attribute dont_touch of G19622: signal is true;
	signal G19623: std_logic; attribute dont_touch of G19623: signal is true;
	signal G19624: std_logic; attribute dont_touch of G19624: signal is true;
	signal G19625: std_logic; attribute dont_touch of G19625: signal is true;
	signal G19626: std_logic; attribute dont_touch of G19626: signal is true;
	signal G19627: std_logic; attribute dont_touch of G19627: signal is true;
	signal G19628: std_logic; attribute dont_touch of G19628: signal is true;
	signal G19629: std_logic; attribute dont_touch of G19629: signal is true;
	signal G19630: std_logic; attribute dont_touch of G19630: signal is true;
	signal G19631: std_logic; attribute dont_touch of G19631: signal is true;
	signal G19632: std_logic; attribute dont_touch of G19632: signal is true;
	signal G19633: std_logic; attribute dont_touch of G19633: signal is true;
	signal G19634: std_logic; attribute dont_touch of G19634: signal is true;
	signal G19635: std_logic; attribute dont_touch of G19635: signal is true;
	signal G19636: std_logic; attribute dont_touch of G19636: signal is true;
	signal G19637: std_logic; attribute dont_touch of G19637: signal is true;
	signal G19638: std_logic; attribute dont_touch of G19638: signal is true;
	signal G19639: std_logic; attribute dont_touch of G19639: signal is true;
	signal G19640: std_logic; attribute dont_touch of G19640: signal is true;
	signal G19641: std_logic; attribute dont_touch of G19641: signal is true;
	signal G19647: std_logic; attribute dont_touch of G19647: signal is true;
	signal G19648: std_logic; attribute dont_touch of G19648: signal is true;
	signal G19649: std_logic; attribute dont_touch of G19649: signal is true;
	signal G19650: std_logic; attribute dont_touch of G19650: signal is true;
	signal G19651: std_logic; attribute dont_touch of G19651: signal is true;
	signal G19652: std_logic; attribute dont_touch of G19652: signal is true;
	signal G19653: std_logic; attribute dont_touch of G19653: signal is true;
	signal G19654: std_logic; attribute dont_touch of G19654: signal is true;
	signal G19655: std_logic; attribute dont_touch of G19655: signal is true;
	signal G19656: std_logic; attribute dont_touch of G19656: signal is true;
	signal G19657: std_logic; attribute dont_touch of G19657: signal is true;
	signal G19660: std_logic; attribute dont_touch of G19660: signal is true;
	signal G19661: std_logic; attribute dont_touch of G19661: signal is true;
	signal G19662: std_logic; attribute dont_touch of G19662: signal is true;
	signal G19663: std_logic; attribute dont_touch of G19663: signal is true;
	signal G19664: std_logic; attribute dont_touch of G19664: signal is true;
	signal G19665: std_logic; attribute dont_touch of G19665: signal is true;
	signal G19666: std_logic; attribute dont_touch of G19666: signal is true;
	signal G19667: std_logic; attribute dont_touch of G19667: signal is true;
	signal G19668: std_logic; attribute dont_touch of G19668: signal is true;
	signal G19669: std_logic; attribute dont_touch of G19669: signal is true;
	signal G19670: std_logic; attribute dont_touch of G19670: signal is true;
	signal G19671: std_logic; attribute dont_touch of G19671: signal is true;
	signal G19672: std_logic; attribute dont_touch of G19672: signal is true;
	signal G19673: std_logic; attribute dont_touch of G19673: signal is true;
	signal G19674: std_logic; attribute dont_touch of G19674: signal is true;
	signal G19675: std_logic; attribute dont_touch of G19675: signal is true;
	signal G19676: std_logic; attribute dont_touch of G19676: signal is true;
	signal G19677: std_logic; attribute dont_touch of G19677: signal is true;
	signal G19678: std_logic; attribute dont_touch of G19678: signal is true;
	signal G19679: std_logic; attribute dont_touch of G19679: signal is true;
	signal G19680: std_logic; attribute dont_touch of G19680: signal is true;
	signal G19681: std_logic; attribute dont_touch of G19681: signal is true;
	signal G19687: std_logic; attribute dont_touch of G19687: signal is true;
	signal G19688: std_logic; attribute dont_touch of G19688: signal is true;
	signal G19689: std_logic; attribute dont_touch of G19689: signal is true;
	signal G19690: std_logic; attribute dont_touch of G19690: signal is true;
	signal G19691: std_logic; attribute dont_touch of G19691: signal is true;
	signal G19692: std_logic; attribute dont_touch of G19692: signal is true;
	signal G19693: std_logic; attribute dont_touch of G19693: signal is true;
	signal G19694: std_logic; attribute dont_touch of G19694: signal is true;
	signal G19695: std_logic; attribute dont_touch of G19695: signal is true;
	signal G19696: std_logic; attribute dont_touch of G19696: signal is true;
	signal G19697: std_logic; attribute dont_touch of G19697: signal is true;
	signal G19698: std_logic; attribute dont_touch of G19698: signal is true;
	signal G19699: std_logic; attribute dont_touch of G19699: signal is true;
	signal G19700: std_logic; attribute dont_touch of G19700: signal is true;
	signal G19701: std_logic; attribute dont_touch of G19701: signal is true;
	signal G19702: std_logic; attribute dont_touch of G19702: signal is true;
	signal G19703: std_logic; attribute dont_touch of G19703: signal is true;
	signal G19704: std_logic; attribute dont_touch of G19704: signal is true;
	signal G19705: std_logic; attribute dont_touch of G19705: signal is true;
	signal G19708: std_logic; attribute dont_touch of G19708: signal is true;
	signal G19709: std_logic; attribute dont_touch of G19709: signal is true;
	signal G19710: std_logic; attribute dont_touch of G19710: signal is true;
	signal G19711: std_logic; attribute dont_touch of G19711: signal is true;
	signal G19712: std_logic; attribute dont_touch of G19712: signal is true;
	signal G19713: std_logic; attribute dont_touch of G19713: signal is true;
	signal G19714: std_logic; attribute dont_touch of G19714: signal is true;
	signal G19715: std_logic; attribute dont_touch of G19715: signal is true;
	signal G19716: std_logic; attribute dont_touch of G19716: signal is true;
	signal G19717: std_logic; attribute dont_touch of G19717: signal is true;
	signal G19718: std_logic; attribute dont_touch of G19718: signal is true;
	signal G19719: std_logic; attribute dont_touch of G19719: signal is true;
	signal G19720: std_logic; attribute dont_touch of G19720: signal is true;
	signal G19721: std_logic; attribute dont_touch of G19721: signal is true;
	signal G19722: std_logic; attribute dont_touch of G19722: signal is true;
	signal G19723: std_logic; attribute dont_touch of G19723: signal is true;
	signal G19724: std_logic; attribute dont_touch of G19724: signal is true;
	signal G19725: std_logic; attribute dont_touch of G19725: signal is true;
	signal G19726: std_logic; attribute dont_touch of G19726: signal is true;
	signal G19727: std_logic; attribute dont_touch of G19727: signal is true;
	signal G19728: std_logic; attribute dont_touch of G19728: signal is true;
	signal G19729: std_logic; attribute dont_touch of G19729: signal is true;
	signal G19730: std_logic; attribute dont_touch of G19730: signal is true;
	signal G19731: std_logic; attribute dont_touch of G19731: signal is true;
	signal G19732: std_logic; attribute dont_touch of G19732: signal is true;
	signal G19733: std_logic; attribute dont_touch of G19733: signal is true;
	signal G19734: std_logic; attribute dont_touch of G19734: signal is true;
	signal G19735: std_logic; attribute dont_touch of G19735: signal is true;
	signal G19736: std_logic; attribute dont_touch of G19736: signal is true;
	signal G19737: std_logic; attribute dont_touch of G19737: signal is true;
	signal G19738: std_logic; attribute dont_touch of G19738: signal is true;
	signal G19739: std_logic; attribute dont_touch of G19739: signal is true;
	signal G19740: std_logic; attribute dont_touch of G19740: signal is true;
	signal G19741: std_logic; attribute dont_touch of G19741: signal is true;
	signal G19742: std_logic; attribute dont_touch of G19742: signal is true;
	signal G19743: std_logic; attribute dont_touch of G19743: signal is true;
	signal G19744: std_logic; attribute dont_touch of G19744: signal is true;
	signal G19745: std_logic; attribute dont_touch of G19745: signal is true;
	signal G19746: std_logic; attribute dont_touch of G19746: signal is true;
	signal G19747: std_logic; attribute dont_touch of G19747: signal is true;
	signal G19748: std_logic; attribute dont_touch of G19748: signal is true;
	signal G19749: std_logic; attribute dont_touch of G19749: signal is true;
	signal G19752: std_logic; attribute dont_touch of G19752: signal is true;
	signal G19753: std_logic; attribute dont_touch of G19753: signal is true;
	signal G19754: std_logic; attribute dont_touch of G19754: signal is true;
	signal G19755: std_logic; attribute dont_touch of G19755: signal is true;
	signal G19756: std_logic; attribute dont_touch of G19756: signal is true;
	signal G19757: std_logic; attribute dont_touch of G19757: signal is true;
	signal G19758: std_logic; attribute dont_touch of G19758: signal is true;
	signal G19759: std_logic; attribute dont_touch of G19759: signal is true;
	signal G19760: std_logic; attribute dont_touch of G19760: signal is true;
	signal G19761: std_logic; attribute dont_touch of G19761: signal is true;
	signal G19762: std_logic; attribute dont_touch of G19762: signal is true;
	signal G19763: std_logic; attribute dont_touch of G19763: signal is true;
	signal G19764: std_logic; attribute dont_touch of G19764: signal is true;
	signal G19765: std_logic; attribute dont_touch of G19765: signal is true;
	signal G19766: std_logic; attribute dont_touch of G19766: signal is true;
	signal G19767: std_logic; attribute dont_touch of G19767: signal is true;
	signal G19768: std_logic; attribute dont_touch of G19768: signal is true;
	signal G19769: std_logic; attribute dont_touch of G19769: signal is true;
	signal G19770: std_logic; attribute dont_touch of G19770: signal is true;
	signal G19771: std_logic; attribute dont_touch of G19771: signal is true;
	signal G19772: std_logic; attribute dont_touch of G19772: signal is true;
	signal G19773: std_logic; attribute dont_touch of G19773: signal is true;
	signal G19774: std_logic; attribute dont_touch of G19774: signal is true;
	signal G19775: std_logic; attribute dont_touch of G19775: signal is true;
	signal G19776: std_logic; attribute dont_touch of G19776: signal is true;
	signal G19777: std_logic; attribute dont_touch of G19777: signal is true;
	signal G19778: std_logic; attribute dont_touch of G19778: signal is true;
	signal G19779: std_logic; attribute dont_touch of G19779: signal is true;
	signal G19780: std_logic; attribute dont_touch of G19780: signal is true;
	signal G19781: std_logic; attribute dont_touch of G19781: signal is true;
	signal G19782: std_logic; attribute dont_touch of G19782: signal is true;
	signal G19783: std_logic; attribute dont_touch of G19783: signal is true;
	signal G19784: std_logic; attribute dont_touch of G19784: signal is true;
	signal G19785: std_logic; attribute dont_touch of G19785: signal is true;
	signal G19786: std_logic; attribute dont_touch of G19786: signal is true;
	signal G19787: std_logic; attribute dont_touch of G19787: signal is true;
	signal G19788: std_logic; attribute dont_touch of G19788: signal is true;
	signal G19789: std_logic; attribute dont_touch of G19789: signal is true;
	signal G19790: std_logic; attribute dont_touch of G19790: signal is true;
	signal G19791: std_logic; attribute dont_touch of G19791: signal is true;
	signal G19792: std_logic; attribute dont_touch of G19792: signal is true;
	signal G19795: std_logic; attribute dont_touch of G19795: signal is true;
	signal G19796: std_logic; attribute dont_touch of G19796: signal is true;
	signal G19797: std_logic; attribute dont_touch of G19797: signal is true;
	signal G19798: std_logic; attribute dont_touch of G19798: signal is true;
	signal G19799: std_logic; attribute dont_touch of G19799: signal is true;
	signal G19802: std_logic; attribute dont_touch of G19802: signal is true;
	signal G19803: std_logic; attribute dont_touch of G19803: signal is true;
	signal G19804: std_logic; attribute dont_touch of G19804: signal is true;
	signal G19805: std_logic; attribute dont_touch of G19805: signal is true;
	signal G19806: std_logic; attribute dont_touch of G19806: signal is true;
	signal G19807: std_logic; attribute dont_touch of G19807: signal is true;
	signal G19808: std_logic; attribute dont_touch of G19808: signal is true;
	signal G19809: std_logic; attribute dont_touch of G19809: signal is true;
	signal G19810: std_logic; attribute dont_touch of G19810: signal is true;
	signal G19811: std_logic; attribute dont_touch of G19811: signal is true;
	signal G19812: std_logic; attribute dont_touch of G19812: signal is true;
	signal G19813: std_logic; attribute dont_touch of G19813: signal is true;
	signal G19814: std_logic; attribute dont_touch of G19814: signal is true;
	signal G19815: std_logic; attribute dont_touch of G19815: signal is true;
	signal G19816: std_logic; attribute dont_touch of G19816: signal is true;
	signal G19817: std_logic; attribute dont_touch of G19817: signal is true;
	signal G19818: std_logic; attribute dont_touch of G19818: signal is true;
	signal G19819: std_logic; attribute dont_touch of G19819: signal is true;
	signal G19820: std_logic; attribute dont_touch of G19820: signal is true;
	signal G19821: std_logic; attribute dont_touch of G19821: signal is true;
	signal G19822: std_logic; attribute dont_touch of G19822: signal is true;
	signal G19823: std_logic; attribute dont_touch of G19823: signal is true;
	signal G19824: std_logic; attribute dont_touch of G19824: signal is true;
	signal G19825: std_logic; attribute dont_touch of G19825: signal is true;
	signal G19826: std_logic; attribute dont_touch of G19826: signal is true;
	signal G19827: std_logic; attribute dont_touch of G19827: signal is true;
	signal G19828: std_logic; attribute dont_touch of G19828: signal is true;
	signal G19829: std_logic; attribute dont_touch of G19829: signal is true;
	signal G19830: std_logic; attribute dont_touch of G19830: signal is true;
	signal G19836: std_logic; attribute dont_touch of G19836: signal is true;
	signal G19837: std_logic; attribute dont_touch of G19837: signal is true;
	signal G19838: std_logic; attribute dont_touch of G19838: signal is true;
	signal G19839: std_logic; attribute dont_touch of G19839: signal is true;
	signal G19840: std_logic; attribute dont_touch of G19840: signal is true;
	signal G19841: std_logic; attribute dont_touch of G19841: signal is true;
	signal G19842: std_logic; attribute dont_touch of G19842: signal is true;
	signal G19843: std_logic; attribute dont_touch of G19843: signal is true;
	signal G19846: std_logic; attribute dont_touch of G19846: signal is true;
	signal G19847: std_logic; attribute dont_touch of G19847: signal is true;
	signal G19848: std_logic; attribute dont_touch of G19848: signal is true;
	signal G19849: std_logic; attribute dont_touch of G19849: signal is true;
	signal G19850: std_logic; attribute dont_touch of G19850: signal is true;
	signal G19851: std_logic; attribute dont_touch of G19851: signal is true;
	signal G19852: std_logic; attribute dont_touch of G19852: signal is true;
	signal G19853: std_logic; attribute dont_touch of G19853: signal is true;
	signal G19854: std_logic; attribute dont_touch of G19854: signal is true;
	signal G19855: std_logic; attribute dont_touch of G19855: signal is true;
	signal G19856: std_logic; attribute dont_touch of G19856: signal is true;
	signal G19857: std_logic; attribute dont_touch of G19857: signal is true;
	signal G19858: std_logic; attribute dont_touch of G19858: signal is true;
	signal G19859: std_logic; attribute dont_touch of G19859: signal is true;
	signal G19860: std_logic; attribute dont_touch of G19860: signal is true;
	signal G19861: std_logic; attribute dont_touch of G19861: signal is true;
	signal G19862: std_logic; attribute dont_touch of G19862: signal is true;
	signal G19863: std_logic; attribute dont_touch of G19863: signal is true;
	signal G19864: std_logic; attribute dont_touch of G19864: signal is true;
	signal G19865: std_logic; attribute dont_touch of G19865: signal is true;
	signal G19868: std_logic; attribute dont_touch of G19868: signal is true;
	signal G19869: std_logic; attribute dont_touch of G19869: signal is true;
	signal G19870: std_logic; attribute dont_touch of G19870: signal is true;
	signal G19871: std_logic; attribute dont_touch of G19871: signal is true;
	signal G19872: std_logic; attribute dont_touch of G19872: signal is true;
	signal G19873: std_logic; attribute dont_touch of G19873: signal is true;
	signal G19874: std_logic; attribute dont_touch of G19874: signal is true;
	signal G19875: std_logic; attribute dont_touch of G19875: signal is true;
	signal G19876: std_logic; attribute dont_touch of G19876: signal is true;
	signal G19879: std_logic; attribute dont_touch of G19879: signal is true;
	signal G19880: std_logic; attribute dont_touch of G19880: signal is true;
	signal G19881: std_logic; attribute dont_touch of G19881: signal is true;
	signal G19882: std_logic; attribute dont_touch of G19882: signal is true;
	signal G19883: std_logic; attribute dont_touch of G19883: signal is true;
	signal G19884: std_logic; attribute dont_touch of G19884: signal is true;
	signal G19885: std_logic; attribute dont_touch of G19885: signal is true;
	signal G19886: std_logic; attribute dont_touch of G19886: signal is true;
	signal G19887: std_logic; attribute dont_touch of G19887: signal is true;
	signal G19888: std_logic; attribute dont_touch of G19888: signal is true;
	signal G19889: std_logic; attribute dont_touch of G19889: signal is true;
	signal G19890: std_logic; attribute dont_touch of G19890: signal is true;
	signal G19893: std_logic; attribute dont_touch of G19893: signal is true;
	signal G19894: std_logic; attribute dont_touch of G19894: signal is true;
	signal G19895: std_logic; attribute dont_touch of G19895: signal is true;
	signal G19896: std_logic; attribute dont_touch of G19896: signal is true;
	signal G19899: std_logic; attribute dont_touch of G19899: signal is true;
	signal G19900: std_logic; attribute dont_touch of G19900: signal is true;
	signal G19901: std_logic; attribute dont_touch of G19901: signal is true;
	signal G19902: std_logic; attribute dont_touch of G19902: signal is true;
	signal G19903: std_logic; attribute dont_touch of G19903: signal is true;
	signal G19904: std_logic; attribute dont_touch of G19904: signal is true;
	signal G19905: std_logic; attribute dont_touch of G19905: signal is true;
	signal G19906: std_logic; attribute dont_touch of G19906: signal is true;
	signal G19907: std_logic; attribute dont_touch of G19907: signal is true;
	signal G19910: std_logic; attribute dont_touch of G19910: signal is true;
	signal G19911: std_logic; attribute dont_touch of G19911: signal is true;
	signal G19912: std_logic; attribute dont_touch of G19912: signal is true;
	signal G19913: std_logic; attribute dont_touch of G19913: signal is true;
	signal G19914: std_logic; attribute dont_touch of G19914: signal is true;
	signal G19915: std_logic; attribute dont_touch of G19915: signal is true;
	signal G19918: std_logic; attribute dont_touch of G19918: signal is true;
	signal G19919: std_logic; attribute dont_touch of G19919: signal is true;
	signal G19920: std_logic; attribute dont_touch of G19920: signal is true;
	signal G19921: std_logic; attribute dont_touch of G19921: signal is true;
	signal G19924: std_logic; attribute dont_touch of G19924: signal is true;
	signal G19925: std_logic; attribute dont_touch of G19925: signal is true;
	signal G19926: std_logic; attribute dont_touch of G19926: signal is true;
	signal G19927: std_logic; attribute dont_touch of G19927: signal is true;
	signal G19928: std_logic; attribute dont_touch of G19928: signal is true;
	signal G19929: std_logic; attribute dont_touch of G19929: signal is true;
	signal G19930: std_logic; attribute dont_touch of G19930: signal is true;
	signal G19931: std_logic; attribute dont_touch of G19931: signal is true;
	signal G19932: std_logic; attribute dont_touch of G19932: signal is true;
	signal G19933: std_logic; attribute dont_touch of G19933: signal is true;
	signal G19934: std_logic; attribute dont_touch of G19934: signal is true;
	signal G19935: std_logic; attribute dont_touch of G19935: signal is true;
	signal G19936: std_logic; attribute dont_touch of G19936: signal is true;
	signal G19939: std_logic; attribute dont_touch of G19939: signal is true;
	signal G19940: std_logic; attribute dont_touch of G19940: signal is true;
	signal G19941: std_logic; attribute dont_touch of G19941: signal is true;
	signal G19942: std_logic; attribute dont_touch of G19942: signal is true;
	signal G19943: std_logic; attribute dont_touch of G19943: signal is true;
	signal G19944: std_logic; attribute dont_touch of G19944: signal is true;
	signal G19945: std_logic; attribute dont_touch of G19945: signal is true;
	signal G19948: std_logic; attribute dont_touch of G19948: signal is true;
	signal G19949: std_logic; attribute dont_touch of G19949: signal is true;
	signal G19950: std_logic; attribute dont_touch of G19950: signal is true;
	signal G19951: std_logic; attribute dont_touch of G19951: signal is true;
	signal G19952: std_logic; attribute dont_touch of G19952: signal is true;
	signal G19953: std_logic; attribute dont_touch of G19953: signal is true;
	signal G19954: std_logic; attribute dont_touch of G19954: signal is true;
	signal G19957: std_logic; attribute dont_touch of G19957: signal is true;
	signal G19970: std_logic; attribute dont_touch of G19970: signal is true;
	signal G19971: std_logic; attribute dont_touch of G19971: signal is true;
	signal G19972: std_logic; attribute dont_touch of G19972: signal is true;
	signal G19975: std_logic; attribute dont_touch of G19975: signal is true;
	signal G19976: std_logic; attribute dont_touch of G19976: signal is true;
	signal G19977: std_logic; attribute dont_touch of G19977: signal is true;
	signal G19978: std_logic; attribute dont_touch of G19978: signal is true;
	signal G19981: std_logic; attribute dont_touch of G19981: signal is true;
	signal G19982: std_logic; attribute dont_touch of G19982: signal is true;
	signal G19983: std_logic; attribute dont_touch of G19983: signal is true;
	signal G19984: std_logic; attribute dont_touch of G19984: signal is true;
	signal G19987: std_logic; attribute dont_touch of G19987: signal is true;
	signal G20000: std_logic; attribute dont_touch of G20000: signal is true;
	signal G20001: std_logic; attribute dont_touch of G20001: signal is true;
	signal G20002: std_logic; attribute dont_touch of G20002: signal is true;
	signal G20005: std_logic; attribute dont_touch of G20005: signal is true;
	signal G20006: std_logic; attribute dont_touch of G20006: signal is true;
	signal G20007: std_logic; attribute dont_touch of G20007: signal is true;
	signal G20008: std_logic; attribute dont_touch of G20008: signal is true;
	signal G20011: std_logic; attribute dont_touch of G20011: signal is true;
	signal G20012: std_logic; attribute dont_touch of G20012: signal is true;
	signal G20013: std_logic; attribute dont_touch of G20013: signal is true;
	signal G20014: std_logic; attribute dont_touch of G20014: signal is true;
	signal G20015: std_logic; attribute dont_touch of G20015: signal is true;
	signal G20016: std_logic; attribute dont_touch of G20016: signal is true;
	signal G20019: std_logic; attribute dont_touch of G20019: signal is true;
	signal G20020: std_logic; attribute dont_touch of G20020: signal is true;
	signal G20021: std_logic; attribute dont_touch of G20021: signal is true;
	signal G20022: std_logic; attribute dont_touch of G20022: signal is true;
	signal G20025: std_logic; attribute dont_touch of G20025: signal is true;
	signal G20038: std_logic; attribute dont_touch of G20038: signal is true;
	signal G20039: std_logic; attribute dont_touch of G20039: signal is true;
	signal G20040: std_logic; attribute dont_touch of G20040: signal is true;
	signal G20043: std_logic; attribute dont_touch of G20043: signal is true;
	signal G20044: std_logic; attribute dont_touch of G20044: signal is true;
	signal G20045: std_logic; attribute dont_touch of G20045: signal is true;
	signal G20048: std_logic; attribute dont_touch of G20048: signal is true;
	signal G20049: std_logic; attribute dont_touch of G20049: signal is true;
	signal G20050: std_logic; attribute dont_touch of G20050: signal is true;
	signal G20051: std_logic; attribute dont_touch of G20051: signal is true;
	signal G20052: std_logic; attribute dont_touch of G20052: signal is true;
	signal G20053: std_logic; attribute dont_touch of G20053: signal is true;
	signal G20054: std_logic; attribute dont_touch of G20054: signal is true;
	signal G20057: std_logic; attribute dont_touch of G20057: signal is true;
	signal G20058: std_logic; attribute dont_touch of G20058: signal is true;
	signal G20061: std_logic; attribute dont_touch of G20061: signal is true;
	signal G20062: std_logic; attribute dont_touch of G20062: signal is true;
	signal G20063: std_logic; attribute dont_touch of G20063: signal is true;
	signal G20064: std_logic; attribute dont_touch of G20064: signal is true;
	signal G20067: std_logic; attribute dont_touch of G20067: signal is true;
	signal G20080: std_logic; attribute dont_touch of G20080: signal is true;
	signal G20081: std_logic; attribute dont_touch of G20081: signal is true;
	signal G20082: std_logic; attribute dont_touch of G20082: signal is true;
	signal G20083: std_logic; attribute dont_touch of G20083: signal is true;
	signal G20084: std_logic; attribute dont_touch of G20084: signal is true;
	signal G20085: std_logic; attribute dont_touch of G20085: signal is true;
	signal G20086: std_logic; attribute dont_touch of G20086: signal is true;
	signal G20087: std_logic; attribute dont_touch of G20087: signal is true;
	signal G20088: std_logic; attribute dont_touch of G20088: signal is true;
	signal G20089: std_logic; attribute dont_touch of G20089: signal is true;
	signal G20090: std_logic; attribute dont_touch of G20090: signal is true;
	signal G20091: std_logic; attribute dont_touch of G20091: signal is true;
	signal G20092: std_logic; attribute dont_touch of G20092: signal is true;
	signal G20093: std_logic; attribute dont_touch of G20093: signal is true;
	signal G20094: std_logic; attribute dont_touch of G20094: signal is true;
	signal G20095: std_logic; attribute dont_touch of G20095: signal is true;
	signal G20098: std_logic; attribute dont_touch of G20098: signal is true;
	signal G20099: std_logic; attribute dont_touch of G20099: signal is true;
	signal G20102: std_logic; attribute dont_touch of G20102: signal is true;
	signal G20103: std_logic; attribute dont_touch of G20103: signal is true;
	signal G20104: std_logic; attribute dont_touch of G20104: signal is true;
	signal G20105: std_logic; attribute dont_touch of G20105: signal is true;
	signal G20106: std_logic; attribute dont_touch of G20106: signal is true;
	signal G20107: std_logic; attribute dont_touch of G20107: signal is true;
	signal G20108: std_logic; attribute dont_touch of G20108: signal is true;
	signal G20109: std_logic; attribute dont_touch of G20109: signal is true;
	signal G20110: std_logic; attribute dont_touch of G20110: signal is true;
	signal G20111: std_logic; attribute dont_touch of G20111: signal is true;
	signal G20112: std_logic; attribute dont_touch of G20112: signal is true;
	signal G20113: std_logic; attribute dont_touch of G20113: signal is true;
	signal G20114: std_logic; attribute dont_touch of G20114: signal is true;
	signal G20115: std_logic; attribute dont_touch of G20115: signal is true;
	signal G20116: std_logic; attribute dont_touch of G20116: signal is true;
	signal G20117: std_logic; attribute dont_touch of G20117: signal is true;
	signal G20118: std_logic; attribute dont_touch of G20118: signal is true;
	signal G20119: std_logic; attribute dont_touch of G20119: signal is true;
	signal G20120: std_logic; attribute dont_touch of G20120: signal is true;
	signal G20123: std_logic; attribute dont_touch of G20123: signal is true;
	signal G20124: std_logic; attribute dont_touch of G20124: signal is true;
	signal G20127: std_logic; attribute dont_touch of G20127: signal is true;
	signal G20131: std_logic; attribute dont_touch of G20131: signal is true;
	signal G20132: std_logic; attribute dont_touch of G20132: signal is true;
	signal G20133: std_logic; attribute dont_touch of G20133: signal is true;
	signal G20134: std_logic; attribute dont_touch of G20134: signal is true;
	signal G20135: std_logic; attribute dont_touch of G20135: signal is true;
	signal G20136: std_logic; attribute dont_touch of G20136: signal is true;
	signal G20137: std_logic; attribute dont_touch of G20137: signal is true;
	signal G20138: std_logic; attribute dont_touch of G20138: signal is true;
	signal G20139: std_logic; attribute dont_touch of G20139: signal is true;
	signal G20140: std_logic; attribute dont_touch of G20140: signal is true;
	signal G20144: std_logic; attribute dont_touch of G20144: signal is true;
	signal G20145: std_logic; attribute dont_touch of G20145: signal is true;
	signal G20146: std_logic; attribute dont_touch of G20146: signal is true;
	signal G20147: std_logic; attribute dont_touch of G20147: signal is true;
	signal G20148: std_logic; attribute dont_touch of G20148: signal is true;
	signal G20149: std_logic; attribute dont_touch of G20149: signal is true;
	signal G20150: std_logic; attribute dont_touch of G20150: signal is true;
	signal G20153: std_logic; attribute dont_touch of G20153: signal is true;
	signal G20156: std_logic; attribute dont_touch of G20156: signal is true;
	signal G20157: std_logic; attribute dont_touch of G20157: signal is true;
	signal G20158: std_logic; attribute dont_touch of G20158: signal is true;
	signal G20159: std_logic; attribute dont_touch of G20159: signal is true;
	signal G20160: std_logic; attribute dont_touch of G20160: signal is true;
	signal G20161: std_logic; attribute dont_touch of G20161: signal is true;
	signal G20162: std_logic; attribute dont_touch of G20162: signal is true;
	signal G20163: std_logic; attribute dont_touch of G20163: signal is true;
	signal G20164: std_logic; attribute dont_touch of G20164: signal is true;
	signal G20177: std_logic; attribute dont_touch of G20177: signal is true;
	signal G20178: std_logic; attribute dont_touch of G20178: signal is true;
	signal G20182: std_logic; attribute dont_touch of G20182: signal is true;
	signal G20183: std_logic; attribute dont_touch of G20183: signal is true;
	signal G20184: std_logic; attribute dont_touch of G20184: signal is true;
	signal G20185: std_logic; attribute dont_touch of G20185: signal is true;
	signal G20186: std_logic; attribute dont_touch of G20186: signal is true;
	signal G20187: std_logic; attribute dont_touch of G20187: signal is true;
	signal G20188: std_logic; attribute dont_touch of G20188: signal is true;
	signal G20189: std_logic; attribute dont_touch of G20189: signal is true;
	signal G20190: std_logic; attribute dont_touch of G20190: signal is true;
	signal G20191: std_logic; attribute dont_touch of G20191: signal is true;
	signal G20192: std_logic; attribute dont_touch of G20192: signal is true;
	signal G20193: std_logic; attribute dont_touch of G20193: signal is true;
	signal G20197: std_logic; attribute dont_touch of G20197: signal is true;
	signal G20198: std_logic; attribute dont_touch of G20198: signal is true;
	signal G20211: std_logic; attribute dont_touch of G20211: signal is true;
	signal G20212: std_logic; attribute dont_touch of G20212: signal is true;
	signal G20216: std_logic; attribute dont_touch of G20216: signal is true;
	signal G20217: std_logic; attribute dont_touch of G20217: signal is true;
	signal G20218: std_logic; attribute dont_touch of G20218: signal is true;
	signal G20219: std_logic; attribute dont_touch of G20219: signal is true;
	signal G20220: std_logic; attribute dont_touch of G20220: signal is true;
	signal G20221: std_logic; attribute dont_touch of G20221: signal is true;
	signal G20222: std_logic; attribute dont_touch of G20222: signal is true;
	signal G20223: std_logic; attribute dont_touch of G20223: signal is true;
	signal G20227: std_logic; attribute dont_touch of G20227: signal is true;
	signal G20228: std_logic; attribute dont_touch of G20228: signal is true;
	signal G20241: std_logic; attribute dont_touch of G20241: signal is true;
	signal G20242: std_logic; attribute dont_touch of G20242: signal is true;
	signal G20246: std_logic; attribute dont_touch of G20246: signal is true;
	signal G20247: std_logic; attribute dont_touch of G20247: signal is true;
	signal G20248: std_logic; attribute dont_touch of G20248: signal is true;
	signal G20249: std_logic; attribute dont_touch of G20249: signal is true;
	signal G20250: std_logic; attribute dont_touch of G20250: signal is true;
	signal G20254: std_logic; attribute dont_touch of G20254: signal is true;
	signal G20255: std_logic; attribute dont_touch of G20255: signal is true;
	signal G20268: std_logic; attribute dont_touch of G20268: signal is true;
	signal G20269: std_logic; attribute dont_touch of G20269: signal is true;
	signal G20270: std_logic; attribute dont_touch of G20270: signal is true;
	signal G20271: std_logic; attribute dont_touch of G20271: signal is true;
	signal G20272: std_logic; attribute dont_touch of G20272: signal is true;
	signal G20273: std_logic; attribute dont_touch of G20273: signal is true;
	signal G20277: std_logic; attribute dont_touch of G20277: signal is true;
	signal G20278: std_logic; attribute dont_touch of G20278: signal is true;
	signal G20279: std_logic; attribute dont_touch of G20279: signal is true;
	signal G20280: std_logic; attribute dont_touch of G20280: signal is true;
	signal G20281: std_logic; attribute dont_touch of G20281: signal is true;
	signal G20282: std_logic; attribute dont_touch of G20282: signal is true;
	signal G20283: std_logic; attribute dont_touch of G20283: signal is true;
	signal G20284: std_logic; attribute dont_touch of G20284: signal is true;
	signal G20285: std_logic; attribute dont_touch of G20285: signal is true;
	signal G20286: std_logic; attribute dont_touch of G20286: signal is true;
	signal G20287: std_logic; attribute dont_touch of G20287: signal is true;
	signal G20288: std_logic; attribute dont_touch of G20288: signal is true;
	signal G20289: std_logic; attribute dont_touch of G20289: signal is true;
	signal G20290: std_logic; attribute dont_touch of G20290: signal is true;
	signal G20291: std_logic; attribute dont_touch of G20291: signal is true;
	signal G20292: std_logic; attribute dont_touch of G20292: signal is true;
	signal G20293: std_logic; attribute dont_touch of G20293: signal is true;
	signal G20294: std_logic; attribute dont_touch of G20294: signal is true;
	signal G20295: std_logic; attribute dont_touch of G20295: signal is true;
	signal G20296: std_logic; attribute dont_touch of G20296: signal is true;
	signal G20297: std_logic; attribute dont_touch of G20297: signal is true;
	signal G20298: std_logic; attribute dont_touch of G20298: signal is true;
	signal G20299: std_logic; attribute dont_touch of G20299: signal is true;
	signal G20302: std_logic; attribute dont_touch of G20302: signal is true;
	signal G20303: std_logic; attribute dont_touch of G20303: signal is true;
	signal G20304: std_logic; attribute dont_touch of G20304: signal is true;
	signal G20305: std_logic; attribute dont_touch of G20305: signal is true;
	signal G20306: std_logic; attribute dont_touch of G20306: signal is true;
	signal G20307: std_logic; attribute dont_touch of G20307: signal is true;
	signal G20308: std_logic; attribute dont_touch of G20308: signal is true;
	signal G20309: std_logic; attribute dont_touch of G20309: signal is true;
	signal G20310: std_logic; attribute dont_touch of G20310: signal is true;
	signal G20311: std_logic; attribute dont_touch of G20311: signal is true;
	signal G20312: std_logic; attribute dont_touch of G20312: signal is true;
	signal G20313: std_logic; attribute dont_touch of G20313: signal is true;
	signal G20314: std_logic; attribute dont_touch of G20314: signal is true;
	signal G20315: std_logic; attribute dont_touch of G20315: signal is true;
	signal G20316: std_logic; attribute dont_touch of G20316: signal is true;
	signal G20317: std_logic; attribute dont_touch of G20317: signal is true;
	signal G20318: std_logic; attribute dont_touch of G20318: signal is true;
	signal G20321: std_logic; attribute dont_touch of G20321: signal is true;
	signal G20322: std_logic; attribute dont_touch of G20322: signal is true;
	signal G20323: std_logic; attribute dont_touch of G20323: signal is true;
	signal G20324: std_logic; attribute dont_touch of G20324: signal is true;
	signal G20325: std_logic; attribute dont_touch of G20325: signal is true;
	signal G20326: std_logic; attribute dont_touch of G20326: signal is true;
	signal G20327: std_logic; attribute dont_touch of G20327: signal is true;
	signal G20328: std_logic; attribute dont_touch of G20328: signal is true;
	signal G20329: std_logic; attribute dont_touch of G20329: signal is true;
	signal G20330: std_logic; attribute dont_touch of G20330: signal is true;
	signal G20331: std_logic; attribute dont_touch of G20331: signal is true;
	signal G20332: std_logic; attribute dont_touch of G20332: signal is true;
	signal G20333: std_logic; attribute dont_touch of G20333: signal is true;
	signal G20334: std_logic; attribute dont_touch of G20334: signal is true;
	signal G20335: std_logic; attribute dont_touch of G20335: signal is true;
	signal G20336: std_logic; attribute dont_touch of G20336: signal is true;
	signal G20337: std_logic; attribute dont_touch of G20337: signal is true;
	signal G20340: std_logic; attribute dont_touch of G20340: signal is true;
	signal G20341: std_logic; attribute dont_touch of G20341: signal is true;
	signal G20342: std_logic; attribute dont_touch of G20342: signal is true;
	signal G20343: std_logic; attribute dont_touch of G20343: signal is true;
	signal G20344: std_logic; attribute dont_touch of G20344: signal is true;
	signal G20345: std_logic; attribute dont_touch of G20345: signal is true;
	signal G20346: std_logic; attribute dont_touch of G20346: signal is true;
	signal G20347: std_logic; attribute dont_touch of G20347: signal is true;
	signal G20348: std_logic; attribute dont_touch of G20348: signal is true;
	signal G20349: std_logic; attribute dont_touch of G20349: signal is true;
	signal G20350: std_logic; attribute dont_touch of G20350: signal is true;
	signal G20351: std_logic; attribute dont_touch of G20351: signal is true;
	signal G20352: std_logic; attribute dont_touch of G20352: signal is true;
	signal G20353: std_logic; attribute dont_touch of G20353: signal is true;
	signal G20354: std_logic; attribute dont_touch of G20354: signal is true;
	signal G20355: std_logic; attribute dont_touch of G20355: signal is true;
	signal G20356: std_logic; attribute dont_touch of G20356: signal is true;
	signal G20357: std_logic; attribute dont_touch of G20357: signal is true;
	signal G20360: std_logic; attribute dont_touch of G20360: signal is true;
	signal G20361: std_logic; attribute dont_touch of G20361: signal is true;
	signal G20362: std_logic; attribute dont_touch of G20362: signal is true;
	signal G20363: std_logic; attribute dont_touch of G20363: signal is true;
	signal G20364: std_logic; attribute dont_touch of G20364: signal is true;
	signal G20365: std_logic; attribute dont_touch of G20365: signal is true;
	signal G20366: std_logic; attribute dont_touch of G20366: signal is true;
	signal G20367: std_logic; attribute dont_touch of G20367: signal is true;
	signal G20368: std_logic; attribute dont_touch of G20368: signal is true;
	signal G20369: std_logic; attribute dont_touch of G20369: signal is true;
	signal G20370: std_logic; attribute dont_touch of G20370: signal is true;
	signal G20371: std_logic; attribute dont_touch of G20371: signal is true;
	signal G20372: std_logic; attribute dont_touch of G20372: signal is true;
	signal G20373: std_logic; attribute dont_touch of G20373: signal is true;
	signal G20374: std_logic; attribute dont_touch of G20374: signal is true;
	signal G20375: std_logic; attribute dont_touch of G20375: signal is true;
	signal G20376: std_logic; attribute dont_touch of G20376: signal is true;
	signal G20377: std_logic; attribute dont_touch of G20377: signal is true;
	signal G20378: std_logic; attribute dont_touch of G20378: signal is true;
	signal G20379: std_logic; attribute dont_touch of G20379: signal is true;
	signal G20380: std_logic; attribute dont_touch of G20380: signal is true;
	signal G20381: std_logic; attribute dont_touch of G20381: signal is true;
	signal G20382: std_logic; attribute dont_touch of G20382: signal is true;
	signal G20383: std_logic; attribute dont_touch of G20383: signal is true;
	signal G20384: std_logic; attribute dont_touch of G20384: signal is true;
	signal G20385: std_logic; attribute dont_touch of G20385: signal is true;
	signal G20386: std_logic; attribute dont_touch of G20386: signal is true;
	signal G20387: std_logic; attribute dont_touch of G20387: signal is true;
	signal G20388: std_logic; attribute dont_touch of G20388: signal is true;
	signal G20389: std_logic; attribute dont_touch of G20389: signal is true;
	signal G20390: std_logic; attribute dont_touch of G20390: signal is true;
	signal G20391: std_logic; attribute dont_touch of G20391: signal is true;
	signal G20392: std_logic; attribute dont_touch of G20392: signal is true;
	signal G20393: std_logic; attribute dont_touch of G20393: signal is true;
	signal G20394: std_logic; attribute dont_touch of G20394: signal is true;
	signal G20395: std_logic; attribute dont_touch of G20395: signal is true;
	signal G20396: std_logic; attribute dont_touch of G20396: signal is true;
	signal G20397: std_logic; attribute dont_touch of G20397: signal is true;
	signal G20398: std_logic; attribute dont_touch of G20398: signal is true;
	signal G20399: std_logic; attribute dont_touch of G20399: signal is true;
	signal G20400: std_logic; attribute dont_touch of G20400: signal is true;
	signal G20401: std_logic; attribute dont_touch of G20401: signal is true;
	signal G20402: std_logic; attribute dont_touch of G20402: signal is true;
	signal G20403: std_logic; attribute dont_touch of G20403: signal is true;
	signal G20404: std_logic; attribute dont_touch of G20404: signal is true;
	signal G20405: std_logic; attribute dont_touch of G20405: signal is true;
	signal G20406: std_logic; attribute dont_touch of G20406: signal is true;
	signal G20407: std_logic; attribute dont_touch of G20407: signal is true;
	signal G20408: std_logic; attribute dont_touch of G20408: signal is true;
	signal G20409: std_logic; attribute dont_touch of G20409: signal is true;
	signal G20410: std_logic; attribute dont_touch of G20410: signal is true;
	signal G20411: std_logic; attribute dont_touch of G20411: signal is true;
	signal G20412: std_logic; attribute dont_touch of G20412: signal is true;
	signal G20413: std_logic; attribute dont_touch of G20413: signal is true;
	signal G20414: std_logic; attribute dont_touch of G20414: signal is true;
	signal G20415: std_logic; attribute dont_touch of G20415: signal is true;
	signal G20416: std_logic; attribute dont_touch of G20416: signal is true;
	signal G20417: std_logic; attribute dont_touch of G20417: signal is true;
	signal G20418: std_logic; attribute dont_touch of G20418: signal is true;
	signal G20419: std_logic; attribute dont_touch of G20419: signal is true;
	signal G20420: std_logic; attribute dont_touch of G20420: signal is true;
	signal G20421: std_logic; attribute dont_touch of G20421: signal is true;
	signal G20422: std_logic; attribute dont_touch of G20422: signal is true;
	signal G20423: std_logic; attribute dont_touch of G20423: signal is true;
	signal G20424: std_logic; attribute dont_touch of G20424: signal is true;
	signal G20425: std_logic; attribute dont_touch of G20425: signal is true;
	signal G20426: std_logic; attribute dont_touch of G20426: signal is true;
	signal G20427: std_logic; attribute dont_touch of G20427: signal is true;
	signal G20428: std_logic; attribute dont_touch of G20428: signal is true;
	signal G20429: std_logic; attribute dont_touch of G20429: signal is true;
	signal G20430: std_logic; attribute dont_touch of G20430: signal is true;
	signal G20431: std_logic; attribute dont_touch of G20431: signal is true;
	signal G20432: std_logic; attribute dont_touch of G20432: signal is true;
	signal G20433: std_logic; attribute dont_touch of G20433: signal is true;
	signal G20434: std_logic; attribute dont_touch of G20434: signal is true;
	signal G20435: std_logic; attribute dont_touch of G20435: signal is true;
	signal G20436: std_logic; attribute dont_touch of G20436: signal is true;
	signal G20437: std_logic; attribute dont_touch of G20437: signal is true;
	signal G20438: std_logic; attribute dont_touch of G20438: signal is true;
	signal G20439: std_logic; attribute dont_touch of G20439: signal is true;
	signal G20440: std_logic; attribute dont_touch of G20440: signal is true;
	signal G20441: std_logic; attribute dont_touch of G20441: signal is true;
	signal G20442: std_logic; attribute dont_touch of G20442: signal is true;
	signal G20443: std_logic; attribute dont_touch of G20443: signal is true;
	signal G20444: std_logic; attribute dont_touch of G20444: signal is true;
	signal G20445: std_logic; attribute dont_touch of G20445: signal is true;
	signal G20446: std_logic; attribute dont_touch of G20446: signal is true;
	signal G20447: std_logic; attribute dont_touch of G20447: signal is true;
	signal G20448: std_logic; attribute dont_touch of G20448: signal is true;
	signal G20449: std_logic; attribute dont_touch of G20449: signal is true;
	signal G20450: std_logic; attribute dont_touch of G20450: signal is true;
	signal G20451: std_logic; attribute dont_touch of G20451: signal is true;
	signal G20452: std_logic; attribute dont_touch of G20452: signal is true;
	signal G20453: std_logic; attribute dont_touch of G20453: signal is true;
	signal G20454: std_logic; attribute dont_touch of G20454: signal is true;
	signal G20455: std_logic; attribute dont_touch of G20455: signal is true;
	signal G20456: std_logic; attribute dont_touch of G20456: signal is true;
	signal G20457: std_logic; attribute dont_touch of G20457: signal is true;
	signal G20458: std_logic; attribute dont_touch of G20458: signal is true;
	signal G20459: std_logic; attribute dont_touch of G20459: signal is true;
	signal G20460: std_logic; attribute dont_touch of G20460: signal is true;
	signal G20461: std_logic; attribute dont_touch of G20461: signal is true;
	signal G20462: std_logic; attribute dont_touch of G20462: signal is true;
	signal G20463: std_logic; attribute dont_touch of G20463: signal is true;
	signal G20464: std_logic; attribute dont_touch of G20464: signal is true;
	signal G20465: std_logic; attribute dont_touch of G20465: signal is true;
	signal G20466: std_logic; attribute dont_touch of G20466: signal is true;
	signal G20467: std_logic; attribute dont_touch of G20467: signal is true;
	signal G20468: std_logic; attribute dont_touch of G20468: signal is true;
	signal G20469: std_logic; attribute dont_touch of G20469: signal is true;
	signal G20470: std_logic; attribute dont_touch of G20470: signal is true;
	signal G20471: std_logic; attribute dont_touch of G20471: signal is true;
	signal G20472: std_logic; attribute dont_touch of G20472: signal is true;
	signal G20473: std_logic; attribute dont_touch of G20473: signal is true;
	signal G20476: std_logic; attribute dont_touch of G20476: signal is true;
	signal G20477: std_logic; attribute dont_touch of G20477: signal is true;
	signal G20478: std_logic; attribute dont_touch of G20478: signal is true;
	signal G20479: std_logic; attribute dont_touch of G20479: signal is true;
	signal G20480: std_logic; attribute dont_touch of G20480: signal is true;
	signal G20481: std_logic; attribute dont_touch of G20481: signal is true;
	signal G20484: std_logic; attribute dont_touch of G20484: signal is true;
	signal G20485: std_logic; attribute dont_touch of G20485: signal is true;
	signal G20486: std_logic; attribute dont_touch of G20486: signal is true;
	signal G20487: std_logic; attribute dont_touch of G20487: signal is true;
	signal G20490: std_logic; attribute dont_touch of G20490: signal is true;
	signal G20491: std_logic; attribute dont_touch of G20491: signal is true;
	signal G20492: std_logic; attribute dont_touch of G20492: signal is true;
	signal G20493: std_logic; attribute dont_touch of G20493: signal is true;
	signal G20496: std_logic; attribute dont_touch of G20496: signal is true;
	signal G20497: std_logic; attribute dont_touch of G20497: signal is true;
	signal G20498: std_logic; attribute dont_touch of G20498: signal is true;
	signal G20499: std_logic; attribute dont_touch of G20499: signal is true;
	signal G20500: std_logic; attribute dont_touch of G20500: signal is true;
	signal G20501: std_logic; attribute dont_touch of G20501: signal is true;
	signal G20502: std_logic; attribute dont_touch of G20502: signal is true;
	signal G20503: std_logic; attribute dont_touch of G20503: signal is true;
	signal G20504: std_logic; attribute dont_touch of G20504: signal is true;
	signal G20505: std_logic; attribute dont_touch of G20505: signal is true;
	signal G20506: std_logic; attribute dont_touch of G20506: signal is true;
	signal G20507: std_logic; attribute dont_touch of G20507: signal is true;
	signal G20512: std_logic; attribute dont_touch of G20512: signal is true;
	signal G20513: std_logic; attribute dont_touch of G20513: signal is true;
	signal G20516: std_logic; attribute dont_touch of G20516: signal is true;
	signal G20517: std_logic; attribute dont_touch of G20517: signal is true;
	signal G20518: std_logic; attribute dont_touch of G20518: signal is true;
	signal G20519: std_logic; attribute dont_touch of G20519: signal is true;
	signal G20522: std_logic; attribute dont_touch of G20522: signal is true;
	signal G20525: std_logic; attribute dont_touch of G20525: signal is true;
	signal G20526: std_logic; attribute dont_touch of G20526: signal is true;
	signal G20531: std_logic; attribute dont_touch of G20531: signal is true;
	signal G20534: std_logic; attribute dont_touch of G20534: signal is true;
	signal G20535: std_logic; attribute dont_touch of G20535: signal is true;
	signal G20536: std_logic; attribute dont_touch of G20536: signal is true;
	signal G20537: std_logic; attribute dont_touch of G20537: signal is true;
	signal G20538: std_logic; attribute dont_touch of G20538: signal is true;
	signal G20539: std_logic; attribute dont_touch of G20539: signal is true;
	signal G20542: std_logic; attribute dont_touch of G20542: signal is true;
	signal G20545: std_logic; attribute dont_touch of G20545: signal is true;
	signal G20550: std_logic; attribute dont_touch of G20550: signal is true;
	signal G20553: std_logic; attribute dont_touch of G20553: signal is true;
	signal G20554: std_logic; attribute dont_touch of G20554: signal is true;
	signal G20555: std_logic; attribute dont_touch of G20555: signal is true;
	signal G20556: std_logic; attribute dont_touch of G20556: signal is true;
	signal G20557: std_logic; attribute dont_touch of G20557: signal is true;
	signal G20558: std_logic; attribute dont_touch of G20558: signal is true;
	signal G20559: std_logic; attribute dont_touch of G20559: signal is true;
	signal G20560: std_logic; attribute dont_touch of G20560: signal is true;
	signal G20561: std_logic; attribute dont_touch of G20561: signal is true;
	signal G20562: std_logic; attribute dont_touch of G20562: signal is true;
	signal G20563: std_logic; attribute dont_touch of G20563: signal is true;
	signal G20564: std_logic; attribute dont_touch of G20564: signal is true;
	signal G20565: std_logic; attribute dont_touch of G20565: signal is true;
	signal G20566: std_logic; attribute dont_touch of G20566: signal is true;
	signal G20567: std_logic; attribute dont_touch of G20567: signal is true;
	signal G20568: std_logic; attribute dont_touch of G20568: signal is true;
	signal G20569: std_logic; attribute dont_touch of G20569: signal is true;
	signal G20570: std_logic; attribute dont_touch of G20570: signal is true;
	signal G20571: std_logic; attribute dont_touch of G20571: signal is true;
	signal G20572: std_logic; attribute dont_touch of G20572: signal is true;
	signal G20573: std_logic; attribute dont_touch of G20573: signal is true;
	signal G20574: std_logic; attribute dont_touch of G20574: signal is true;
	signal G20575: std_logic; attribute dont_touch of G20575: signal is true;
	signal G20576: std_logic; attribute dont_touch of G20576: signal is true;
	signal G20577: std_logic; attribute dont_touch of G20577: signal is true;
	signal G20578: std_logic; attribute dont_touch of G20578: signal is true;
	signal G20579: std_logic; attribute dont_touch of G20579: signal is true;
	signal G20580: std_logic; attribute dont_touch of G20580: signal is true;
	signal G20581: std_logic; attribute dont_touch of G20581: signal is true;
	signal G20582: std_logic; attribute dont_touch of G20582: signal is true;
	signal G20583: std_logic; attribute dont_touch of G20583: signal is true;
	signal G20584: std_logic; attribute dont_touch of G20584: signal is true;
	signal G20585: std_logic; attribute dont_touch of G20585: signal is true;
	signal G20586: std_logic; attribute dont_touch of G20586: signal is true;
	signal G20587: std_logic; attribute dont_touch of G20587: signal is true;
	signal G20588: std_logic; attribute dont_touch of G20588: signal is true;
	signal G20589: std_logic; attribute dont_touch of G20589: signal is true;
	signal G20590: std_logic; attribute dont_touch of G20590: signal is true;
	signal G20591: std_logic; attribute dont_touch of G20591: signal is true;
	signal G20592: std_logic; attribute dont_touch of G20592: signal is true;
	signal G20593: std_logic; attribute dont_touch of G20593: signal is true;
	signal G20594: std_logic; attribute dont_touch of G20594: signal is true;
	signal G20595: std_logic; attribute dont_touch of G20595: signal is true;
	signal G20596: std_logic; attribute dont_touch of G20596: signal is true;
	signal G20597: std_logic; attribute dont_touch of G20597: signal is true;
	signal G20598: std_logic; attribute dont_touch of G20598: signal is true;
	signal G20599: std_logic; attribute dont_touch of G20599: signal is true;
	signal G20600: std_logic; attribute dont_touch of G20600: signal is true;
	signal G20601: std_logic; attribute dont_touch of G20601: signal is true;
	signal G20602: std_logic; attribute dont_touch of G20602: signal is true;
	signal G20603: std_logic; attribute dont_touch of G20603: signal is true;
	signal G20604: std_logic; attribute dont_touch of G20604: signal is true;
	signal G20605: std_logic; attribute dont_touch of G20605: signal is true;
	signal G20606: std_logic; attribute dont_touch of G20606: signal is true;
	signal G20607: std_logic; attribute dont_touch of G20607: signal is true;
	signal G20608: std_logic; attribute dont_touch of G20608: signal is true;
	signal G20609: std_logic; attribute dont_touch of G20609: signal is true;
	signal G20610: std_logic; attribute dont_touch of G20610: signal is true;
	signal G20611: std_logic; attribute dont_touch of G20611: signal is true;
	signal G20612: std_logic; attribute dont_touch of G20612: signal is true;
	signal G20613: std_logic; attribute dont_touch of G20613: signal is true;
	signal G20614: std_logic; attribute dont_touch of G20614: signal is true;
	signal G20615: std_logic; attribute dont_touch of G20615: signal is true;
	signal G20616: std_logic; attribute dont_touch of G20616: signal is true;
	signal G20617: std_logic; attribute dont_touch of G20617: signal is true;
	signal G20618: std_logic; attribute dont_touch of G20618: signal is true;
	signal G20619: std_logic; attribute dont_touch of G20619: signal is true;
	signal G20620: std_logic; attribute dont_touch of G20620: signal is true;
	signal G20621: std_logic; attribute dont_touch of G20621: signal is true;
	signal G20622: std_logic; attribute dont_touch of G20622: signal is true;
	signal G20623: std_logic; attribute dont_touch of G20623: signal is true;
	signal G20624: std_logic; attribute dont_touch of G20624: signal is true;
	signal G20625: std_logic; attribute dont_touch of G20625: signal is true;
	signal G20626: std_logic; attribute dont_touch of G20626: signal is true;
	signal G20627: std_logic; attribute dont_touch of G20627: signal is true;
	signal G20628: std_logic; attribute dont_touch of G20628: signal is true;
	signal G20629: std_logic; attribute dont_touch of G20629: signal is true;
	signal G20630: std_logic; attribute dont_touch of G20630: signal is true;
	signal G20631: std_logic; attribute dont_touch of G20631: signal is true;
	signal G20632: std_logic; attribute dont_touch of G20632: signal is true;
	signal G20633: std_logic; attribute dont_touch of G20633: signal is true;
	signal G20634: std_logic; attribute dont_touch of G20634: signal is true;
	signal G20637: std_logic; attribute dont_touch of G20637: signal is true;
	signal G20640: std_logic; attribute dont_touch of G20640: signal is true;
	signal G20641: std_logic; attribute dont_touch of G20641: signal is true;
	signal G20644: std_logic; attribute dont_touch of G20644: signal is true;
	signal G20647: std_logic; attribute dont_touch of G20647: signal is true;
	signal G20648: std_logic; attribute dont_touch of G20648: signal is true;
	signal G20649: std_logic; attribute dont_touch of G20649: signal is true;
	signal G20652: std_logic; attribute dont_touch of G20652: signal is true;
	signal G20655: std_logic; attribute dont_touch of G20655: signal is true;
	signal G20658: std_logic; attribute dont_touch of G20658: signal is true;
	signal G20659: std_logic; attribute dont_touch of G20659: signal is true;
	signal G20662: std_logic; attribute dont_touch of G20662: signal is true;
	signal G20665: std_logic; attribute dont_touch of G20665: signal is true;
	signal G20666: std_logic; attribute dont_touch of G20666: signal is true;
	signal G20669: std_logic; attribute dont_touch of G20669: signal is true;
	signal G20672: std_logic; attribute dont_touch of G20672: signal is true;
	signal G20673: std_logic; attribute dont_touch of G20673: signal is true;
	signal G20676: std_logic; attribute dont_touch of G20676: signal is true;
	signal G20679: std_logic; attribute dont_touch of G20679: signal is true;
	signal G20682: std_logic; attribute dont_touch of G20682: signal is true;
	signal G20683: std_logic; attribute dont_touch of G20683: signal is true;
	signal G20684: std_logic; attribute dont_touch of G20684: signal is true;
	signal G20687: std_logic; attribute dont_touch of G20687: signal is true;
	signal G20690: std_logic; attribute dont_touch of G20690: signal is true;
	signal G20693: std_logic; attribute dont_touch of G20693: signal is true;
	signal G20694: std_logic; attribute dont_touch of G20694: signal is true;
	signal G20697: std_logic; attribute dont_touch of G20697: signal is true;
	signal G20700: std_logic; attribute dont_touch of G20700: signal is true;
	signal G20703: std_logic; attribute dont_touch of G20703: signal is true;
	signal G20704: std_logic; attribute dont_touch of G20704: signal is true;
	signal G20707: std_logic; attribute dont_touch of G20707: signal is true;
	signal G20708: std_logic; attribute dont_touch of G20708: signal is true;
	signal G20711: std_logic; attribute dont_touch of G20711: signal is true;
	signal G20714: std_logic; attribute dont_touch of G20714: signal is true;
	signal G20717: std_logic; attribute dont_touch of G20717: signal is true;
	signal G20718: std_logic; attribute dont_touch of G20718: signal is true;
	signal G20719: std_logic; attribute dont_touch of G20719: signal is true;
	signal G20722: std_logic; attribute dont_touch of G20722: signal is true;
	signal G20725: std_logic; attribute dont_touch of G20725: signal is true;
	signal G20728: std_logic; attribute dont_touch of G20728: signal is true;
	signal G20729: std_logic; attribute dont_touch of G20729: signal is true;
	signal G20732: std_logic; attribute dont_touch of G20732: signal is true;
	signal G20735: std_logic; attribute dont_touch of G20735: signal is true;
	signal G20738: std_logic; attribute dont_touch of G20738: signal is true;
	signal G20739: std_logic; attribute dont_touch of G20739: signal is true;
	signal G20742: std_logic; attribute dont_touch of G20742: signal is true;
	signal G20743: std_logic; attribute dont_touch of G20743: signal is true;
	signal G20746: std_logic; attribute dont_touch of G20746: signal is true;
	signal G20749: std_logic; attribute dont_touch of G20749: signal is true;
	signal G20752: std_logic; attribute dont_touch of G20752: signal is true;
	signal G20753: std_logic; attribute dont_touch of G20753: signal is true;
	signal G20754: std_logic; attribute dont_touch of G20754: signal is true;
	signal G20757: std_logic; attribute dont_touch of G20757: signal is true;
	signal G20760: std_logic; attribute dont_touch of G20760: signal is true;
	signal G20763: std_logic; attribute dont_touch of G20763: signal is true;
	signal G20766: std_logic; attribute dont_touch of G20766: signal is true;
	signal G20769: std_logic; attribute dont_touch of G20769: signal is true;
	signal G20772: std_logic; attribute dont_touch of G20772: signal is true;
	signal G20775: std_logic; attribute dont_touch of G20775: signal is true;
	signal G20776: std_logic; attribute dont_touch of G20776: signal is true;
	signal G20779: std_logic; attribute dont_touch of G20779: signal is true;
	signal G20780: std_logic; attribute dont_touch of G20780: signal is true;
	signal G20783: std_logic; attribute dont_touch of G20783: signal is true;
	signal G20786: std_logic; attribute dont_touch of G20786: signal is true;
	signal G20789: std_logic; attribute dont_touch of G20789: signal is true;
	signal G20790: std_logic; attribute dont_touch of G20790: signal is true;
	signal G20793: std_logic; attribute dont_touch of G20793: signal is true;
	signal G20796: std_logic; attribute dont_touch of G20796: signal is true;
	signal G20799: std_logic; attribute dont_touch of G20799: signal is true;
	signal G20802: std_logic; attribute dont_touch of G20802: signal is true;
	signal G20805: std_logic; attribute dont_touch of G20805: signal is true;
	signal G20806: std_logic; attribute dont_touch of G20806: signal is true;
	signal G20809: std_logic; attribute dont_touch of G20809: signal is true;
	signal G20810: std_logic; attribute dont_touch of G20810: signal is true;
	signal G20813: std_logic; attribute dont_touch of G20813: signal is true;
	signal G20816: std_logic; attribute dont_touch of G20816: signal is true;
	signal G20819: std_logic; attribute dont_touch of G20819: signal is true;
	signal G20822: std_logic; attribute dont_touch of G20822: signal is true;
	signal G20825: std_logic; attribute dont_touch of G20825: signal is true;
	signal G20826: std_logic; attribute dont_touch of G20826: signal is true;
	signal G20827: std_logic; attribute dont_touch of G20827: signal is true;
	signal G20830: std_logic; attribute dont_touch of G20830: signal is true;
	signal G20833: std_logic; attribute dont_touch of G20833: signal is true;
	signal G20836: std_logic; attribute dont_touch of G20836: signal is true;
	signal G20837: std_logic; attribute dont_touch of G20837: signal is true;
	signal G20840: std_logic; attribute dont_touch of G20840: signal is true;
	signal G20841: std_logic; attribute dont_touch of G20841: signal is true;
	signal G20842: std_logic; attribute dont_touch of G20842: signal is true;
	signal G20850: std_logic; attribute dont_touch of G20850: signal is true;
	signal G20858: std_logic; attribute dont_touch of G20858: signal is true;
	signal G20866: std_logic; attribute dont_touch of G20866: signal is true;
	signal G20874: std_logic; attribute dont_touch of G20874: signal is true;
	signal G20875: std_logic; attribute dont_touch of G20875: signal is true;
	signal G20876: std_logic; attribute dont_touch of G20876: signal is true;
	signal G20877: std_logic; attribute dont_touch of G20877: signal is true;
	signal G20878: std_logic; attribute dont_touch of G20878: signal is true;
	signal G20879: std_logic; attribute dont_touch of G20879: signal is true;
	signal G20880: std_logic; attribute dont_touch of G20880: signal is true;
	signal G20881: std_logic; attribute dont_touch of G20881: signal is true;
	signal G20882: std_logic; attribute dont_touch of G20882: signal is true;
	signal G20883: std_logic; attribute dont_touch of G20883: signal is true;
	signal G20884: std_logic; attribute dont_touch of G20884: signal is true;
	signal G20885: std_logic; attribute dont_touch of G20885: signal is true;
	signal G20891: std_logic; attribute dont_touch of G20891: signal is true;
	signal G20892: std_logic; attribute dont_touch of G20892: signal is true;
	signal G20893: std_logic; attribute dont_touch of G20893: signal is true;
	signal G20894: std_logic; attribute dont_touch of G20894: signal is true;
	signal G20895: std_logic; attribute dont_touch of G20895: signal is true;
	signal G20896: std_logic; attribute dont_touch of G20896: signal is true;
	signal G20897: std_logic; attribute dont_touch of G20897: signal is true;
	signal G20898: std_logic; attribute dont_touch of G20898: signal is true;
	signal G20899: std_logic; attribute dont_touch of G20899: signal is true;
	signal G20900: std_logic; attribute dont_touch of G20900: signal is true;
	signal G20901: std_logic; attribute dont_touch of G20901: signal is true;
	signal G20902: std_logic; attribute dont_touch of G20902: signal is true;
	signal G20903: std_logic; attribute dont_touch of G20903: signal is true;
	signal G20904: std_logic; attribute dont_touch of G20904: signal is true;
	signal G20910: std_logic; attribute dont_touch of G20910: signal is true;
	signal G20911: std_logic; attribute dont_touch of G20911: signal is true;
	signal G20912: std_logic; attribute dont_touch of G20912: signal is true;
	signal G20913: std_logic; attribute dont_touch of G20913: signal is true;
	signal G20914: std_logic; attribute dont_touch of G20914: signal is true;
	signal G20915: std_logic; attribute dont_touch of G20915: signal is true;
	signal G20916: std_logic; attribute dont_touch of G20916: signal is true;
	signal G20917: std_logic; attribute dont_touch of G20917: signal is true;
	signal G20918: std_logic; attribute dont_touch of G20918: signal is true;
	signal G20919: std_logic; attribute dont_touch of G20919: signal is true;
	signal G20920: std_logic; attribute dont_touch of G20920: signal is true;
	signal G20921: std_logic; attribute dont_touch of G20921: signal is true;
	signal G20922: std_logic; attribute dont_touch of G20922: signal is true;
	signal G20923: std_logic; attribute dont_touch of G20923: signal is true;
	signal G20924: std_logic; attribute dont_touch of G20924: signal is true;
	signal G20925: std_logic; attribute dont_touch of G20925: signal is true;
	signal G20926: std_logic; attribute dont_touch of G20926: signal is true;
	signal G20927: std_logic; attribute dont_touch of G20927: signal is true;
	signal G20928: std_logic; attribute dont_touch of G20928: signal is true;
	signal G20934: std_logic; attribute dont_touch of G20934: signal is true;
	signal G20935: std_logic; attribute dont_touch of G20935: signal is true;
	signal G20936: std_logic; attribute dont_touch of G20936: signal is true;
	signal G20937: std_logic; attribute dont_touch of G20937: signal is true;
	signal G20938: std_logic; attribute dont_touch of G20938: signal is true;
	signal G20939: std_logic; attribute dont_touch of G20939: signal is true;
	signal G20940: std_logic; attribute dont_touch of G20940: signal is true;
	signal G20941: std_logic; attribute dont_touch of G20941: signal is true;
	signal G20942: std_logic; attribute dont_touch of G20942: signal is true;
	signal G20943: std_logic; attribute dont_touch of G20943: signal is true;
	signal G20944: std_logic; attribute dont_touch of G20944: signal is true;
	signal G20945: std_logic; attribute dont_touch of G20945: signal is true;
	signal G20946: std_logic; attribute dont_touch of G20946: signal is true;
	signal G20947: std_logic; attribute dont_touch of G20947: signal is true;
	signal G20948: std_logic; attribute dont_touch of G20948: signal is true;
	signal G20949: std_logic; attribute dont_touch of G20949: signal is true;
	signal G20950: std_logic; attribute dont_touch of G20950: signal is true;
	signal G20951: std_logic; attribute dont_touch of G20951: signal is true;
	signal G20952: std_logic; attribute dont_touch of G20952: signal is true;
	signal G20953: std_logic; attribute dont_touch of G20953: signal is true;
	signal G20954: std_logic; attribute dont_touch of G20954: signal is true;
	signal G20955: std_logic; attribute dont_touch of G20955: signal is true;
	signal G20956: std_logic; attribute dont_touch of G20956: signal is true;
	signal G20962: std_logic; attribute dont_touch of G20962: signal is true;
	signal G20963: std_logic; attribute dont_touch of G20963: signal is true;
	signal G20964: std_logic; attribute dont_touch of G20964: signal is true;
	signal G20965: std_logic; attribute dont_touch of G20965: signal is true;
	signal G20966: std_logic; attribute dont_touch of G20966: signal is true;
	signal G20967: std_logic; attribute dont_touch of G20967: signal is true;
	signal G20968: std_logic; attribute dont_touch of G20968: signal is true;
	signal G20969: std_logic; attribute dont_touch of G20969: signal is true;
	signal G20970: std_logic; attribute dont_touch of G20970: signal is true;
	signal G20971: std_logic; attribute dont_touch of G20971: signal is true;
	signal G20972: std_logic; attribute dont_touch of G20972: signal is true;
	signal G20973: std_logic; attribute dont_touch of G20973: signal is true;
	signal G20974: std_logic; attribute dont_touch of G20974: signal is true;
	signal G20975: std_logic; attribute dont_touch of G20975: signal is true;
	signal G20976: std_logic; attribute dont_touch of G20976: signal is true;
	signal G20977: std_logic; attribute dont_touch of G20977: signal is true;
	signal G20978: std_logic; attribute dont_touch of G20978: signal is true;
	signal G20979: std_logic; attribute dont_touch of G20979: signal is true;
	signal G20980: std_logic; attribute dont_touch of G20980: signal is true;
	signal G20981: std_logic; attribute dont_touch of G20981: signal is true;
	signal G20982: std_logic; attribute dont_touch of G20982: signal is true;
	signal G20983: std_logic; attribute dont_touch of G20983: signal is true;
	signal G20984: std_logic; attribute dont_touch of G20984: signal is true;
	signal G20985: std_logic; attribute dont_touch of G20985: signal is true;
	signal G20986: std_logic; attribute dont_touch of G20986: signal is true;
	signal G20989: std_logic; attribute dont_touch of G20989: signal is true;
	signal G20990: std_logic; attribute dont_touch of G20990: signal is true;
	signal G20991: std_logic; attribute dont_touch of G20991: signal is true;
	signal G20992: std_logic; attribute dont_touch of G20992: signal is true;
	signal G20993: std_logic; attribute dont_touch of G20993: signal is true;
	signal G20994: std_logic; attribute dont_touch of G20994: signal is true;
	signal G20995: std_logic; attribute dont_touch of G20995: signal is true;
	signal G20996: std_logic; attribute dont_touch of G20996: signal is true;
	signal G20997: std_logic; attribute dont_touch of G20997: signal is true;
	signal G20998: std_logic; attribute dont_touch of G20998: signal is true;
	signal G20999: std_logic; attribute dont_touch of G20999: signal is true;
	signal G21000: std_logic; attribute dont_touch of G21000: signal is true;
	signal G21001: std_logic; attribute dont_touch of G21001: signal is true;
	signal G21002: std_logic; attribute dont_touch of G21002: signal is true;
	signal G21003: std_logic; attribute dont_touch of G21003: signal is true;
	signal G21004: std_logic; attribute dont_touch of G21004: signal is true;
	signal G21005: std_logic; attribute dont_touch of G21005: signal is true;
	signal G21006: std_logic; attribute dont_touch of G21006: signal is true;
	signal G21007: std_logic; attribute dont_touch of G21007: signal is true;
	signal G21008: std_logic; attribute dont_touch of G21008: signal is true;
	signal G21009: std_logic; attribute dont_touch of G21009: signal is true;
	signal G21010: std_logic; attribute dont_touch of G21010: signal is true;
	signal G21011: std_logic; attribute dont_touch of G21011: signal is true;
	signal G21012: std_logic; attribute dont_touch of G21012: signal is true;
	signal G21015: std_logic; attribute dont_touch of G21015: signal is true;
	signal G21016: std_logic; attribute dont_touch of G21016: signal is true;
	signal G21017: std_logic; attribute dont_touch of G21017: signal is true;
	signal G21018: std_logic; attribute dont_touch of G21018: signal is true;
	signal G21019: std_logic; attribute dont_touch of G21019: signal is true;
	signal G21020: std_logic; attribute dont_touch of G21020: signal is true;
	signal G21021: std_logic; attribute dont_touch of G21021: signal is true;
	signal G21022: std_logic; attribute dont_touch of G21022: signal is true;
	signal G21023: std_logic; attribute dont_touch of G21023: signal is true;
	signal G21024: std_logic; attribute dont_touch of G21024: signal is true;
	signal G21025: std_logic; attribute dont_touch of G21025: signal is true;
	signal G21026: std_logic; attribute dont_touch of G21026: signal is true;
	signal G21027: std_logic; attribute dont_touch of G21027: signal is true;
	signal G21028: std_logic; attribute dont_touch of G21028: signal is true;
	signal G21029: std_logic; attribute dont_touch of G21029: signal is true;
	signal G21030: std_logic; attribute dont_touch of G21030: signal is true;
	signal G21031: std_logic; attribute dont_touch of G21031: signal is true;
	signal G21032: std_logic; attribute dont_touch of G21032: signal is true;
	signal G21033: std_logic; attribute dont_touch of G21033: signal is true;
	signal G21034: std_logic; attribute dont_touch of G21034: signal is true;
	signal G21035: std_logic; attribute dont_touch of G21035: signal is true;
	signal G21036: std_logic; attribute dont_touch of G21036: signal is true;
	signal G21039: std_logic; attribute dont_touch of G21039: signal is true;
	signal G21040: std_logic; attribute dont_touch of G21040: signal is true;
	signal G21041: std_logic; attribute dont_touch of G21041: signal is true;
	signal G21042: std_logic; attribute dont_touch of G21042: signal is true;
	signal G21043: std_logic; attribute dont_touch of G21043: signal is true;
	signal G21044: std_logic; attribute dont_touch of G21044: signal is true;
	signal G21045: std_logic; attribute dont_touch of G21045: signal is true;
	signal G21046: std_logic; attribute dont_touch of G21046: signal is true;
	signal G21047: std_logic; attribute dont_touch of G21047: signal is true;
	signal G21048: std_logic; attribute dont_touch of G21048: signal is true;
	signal G21049: std_logic; attribute dont_touch of G21049: signal is true;
	signal G21050: std_logic; attribute dont_touch of G21050: signal is true;
	signal G21051: std_logic; attribute dont_touch of G21051: signal is true;
	signal G21052: std_logic; attribute dont_touch of G21052: signal is true;
	signal G21053: std_logic; attribute dont_touch of G21053: signal is true;
	signal G21054: std_logic; attribute dont_touch of G21054: signal is true;
	signal G21055: std_logic; attribute dont_touch of G21055: signal is true;
	signal G21056: std_logic; attribute dont_touch of G21056: signal is true;
	signal G21057: std_logic; attribute dont_touch of G21057: signal is true;
	signal G21060: std_logic; attribute dont_touch of G21060: signal is true;
	signal G21061: std_logic; attribute dont_touch of G21061: signal is true;
	signal G21062: std_logic; attribute dont_touch of G21062: signal is true;
	signal G21063: std_logic; attribute dont_touch of G21063: signal is true;
	signal G21064: std_logic; attribute dont_touch of G21064: signal is true;
	signal G21065: std_logic; attribute dont_touch of G21065: signal is true;
	signal G21066: std_logic; attribute dont_touch of G21066: signal is true;
	signal G21067: std_logic; attribute dont_touch of G21067: signal is true;
	signal G21068: std_logic; attribute dont_touch of G21068: signal is true;
	signal G21069: std_logic; attribute dont_touch of G21069: signal is true;
	signal G21070: std_logic; attribute dont_touch of G21070: signal is true;
	signal G21071: std_logic; attribute dont_touch of G21071: signal is true;
	signal G21072: std_logic; attribute dont_touch of G21072: signal is true;
	signal G21073: std_logic; attribute dont_touch of G21073: signal is true;
	signal G21074: std_logic; attribute dont_touch of G21074: signal is true;
	signal G21075: std_logic; attribute dont_touch of G21075: signal is true;
	signal G21076: std_logic; attribute dont_touch of G21076: signal is true;
	signal G21077: std_logic; attribute dont_touch of G21077: signal is true;
	signal G21078: std_logic; attribute dont_touch of G21078: signal is true;
	signal G21079: std_logic; attribute dont_touch of G21079: signal is true;
	signal G21080: std_logic; attribute dont_touch of G21080: signal is true;
	signal G21081: std_logic; attribute dont_touch of G21081: signal is true;
	signal G21082: std_logic; attribute dont_touch of G21082: signal is true;
	signal G21083: std_logic; attribute dont_touch of G21083: signal is true;
	signal G21084: std_logic; attribute dont_touch of G21084: signal is true;
	signal G21085: std_logic; attribute dont_touch of G21085: signal is true;
	signal G21086: std_logic; attribute dont_touch of G21086: signal is true;
	signal G21087: std_logic; attribute dont_touch of G21087: signal is true;
	signal G21090: std_logic; attribute dont_touch of G21090: signal is true;
	signal G21091: std_logic; attribute dont_touch of G21091: signal is true;
	signal G21092: std_logic; attribute dont_touch of G21092: signal is true;
	signal G21093: std_logic; attribute dont_touch of G21093: signal is true;
	signal G21094: std_logic; attribute dont_touch of G21094: signal is true;
	signal G21095: std_logic; attribute dont_touch of G21095: signal is true;
	signal G21096: std_logic; attribute dont_touch of G21096: signal is true;
	signal G21097: std_logic; attribute dont_touch of G21097: signal is true;
	signal G21098: std_logic; attribute dont_touch of G21098: signal is true;
	signal G21099: std_logic; attribute dont_touch of G21099: signal is true;
	signal G21102: std_logic; attribute dont_touch of G21102: signal is true;
	signal G21103: std_logic; attribute dont_touch of G21103: signal is true;
	signal G21104: std_logic; attribute dont_touch of G21104: signal is true;
	signal G21105: std_logic; attribute dont_touch of G21105: signal is true;
	signal G21106: std_logic; attribute dont_touch of G21106: signal is true;
	signal G21107: std_logic; attribute dont_touch of G21107: signal is true;
	signal G21108: std_logic; attribute dont_touch of G21108: signal is true;
	signal G21111: std_logic; attribute dont_touch of G21111: signal is true;
	signal G21112: std_logic; attribute dont_touch of G21112: signal is true;
	signal G21113: std_logic; attribute dont_touch of G21113: signal is true;
	signal G21116: std_logic; attribute dont_touch of G21116: signal is true;
	signal G21117: std_logic; attribute dont_touch of G21117: signal is true;
	signal G21118: std_logic; attribute dont_touch of G21118: signal is true;
	signal G21119: std_logic; attribute dont_touch of G21119: signal is true;
	signal G21120: std_logic; attribute dont_touch of G21120: signal is true;
	signal G21121: std_logic; attribute dont_touch of G21121: signal is true;
	signal G21122: std_logic; attribute dont_touch of G21122: signal is true;
	signal G21123: std_logic; attribute dont_touch of G21123: signal is true;
	signal G21124: std_logic; attribute dont_touch of G21124: signal is true;
	signal G21125: std_logic; attribute dont_touch of G21125: signal is true;
	signal G21128: std_logic; attribute dont_touch of G21128: signal is true;
	signal G21129: std_logic; attribute dont_touch of G21129: signal is true;
	signal G21130: std_logic; attribute dont_touch of G21130: signal is true;
	signal G21133: std_logic; attribute dont_touch of G21133: signal is true;
	signal G21134: std_logic; attribute dont_touch of G21134: signal is true;
	signal G21135: std_logic; attribute dont_touch of G21135: signal is true;
	signal G21136: std_logic; attribute dont_touch of G21136: signal is true;
	signal G21137: std_logic; attribute dont_touch of G21137: signal is true;
	signal G21138: std_logic; attribute dont_touch of G21138: signal is true;
	signal G21139: std_logic; attribute dont_touch of G21139: signal is true;
	signal G21140: std_logic; attribute dont_touch of G21140: signal is true;
	signal G21141: std_logic; attribute dont_touch of G21141: signal is true;
	signal G21142: std_logic; attribute dont_touch of G21142: signal is true;
	signal G21143: std_logic; attribute dont_touch of G21143: signal is true;
	signal G21144: std_logic; attribute dont_touch of G21144: signal is true;
	signal G21147: std_logic; attribute dont_touch of G21147: signal is true;
	signal G21148: std_logic; attribute dont_touch of G21148: signal is true;
	signal G21149: std_logic; attribute dont_touch of G21149: signal is true;
	signal G21152: std_logic; attribute dont_touch of G21152: signal is true;
	signal G21153: std_logic; attribute dont_touch of G21153: signal is true;
	signal G21154: std_logic; attribute dont_touch of G21154: signal is true;
	signal G21155: std_logic; attribute dont_touch of G21155: signal is true;
	signal G21156: std_logic; attribute dont_touch of G21156: signal is true;
	signal G21157: std_logic; attribute dont_touch of G21157: signal is true;
	signal G21158: std_logic; attribute dont_touch of G21158: signal is true;
	signal G21159: std_logic; attribute dont_touch of G21159: signal is true;
	signal G21160: std_logic; attribute dont_touch of G21160: signal is true;
	signal G21161: std_logic; attribute dont_touch of G21161: signal is true;
	signal G21162: std_logic; attribute dont_touch of G21162: signal is true;
	signal G21163: std_logic; attribute dont_touch of G21163: signal is true;
	signal G21164: std_logic; attribute dont_touch of G21164: signal is true;
	signal G21167: std_logic; attribute dont_touch of G21167: signal is true;
	signal G21168: std_logic; attribute dont_touch of G21168: signal is true;
	signal G21169: std_logic; attribute dont_touch of G21169: signal is true;
	signal G21172: std_logic; attribute dont_touch of G21172: signal is true;
	signal G21173: std_logic; attribute dont_touch of G21173: signal is true;
	signal G21174: std_logic; attribute dont_touch of G21174: signal is true;
	signal G21175: std_logic; attribute dont_touch of G21175: signal is true;
	signal G21176: std_logic; attribute dont_touch of G21176: signal is true;
	signal G21177: std_logic; attribute dont_touch of G21177: signal is true;
	signal G21178: std_logic; attribute dont_touch of G21178: signal is true;
	signal G21179: std_logic; attribute dont_touch of G21179: signal is true;
	signal G21180: std_logic; attribute dont_touch of G21180: signal is true;
	signal G21181: std_logic; attribute dont_touch of G21181: signal is true;
	signal G21182: std_logic; attribute dont_touch of G21182: signal is true;
	signal G21183: std_logic; attribute dont_touch of G21183: signal is true;
	signal G21184: std_logic; attribute dont_touch of G21184: signal is true;
	signal G21187: std_logic; attribute dont_touch of G21187: signal is true;
	signal G21188: std_logic; attribute dont_touch of G21188: signal is true;
	signal G21189: std_logic; attribute dont_touch of G21189: signal is true;
	signal G21192: std_logic; attribute dont_touch of G21192: signal is true;
	signal G21193: std_logic; attribute dont_touch of G21193: signal is true;
	signal G21194: std_logic; attribute dont_touch of G21194: signal is true;
	signal G21195: std_logic; attribute dont_touch of G21195: signal is true;
	signal G21196: std_logic; attribute dont_touch of G21196: signal is true;
	signal G21197: std_logic; attribute dont_touch of G21197: signal is true;
	signal G21198: std_logic; attribute dont_touch of G21198: signal is true;
	signal G21199: std_logic; attribute dont_touch of G21199: signal is true;
	signal G21202: std_logic; attribute dont_touch of G21202: signal is true;
	signal G21203: std_logic; attribute dont_touch of G21203: signal is true;
	signal G21204: std_logic; attribute dont_touch of G21204: signal is true;
	signal G21207: std_logic; attribute dont_touch of G21207: signal is true;
	signal G21208: std_logic; attribute dont_touch of G21208: signal is true;
	signal G21209: std_logic; attribute dont_touch of G21209: signal is true;
	signal G21210: std_logic; attribute dont_touch of G21210: signal is true;
	signal G21211: std_logic; attribute dont_touch of G21211: signal is true;
	signal G21214: std_logic; attribute dont_touch of G21214: signal is true;
	signal G21217: std_logic; attribute dont_touch of G21217: signal is true;
	signal G21218: std_logic; attribute dont_touch of G21218: signal is true;
	signal G21219: std_logic; attribute dont_touch of G21219: signal is true;
	signal G21222: std_logic; attribute dont_touch of G21222: signal is true;
	signal G21225: std_logic; attribute dont_touch of G21225: signal is true;
	signal G21226: std_logic; attribute dont_touch of G21226: signal is true;
	signal G21227: std_logic; attribute dont_touch of G21227: signal is true;
	signal G21228: std_logic; attribute dont_touch of G21228: signal is true;
	signal G21229: std_logic; attribute dont_touch of G21229: signal is true;
	signal G21230: std_logic; attribute dont_touch of G21230: signal is true;
	signal G21233: std_logic; attribute dont_touch of G21233: signal is true;
	signal G21234: std_logic; attribute dont_touch of G21234: signal is true;
	signal G21235: std_logic; attribute dont_touch of G21235: signal is true;
	signal G21238: std_logic; attribute dont_touch of G21238: signal is true;
	signal G21241: std_logic; attribute dont_touch of G21241: signal is true;
	signal G21242: std_logic; attribute dont_touch of G21242: signal is true;
	signal G21243: std_logic; attribute dont_touch of G21243: signal is true;
	signal G21244: std_logic; attribute dont_touch of G21244: signal is true;
	signal G21245: std_logic; attribute dont_touch of G21245: signal is true;
	signal G21246: std_logic; attribute dont_touch of G21246: signal is true;
	signal G21249: std_logic; attribute dont_touch of G21249: signal is true;
	signal G21250: std_logic; attribute dont_touch of G21250: signal is true;
	signal G21251: std_logic; attribute dont_touch of G21251: signal is true;
	signal G21252: std_logic; attribute dont_touch of G21252: signal is true;
	signal G21253: std_logic; attribute dont_touch of G21253: signal is true;
	signal G21254: std_logic; attribute dont_touch of G21254: signal is true;
	signal G21255: std_logic; attribute dont_touch of G21255: signal is true;
	signal G21258: std_logic; attribute dont_touch of G21258: signal is true;
	signal G21259: std_logic; attribute dont_touch of G21259: signal is true;
	signal G21260: std_logic; attribute dont_touch of G21260: signal is true;
	signal G21261: std_logic; attribute dont_touch of G21261: signal is true;
	signal G21262: std_logic; attribute dont_touch of G21262: signal is true;
	signal G21263: std_logic; attribute dont_touch of G21263: signal is true;
	signal G21266: std_logic; attribute dont_touch of G21266: signal is true;
	signal G21267: std_logic; attribute dont_touch of G21267: signal is true;
	signal G21268: std_logic; attribute dont_touch of G21268: signal is true;
	signal G21269: std_logic; attribute dont_touch of G21269: signal is true;
	signal G21270: std_logic; attribute dont_touch of G21270: signal is true;
	signal G21271: std_logic; attribute dont_touch of G21271: signal is true;
	signal G21276: std_logic; attribute dont_touch of G21276: signal is true;
	signal G21277: std_logic; attribute dont_touch of G21277: signal is true;
	signal G21278: std_logic; attribute dont_touch of G21278: signal is true;
	signal G21283: std_logic; attribute dont_touch of G21283: signal is true;
	signal G21284: std_logic; attribute dont_touch of G21284: signal is true;
	signal G21285: std_logic; attribute dont_touch of G21285: signal is true;
	signal G21290: std_logic; attribute dont_touch of G21290: signal is true;
	signal G21291: std_logic; attribute dont_touch of G21291: signal is true;
	signal G21292: std_logic; attribute dont_touch of G21292: signal is true;
	signal G21293: std_logic; attribute dont_touch of G21293: signal is true;
	signal G21298: std_logic; attribute dont_touch of G21298: signal is true;
	signal G21299: std_logic; attribute dont_touch of G21299: signal is true;
	signal G21300: std_logic; attribute dont_touch of G21300: signal is true;
	signal G21301: std_logic; attribute dont_touch of G21301: signal is true;
	signal G21302: std_logic; attribute dont_touch of G21302: signal is true;
	signal G21303: std_logic; attribute dont_touch of G21303: signal is true;
	signal G21304: std_logic; attribute dont_touch of G21304: signal is true;
	signal G21305: std_logic; attribute dont_touch of G21305: signal is true;
	signal G21306: std_logic; attribute dont_touch of G21306: signal is true;
	signal G21307: std_logic; attribute dont_touch of G21307: signal is true;
	signal G21308: std_logic; attribute dont_touch of G21308: signal is true;
	signal G21309: std_logic; attribute dont_touch of G21309: signal is true;
	signal G21310: std_logic; attribute dont_touch of G21310: signal is true;
	signal G21311: std_logic; attribute dont_touch of G21311: signal is true;
	signal G21312: std_logic; attribute dont_touch of G21312: signal is true;
	signal G21313: std_logic; attribute dont_touch of G21313: signal is true;
	signal G21314: std_logic; attribute dont_touch of G21314: signal is true;
	signal G21315: std_logic; attribute dont_touch of G21315: signal is true;
	signal G21316: std_logic; attribute dont_touch of G21316: signal is true;
	signal G21319: std_logic; attribute dont_touch of G21319: signal is true;
	signal G21320: std_logic; attribute dont_touch of G21320: signal is true;
	signal G21321: std_logic; attribute dont_touch of G21321: signal is true;
	signal G21322: std_logic; attribute dont_touch of G21322: signal is true;
	signal G21323: std_logic; attribute dont_touch of G21323: signal is true;
	signal G21324: std_logic; attribute dont_touch of G21324: signal is true;
	signal G21325: std_logic; attribute dont_touch of G21325: signal is true;
	signal G21326: std_logic; attribute dont_touch of G21326: signal is true;
	signal G21327: std_logic; attribute dont_touch of G21327: signal is true;
	signal G21328: std_logic; attribute dont_touch of G21328: signal is true;
	signal G21329: std_logic; attribute dont_touch of G21329: signal is true;
	signal G21330: std_logic; attribute dont_touch of G21330: signal is true;
	signal G21331: std_logic; attribute dont_touch of G21331: signal is true;
	signal G21334: std_logic; attribute dont_touch of G21334: signal is true;
	signal G21335: std_logic; attribute dont_touch of G21335: signal is true;
	signal G21336: std_logic; attribute dont_touch of G21336: signal is true;
	signal G21337: std_logic; attribute dont_touch of G21337: signal is true;
	signal G21338: std_logic; attribute dont_touch of G21338: signal is true;
	signal G21339: std_logic; attribute dont_touch of G21339: signal is true;
	signal G21340: std_logic; attribute dont_touch of G21340: signal is true;
	signal G21341: std_logic; attribute dont_touch of G21341: signal is true;
	signal G21342: std_logic; attribute dont_touch of G21342: signal is true;
	signal G21343: std_logic; attribute dont_touch of G21343: signal is true;
	signal G21344: std_logic; attribute dont_touch of G21344: signal is true;
	signal G21345: std_logic; attribute dont_touch of G21345: signal is true;
	signal G21346: std_logic; attribute dont_touch of G21346: signal is true;
	signal G21349: std_logic; attribute dont_touch of G21349: signal is true;
	signal G21350: std_logic; attribute dont_touch of G21350: signal is true;
	signal G21351: std_logic; attribute dont_touch of G21351: signal is true;
	signal G21352: std_logic; attribute dont_touch of G21352: signal is true;
	signal G21353: std_logic; attribute dont_touch of G21353: signal is true;
	signal G21354: std_logic; attribute dont_touch of G21354: signal is true;
	signal G21355: std_logic; attribute dont_touch of G21355: signal is true;
	signal G21356: std_logic; attribute dont_touch of G21356: signal is true;
	signal G21357: std_logic; attribute dont_touch of G21357: signal is true;
	signal G21358: std_logic; attribute dont_touch of G21358: signal is true;
	signal G21359: std_logic; attribute dont_touch of G21359: signal is true;
	signal G21360: std_logic; attribute dont_touch of G21360: signal is true;
	signal G21361: std_logic; attribute dont_touch of G21361: signal is true;
	signal G21362: std_logic; attribute dont_touch of G21362: signal is true;
	signal G21363: std_logic; attribute dont_touch of G21363: signal is true;
	signal G21364: std_logic; attribute dont_touch of G21364: signal is true;
	signal G21367: std_logic; attribute dont_touch of G21367: signal is true;
	signal G21368: std_logic; attribute dont_touch of G21368: signal is true;
	signal G21369: std_logic; attribute dont_touch of G21369: signal is true;
	signal G21370: std_logic; attribute dont_touch of G21370: signal is true;
	signal G21371: std_logic; attribute dont_touch of G21371: signal is true;
	signal G21372: std_logic; attribute dont_touch of G21372: signal is true;
	signal G21373: std_logic; attribute dont_touch of G21373: signal is true;
	signal G21374: std_logic; attribute dont_touch of G21374: signal is true;
	signal G21375: std_logic; attribute dont_touch of G21375: signal is true;
	signal G21376: std_logic; attribute dont_touch of G21376: signal is true;
	signal G21377: std_logic; attribute dont_touch of G21377: signal is true;
	signal G21378: std_logic; attribute dont_touch of G21378: signal is true;
	signal G21379: std_logic; attribute dont_touch of G21379: signal is true;
	signal G21380: std_logic; attribute dont_touch of G21380: signal is true;
	signal G21381: std_logic; attribute dont_touch of G21381: signal is true;
	signal G21382: std_logic; attribute dont_touch of G21382: signal is true;
	signal G21385: std_logic; attribute dont_touch of G21385: signal is true;
	signal G21388: std_logic; attribute dont_touch of G21388: signal is true;
	signal G21389: std_logic; attribute dont_touch of G21389: signal is true;
	signal G21390: std_logic; attribute dont_touch of G21390: signal is true;
	signal G21391: std_logic; attribute dont_touch of G21391: signal is true;
	signal G21392: std_logic; attribute dont_touch of G21392: signal is true;
	signal G21393: std_logic; attribute dont_touch of G21393: signal is true;
	signal G21394: std_logic; attribute dont_touch of G21394: signal is true;
	signal G21395: std_logic; attribute dont_touch of G21395: signal is true;
	signal G21396: std_logic; attribute dont_touch of G21396: signal is true;
	signal G21397: std_logic; attribute dont_touch of G21397: signal is true;
	signal G21398: std_logic; attribute dont_touch of G21398: signal is true;
	signal G21399: std_logic; attribute dont_touch of G21399: signal is true;
	signal G21400: std_logic; attribute dont_touch of G21400: signal is true;
	signal G21401: std_logic; attribute dont_touch of G21401: signal is true;
	signal G21402: std_logic; attribute dont_touch of G21402: signal is true;
	signal G21403: std_logic; attribute dont_touch of G21403: signal is true;
	signal G21404: std_logic; attribute dont_touch of G21404: signal is true;
	signal G21407: std_logic; attribute dont_touch of G21407: signal is true;
	signal G21410: std_logic; attribute dont_touch of G21410: signal is true;
	signal G21411: std_logic; attribute dont_touch of G21411: signal is true;
	signal G21412: std_logic; attribute dont_touch of G21412: signal is true;
	signal G21413: std_logic; attribute dont_touch of G21413: signal is true;
	signal G21414: std_logic; attribute dont_touch of G21414: signal is true;
	signal G21415: std_logic; attribute dont_touch of G21415: signal is true;
	signal G21418: std_logic; attribute dont_touch of G21418: signal is true;
	signal G21419: std_logic; attribute dont_touch of G21419: signal is true;
	signal G21420: std_logic; attribute dont_touch of G21420: signal is true;
	signal G21421: std_logic; attribute dont_touch of G21421: signal is true;
	signal G21422: std_logic; attribute dont_touch of G21422: signal is true;
	signal G21423: std_logic; attribute dont_touch of G21423: signal is true;
	signal G21424: std_logic; attribute dont_touch of G21424: signal is true;
	signal G21425: std_logic; attribute dont_touch of G21425: signal is true;
	signal G21426: std_logic; attribute dont_touch of G21426: signal is true;
	signal G21427: std_logic; attribute dont_touch of G21427: signal is true;
	signal G21428: std_logic; attribute dont_touch of G21428: signal is true;
	signal G21429: std_logic; attribute dont_touch of G21429: signal is true;
	signal G21432: std_logic; attribute dont_touch of G21432: signal is true;
	signal G21435: std_logic; attribute dont_touch of G21435: signal is true;
	signal G21438: std_logic; attribute dont_touch of G21438: signal is true;
	signal G21439: std_logic; attribute dont_touch of G21439: signal is true;
	signal G21440: std_logic; attribute dont_touch of G21440: signal is true;
	signal G21441: std_logic; attribute dont_touch of G21441: signal is true;
	signal G21444: std_logic; attribute dont_touch of G21444: signal is true;
	signal G21445: std_logic; attribute dont_touch of G21445: signal is true;
	signal G21446: std_logic; attribute dont_touch of G21446: signal is true;
	signal G21447: std_logic; attribute dont_touch of G21447: signal is true;
	signal G21448: std_logic; attribute dont_touch of G21448: signal is true;
	signal G21449: std_logic; attribute dont_touch of G21449: signal is true;
	signal G21452: std_logic; attribute dont_touch of G21452: signal is true;
	signal G21453: std_logic; attribute dont_touch of G21453: signal is true;
	signal G21454: std_logic; attribute dont_touch of G21454: signal is true;
	signal G21455: std_logic; attribute dont_touch of G21455: signal is true;
	signal G21456: std_logic; attribute dont_touch of G21456: signal is true;
	signal G21457: std_logic; attribute dont_touch of G21457: signal is true;
	signal G21458: std_logic; attribute dont_touch of G21458: signal is true;
	signal G21461: std_logic; attribute dont_touch of G21461: signal is true;
	signal G21467: std_logic; attribute dont_touch of G21467: signal is true;
	signal G21470: std_logic; attribute dont_touch of G21470: signal is true;
	signal G21473: std_logic; attribute dont_touch of G21473: signal is true;
	signal G21476: std_logic; attribute dont_touch of G21476: signal is true;
	signal G21477: std_logic; attribute dont_touch of G21477: signal is true;
	signal G21480: std_logic; attribute dont_touch of G21480: signal is true;
	signal G21481: std_logic; attribute dont_touch of G21481: signal is true;
	signal G21482: std_logic; attribute dont_touch of G21482: signal is true;
	signal G21483: std_logic; attribute dont_touch of G21483: signal is true;
	signal G21486: std_logic; attribute dont_touch of G21486: signal is true;
	signal G21487: std_logic; attribute dont_touch of G21487: signal is true;
	signal G21488: std_logic; attribute dont_touch of G21488: signal is true;
	signal G21489: std_logic; attribute dont_touch of G21489: signal is true;
	signal G21490: std_logic; attribute dont_touch of G21490: signal is true;
	signal G21491: std_logic; attribute dont_touch of G21491: signal is true;
	signal G21494: std_logic; attribute dont_touch of G21494: signal is true;
	signal G21495: std_logic; attribute dont_touch of G21495: signal is true;
	signal G21496: std_logic; attribute dont_touch of G21496: signal is true;
	signal G21497: std_logic; attribute dont_touch of G21497: signal is true;
	signal G21498: std_logic; attribute dont_touch of G21498: signal is true;
	signal G21501: std_logic; attribute dont_touch of G21501: signal is true;
	signal G21502: std_logic; attribute dont_touch of G21502: signal is true;
	signal G21505: std_logic; attribute dont_touch of G21505: signal is true;
	signal G21508: std_logic; attribute dont_touch of G21508: signal is true;
	signal G21514: std_logic; attribute dont_touch of G21514: signal is true;
	signal G21517: std_logic; attribute dont_touch of G21517: signal is true;
	signal G21518: std_logic; attribute dont_touch of G21518: signal is true;
	signal G21521: std_logic; attribute dont_touch of G21521: signal is true;
	signal G21522: std_logic; attribute dont_touch of G21522: signal is true;
	signal G21523: std_logic; attribute dont_touch of G21523: signal is true;
	signal G21524: std_logic; attribute dont_touch of G21524: signal is true;
	signal G21527: std_logic; attribute dont_touch of G21527: signal is true;
	signal G21528: std_logic; attribute dont_touch of G21528: signal is true;
	signal G21529: std_logic; attribute dont_touch of G21529: signal is true;
	signal G21530: std_logic; attribute dont_touch of G21530: signal is true;
	signal G21533: std_logic; attribute dont_touch of G21533: signal is true;
	signal G21536: std_logic; attribute dont_touch of G21536: signal is true;
	signal G21537: std_logic; attribute dont_touch of G21537: signal is true;
	signal G21540: std_logic; attribute dont_touch of G21540: signal is true;
	signal G21541: std_logic; attribute dont_touch of G21541: signal is true;
	signal G21544: std_logic; attribute dont_touch of G21544: signal is true;
	signal G21550: std_logic; attribute dont_touch of G21550: signal is true;
	signal G21553: std_logic; attribute dont_touch of G21553: signal is true;
	signal G21554: std_logic; attribute dont_touch of G21554: signal is true;
	signal G21557: std_logic; attribute dont_touch of G21557: signal is true;
	signal G21558: std_logic; attribute dont_touch of G21558: signal is true;
	signal G21561: std_logic; attribute dont_touch of G21561: signal is true;
	signal G21564: std_logic; attribute dont_touch of G21564: signal is true;
	signal G21565: std_logic; attribute dont_touch of G21565: signal is true;
	signal G21566: std_logic; attribute dont_touch of G21566: signal is true;
	signal G21569: std_logic; attribute dont_touch of G21569: signal is true;
	signal G21572: std_logic; attribute dont_touch of G21572: signal is true;
	signal G21573: std_logic; attribute dont_touch of G21573: signal is true;
	signal G21576: std_logic; attribute dont_touch of G21576: signal is true;
	signal G21577: std_logic; attribute dont_touch of G21577: signal is true;
	signal G21580: std_logic; attribute dont_touch of G21580: signal is true;
	signal G21586: std_logic; attribute dont_touch of G21586: signal is true;
	signal G21589: std_logic; attribute dont_touch of G21589: signal is true;
	signal G21590: std_logic; attribute dont_touch of G21590: signal is true;
	signal G21593: std_logic; attribute dont_touch of G21593: signal is true;
	signal G21594: std_logic; attribute dont_touch of G21594: signal is true;
	signal G21597: std_logic; attribute dont_touch of G21597: signal is true;
	signal G21598: std_logic; attribute dont_touch of G21598: signal is true;
	signal G21599: std_logic; attribute dont_touch of G21599: signal is true;
	signal G21602: std_logic; attribute dont_touch of G21602: signal is true;
	signal G21605: std_logic; attribute dont_touch of G21605: signal is true;
	signal G21606: std_logic; attribute dont_touch of G21606: signal is true;
	signal G21609: std_logic; attribute dont_touch of G21609: signal is true;
	signal G21610: std_logic; attribute dont_touch of G21610: signal is true;
	signal G21611: std_logic; attribute dont_touch of G21611: signal is true;
	signal G21612: std_logic; attribute dont_touch of G21612: signal is true;
	signal G21615: std_logic; attribute dont_touch of G21615: signal is true;
	signal G21618: std_logic; attribute dont_touch of G21618: signal is true;
	signal G21619: std_logic; attribute dont_touch of G21619: signal is true;
	signal G21622: std_logic; attribute dont_touch of G21622: signal is true;
	signal G21623: std_logic; attribute dont_touch of G21623: signal is true;
	signal G21626: std_logic; attribute dont_touch of G21626: signal is true;
	signal G21627: std_logic; attribute dont_touch of G21627: signal is true;
	signal G21628: std_logic; attribute dont_touch of G21628: signal is true;
	signal G21631: std_logic; attribute dont_touch of G21631: signal is true;
	signal G21634: std_logic; attribute dont_touch of G21634: signal is true;
	signal G21635: std_logic; attribute dont_touch of G21635: signal is true;
	signal G21636: std_logic; attribute dont_touch of G21636: signal is true;
	signal G21639: std_logic; attribute dont_touch of G21639: signal is true;
	signal G21640: std_logic; attribute dont_touch of G21640: signal is true;
	signal G21643: std_logic; attribute dont_touch of G21643: signal is true;
	signal G21646: std_logic; attribute dont_touch of G21646: signal is true;
	signal G21647: std_logic; attribute dont_touch of G21647: signal is true;
	signal G21650: std_logic; attribute dont_touch of G21650: signal is true;
	signal G21651: std_logic; attribute dont_touch of G21651: signal is true;
	signal G21654: std_logic; attribute dont_touch of G21654: signal is true;
	signal G21655: std_logic; attribute dont_touch of G21655: signal is true;
	signal G21658: std_logic; attribute dont_touch of G21658: signal is true;
	signal G21659: std_logic; attribute dont_touch of G21659: signal is true;
	signal G21660: std_logic; attribute dont_touch of G21660: signal is true;
	signal G21661: std_logic; attribute dont_touch of G21661: signal is true;
	signal G21665: std_logic; attribute dont_touch of G21665: signal is true;
	signal G21666: std_logic; attribute dont_touch of G21666: signal is true;
	signal G21667: std_logic; attribute dont_touch of G21667: signal is true;
	signal G21670: std_logic; attribute dont_touch of G21670: signal is true;
	signal G21671: std_logic; attribute dont_touch of G21671: signal is true;
	signal G21674: std_logic; attribute dont_touch of G21674: signal is true;
	signal G21677: std_logic; attribute dont_touch of G21677: signal is true;
	signal G21678: std_logic; attribute dont_touch of G21678: signal is true;
	signal G21681: std_logic; attribute dont_touch of G21681: signal is true;
	signal G21682: std_logic; attribute dont_touch of G21682: signal is true;
	signal G21685: std_logic; attribute dont_touch of G21685: signal is true;
	signal G21686: std_logic; attribute dont_touch of G21686: signal is true;
	signal G21687: std_logic; attribute dont_touch of G21687: signal is true;
	signal G21688: std_logic; attribute dont_touch of G21688: signal is true;
	signal G21689: std_logic; attribute dont_touch of G21689: signal is true;
	signal G21690: std_logic; attribute dont_touch of G21690: signal is true;
	signal G21694: std_logic; attribute dont_touch of G21694: signal is true;
	signal G21695: std_logic; attribute dont_touch of G21695: signal is true;
	signal G21696: std_logic; attribute dont_touch of G21696: signal is true;
	signal G21699: std_logic; attribute dont_touch of G21699: signal is true;
	signal G21700: std_logic; attribute dont_touch of G21700: signal is true;
	signal G21703: std_logic; attribute dont_touch of G21703: signal is true;
	signal G21706: std_logic; attribute dont_touch of G21706: signal is true;
	signal G21707: std_logic; attribute dont_touch of G21707: signal is true;
	signal G21708: std_logic; attribute dont_touch of G21708: signal is true;
	signal G21711: std_logic; attribute dont_touch of G21711: signal is true;
	signal G21714: std_logic; attribute dont_touch of G21714: signal is true;
	signal G21715: std_logic; attribute dont_touch of G21715: signal is true;
	signal G21716: std_logic; attribute dont_touch of G21716: signal is true;
	signal G21720: std_logic; attribute dont_touch of G21720: signal is true;
	signal G21721: std_logic; attribute dont_touch of G21721: signal is true;
	signal G21722: std_logic; attribute dont_touch of G21722: signal is true;
	signal G21723: std_logic; attribute dont_touch of G21723: signal is true;
	signal G21724: std_logic; attribute dont_touch of G21724: signal is true;
	signal G21725: std_logic; attribute dont_touch of G21725: signal is true;
	signal G21726: std_logic; attribute dont_touch of G21726: signal is true;
	signal G21730: std_logic; attribute dont_touch of G21730: signal is true;
	signal G21731: std_logic; attribute dont_touch of G21731: signal is true;
	signal G21732: std_logic; attribute dont_touch of G21732: signal is true;
	signal G21735: std_logic; attribute dont_touch of G21735: signal is true;
	signal G21736: std_logic; attribute dont_touch of G21736: signal is true;
	signal G21737: std_logic; attribute dont_touch of G21737: signal is true;
	signal G21738: std_logic; attribute dont_touch of G21738: signal is true;
	signal G21739: std_logic; attribute dont_touch of G21739: signal is true;
	signal G21740: std_logic; attribute dont_touch of G21740: signal is true;
	signal G21741: std_logic; attribute dont_touch of G21741: signal is true;
	signal G21742: std_logic; attribute dont_touch of G21742: signal is true;
	signal G21746: std_logic; attribute dont_touch of G21746: signal is true;
	signal G21747: std_logic; attribute dont_touch of G21747: signal is true;
	signal G21748: std_logic; attribute dont_touch of G21748: signal is true;
	signal G21749: std_logic; attribute dont_touch of G21749: signal is true;
	signal G21750: std_logic; attribute dont_touch of G21750: signal is true;
	signal G21751: std_logic; attribute dont_touch of G21751: signal is true;
	signal G21752: std_logic; attribute dont_touch of G21752: signal is true;
	signal G21756: std_logic; attribute dont_touch of G21756: signal is true;
	signal G21757: std_logic; attribute dont_touch of G21757: signal is true;
	signal G21758: std_logic; attribute dont_touch of G21758: signal is true;
	signal G21759: std_logic; attribute dont_touch of G21759: signal is true;
	signal G21760: std_logic; attribute dont_touch of G21760: signal is true;
	signal G21761: std_logic; attribute dont_touch of G21761: signal is true;
	signal G21762: std_logic; attribute dont_touch of G21762: signal is true;
	signal G21763: std_logic; attribute dont_touch of G21763: signal is true;
	signal G21764: std_logic; attribute dont_touch of G21764: signal is true;
	signal G21765: std_logic; attribute dont_touch of G21765: signal is true;
	signal G21766: std_logic; attribute dont_touch of G21766: signal is true;
	signal G21770: std_logic; attribute dont_touch of G21770: signal is true;
	signal G21771: std_logic; attribute dont_touch of G21771: signal is true;
	signal G21772: std_logic; attribute dont_touch of G21772: signal is true;
	signal G21773: std_logic; attribute dont_touch of G21773: signal is true;
	signal G21774: std_logic; attribute dont_touch of G21774: signal is true;
	signal G21775: std_logic; attribute dont_touch of G21775: signal is true;
	signal G21776: std_logic; attribute dont_touch of G21776: signal is true;
	signal G21777: std_logic; attribute dont_touch of G21777: signal is true;
	signal G21778: std_logic; attribute dont_touch of G21778: signal is true;
	signal G21779: std_logic; attribute dont_touch of G21779: signal is true;
	signal G21780: std_logic; attribute dont_touch of G21780: signal is true;
	signal G21781: std_logic; attribute dont_touch of G21781: signal is true;
	signal G21782: std_logic; attribute dont_touch of G21782: signal is true;
	signal G21786: std_logic; attribute dont_touch of G21786: signal is true;
	signal G21787: std_logic; attribute dont_touch of G21787: signal is true;
	signal G21788: std_logic; attribute dont_touch of G21788: signal is true;
	signal G21789: std_logic; attribute dont_touch of G21789: signal is true;
	signal G21790: std_logic; attribute dont_touch of G21790: signal is true;
	signal G21791: std_logic; attribute dont_touch of G21791: signal is true;
	signal G21792: std_logic; attribute dont_touch of G21792: signal is true;
	signal G21793: std_logic; attribute dont_touch of G21793: signal is true;
	signal G21794: std_logic; attribute dont_touch of G21794: signal is true;
	signal G21795: std_logic; attribute dont_touch of G21795: signal is true;
	signal G21796: std_logic; attribute dont_touch of G21796: signal is true;
	signal G21799: std_logic; attribute dont_touch of G21799: signal is true;
	signal G21800: std_logic; attribute dont_touch of G21800: signal is true;
	signal G21801: std_logic; attribute dont_touch of G21801: signal is true;
	signal G21802: std_logic; attribute dont_touch of G21802: signal is true;
	signal G21803: std_logic; attribute dont_touch of G21803: signal is true;
	signal G21804: std_logic; attribute dont_touch of G21804: signal is true;
	signal G21805: std_logic; attribute dont_touch of G21805: signal is true;
	signal G21806: std_logic; attribute dont_touch of G21806: signal is true;
	signal G21807: std_logic; attribute dont_touch of G21807: signal is true;
	signal G21808: std_logic; attribute dont_touch of G21808: signal is true;
	signal G21809: std_logic; attribute dont_touch of G21809: signal is true;
	signal G21810: std_logic; attribute dont_touch of G21810: signal is true;
	signal G21811: std_logic; attribute dont_touch of G21811: signal is true;
	signal G21812: std_logic; attribute dont_touch of G21812: signal is true;
	signal G21813: std_logic; attribute dont_touch of G21813: signal is true;
	signal G21814: std_logic; attribute dont_touch of G21814: signal is true;
	signal G21815: std_logic; attribute dont_touch of G21815: signal is true;
	signal G21816: std_logic; attribute dont_touch of G21816: signal is true;
	signal G21817: std_logic; attribute dont_touch of G21817: signal is true;
	signal G21818: std_logic; attribute dont_touch of G21818: signal is true;
	signal G21819: std_logic; attribute dont_touch of G21819: signal is true;
	signal G21820: std_logic; attribute dont_touch of G21820: signal is true;
	signal G21821: std_logic; attribute dont_touch of G21821: signal is true;
	signal G21822: std_logic; attribute dont_touch of G21822: signal is true;
	signal G21823: std_logic; attribute dont_touch of G21823: signal is true;
	signal G21824: std_logic; attribute dont_touch of G21824: signal is true;
	signal G21825: std_logic; attribute dont_touch of G21825: signal is true;
	signal G21842: std_logic; attribute dont_touch of G21842: signal is true;
	signal G21843: std_logic; attribute dont_touch of G21843: signal is true;
	signal G21844: std_logic; attribute dont_touch of G21844: signal is true;
	signal G21845: std_logic; attribute dont_touch of G21845: signal is true;
	signal G21846: std_logic; attribute dont_touch of G21846: signal is true;
	signal G21847: std_logic; attribute dont_touch of G21847: signal is true;
	signal G21848: std_logic; attribute dont_touch of G21848: signal is true;
	signal G21849: std_logic; attribute dont_touch of G21849: signal is true;
	signal G21850: std_logic; attribute dont_touch of G21850: signal is true;
	signal G21851: std_logic; attribute dont_touch of G21851: signal is true;
	signal G21855: std_logic; attribute dont_touch of G21855: signal is true;
	signal G21856: std_logic; attribute dont_touch of G21856: signal is true;
	signal G21857: std_logic; attribute dont_touch of G21857: signal is true;
	signal G21858: std_logic; attribute dont_touch of G21858: signal is true;
	signal G21859: std_logic; attribute dont_touch of G21859: signal is true;
	signal G21860: std_logic; attribute dont_touch of G21860: signal is true;
	signal G21861: std_logic; attribute dont_touch of G21861: signal is true;
	signal G21862: std_logic; attribute dont_touch of G21862: signal is true;
	signal G21863: std_logic; attribute dont_touch of G21863: signal is true;
	signal G21864: std_logic; attribute dont_touch of G21864: signal is true;
	signal G21865: std_logic; attribute dont_touch of G21865: signal is true;
	signal G21866: std_logic; attribute dont_touch of G21866: signal is true;
	signal G21867: std_logic; attribute dont_touch of G21867: signal is true;
	signal G21868: std_logic; attribute dont_touch of G21868: signal is true;
	signal G21869: std_logic; attribute dont_touch of G21869: signal is true;
	signal G21870: std_logic; attribute dont_touch of G21870: signal is true;
	signal G21871: std_logic; attribute dont_touch of G21871: signal is true;
	signal G21872: std_logic; attribute dont_touch of G21872: signal is true;
	signal G21873: std_logic; attribute dont_touch of G21873: signal is true;
	signal G21874: std_logic; attribute dont_touch of G21874: signal is true;
	signal G21875: std_logic; attribute dont_touch of G21875: signal is true;
	signal G21876: std_logic; attribute dont_touch of G21876: signal is true;
	signal G21877: std_logic; attribute dont_touch of G21877: signal is true;
	signal G21878: std_logic; attribute dont_touch of G21878: signal is true;
	signal G21879: std_logic; attribute dont_touch of G21879: signal is true;
	signal G21880: std_logic; attribute dont_touch of G21880: signal is true;
	signal G21881: std_logic; attribute dont_touch of G21881: signal is true;
	signal G21882: std_logic; attribute dont_touch of G21882: signal is true;
	signal G21883: std_logic; attribute dont_touch of G21883: signal is true;
	signal G21884: std_logic; attribute dont_touch of G21884: signal is true;
	signal G21885: std_logic; attribute dont_touch of G21885: signal is true;
	signal G21886: std_logic; attribute dont_touch of G21886: signal is true;
	signal G21887: std_logic; attribute dont_touch of G21887: signal is true;
	signal G21888: std_logic; attribute dont_touch of G21888: signal is true;
	signal G21889: std_logic; attribute dont_touch of G21889: signal is true;
	signal G21890: std_logic; attribute dont_touch of G21890: signal is true;
	signal G21891: std_logic; attribute dont_touch of G21891: signal is true;
	signal G21892: std_logic; attribute dont_touch of G21892: signal is true;
	signal G21893: std_logic; attribute dont_touch of G21893: signal is true;
	signal G21894: std_logic; attribute dont_touch of G21894: signal is true;
	signal G21895: std_logic; attribute dont_touch of G21895: signal is true;
	signal G21899: std_logic; attribute dont_touch of G21899: signal is true;
	signal G21900: std_logic; attribute dont_touch of G21900: signal is true;
	signal G21901: std_logic; attribute dont_touch of G21901: signal is true;
	signal G21902: std_logic; attribute dont_touch of G21902: signal is true;
	signal G21903: std_logic; attribute dont_touch of G21903: signal is true;
	signal G21906: std_logic; attribute dont_touch of G21906: signal is true;
	signal G21907: std_logic; attribute dont_touch of G21907: signal is true;
	signal G21911: std_logic; attribute dont_touch of G21911: signal is true;
	signal G21912: std_logic; attribute dont_touch of G21912: signal is true;
	signal G21913: std_logic; attribute dont_touch of G21913: signal is true;
	signal G21914: std_logic; attribute dont_touch of G21914: signal is true;
	signal G21917: std_logic; attribute dont_touch of G21917: signal is true;
	signal G21920: std_logic; attribute dont_touch of G21920: signal is true;
	signal G21921: std_logic; attribute dont_touch of G21921: signal is true;
	signal G21925: std_logic; attribute dont_touch of G21925: signal is true;
	signal G21926: std_logic; attribute dont_touch of G21926: signal is true;
	signal G21927: std_logic; attribute dont_touch of G21927: signal is true;
	signal G21928: std_logic; attribute dont_touch of G21928: signal is true;
	signal G21931: std_logic; attribute dont_touch of G21931: signal is true;
	signal G21932: std_logic; attribute dont_touch of G21932: signal is true;
	signal G21935: std_logic; attribute dont_touch of G21935: signal is true;
	signal G21938: std_logic; attribute dont_touch of G21938: signal is true;
	signal G21939: std_logic; attribute dont_touch of G21939: signal is true;
	signal G21943: std_logic; attribute dont_touch of G21943: signal is true;
	signal G21944: std_logic; attribute dont_touch of G21944: signal is true;
	signal G21945: std_logic; attribute dont_touch of G21945: signal is true;
	signal G21946: std_logic; attribute dont_touch of G21946: signal is true;
	signal G21947: std_logic; attribute dont_touch of G21947: signal is true;
	signal G21948: std_logic; attribute dont_touch of G21948: signal is true;
	signal G21949: std_logic; attribute dont_touch of G21949: signal is true;
	signal G21950: std_logic; attribute dont_touch of G21950: signal is true;
	signal G21951: std_logic; attribute dont_touch of G21951: signal is true;
	signal G21952: std_logic; attribute dont_touch of G21952: signal is true;
	signal G21953: std_logic; attribute dont_touch of G21953: signal is true;
	signal G21954: std_logic; attribute dont_touch of G21954: signal is true;
	signal G21955: std_logic; attribute dont_touch of G21955: signal is true;
	signal G21956: std_logic; attribute dont_touch of G21956: signal is true;
	signal G21957: std_logic; attribute dont_touch of G21957: signal is true;
	signal G21958: std_logic; attribute dont_touch of G21958: signal is true;
	signal G21959: std_logic; attribute dont_touch of G21959: signal is true;
	signal G21960: std_logic; attribute dont_touch of G21960: signal is true;
	signal G21961: std_logic; attribute dont_touch of G21961: signal is true;
	signal G21962: std_logic; attribute dont_touch of G21962: signal is true;
	signal G21963: std_logic; attribute dont_touch of G21963: signal is true;
	signal G21964: std_logic; attribute dont_touch of G21964: signal is true;
	signal G21965: std_logic; attribute dont_touch of G21965: signal is true;
	signal G21966: std_logic; attribute dont_touch of G21966: signal is true;
	signal G21967: std_logic; attribute dont_touch of G21967: signal is true;
	signal G21968: std_logic; attribute dont_touch of G21968: signal is true;
	signal G21969: std_logic; attribute dont_touch of G21969: signal is true;
	signal G21970: std_logic; attribute dont_touch of G21970: signal is true;
	signal G21971: std_logic; attribute dont_touch of G21971: signal is true;
	signal G21972: std_logic; attribute dont_touch of G21972: signal is true;
	signal G21973: std_logic; attribute dont_touch of G21973: signal is true;
	signal G21974: std_logic; attribute dont_touch of G21974: signal is true;
	signal G21975: std_logic; attribute dont_touch of G21975: signal is true;
	signal G21976: std_logic; attribute dont_touch of G21976: signal is true;
	signal G21980: std_logic; attribute dont_touch of G21980: signal is true;
	signal G21981: std_logic; attribute dont_touch of G21981: signal is true;
	signal G21982: std_logic; attribute dont_touch of G21982: signal is true;
	signal G21983: std_logic; attribute dont_touch of G21983: signal is true;
	signal G21987: std_logic; attribute dont_touch of G21987: signal is true;
	signal G21988: std_logic; attribute dont_touch of G21988: signal is true;
	signal G21989: std_logic; attribute dont_touch of G21989: signal is true;
	signal G21990: std_logic; attribute dont_touch of G21990: signal is true;
	signal G21991: std_logic; attribute dont_touch of G21991: signal is true;
	signal G21995: std_logic; attribute dont_touch of G21995: signal is true;
	signal G21996: std_logic; attribute dont_touch of G21996: signal is true;
	signal G22000: std_logic; attribute dont_touch of G22000: signal is true;
	signal G22001: std_logic; attribute dont_touch of G22001: signal is true;
	signal G22002: std_logic; attribute dont_touch of G22002: signal is true;
	signal G22003: std_logic; attribute dont_touch of G22003: signal is true;
	signal G22004: std_logic; attribute dont_touch of G22004: signal is true;
	signal G22005: std_logic; attribute dont_touch of G22005: signal is true;
	signal G22009: std_logic; attribute dont_touch of G22009: signal is true;
	signal G22013: std_logic; attribute dont_touch of G22013: signal is true;
	signal G22014: std_logic; attribute dont_touch of G22014: signal is true;
	signal G22015: std_logic; attribute dont_touch of G22015: signal is true;
	signal G22016: std_logic; attribute dont_touch of G22016: signal is true;
	signal G22020: std_logic; attribute dont_touch of G22020: signal is true;
	signal G22021: std_logic; attribute dont_touch of G22021: signal is true;
	signal G22025: std_logic; attribute dont_touch of G22025: signal is true;
	signal G22026: std_logic; attribute dont_touch of G22026: signal is true;
	signal G22027: std_logic; attribute dont_touch of G22027: signal is true;
	signal G22028: std_logic; attribute dont_touch of G22028: signal is true;
	signal G22029: std_logic; attribute dont_touch of G22029: signal is true;
	signal G22030: std_logic; attribute dont_touch of G22030: signal is true;
	signal G22031: std_logic; attribute dont_touch of G22031: signal is true;
	signal G22032: std_logic; attribute dont_touch of G22032: signal is true;
	signal G22033: std_logic; attribute dont_touch of G22033: signal is true;
	signal G22034: std_logic; attribute dont_touch of G22034: signal is true;
	signal G22035: std_logic; attribute dont_touch of G22035: signal is true;
	signal G22036: std_logic; attribute dont_touch of G22036: signal is true;
	signal G22037: std_logic; attribute dont_touch of G22037: signal is true;
	signal G22038: std_logic; attribute dont_touch of G22038: signal is true;
	signal G22039: std_logic; attribute dont_touch of G22039: signal is true;
	signal G22040: std_logic; attribute dont_touch of G22040: signal is true;
	signal G22041: std_logic; attribute dont_touch of G22041: signal is true;
	signal G22042: std_logic; attribute dont_touch of G22042: signal is true;
	signal G22043: std_logic; attribute dont_touch of G22043: signal is true;
	signal G22044: std_logic; attribute dont_touch of G22044: signal is true;
	signal G22045: std_logic; attribute dont_touch of G22045: signal is true;
	signal G22046: std_logic; attribute dont_touch of G22046: signal is true;
	signal G22047: std_logic; attribute dont_touch of G22047: signal is true;
	signal G22048: std_logic; attribute dont_touch of G22048: signal is true;
	signal G22049: std_logic; attribute dont_touch of G22049: signal is true;
	signal G22050: std_logic; attribute dont_touch of G22050: signal is true;
	signal G22054: std_logic; attribute dont_touch of G22054: signal is true;
	signal G22055: std_logic; attribute dont_touch of G22055: signal is true;
	signal G22056: std_logic; attribute dont_touch of G22056: signal is true;
	signal G22057: std_logic; attribute dont_touch of G22057: signal is true;
	signal G22058: std_logic; attribute dont_touch of G22058: signal is true;
	signal G22059: std_logic; attribute dont_touch of G22059: signal is true;
	signal G22060: std_logic; attribute dont_touch of G22060: signal is true;
	signal G22061: std_logic; attribute dont_touch of G22061: signal is true;
	signal G22062: std_logic; attribute dont_touch of G22062: signal is true;
	signal G22063: std_logic; attribute dont_touch of G22063: signal is true;
	signal G22064: std_logic; attribute dont_touch of G22064: signal is true;
	signal G22065: std_logic; attribute dont_touch of G22065: signal is true;
	signal G22066: std_logic; attribute dont_touch of G22066: signal is true;
	signal G22067: std_logic; attribute dont_touch of G22067: signal is true;
	signal G22068: std_logic; attribute dont_touch of G22068: signal is true;
	signal G22069: std_logic; attribute dont_touch of G22069: signal is true;
	signal G22073: std_logic; attribute dont_touch of G22073: signal is true;
	signal G22074: std_logic; attribute dont_touch of G22074: signal is true;
	signal G22075: std_logic; attribute dont_touch of G22075: signal is true;
	signal G22076: std_logic; attribute dont_touch of G22076: signal is true;
	signal G22077: std_logic; attribute dont_touch of G22077: signal is true;
	signal G22078: std_logic; attribute dont_touch of G22078: signal is true;
	signal G22079: std_logic; attribute dont_touch of G22079: signal is true;
	signal G22080: std_logic; attribute dont_touch of G22080: signal is true;
	signal G22081: std_logic; attribute dont_touch of G22081: signal is true;
	signal G22082: std_logic; attribute dont_touch of G22082: signal is true;
	signal G22083: std_logic; attribute dont_touch of G22083: signal is true;
	signal G22087: std_logic; attribute dont_touch of G22087: signal is true;
	signal G22088: std_logic; attribute dont_touch of G22088: signal is true;
	signal G22089: std_logic; attribute dont_touch of G22089: signal is true;
	signal G22090: std_logic; attribute dont_touch of G22090: signal is true;
	signal G22091: std_logic; attribute dont_touch of G22091: signal is true;
	signal G22092: std_logic; attribute dont_touch of G22092: signal is true;
	signal G22093: std_logic; attribute dont_touch of G22093: signal is true;
	signal G22097: std_logic; attribute dont_touch of G22097: signal is true;
	signal G22098: std_logic; attribute dont_touch of G22098: signal is true;
	signal G22099: std_logic; attribute dont_touch of G22099: signal is true;
	signal G22100: std_logic; attribute dont_touch of G22100: signal is true;
	signal G22101: std_logic; attribute dont_touch of G22101: signal is true;
	signal G22102: std_logic; attribute dont_touch of G22102: signal is true;
	signal G22103: std_logic; attribute dont_touch of G22103: signal is true;
	signal G22104: std_logic; attribute dont_touch of G22104: signal is true;
	signal G22105: std_logic; attribute dont_touch of G22105: signal is true;
	signal G22106: std_logic; attribute dont_touch of G22106: signal is true;
	signal G22107: std_logic; attribute dont_touch of G22107: signal is true;
	signal G22108: std_logic; attribute dont_touch of G22108: signal is true;
	signal G22112: std_logic; attribute dont_touch of G22112: signal is true;
	signal G22113: std_logic; attribute dont_touch of G22113: signal is true;
	signal G22114: std_logic; attribute dont_touch of G22114: signal is true;
	signal G22115: std_logic; attribute dont_touch of G22115: signal is true;
	signal G22116: std_logic; attribute dont_touch of G22116: signal is true;
	signal G22117: std_logic; attribute dont_touch of G22117: signal is true;
	signal G22118: std_logic; attribute dont_touch of G22118: signal is true;
	signal G22122: std_logic; attribute dont_touch of G22122: signal is true;
	signal G22123: std_logic; attribute dont_touch of G22123: signal is true;
	signal G22124: std_logic; attribute dont_touch of G22124: signal is true;
	signal G22125: std_logic; attribute dont_touch of G22125: signal is true;
	signal G22126: std_logic; attribute dont_touch of G22126: signal is true;
	signal G22127: std_logic; attribute dont_touch of G22127: signal is true;
	signal G22128: std_logic; attribute dont_touch of G22128: signal is true;
	signal G22129: std_logic; attribute dont_touch of G22129: signal is true;
	signal G22130: std_logic; attribute dont_touch of G22130: signal is true;
	signal G22131: std_logic; attribute dont_touch of G22131: signal is true;
	signal G22132: std_logic; attribute dont_touch of G22132: signal is true;
	signal G22133: std_logic; attribute dont_touch of G22133: signal is true;
	signal G22134: std_logic; attribute dont_touch of G22134: signal is true;
	signal G22138: std_logic; attribute dont_touch of G22138: signal is true;
	signal G22139: std_logic; attribute dont_touch of G22139: signal is true;
	signal G22140: std_logic; attribute dont_touch of G22140: signal is true;
	signal G22141: std_logic; attribute dont_touch of G22141: signal is true;
	signal G22142: std_logic; attribute dont_touch of G22142: signal is true;
	signal G22143: std_logic; attribute dont_touch of G22143: signal is true;
	signal G22144: std_logic; attribute dont_touch of G22144: signal is true;
	signal G22145: std_logic; attribute dont_touch of G22145: signal is true;
	signal G22146: std_logic; attribute dont_touch of G22146: signal is true;
	signal G22147: std_logic; attribute dont_touch of G22147: signal is true;
	signal G22148: std_logic; attribute dont_touch of G22148: signal is true;
	signal G22149: std_logic; attribute dont_touch of G22149: signal is true;
	signal G22150: std_logic; attribute dont_touch of G22150: signal is true;
	signal G22151: std_logic; attribute dont_touch of G22151: signal is true;
	signal G22152: std_logic; attribute dont_touch of G22152: signal is true;
	signal G22153: std_logic; attribute dont_touch of G22153: signal is true;
	signal G22154: std_logic; attribute dont_touch of G22154: signal is true;
	signal G22155: std_logic; attribute dont_touch of G22155: signal is true;
	signal G22156: std_logic; attribute dont_touch of G22156: signal is true;
	signal G22157: std_logic; attribute dont_touch of G22157: signal is true;
	signal G22161: std_logic; attribute dont_touch of G22161: signal is true;
	signal G22162: std_logic; attribute dont_touch of G22162: signal is true;
	signal G22163: std_logic; attribute dont_touch of G22163: signal is true;
	signal G22164: std_logic; attribute dont_touch of G22164: signal is true;
	signal G22165: std_logic; attribute dont_touch of G22165: signal is true;
	signal G22166: std_logic; attribute dont_touch of G22166: signal is true;
	signal G22167: std_logic; attribute dont_touch of G22167: signal is true;
	signal G22168: std_logic; attribute dont_touch of G22168: signal is true;
	signal G22169: std_logic; attribute dont_touch of G22169: signal is true;
	signal G22170: std_logic; attribute dont_touch of G22170: signal is true;
	signal G22171: std_logic; attribute dont_touch of G22171: signal is true;
	signal G22172: std_logic; attribute dont_touch of G22172: signal is true;
	signal G22173: std_logic; attribute dont_touch of G22173: signal is true;
	signal G22174: std_logic; attribute dont_touch of G22174: signal is true;
	signal G22175: std_logic; attribute dont_touch of G22175: signal is true;
	signal G22176: std_logic; attribute dont_touch of G22176: signal is true;
	signal G22177: std_logic; attribute dont_touch of G22177: signal is true;
	signal G22178: std_logic; attribute dont_touch of G22178: signal is true;
	signal G22179: std_logic; attribute dont_touch of G22179: signal is true;
	signal G22180: std_logic; attribute dont_touch of G22180: signal is true;
	signal G22181: std_logic; attribute dont_touch of G22181: signal is true;
	signal G22182: std_logic; attribute dont_touch of G22182: signal is true;
	signal G22183: std_logic; attribute dont_touch of G22183: signal is true;
	signal G22184: std_logic; attribute dont_touch of G22184: signal is true;
	signal G22185: std_logic; attribute dont_touch of G22185: signal is true;
	signal G22186: std_logic; attribute dont_touch of G22186: signal is true;
	signal G22187: std_logic; attribute dont_touch of G22187: signal is true;
	signal G22188: std_logic; attribute dont_touch of G22188: signal is true;
	signal G22189: std_logic; attribute dont_touch of G22189: signal is true;
	signal G22190: std_logic; attribute dont_touch of G22190: signal is true;
	signal G22191: std_logic; attribute dont_touch of G22191: signal is true;
	signal G22192: std_logic; attribute dont_touch of G22192: signal is true;
	signal G22193: std_logic; attribute dont_touch of G22193: signal is true;
	signal G22194: std_logic; attribute dont_touch of G22194: signal is true;
	signal G22195: std_logic; attribute dont_touch of G22195: signal is true;
	signal G22196: std_logic; attribute dont_touch of G22196: signal is true;
	signal G22197: std_logic; attribute dont_touch of G22197: signal is true;
	signal G22198: std_logic; attribute dont_touch of G22198: signal is true;
	signal G22199: std_logic; attribute dont_touch of G22199: signal is true;
	signal G22200: std_logic; attribute dont_touch of G22200: signal is true;
	signal G22201: std_logic; attribute dont_touch of G22201: signal is true;
	signal G22202: std_logic; attribute dont_touch of G22202: signal is true;
	signal G22203: std_logic; attribute dont_touch of G22203: signal is true;
	signal G22204: std_logic; attribute dont_touch of G22204: signal is true;
	signal G22205: std_logic; attribute dont_touch of G22205: signal is true;
	signal G22206: std_logic; attribute dont_touch of G22206: signal is true;
	signal G22207: std_logic; attribute dont_touch of G22207: signal is true;
	signal G22208: std_logic; attribute dont_touch of G22208: signal is true;
	signal G22209: std_logic; attribute dont_touch of G22209: signal is true;
	signal G22210: std_logic; attribute dont_touch of G22210: signal is true;
	signal G22211: std_logic; attribute dont_touch of G22211: signal is true;
	signal G22212: std_logic; attribute dont_touch of G22212: signal is true;
	signal G22213: std_logic; attribute dont_touch of G22213: signal is true;
	signal G22214: std_logic; attribute dont_touch of G22214: signal is true;
	signal G22215: std_logic; attribute dont_touch of G22215: signal is true;
	signal G22216: std_logic; attribute dont_touch of G22216: signal is true;
	signal G22217: std_logic; attribute dont_touch of G22217: signal is true;
	signal G22218: std_logic; attribute dont_touch of G22218: signal is true;
	signal G22219: std_logic; attribute dont_touch of G22219: signal is true;
	signal G22220: std_logic; attribute dont_touch of G22220: signal is true;
	signal G22221: std_logic; attribute dont_touch of G22221: signal is true;
	signal G22222: std_logic; attribute dont_touch of G22222: signal is true;
	signal G22223: std_logic; attribute dont_touch of G22223: signal is true;
	signal G22224: std_logic; attribute dont_touch of G22224: signal is true;
	signal G22225: std_logic; attribute dont_touch of G22225: signal is true;
	signal G22226: std_logic; attribute dont_touch of G22226: signal is true;
	signal G22227: std_logic; attribute dont_touch of G22227: signal is true;
	signal G22228: std_logic; attribute dont_touch of G22228: signal is true;
	signal G22229: std_logic; attribute dont_touch of G22229: signal is true;
	signal G22230: std_logic; attribute dont_touch of G22230: signal is true;
	signal G22231: std_logic; attribute dont_touch of G22231: signal is true;
	signal G22232: std_logic; attribute dont_touch of G22232: signal is true;
	signal G22233: std_logic; attribute dont_touch of G22233: signal is true;
	signal G22234: std_logic; attribute dont_touch of G22234: signal is true;
	signal G22235: std_logic; attribute dont_touch of G22235: signal is true;
	signal G22236: std_logic; attribute dont_touch of G22236: signal is true;
	signal G22237: std_logic; attribute dont_touch of G22237: signal is true;
	signal G22238: std_logic; attribute dont_touch of G22238: signal is true;
	signal G22239: std_logic; attribute dont_touch of G22239: signal is true;
	signal G22240: std_logic; attribute dont_touch of G22240: signal is true;
	signal G22241: std_logic; attribute dont_touch of G22241: signal is true;
	signal G22242: std_logic; attribute dont_touch of G22242: signal is true;
	signal G22243: std_logic; attribute dont_touch of G22243: signal is true;
	signal G22244: std_logic; attribute dont_touch of G22244: signal is true;
	signal G22245: std_logic; attribute dont_touch of G22245: signal is true;
	signal G22246: std_logic; attribute dont_touch of G22246: signal is true;
	signal G22247: std_logic; attribute dont_touch of G22247: signal is true;
	signal G22248: std_logic; attribute dont_touch of G22248: signal is true;
	signal G22249: std_logic; attribute dont_touch of G22249: signal is true;
	signal G22250: std_logic; attribute dont_touch of G22250: signal is true;
	signal G22251: std_logic; attribute dont_touch of G22251: signal is true;
	signal G22252: std_logic; attribute dont_touch of G22252: signal is true;
	signal G22253: std_logic; attribute dont_touch of G22253: signal is true;
	signal G22254: std_logic; attribute dont_touch of G22254: signal is true;
	signal G22255: std_logic; attribute dont_touch of G22255: signal is true;
	signal G22256: std_logic; attribute dont_touch of G22256: signal is true;
	signal G22257: std_logic; attribute dont_touch of G22257: signal is true;
	signal G22258: std_logic; attribute dont_touch of G22258: signal is true;
	signal G22259: std_logic; attribute dont_touch of G22259: signal is true;
	signal G22260: std_logic; attribute dont_touch of G22260: signal is true;
	signal G22261: std_logic; attribute dont_touch of G22261: signal is true;
	signal G22262: std_logic; attribute dont_touch of G22262: signal is true;
	signal G22263: std_logic; attribute dont_touch of G22263: signal is true;
	signal G22264: std_logic; attribute dont_touch of G22264: signal is true;
	signal G22265: std_logic; attribute dont_touch of G22265: signal is true;
	signal G22266: std_logic; attribute dont_touch of G22266: signal is true;
	signal G22267: std_logic; attribute dont_touch of G22267: signal is true;
	signal G22268: std_logic; attribute dont_touch of G22268: signal is true;
	signal G22269: std_logic; attribute dont_touch of G22269: signal is true;
	signal G22270: std_logic; attribute dont_touch of G22270: signal is true;
	signal G22271: std_logic; attribute dont_touch of G22271: signal is true;
	signal G22272: std_logic; attribute dont_touch of G22272: signal is true;
	signal G22273: std_logic; attribute dont_touch of G22273: signal is true;
	signal G22274: std_logic; attribute dont_touch of G22274: signal is true;
	signal G22275: std_logic; attribute dont_touch of G22275: signal is true;
	signal G22276: std_logic; attribute dont_touch of G22276: signal is true;
	signal G22277: std_logic; attribute dont_touch of G22277: signal is true;
	signal G22278: std_logic; attribute dont_touch of G22278: signal is true;
	signal G22279: std_logic; attribute dont_touch of G22279: signal is true;
	signal G22280: std_logic; attribute dont_touch of G22280: signal is true;
	signal G22281: std_logic; attribute dont_touch of G22281: signal is true;
	signal G22282: std_logic; attribute dont_touch of G22282: signal is true;
	signal G22283: std_logic; attribute dont_touch of G22283: signal is true;
	signal G22284: std_logic; attribute dont_touch of G22284: signal is true;
	signal G22285: std_logic; attribute dont_touch of G22285: signal is true;
	signal G22286: std_logic; attribute dont_touch of G22286: signal is true;
	signal G22287: std_logic; attribute dont_touch of G22287: signal is true;
	signal G22288: std_logic; attribute dont_touch of G22288: signal is true;
	signal G22289: std_logic; attribute dont_touch of G22289: signal is true;
	signal G22290: std_logic; attribute dont_touch of G22290: signal is true;
	signal G22291: std_logic; attribute dont_touch of G22291: signal is true;
	signal G22292: std_logic; attribute dont_touch of G22292: signal is true;
	signal G22293: std_logic; attribute dont_touch of G22293: signal is true;
	signal G22294: std_logic; attribute dont_touch of G22294: signal is true;
	signal G22295: std_logic; attribute dont_touch of G22295: signal is true;
	signal G22296: std_logic; attribute dont_touch of G22296: signal is true;
	signal G22297: std_logic; attribute dont_touch of G22297: signal is true;
	signal G22298: std_logic; attribute dont_touch of G22298: signal is true;
	signal G22299: std_logic; attribute dont_touch of G22299: signal is true;
	signal G22300: std_logic; attribute dont_touch of G22300: signal is true;
	signal G22303: std_logic; attribute dont_touch of G22303: signal is true;
	signal G22304: std_logic; attribute dont_touch of G22304: signal is true;
	signal G22305: std_logic; attribute dont_touch of G22305: signal is true;
	signal G22306: std_logic; attribute dont_touch of G22306: signal is true;
	signal G22307: std_logic; attribute dont_touch of G22307: signal is true;
	signal G22308: std_logic; attribute dont_touch of G22308: signal is true;
	signal G22309: std_logic; attribute dont_touch of G22309: signal is true;
	signal G22310: std_logic; attribute dont_touch of G22310: signal is true;
	signal G22311: std_logic; attribute dont_touch of G22311: signal is true;
	signal G22312: std_logic; attribute dont_touch of G22312: signal is true;
	signal G22313: std_logic; attribute dont_touch of G22313: signal is true;
	signal G22314: std_logic; attribute dont_touch of G22314: signal is true;
	signal G22315: std_logic; attribute dont_touch of G22315: signal is true;
	signal G22316: std_logic; attribute dont_touch of G22316: signal is true;
	signal G22317: std_logic; attribute dont_touch of G22317: signal is true;
	signal G22318: std_logic; attribute dont_touch of G22318: signal is true;
	signal G22319: std_logic; attribute dont_touch of G22319: signal is true;
	signal G22328: std_logic; attribute dont_touch of G22328: signal is true;
	signal G22331: std_logic; attribute dont_touch of G22331: signal is true;
	signal G22332: std_logic; attribute dont_touch of G22332: signal is true;
	signal G22333: std_logic; attribute dont_touch of G22333: signal is true;
	signal G22334: std_logic; attribute dont_touch of G22334: signal is true;
	signal G22335: std_logic; attribute dont_touch of G22335: signal is true;
	signal G22336: std_logic; attribute dont_touch of G22336: signal is true;
	signal G22337: std_logic; attribute dont_touch of G22337: signal is true;
	signal G22338: std_logic; attribute dont_touch of G22338: signal is true;
	signal G22339: std_logic; attribute dont_touch of G22339: signal is true;
	signal G22340: std_logic; attribute dont_touch of G22340: signal is true;
	signal G22341: std_logic; attribute dont_touch of G22341: signal is true;
	signal G22342: std_logic; attribute dont_touch of G22342: signal is true;
	signal G22343: std_logic; attribute dont_touch of G22343: signal is true;
	signal G22344: std_logic; attribute dont_touch of G22344: signal is true;
	signal G22353: std_logic; attribute dont_touch of G22353: signal is true;
	signal G22356: std_logic; attribute dont_touch of G22356: signal is true;
	signal G22357: std_logic; attribute dont_touch of G22357: signal is true;
	signal G22358: std_logic; attribute dont_touch of G22358: signal is true;
	signal G22359: std_logic; attribute dont_touch of G22359: signal is true;
	signal G22360: std_logic; attribute dont_touch of G22360: signal is true;
	signal G22361: std_logic; attribute dont_touch of G22361: signal is true;
	signal G22362: std_logic; attribute dont_touch of G22362: signal is true;
	signal G22363: std_logic; attribute dont_touch of G22363: signal is true;
	signal G22364: std_logic; attribute dont_touch of G22364: signal is true;
	signal G22365: std_logic; attribute dont_touch of G22365: signal is true;
	signal G22366: std_logic; attribute dont_touch of G22366: signal is true;
	signal G22367: std_logic; attribute dont_touch of G22367: signal is true;
	signal G22376: std_logic; attribute dont_touch of G22376: signal is true;
	signal G22379: std_logic; attribute dont_touch of G22379: signal is true;
	signal G22380: std_logic; attribute dont_touch of G22380: signal is true;
	signal G22381: std_logic; attribute dont_touch of G22381: signal is true;
	signal G22382: std_logic; attribute dont_touch of G22382: signal is true;
	signal G22383: std_logic; attribute dont_touch of G22383: signal is true;
	signal G22384: std_logic; attribute dont_touch of G22384: signal is true;
	signal G22385: std_logic; attribute dont_touch of G22385: signal is true;
	signal G22386: std_logic; attribute dont_touch of G22386: signal is true;
	signal G22387: std_logic; attribute dont_touch of G22387: signal is true;
	signal G22396: std_logic; attribute dont_touch of G22396: signal is true;
	signal G22397: std_logic; attribute dont_touch of G22397: signal is true;
	signal G22398: std_logic; attribute dont_touch of G22398: signal is true;
	signal G22399: std_logic; attribute dont_touch of G22399: signal is true;
	signal G22400: std_logic; attribute dont_touch of G22400: signal is true;
	signal G22401: std_logic; attribute dont_touch of G22401: signal is true;
	signal G22402: std_logic; attribute dont_touch of G22402: signal is true;
	signal G22403: std_logic; attribute dont_touch of G22403: signal is true;
	signal G22404: std_logic; attribute dont_touch of G22404: signal is true;
	signal G22405: std_logic; attribute dont_touch of G22405: signal is true;
	signal G22408: std_logic; attribute dont_touch of G22408: signal is true;
	signal G22409: std_logic; attribute dont_touch of G22409: signal is true;
	signal G22412: std_logic; attribute dont_touch of G22412: signal is true;
	signal G22415: std_logic; attribute dont_touch of G22415: signal is true;
	signal G22418: std_logic; attribute dont_touch of G22418: signal is true;
	signal G22421: std_logic; attribute dont_touch of G22421: signal is true;
	signal G22422: std_logic; attribute dont_touch of G22422: signal is true;
	signal G22425: std_logic; attribute dont_touch of G22425: signal is true;
	signal G22428: std_logic; attribute dont_touch of G22428: signal is true;
	signal G22431: std_logic; attribute dont_touch of G22431: signal is true;
	signal G22434: std_logic; attribute dont_touch of G22434: signal is true;
	signal G22437: std_logic; attribute dont_touch of G22437: signal is true;
	signal G22440: std_logic; attribute dont_touch of G22440: signal is true;
	signal G22443: std_logic; attribute dont_touch of G22443: signal is true;
	signal G22444: std_logic; attribute dont_touch of G22444: signal is true;
	signal G22445: std_logic; attribute dont_touch of G22445: signal is true;
	signal G22448: std_logic; attribute dont_touch of G22448: signal is true;
	signal G22451: std_logic; attribute dont_touch of G22451: signal is true;
	signal G22454: std_logic; attribute dont_touch of G22454: signal is true;
	signal G22455: std_logic; attribute dont_touch of G22455: signal is true;
	signal G22458: std_logic; attribute dont_touch of G22458: signal is true;
	signal G22461: std_logic; attribute dont_touch of G22461: signal is true;
	signal G22464: std_logic; attribute dont_touch of G22464: signal is true;
	signal G22467: std_logic; attribute dont_touch of G22467: signal is true;
	signal G22470: std_logic; attribute dont_touch of G22470: signal is true;
	signal G22473: std_logic; attribute dont_touch of G22473: signal is true;
	signal G22476: std_logic; attribute dont_touch of G22476: signal is true;
	signal G22477: std_logic; attribute dont_touch of G22477: signal is true;
	signal G22480: std_logic; attribute dont_touch of G22480: signal is true;
	signal G22483: std_logic; attribute dont_touch of G22483: signal is true;
	signal G22484: std_logic; attribute dont_touch of G22484: signal is true;
	signal G22487: std_logic; attribute dont_touch of G22487: signal is true;
	signal G22490: std_logic; attribute dont_touch of G22490: signal is true;
	signal G22493: std_logic; attribute dont_touch of G22493: signal is true;
	signal G22494: std_logic; attribute dont_touch of G22494: signal is true;
	signal G22497: std_logic; attribute dont_touch of G22497: signal is true;
	signal G22500: std_logic; attribute dont_touch of G22500: signal is true;
	signal G22503: std_logic; attribute dont_touch of G22503: signal is true;
	signal G22506: std_logic; attribute dont_touch of G22506: signal is true;
	signal G22509: std_logic; attribute dont_touch of G22509: signal is true;
	signal G22512: std_logic; attribute dont_touch of G22512: signal is true;
	signal G22515: std_logic; attribute dont_touch of G22515: signal is true;
	signal G22516: std_logic; attribute dont_touch of G22516: signal is true;
	signal G22517: std_logic; attribute dont_touch of G22517: signal is true;
	signal G22518: std_logic; attribute dont_touch of G22518: signal is true;
	signal G22519: std_logic; attribute dont_touch of G22519: signal is true;
	signal G22520: std_logic; attribute dont_touch of G22520: signal is true;
	signal G22523: std_logic; attribute dont_touch of G22523: signal is true;
	signal G22526: std_logic; attribute dont_touch of G22526: signal is true;
	signal G22527: std_logic; attribute dont_touch of G22527: signal is true;
	signal G22530: std_logic; attribute dont_touch of G22530: signal is true;
	signal G22533: std_logic; attribute dont_touch of G22533: signal is true;
	signal G22536: std_logic; attribute dont_touch of G22536: signal is true;
	signal G22537: std_logic; attribute dont_touch of G22537: signal is true;
	signal G22540: std_logic; attribute dont_touch of G22540: signal is true;
	signal G22543: std_logic; attribute dont_touch of G22543: signal is true;
	signal G22546: std_logic; attribute dont_touch of G22546: signal is true;
	signal G22547: std_logic; attribute dont_touch of G22547: signal is true;
	signal G22548: std_logic; attribute dont_touch of G22548: signal is true;
	signal G22549: std_logic; attribute dont_touch of G22549: signal is true;
	signal G22550: std_logic; attribute dont_touch of G22550: signal is true;
	signal G22551: std_logic; attribute dont_touch of G22551: signal is true;
	signal G22552: std_logic; attribute dont_touch of G22552: signal is true;
	signal G22555: std_logic; attribute dont_touch of G22555: signal is true;
	signal G22556: std_logic; attribute dont_touch of G22556: signal is true;
	signal G22557: std_logic; attribute dont_touch of G22557: signal is true;
	signal G22558: std_logic; attribute dont_touch of G22558: signal is true;
	signal G22559: std_logic; attribute dont_touch of G22559: signal is true;
	signal G22560: std_logic; attribute dont_touch of G22560: signal is true;
	signal G22563: std_logic; attribute dont_touch of G22563: signal is true;
	signal G22566: std_logic; attribute dont_touch of G22566: signal is true;
	signal G22567: std_logic; attribute dont_touch of G22567: signal is true;
	signal G22570: std_logic; attribute dont_touch of G22570: signal is true;
	signal G22573: std_logic; attribute dont_touch of G22573: signal is true;
	signal G22576: std_logic; attribute dont_touch of G22576: signal is true;
	signal G22577: std_logic; attribute dont_touch of G22577: signal is true;
	signal G22578: std_logic; attribute dont_touch of G22578: signal is true;
	signal G22581: std_logic; attribute dont_touch of G22581: signal is true;
	signal G22582: std_logic; attribute dont_touch of G22582: signal is true;
	signal G22583: std_logic; attribute dont_touch of G22583: signal is true;
	signal G22584: std_logic; attribute dont_touch of G22584: signal is true;
	signal G22585: std_logic; attribute dont_touch of G22585: signal is true;
	signal G22586: std_logic; attribute dont_touch of G22586: signal is true;
	signal G22587: std_logic; attribute dont_touch of G22587: signal is true;
	signal G22588: std_logic; attribute dont_touch of G22588: signal is true;
	signal G22589: std_logic; attribute dont_touch of G22589: signal is true;
	signal G22590: std_logic; attribute dont_touch of G22590: signal is true;
	signal G22591: std_logic; attribute dont_touch of G22591: signal is true;
	signal G22592: std_logic; attribute dont_touch of G22592: signal is true;
	signal G22595: std_logic; attribute dont_touch of G22595: signal is true;
	signal G22596: std_logic; attribute dont_touch of G22596: signal is true;
	signal G22597: std_logic; attribute dont_touch of G22597: signal is true;
	signal G22598: std_logic; attribute dont_touch of G22598: signal is true;
	signal G22599: std_logic; attribute dont_touch of G22599: signal is true;
	signal G22600: std_logic; attribute dont_touch of G22600: signal is true;
	signal G22603: std_logic; attribute dont_touch of G22603: signal is true;
	signal G22606: std_logic; attribute dont_touch of G22606: signal is true;
	signal G22607: std_logic; attribute dont_touch of G22607: signal is true;
	signal G22608: std_logic; attribute dont_touch of G22608: signal is true;
	signal G22609: std_logic; attribute dont_touch of G22609: signal is true;
	signal G22610: std_logic; attribute dont_touch of G22610: signal is true;
	signal G22611: std_logic; attribute dont_touch of G22611: signal is true;
	signal G22612: std_logic; attribute dont_touch of G22612: signal is true;
	signal G22613: std_logic; attribute dont_touch of G22613: signal is true;
	signal G22614: std_logic; attribute dont_touch of G22614: signal is true;
	signal G22615: std_logic; attribute dont_touch of G22615: signal is true;
	signal G22618: std_logic; attribute dont_touch of G22618: signal is true;
	signal G22619: std_logic; attribute dont_touch of G22619: signal is true;
	signal G22620: std_logic; attribute dont_touch of G22620: signal is true;
	signal G22621: std_logic; attribute dont_touch of G22621: signal is true;
	signal G22622: std_logic; attribute dont_touch of G22622: signal is true;
	signal G22623: std_logic; attribute dont_touch of G22623: signal is true;
	signal G22624: std_logic; attribute dont_touch of G22624: signal is true;
	signal G22625: std_logic; attribute dont_touch of G22625: signal is true;
	signal G22626: std_logic; attribute dont_touch of G22626: signal is true;
	signal G22627: std_logic; attribute dont_touch of G22627: signal is true;
	signal G22628: std_logic; attribute dont_touch of G22628: signal is true;
	signal G22629: std_logic; attribute dont_touch of G22629: signal is true;
	signal G22632: std_logic; attribute dont_touch of G22632: signal is true;
	signal G22633: std_logic; attribute dont_touch of G22633: signal is true;
	signal G22634: std_logic; attribute dont_touch of G22634: signal is true;
	signal G22635: std_logic; attribute dont_touch of G22635: signal is true;
	signal G22636: std_logic; attribute dont_touch of G22636: signal is true;
	signal G22637: std_logic; attribute dont_touch of G22637: signal is true;
	signal G22638: std_logic; attribute dont_touch of G22638: signal is true;
	signal G22639: std_logic; attribute dont_touch of G22639: signal is true;
	signal G22640: std_logic; attribute dont_touch of G22640: signal is true;
	signal G22641: std_logic; attribute dont_touch of G22641: signal is true;
	signal G22642: std_logic; attribute dont_touch of G22642: signal is true;
	signal G22643: std_logic; attribute dont_touch of G22643: signal is true;
	signal G22644: std_logic; attribute dont_touch of G22644: signal is true;
	signal G22645: std_logic; attribute dont_touch of G22645: signal is true;
	signal G22646: std_logic; attribute dont_touch of G22646: signal is true;
	signal G22647: std_logic; attribute dont_touch of G22647: signal is true;
	signal G22648: std_logic; attribute dont_touch of G22648: signal is true;
	signal G22649: std_logic; attribute dont_touch of G22649: signal is true;
	signal G22650: std_logic; attribute dont_touch of G22650: signal is true;
	signal G22651: std_logic; attribute dont_touch of G22651: signal is true;
	signal G22654: std_logic; attribute dont_touch of G22654: signal is true;
	signal G22655: std_logic; attribute dont_touch of G22655: signal is true;
	signal G22656: std_logic; attribute dont_touch of G22656: signal is true;
	signal G22657: std_logic; attribute dont_touch of G22657: signal is true;
	signal G22658: std_logic; attribute dont_touch of G22658: signal is true;
	signal G22659: std_logic; attribute dont_touch of G22659: signal is true;
	signal G22660: std_logic; attribute dont_touch of G22660: signal is true;
	signal G22661: std_logic; attribute dont_touch of G22661: signal is true;
	signal G22662: std_logic; attribute dont_touch of G22662: signal is true;
	signal G22663: std_logic; attribute dont_touch of G22663: signal is true;
	signal G22664: std_logic; attribute dont_touch of G22664: signal is true;
	signal G22665: std_logic; attribute dont_touch of G22665: signal is true;
	signal G22666: std_logic; attribute dont_touch of G22666: signal is true;
	signal G22667: std_logic; attribute dont_touch of G22667: signal is true;
	signal G22668: std_logic; attribute dont_touch of G22668: signal is true;
	signal G22669: std_logic; attribute dont_touch of G22669: signal is true;
	signal G22670: std_logic; attribute dont_touch of G22670: signal is true;
	signal G22671: std_logic; attribute dont_touch of G22671: signal is true;
	signal G22672: std_logic; attribute dont_touch of G22672: signal is true;
	signal G22673: std_logic; attribute dont_touch of G22673: signal is true;
	signal G22674: std_logic; attribute dont_touch of G22674: signal is true;
	signal G22675: std_logic; attribute dont_touch of G22675: signal is true;
	signal G22676: std_logic; attribute dont_touch of G22676: signal is true;
	signal G22677: std_logic; attribute dont_touch of G22677: signal is true;
	signal G22678: std_logic; attribute dont_touch of G22678: signal is true;
	signal G22679: std_logic; attribute dont_touch of G22679: signal is true;
	signal G22680: std_logic; attribute dont_touch of G22680: signal is true;
	signal G22681: std_logic; attribute dont_touch of G22681: signal is true;
	signal G22682: std_logic; attribute dont_touch of G22682: signal is true;
	signal G22683: std_logic; attribute dont_touch of G22683: signal is true;
	signal G22684: std_logic; attribute dont_touch of G22684: signal is true;
	signal G22685: std_logic; attribute dont_touch of G22685: signal is true;
	signal G22686: std_logic; attribute dont_touch of G22686: signal is true;
	signal G22687: std_logic; attribute dont_touch of G22687: signal is true;
	signal G22690: std_logic; attribute dont_touch of G22690: signal is true;
	signal G22691: std_logic; attribute dont_touch of G22691: signal is true;
	signal G22692: std_logic; attribute dont_touch of G22692: signal is true;
	signal G22693: std_logic; attribute dont_touch of G22693: signal is true;
	signal G22694: std_logic; attribute dont_touch of G22694: signal is true;
	signal G22695: std_logic; attribute dont_touch of G22695: signal is true;
	signal G22696: std_logic; attribute dont_touch of G22696: signal is true;
	signal G22699: std_logic; attribute dont_touch of G22699: signal is true;
	signal G22700: std_logic; attribute dont_touch of G22700: signal is true;
	signal G22701: std_logic; attribute dont_touch of G22701: signal is true;
	signal G22702: std_logic; attribute dont_touch of G22702: signal is true;
	signal G22703: std_logic; attribute dont_touch of G22703: signal is true;
	signal G22704: std_logic; attribute dont_touch of G22704: signal is true;
	signal G22705: std_logic; attribute dont_touch of G22705: signal is true;
	signal G22706: std_logic; attribute dont_touch of G22706: signal is true;
	signal G22707: std_logic; attribute dont_touch of G22707: signal is true;
	signal G22708: std_logic; attribute dont_touch of G22708: signal is true;
	signal G22709: std_logic; attribute dont_touch of G22709: signal is true;
	signal G22710: std_logic; attribute dont_touch of G22710: signal is true;
	signal G22711: std_logic; attribute dont_touch of G22711: signal is true;
	signal G22712: std_logic; attribute dont_touch of G22712: signal is true;
	signal G22713: std_logic; attribute dont_touch of G22713: signal is true;
	signal G22714: std_logic; attribute dont_touch of G22714: signal is true;
	signal G22715: std_logic; attribute dont_touch of G22715: signal is true;
	signal G22716: std_logic; attribute dont_touch of G22716: signal is true;
	signal G22717: std_logic; attribute dont_touch of G22717: signal is true;
	signal G22718: std_logic; attribute dont_touch of G22718: signal is true;
	signal G22719: std_logic; attribute dont_touch of G22719: signal is true;
	signal G22720: std_logic; attribute dont_touch of G22720: signal is true;
	signal G22721: std_logic; attribute dont_touch of G22721: signal is true;
	signal G22722: std_logic; attribute dont_touch of G22722: signal is true;
	signal G22723: std_logic; attribute dont_touch of G22723: signal is true;
	signal G22724: std_logic; attribute dont_touch of G22724: signal is true;
	signal G22725: std_logic; attribute dont_touch of G22725: signal is true;
	signal G22726: std_logic; attribute dont_touch of G22726: signal is true;
	signal G22727: std_logic; attribute dont_touch of G22727: signal is true;
	signal G22728: std_logic; attribute dont_touch of G22728: signal is true;
	signal G22729: std_logic; attribute dont_touch of G22729: signal is true;
	signal G22730: std_logic; attribute dont_touch of G22730: signal is true;
	signal G22731: std_logic; attribute dont_touch of G22731: signal is true;
	signal G22732: std_logic; attribute dont_touch of G22732: signal is true;
	signal G22733: std_logic; attribute dont_touch of G22733: signal is true;
	signal G22734: std_logic; attribute dont_touch of G22734: signal is true;
	signal G22735: std_logic; attribute dont_touch of G22735: signal is true;
	signal G22736: std_logic; attribute dont_touch of G22736: signal is true;
	signal G22737: std_logic; attribute dont_touch of G22737: signal is true;
	signal G22738: std_logic; attribute dont_touch of G22738: signal is true;
	signal G22739: std_logic; attribute dont_touch of G22739: signal is true;
	signal G22740: std_logic; attribute dont_touch of G22740: signal is true;
	signal G22741: std_logic; attribute dont_touch of G22741: signal is true;
	signal G22742: std_logic; attribute dont_touch of G22742: signal is true;
	signal G22743: std_logic; attribute dont_touch of G22743: signal is true;
	signal G22744: std_logic; attribute dont_touch of G22744: signal is true;
	signal G22745: std_logic; attribute dont_touch of G22745: signal is true;
	signal G22746: std_logic; attribute dont_touch of G22746: signal is true;
	signal G22747: std_logic; attribute dont_touch of G22747: signal is true;
	signal G22748: std_logic; attribute dont_touch of G22748: signal is true;
	signal G22749: std_logic; attribute dont_touch of G22749: signal is true;
	signal G22750: std_logic; attribute dont_touch of G22750: signal is true;
	signal G22753: std_logic; attribute dont_touch of G22753: signal is true;
	signal G22754: std_logic; attribute dont_touch of G22754: signal is true;
	signal G22755: std_logic; attribute dont_touch of G22755: signal is true;
	signal G22756: std_logic; attribute dont_touch of G22756: signal is true;
	signal G22757: std_logic; attribute dont_touch of G22757: signal is true;
	signal G22758: std_logic; attribute dont_touch of G22758: signal is true;
	signal G22759: std_logic; attribute dont_touch of G22759: signal is true;
	signal G22760: std_logic; attribute dont_touch of G22760: signal is true;
	signal G22761: std_logic; attribute dont_touch of G22761: signal is true;
	signal G22762: std_logic; attribute dont_touch of G22762: signal is true;
	signal G22763: std_logic; attribute dont_touch of G22763: signal is true;
	signal G22764: std_logic; attribute dont_touch of G22764: signal is true;
	signal G22765: std_logic; attribute dont_touch of G22765: signal is true;
	signal G22766: std_logic; attribute dont_touch of G22766: signal is true;
	signal G22767: std_logic; attribute dont_touch of G22767: signal is true;
	signal G22768: std_logic; attribute dont_touch of G22768: signal is true;
	signal G22769: std_logic; attribute dont_touch of G22769: signal is true;
	signal G22770: std_logic; attribute dont_touch of G22770: signal is true;
	signal G22771: std_logic; attribute dont_touch of G22771: signal is true;
	signal G22772: std_logic; attribute dont_touch of G22772: signal is true;
	signal G22773: std_logic; attribute dont_touch of G22773: signal is true;
	signal G22774: std_logic; attribute dont_touch of G22774: signal is true;
	signal G22775: std_logic; attribute dont_touch of G22775: signal is true;
	signal G22776: std_logic; attribute dont_touch of G22776: signal is true;
	signal G22777: std_logic; attribute dont_touch of G22777: signal is true;
	signal G22784: std_logic; attribute dont_touch of G22784: signal is true;
	signal G22785: std_logic; attribute dont_touch of G22785: signal is true;
	signal G22786: std_logic; attribute dont_touch of G22786: signal is true;
	signal G22787: std_logic; attribute dont_touch of G22787: signal is true;
	signal G22788: std_logic; attribute dont_touch of G22788: signal is true;
	signal G22789: std_logic; attribute dont_touch of G22789: signal is true;
	signal G22790: std_logic; attribute dont_touch of G22790: signal is true;
	signal G22791: std_logic; attribute dont_touch of G22791: signal is true;
	signal G22792: std_logic; attribute dont_touch of G22792: signal is true;
	signal G22793: std_logic; attribute dont_touch of G22793: signal is true;
	signal G22794: std_logic; attribute dont_touch of G22794: signal is true;
	signal G22795: std_logic; attribute dont_touch of G22795: signal is true;
	signal G22796: std_logic; attribute dont_touch of G22796: signal is true;
	signal G22797: std_logic; attribute dont_touch of G22797: signal is true;
	signal G22798: std_logic; attribute dont_touch of G22798: signal is true;
	signal G22799: std_logic; attribute dont_touch of G22799: signal is true;
	signal G22800: std_logic; attribute dont_touch of G22800: signal is true;
	signal G22801: std_logic; attribute dont_touch of G22801: signal is true;
	signal G22802: std_logic; attribute dont_touch of G22802: signal is true;
	signal G22803: std_logic; attribute dont_touch of G22803: signal is true;
	signal G22804: std_logic; attribute dont_touch of G22804: signal is true;
	signal G22805: std_logic; attribute dont_touch of G22805: signal is true;
	signal G22806: std_logic; attribute dont_touch of G22806: signal is true;
	signal G22809: std_logic; attribute dont_touch of G22809: signal is true;
	signal G22810: std_logic; attribute dont_touch of G22810: signal is true;
	signal G22811: std_logic; attribute dont_touch of G22811: signal is true;
	signal G22812: std_logic; attribute dont_touch of G22812: signal is true;
	signal G22824: std_logic; attribute dont_touch of G22824: signal is true;
	signal G22825: std_logic; attribute dont_touch of G22825: signal is true;
	signal G22826: std_logic; attribute dont_touch of G22826: signal is true;
	signal G22827: std_logic; attribute dont_touch of G22827: signal is true;
	signal G22828: std_logic; attribute dont_touch of G22828: signal is true;
	signal G22829: std_logic; attribute dont_touch of G22829: signal is true;
	signal G22830: std_logic; attribute dont_touch of G22830: signal is true;
	signal G22831: std_logic; attribute dont_touch of G22831: signal is true;
	signal G22832: std_logic; attribute dont_touch of G22832: signal is true;
	signal G22833: std_logic; attribute dont_touch of G22833: signal is true;
	signal G22834: std_logic; attribute dont_touch of G22834: signal is true;
	signal G22835: std_logic; attribute dont_touch of G22835: signal is true;
	signal G22836: std_logic; attribute dont_touch of G22836: signal is true;
	signal G22837: std_logic; attribute dont_touch of G22837: signal is true;
	signal G22838: std_logic; attribute dont_touch of G22838: signal is true;
	signal G22839: std_logic; attribute dont_touch of G22839: signal is true;
	signal G22840: std_logic; attribute dont_touch of G22840: signal is true;
	signal G22841: std_logic; attribute dont_touch of G22841: signal is true;
	signal G22842: std_logic; attribute dont_touch of G22842: signal is true;
	signal G22843: std_logic; attribute dont_touch of G22843: signal is true;
	signal G22844: std_logic; attribute dont_touch of G22844: signal is true;
	signal G22845: std_logic; attribute dont_touch of G22845: signal is true;
	signal G22846: std_logic; attribute dont_touch of G22846: signal is true;
	signal G22847: std_logic; attribute dont_touch of G22847: signal is true;
	signal G22850: std_logic; attribute dont_touch of G22850: signal is true;
	signal G22851: std_logic; attribute dont_touch of G22851: signal is true;
	signal G22852: std_logic; attribute dont_touch of G22852: signal is true;
	signal G22864: std_logic; attribute dont_touch of G22864: signal is true;
	signal G22865: std_logic; attribute dont_touch of G22865: signal is true;
	signal G22866: std_logic; attribute dont_touch of G22866: signal is true;
	signal G22867: std_logic; attribute dont_touch of G22867: signal is true;
	signal G22868: std_logic; attribute dont_touch of G22868: signal is true;
	signal G22869: std_logic; attribute dont_touch of G22869: signal is true;
	signal G22870: std_logic; attribute dont_touch of G22870: signal is true;
	signal G22871: std_logic; attribute dont_touch of G22871: signal is true;
	signal G22872: std_logic; attribute dont_touch of G22872: signal is true;
	signal G22873: std_logic; attribute dont_touch of G22873: signal is true;
	signal G22874: std_logic; attribute dont_touch of G22874: signal is true;
	signal G22875: std_logic; attribute dont_touch of G22875: signal is true;
	signal G22876: std_logic; attribute dont_touch of G22876: signal is true;
	signal G22879: std_logic; attribute dont_touch of G22879: signal is true;
	signal G22880: std_logic; attribute dont_touch of G22880: signal is true;
	signal G22881: std_logic; attribute dont_touch of G22881: signal is true;
	signal G22882: std_logic; attribute dont_touch of G22882: signal is true;
	signal G22885: std_logic; attribute dont_touch of G22885: signal is true;
	signal G22886: std_logic; attribute dont_touch of G22886: signal is true;
	signal G22887: std_logic; attribute dont_touch of G22887: signal is true;
	signal G22899: std_logic; attribute dont_touch of G22899: signal is true;
	signal G22900: std_logic; attribute dont_touch of G22900: signal is true;
	signal G22901: std_logic; attribute dont_touch of G22901: signal is true;
	signal G22902: std_logic; attribute dont_touch of G22902: signal is true;
	signal G22903: std_logic; attribute dont_touch of G22903: signal is true;
	signal G22906: std_logic; attribute dont_touch of G22906: signal is true;
	signal G22907: std_logic; attribute dont_touch of G22907: signal is true;
	signal G22911: std_logic; attribute dont_touch of G22911: signal is true;
	signal G22914: std_logic; attribute dont_touch of G22914: signal is true;
	signal G22915: std_logic; attribute dont_touch of G22915: signal is true;
	signal G22916: std_logic; attribute dont_touch of G22916: signal is true;
	signal G22917: std_logic; attribute dont_touch of G22917: signal is true;
	signal G22920: std_logic; attribute dont_touch of G22920: signal is true;
	signal G22921: std_logic; attribute dont_touch of G22921: signal is true;
	signal G22922: std_logic; attribute dont_touch of G22922: signal is true;
	signal G22934: std_logic; attribute dont_touch of G22934: signal is true;
	signal G22935: std_logic; attribute dont_touch of G22935: signal is true;
	signal G22936: std_logic; attribute dont_touch of G22936: signal is true;
	signal G22939: std_logic; attribute dont_touch of G22939: signal is true;
	signal G22940: std_logic; attribute dont_touch of G22940: signal is true;
	signal G22941: std_logic; attribute dont_touch of G22941: signal is true;
	signal G22942: std_logic; attribute dont_touch of G22942: signal is true;
	signal G22945: std_logic; attribute dont_touch of G22945: signal is true;
	signal G22948: std_logic; attribute dont_touch of G22948: signal is true;
	signal G22949: std_logic; attribute dont_touch of G22949: signal is true;
	signal G22953: std_logic; attribute dont_touch of G22953: signal is true;
	signal G22954: std_logic; attribute dont_touch of G22954: signal is true;
	signal G22958: std_logic; attribute dont_touch of G22958: signal is true;
	signal G22962: std_logic; attribute dont_touch of G22962: signal is true;
	signal G22966: std_logic; attribute dont_touch of G22966: signal is true;
	signal G22970: std_logic; attribute dont_touch of G22970: signal is true;
	signal G22971: std_logic; attribute dont_touch of G22971: signal is true;
	signal G22975: std_logic; attribute dont_touch of G22975: signal is true;
	signal G22979: std_logic; attribute dont_touch of G22979: signal is true;
	signal G22980: std_logic; attribute dont_touch of G22980: signal is true;
	signal G22984: std_logic; attribute dont_touch of G22984: signal is true;
	signal G22985: std_logic; attribute dont_touch of G22985: signal is true;
	signal G22986: std_logic; attribute dont_touch of G22986: signal is true;
	signal G22987: std_logic; attribute dont_touch of G22987: signal is true;
	signal G22988: std_logic; attribute dont_touch of G22988: signal is true;
	signal G22989: std_logic; attribute dont_touch of G22989: signal is true;
	signal G22990: std_logic; attribute dont_touch of G22990: signal is true;
	signal G22991: std_logic; attribute dont_touch of G22991: signal is true;
	signal G22992: std_logic; attribute dont_touch of G22992: signal is true;
	signal G22995: std_logic; attribute dont_touch of G22995: signal is true;
	signal G22996: std_logic; attribute dont_touch of G22996: signal is true;
	signal G22997: std_logic; attribute dont_touch of G22997: signal is true;
	signal G22998: std_logic; attribute dont_touch of G22998: signal is true;
	signal G22999: std_logic; attribute dont_touch of G22999: signal is true;
	signal G23000: std_logic; attribute dont_touch of G23000: signal is true;
	signal G23001: std_logic; attribute dont_touch of G23001: signal is true;
	signal G23002: std_logic; attribute dont_touch of G23002: signal is true;
	signal G23003: std_logic; attribute dont_touch of G23003: signal is true;
	signal G23006: std_logic; attribute dont_touch of G23006: signal is true;
	signal G23007: std_logic; attribute dont_touch of G23007: signal is true;
	signal G23008: std_logic; attribute dont_touch of G23008: signal is true;
	signal G23009: std_logic; attribute dont_touch of G23009: signal is true;
	signal G23012: std_logic; attribute dont_touch of G23012: signal is true;
	signal G23013: std_logic; attribute dont_touch of G23013: signal is true;
	signal G23014: std_logic; attribute dont_touch of G23014: signal is true;
	signal G23015: std_logic; attribute dont_touch of G23015: signal is true;
	signal G23016: std_logic; attribute dont_touch of G23016: signal is true;
	signal G23017: std_logic; attribute dont_touch of G23017: signal is true;
	signal G23020: std_logic; attribute dont_touch of G23020: signal is true;
	signal G23021: std_logic; attribute dont_touch of G23021: signal is true;
	signal G23022: std_logic; attribute dont_touch of G23022: signal is true;
	signal G23023: std_logic; attribute dont_touch of G23023: signal is true;
	signal G23024: std_logic; attribute dont_touch of G23024: signal is true;
	signal G23025: std_logic; attribute dont_touch of G23025: signal is true;
	signal G23028: std_logic; attribute dont_touch of G23028: signal is true;
	signal G23029: std_logic; attribute dont_touch of G23029: signal is true;
	signal G23030: std_logic; attribute dont_touch of G23030: signal is true;
	signal G23031: std_logic; attribute dont_touch of G23031: signal is true;
	signal G23032: std_logic; attribute dont_touch of G23032: signal is true;
	signal G23033: std_logic; attribute dont_touch of G23033: signal is true;
	signal G23036: std_logic; attribute dont_touch of G23036: signal is true;
	signal G23037: std_logic; attribute dont_touch of G23037: signal is true;
	signal G23038: std_logic; attribute dont_touch of G23038: signal is true;
	signal G23039: std_logic; attribute dont_touch of G23039: signal is true;
	signal G23040: std_logic; attribute dont_touch of G23040: signal is true;
	signal G23041: std_logic; attribute dont_touch of G23041: signal is true;
	signal G23042: std_logic; attribute dont_touch of G23042: signal is true;
	signal G23045: std_logic; attribute dont_touch of G23045: signal is true;
	signal G23046: std_logic; attribute dont_touch of G23046: signal is true;
	signal G23047: std_logic; attribute dont_touch of G23047: signal is true;
	signal G23048: std_logic; attribute dont_touch of G23048: signal is true;
	signal G23049: std_logic; attribute dont_touch of G23049: signal is true;
	signal G23050: std_logic; attribute dont_touch of G23050: signal is true;
	signal G23051: std_logic; attribute dont_touch of G23051: signal is true;
	signal G23052: std_logic; attribute dont_touch of G23052: signal is true;
	signal G23055: std_logic; attribute dont_touch of G23055: signal is true;
	signal G23056: std_logic; attribute dont_touch of G23056: signal is true;
	signal G23057: std_logic; attribute dont_touch of G23057: signal is true;
	signal G23058: std_logic; attribute dont_touch of G23058: signal is true;
	signal G23059: std_logic; attribute dont_touch of G23059: signal is true;
	signal G23060: std_logic; attribute dont_touch of G23060: signal is true;
	signal G23061: std_logic; attribute dont_touch of G23061: signal is true;
	signal G23064: std_logic; attribute dont_touch of G23064: signal is true;
	signal G23065: std_logic; attribute dont_touch of G23065: signal is true;
	signal G23066: std_logic; attribute dont_touch of G23066: signal is true;
	signal G23067: std_logic; attribute dont_touch of G23067: signal is true;
	signal G23068: std_logic; attribute dont_touch of G23068: signal is true;
	signal G23069: std_logic; attribute dont_touch of G23069: signal is true;
	signal G23070: std_logic; attribute dont_touch of G23070: signal is true;
	signal G23071: std_logic; attribute dont_touch of G23071: signal is true;
	signal G23074: std_logic; attribute dont_touch of G23074: signal is true;
	signal G23075: std_logic; attribute dont_touch of G23075: signal is true;
	signal G23076: std_logic; attribute dont_touch of G23076: signal is true;
	signal G23077: std_logic; attribute dont_touch of G23077: signal is true;
	signal G23078: std_logic; attribute dont_touch of G23078: signal is true;
	signal G23079: std_logic; attribute dont_touch of G23079: signal is true;
	signal G23080: std_logic; attribute dont_touch of G23080: signal is true;
	signal G23081: std_logic; attribute dont_touch of G23081: signal is true;
	signal G23082: std_logic; attribute dont_touch of G23082: signal is true;
	signal G23083: std_logic; attribute dont_touch of G23083: signal is true;
	signal G23084: std_logic; attribute dont_touch of G23084: signal is true;
	signal G23087: std_logic; attribute dont_touch of G23087: signal is true;
	signal G23088: std_logic; attribute dont_touch of G23088: signal is true;
	signal G23089: std_logic; attribute dont_touch of G23089: signal is true;
	signal G23092: std_logic; attribute dont_touch of G23092: signal is true;
	signal G23093: std_logic; attribute dont_touch of G23093: signal is true;
	signal G23094: std_logic; attribute dont_touch of G23094: signal is true;
	signal G23095: std_logic; attribute dont_touch of G23095: signal is true;
	signal G23096: std_logic; attribute dont_touch of G23096: signal is true;
	signal G23097: std_logic; attribute dont_touch of G23097: signal is true;
	signal G23098: std_logic; attribute dont_touch of G23098: signal is true;
	signal G23099: std_logic; attribute dont_touch of G23099: signal is true;
	signal G23100: std_logic; attribute dont_touch of G23100: signal is true;
	signal G23103: std_logic; attribute dont_touch of G23103: signal is true;
	signal G23104: std_logic; attribute dont_touch of G23104: signal is true;
	signal G23105: std_logic; attribute dont_touch of G23105: signal is true;
	signal G23106: std_logic; attribute dont_touch of G23106: signal is true;
	signal G23107: std_logic; attribute dont_touch of G23107: signal is true;
	signal G23110: std_logic; attribute dont_touch of G23110: signal is true;
	signal G23111: std_logic; attribute dont_touch of G23111: signal is true;
	signal G23112: std_logic; attribute dont_touch of G23112: signal is true;
	signal G23113: std_logic; attribute dont_touch of G23113: signal is true;
	signal G23114: std_logic; attribute dont_touch of G23114: signal is true;
	signal G23115: std_logic; attribute dont_touch of G23115: signal is true;
	signal G23116: std_logic; attribute dont_touch of G23116: signal is true;
	signal G23117: std_logic; attribute dont_touch of G23117: signal is true;
	signal G23118: std_logic; attribute dont_touch of G23118: signal is true;
	signal G23119: std_logic; attribute dont_touch of G23119: signal is true;
	signal G23120: std_logic; attribute dont_touch of G23120: signal is true;
	signal G23123: std_logic; attribute dont_touch of G23123: signal is true;
	signal G23124: std_logic; attribute dont_touch of G23124: signal is true;
	signal G23125: std_logic; attribute dont_touch of G23125: signal is true;
	signal G23126: std_logic; attribute dont_touch of G23126: signal is true;
	signal G23127: std_logic; attribute dont_touch of G23127: signal is true;
	signal G23128: std_logic; attribute dont_touch of G23128: signal is true;
	signal G23129: std_logic; attribute dont_touch of G23129: signal is true;
	signal G23132: std_logic; attribute dont_touch of G23132: signal is true;
	signal G23133: std_logic; attribute dont_touch of G23133: signal is true;
	signal G23134: std_logic; attribute dont_touch of G23134: signal is true;
	signal G23135: std_logic; attribute dont_touch of G23135: signal is true;
	signal G23136: std_logic; attribute dont_touch of G23136: signal is true;
	signal G23137: std_logic; attribute dont_touch of G23137: signal is true;
	signal G23138: std_logic; attribute dont_touch of G23138: signal is true;
	signal G23139: std_logic; attribute dont_touch of G23139: signal is true;
	signal G23140: std_logic; attribute dont_touch of G23140: signal is true;
	signal G23141: std_logic; attribute dont_touch of G23141: signal is true;
	signal G23142: std_logic; attribute dont_touch of G23142: signal is true;
	signal G23143: std_logic; attribute dont_touch of G23143: signal is true;
	signal G23144: std_logic; attribute dont_touch of G23144: signal is true;
	signal G23145: std_logic; attribute dont_touch of G23145: signal is true;
	signal G23146: std_logic; attribute dont_touch of G23146: signal is true;
	signal G23147: std_logic; attribute dont_touch of G23147: signal is true;
	signal G23148: std_logic; attribute dont_touch of G23148: signal is true;
	signal G23149: std_logic; attribute dont_touch of G23149: signal is true;
	signal G23150: std_logic; attribute dont_touch of G23150: signal is true;
	signal G23151: std_logic; attribute dont_touch of G23151: signal is true;
	signal G23152: std_logic; attribute dont_touch of G23152: signal is true;
	signal G23153: std_logic; attribute dont_touch of G23153: signal is true;
	signal G23154: std_logic; attribute dont_touch of G23154: signal is true;
	signal G23155: std_logic; attribute dont_touch of G23155: signal is true;
	signal G23156: std_logic; attribute dont_touch of G23156: signal is true;
	signal G23157: std_logic; attribute dont_touch of G23157: signal is true;
	signal G23158: std_logic; attribute dont_touch of G23158: signal is true;
	signal G23159: std_logic; attribute dont_touch of G23159: signal is true;
	signal G23160: std_logic; attribute dont_touch of G23160: signal is true;
	signal G23161: std_logic; attribute dont_touch of G23161: signal is true;
	signal G23162: std_logic; attribute dont_touch of G23162: signal is true;
	signal G23163: std_logic; attribute dont_touch of G23163: signal is true;
	signal G23164: std_logic; attribute dont_touch of G23164: signal is true;
	signal G23165: std_logic; attribute dont_touch of G23165: signal is true;
	signal G23166: std_logic; attribute dont_touch of G23166: signal is true;
	signal G23167: std_logic; attribute dont_touch of G23167: signal is true;
	signal G23168: std_logic; attribute dont_touch of G23168: signal is true;
	signal G23169: std_logic; attribute dont_touch of G23169: signal is true;
	signal G23170: std_logic; attribute dont_touch of G23170: signal is true;
	signal G23171: std_logic; attribute dont_touch of G23171: signal is true;
	signal G23172: std_logic; attribute dont_touch of G23172: signal is true;
	signal G23173: std_logic; attribute dont_touch of G23173: signal is true;
	signal G23174: std_logic; attribute dont_touch of G23174: signal is true;
	signal G23175: std_logic; attribute dont_touch of G23175: signal is true;
	signal G23176: std_logic; attribute dont_touch of G23176: signal is true;
	signal G23177: std_logic; attribute dont_touch of G23177: signal is true;
	signal G23178: std_logic; attribute dont_touch of G23178: signal is true;
	signal G23179: std_logic; attribute dont_touch of G23179: signal is true;
	signal G23180: std_logic; attribute dont_touch of G23180: signal is true;
	signal G23181: std_logic; attribute dont_touch of G23181: signal is true;
	signal G23182: std_logic; attribute dont_touch of G23182: signal is true;
	signal G23183: std_logic; attribute dont_touch of G23183: signal is true;
	signal G23184: std_logic; attribute dont_touch of G23184: signal is true;
	signal G23185: std_logic; attribute dont_touch of G23185: signal is true;
	signal G23186: std_logic; attribute dont_touch of G23186: signal is true;
	signal G23187: std_logic; attribute dont_touch of G23187: signal is true;
	signal G23188: std_logic; attribute dont_touch of G23188: signal is true;
	signal G23189: std_logic; attribute dont_touch of G23189: signal is true;
	signal G23190: std_logic; attribute dont_touch of G23190: signal is true;
	signal G23191: std_logic; attribute dont_touch of G23191: signal is true;
	signal G23192: std_logic; attribute dont_touch of G23192: signal is true;
	signal G23193: std_logic; attribute dont_touch of G23193: signal is true;
	signal G23194: std_logic; attribute dont_touch of G23194: signal is true;
	signal G23195: std_logic; attribute dont_touch of G23195: signal is true;
	signal G23196: std_logic; attribute dont_touch of G23196: signal is true;
	signal G23197: std_logic; attribute dont_touch of G23197: signal is true;
	signal G23198: std_logic; attribute dont_touch of G23198: signal is true;
	signal G23199: std_logic; attribute dont_touch of G23199: signal is true;
	signal G23200: std_logic; attribute dont_touch of G23200: signal is true;
	signal G23201: std_logic; attribute dont_touch of G23201: signal is true;
	signal G23202: std_logic; attribute dont_touch of G23202: signal is true;
	signal G23203: std_logic; attribute dont_touch of G23203: signal is true;
	signal G23204: std_logic; attribute dont_touch of G23204: signal is true;
	signal G23205: std_logic; attribute dont_touch of G23205: signal is true;
	signal G23206: std_logic; attribute dont_touch of G23206: signal is true;
	signal G23207: std_logic; attribute dont_touch of G23207: signal is true;
	signal G23208: std_logic; attribute dont_touch of G23208: signal is true;
	signal G23209: std_logic; attribute dont_touch of G23209: signal is true;
	signal G23210: std_logic; attribute dont_touch of G23210: signal is true;
	signal G23211: std_logic; attribute dont_touch of G23211: signal is true;
	signal G23212: std_logic; attribute dont_touch of G23212: signal is true;
	signal G23213: std_logic; attribute dont_touch of G23213: signal is true;
	signal G23214: std_logic; attribute dont_touch of G23214: signal is true;
	signal G23215: std_logic; attribute dont_touch of G23215: signal is true;
	signal G23216: std_logic; attribute dont_touch of G23216: signal is true;
	signal G23217: std_logic; attribute dont_touch of G23217: signal is true;
	signal G23218: std_logic; attribute dont_touch of G23218: signal is true;
	signal G23219: std_logic; attribute dont_touch of G23219: signal is true;
	signal G23220: std_logic; attribute dont_touch of G23220: signal is true;
	signal G23221: std_logic; attribute dont_touch of G23221: signal is true;
	signal G23222: std_logic; attribute dont_touch of G23222: signal is true;
	signal G23223: std_logic; attribute dont_touch of G23223: signal is true;
	signal G23224: std_logic; attribute dont_touch of G23224: signal is true;
	signal G23225: std_logic; attribute dont_touch of G23225: signal is true;
	signal G23226: std_logic; attribute dont_touch of G23226: signal is true;
	signal G23227: std_logic; attribute dont_touch of G23227: signal is true;
	signal G23228: std_logic; attribute dont_touch of G23228: signal is true;
	signal G23229: std_logic; attribute dont_touch of G23229: signal is true;
	signal G23230: std_logic; attribute dont_touch of G23230: signal is true;
	signal G23231: std_logic; attribute dont_touch of G23231: signal is true;
	signal G23232: std_logic; attribute dont_touch of G23232: signal is true;
	signal G23233: std_logic; attribute dont_touch of G23233: signal is true;
	signal G23234: std_logic; attribute dont_touch of G23234: signal is true;
	signal G23235: std_logic; attribute dont_touch of G23235: signal is true;
	signal G23236: std_logic; attribute dont_touch of G23236: signal is true;
	signal G23237: std_logic; attribute dont_touch of G23237: signal is true;
	signal G23238: std_logic; attribute dont_touch of G23238: signal is true;
	signal G23239: std_logic; attribute dont_touch of G23239: signal is true;
	signal G23240: std_logic; attribute dont_touch of G23240: signal is true;
	signal G23241: std_logic; attribute dont_touch of G23241: signal is true;
	signal G23242: std_logic; attribute dont_touch of G23242: signal is true;
	signal G23243: std_logic; attribute dont_touch of G23243: signal is true;
	signal G23244: std_logic; attribute dont_touch of G23244: signal is true;
	signal G23245: std_logic; attribute dont_touch of G23245: signal is true;
	signal G23246: std_logic; attribute dont_touch of G23246: signal is true;
	signal G23247: std_logic; attribute dont_touch of G23247: signal is true;
	signal G23248: std_logic; attribute dont_touch of G23248: signal is true;
	signal G23249: std_logic; attribute dont_touch of G23249: signal is true;
	signal G23250: std_logic; attribute dont_touch of G23250: signal is true;
	signal G23251: std_logic; attribute dont_touch of G23251: signal is true;
	signal G23252: std_logic; attribute dont_touch of G23252: signal is true;
	signal G23253: std_logic; attribute dont_touch of G23253: signal is true;
	signal G23254: std_logic; attribute dont_touch of G23254: signal is true;
	signal G23255: std_logic; attribute dont_touch of G23255: signal is true;
	signal G23256: std_logic; attribute dont_touch of G23256: signal is true;
	signal G23257: std_logic; attribute dont_touch of G23257: signal is true;
	signal G23258: std_logic; attribute dont_touch of G23258: signal is true;
	signal G23259: std_logic; attribute dont_touch of G23259: signal is true;
	signal G23260: std_logic; attribute dont_touch of G23260: signal is true;
	signal G23261: std_logic; attribute dont_touch of G23261: signal is true;
	signal G23262: std_logic; attribute dont_touch of G23262: signal is true;
	signal G23263: std_logic; attribute dont_touch of G23263: signal is true;
	signal G23264: std_logic; attribute dont_touch of G23264: signal is true;
	signal G23265: std_logic; attribute dont_touch of G23265: signal is true;
	signal G23266: std_logic; attribute dont_touch of G23266: signal is true;
	signal G23267: std_logic; attribute dont_touch of G23267: signal is true;
	signal G23268: std_logic; attribute dont_touch of G23268: signal is true;
	signal G23269: std_logic; attribute dont_touch of G23269: signal is true;
	signal G23270: std_logic; attribute dont_touch of G23270: signal is true;
	signal G23271: std_logic; attribute dont_touch of G23271: signal is true;
	signal G23272: std_logic; attribute dont_touch of G23272: signal is true;
	signal G23273: std_logic; attribute dont_touch of G23273: signal is true;
	signal G23274: std_logic; attribute dont_touch of G23274: signal is true;
	signal G23275: std_logic; attribute dont_touch of G23275: signal is true;
	signal G23276: std_logic; attribute dont_touch of G23276: signal is true;
	signal G23277: std_logic; attribute dont_touch of G23277: signal is true;
	signal G23278: std_logic; attribute dont_touch of G23278: signal is true;
	signal G23279: std_logic; attribute dont_touch of G23279: signal is true;
	signal G23280: std_logic; attribute dont_touch of G23280: signal is true;
	signal G23281: std_logic; attribute dont_touch of G23281: signal is true;
	signal G23282: std_logic; attribute dont_touch of G23282: signal is true;
	signal G23283: std_logic; attribute dont_touch of G23283: signal is true;
	signal G23284: std_logic; attribute dont_touch of G23284: signal is true;
	signal G23285: std_logic; attribute dont_touch of G23285: signal is true;
	signal G23286: std_logic; attribute dont_touch of G23286: signal is true;
	signal G23287: std_logic; attribute dont_touch of G23287: signal is true;
	signal G23288: std_logic; attribute dont_touch of G23288: signal is true;
	signal G23289: std_logic; attribute dont_touch of G23289: signal is true;
	signal G23290: std_logic; attribute dont_touch of G23290: signal is true;
	signal G23291: std_logic; attribute dont_touch of G23291: signal is true;
	signal G23292: std_logic; attribute dont_touch of G23292: signal is true;
	signal G23293: std_logic; attribute dont_touch of G23293: signal is true;
	signal G23294: std_logic; attribute dont_touch of G23294: signal is true;
	signal G23295: std_logic; attribute dont_touch of G23295: signal is true;
	signal G23296: std_logic; attribute dont_touch of G23296: signal is true;
	signal G23297: std_logic; attribute dont_touch of G23297: signal is true;
	signal G23298: std_logic; attribute dont_touch of G23298: signal is true;
	signal G23299: std_logic; attribute dont_touch of G23299: signal is true;
	signal G23300: std_logic; attribute dont_touch of G23300: signal is true;
	signal G23301: std_logic; attribute dont_touch of G23301: signal is true;
	signal G23302: std_logic; attribute dont_touch of G23302: signal is true;
	signal G23303: std_logic; attribute dont_touch of G23303: signal is true;
	signal G23304: std_logic; attribute dont_touch of G23304: signal is true;
	signal G23305: std_logic; attribute dont_touch of G23305: signal is true;
	signal G23306: std_logic; attribute dont_touch of G23306: signal is true;
	signal G23307: std_logic; attribute dont_touch of G23307: signal is true;
	signal G23308: std_logic; attribute dont_touch of G23308: signal is true;
	signal G23309: std_logic; attribute dont_touch of G23309: signal is true;
	signal G23310: std_logic; attribute dont_touch of G23310: signal is true;
	signal G23311: std_logic; attribute dont_touch of G23311: signal is true;
	signal G23312: std_logic; attribute dont_touch of G23312: signal is true;
	signal G23313: std_logic; attribute dont_touch of G23313: signal is true;
	signal G23314: std_logic; attribute dont_touch of G23314: signal is true;
	signal G23315: std_logic; attribute dont_touch of G23315: signal is true;
	signal G23316: std_logic; attribute dont_touch of G23316: signal is true;
	signal G23317: std_logic; attribute dont_touch of G23317: signal is true;
	signal G23318: std_logic; attribute dont_touch of G23318: signal is true;
	signal G23319: std_logic; attribute dont_touch of G23319: signal is true;
	signal G23320: std_logic; attribute dont_touch of G23320: signal is true;
	signal G23324: std_logic; attribute dont_touch of G23324: signal is true;
	signal G23325: std_logic; attribute dont_touch of G23325: signal is true;
	signal G23329: std_logic; attribute dont_touch of G23329: signal is true;
	signal G23330: std_logic; attribute dont_touch of G23330: signal is true;
	signal G23331: std_logic; attribute dont_touch of G23331: signal is true;
	signal G23335: std_logic; attribute dont_touch of G23335: signal is true;
	signal G23339: std_logic; attribute dont_touch of G23339: signal is true;
	signal G23340: std_logic; attribute dont_touch of G23340: signal is true;
	signal G23344: std_logic; attribute dont_touch of G23344: signal is true;
	signal G23348: std_logic; attribute dont_touch of G23348: signal is true;
	signal G23349: std_logic; attribute dont_touch of G23349: signal is true;
	signal G23353: std_logic; attribute dont_touch of G23353: signal is true;
	signal G23357: std_logic; attribute dont_touch of G23357: signal is true;
	signal G23358: std_logic; attribute dont_touch of G23358: signal is true;
	signal G23359: std_logic; attribute dont_touch of G23359: signal is true;
	signal G23360: std_logic; attribute dont_touch of G23360: signal is true;
	signal G23364: std_logic; attribute dont_touch of G23364: signal is true;
	signal G23368: std_logic; attribute dont_touch of G23368: signal is true;
	signal G23372: std_logic; attribute dont_touch of G23372: signal is true;
	signal G23376: std_logic; attribute dont_touch of G23376: signal is true;
	signal G23377: std_logic; attribute dont_touch of G23377: signal is true;
	signal G23381: std_logic; attribute dont_touch of G23381: signal is true;
	signal G23385: std_logic; attribute dont_touch of G23385: signal is true;
	signal G23386: std_logic; attribute dont_touch of G23386: signal is true;
	signal G23387: std_logic; attribute dont_touch of G23387: signal is true;
	signal G23388: std_logic; attribute dont_touch of G23388: signal is true;
	signal G23392: std_logic; attribute dont_touch of G23392: signal is true;
	signal G23393: std_logic; attribute dont_touch of G23393: signal is true;
	signal G23394: std_logic; attribute dont_touch of G23394: signal is true;
	signal G23395: std_logic; attribute dont_touch of G23395: signal is true;
	signal G23399: std_logic; attribute dont_touch of G23399: signal is true;
	signal G23400: std_logic; attribute dont_touch of G23400: signal is true;
	signal G23401: std_logic; attribute dont_touch of G23401: signal is true;
	signal G23402: std_logic; attribute dont_touch of G23402: signal is true;
	signal G23403: std_logic; attribute dont_touch of G23403: signal is true;
	signal G23406: std_logic; attribute dont_touch of G23406: signal is true;
	signal G23407: std_logic; attribute dont_touch of G23407: signal is true;
	signal G23408: std_logic; attribute dont_touch of G23408: signal is true;
	signal G23409: std_logic; attribute dont_touch of G23409: signal is true;
	signal G23410: std_logic; attribute dont_touch of G23410: signal is true;
	signal G23413: std_logic; attribute dont_touch of G23413: signal is true;
	signal G23414: std_logic; attribute dont_touch of G23414: signal is true;
	signal G23415: std_logic; attribute dont_touch of G23415: signal is true;
	signal G23418: std_logic; attribute dont_touch of G23418: signal is true;
	signal G23419: std_logic; attribute dont_touch of G23419: signal is true;
	signal G23420: std_logic; attribute dont_touch of G23420: signal is true;
	signal G23423: std_logic; attribute dont_touch of G23423: signal is true;
	signal G23424: std_logic; attribute dont_touch of G23424: signal is true;
	signal G23427: std_logic; attribute dont_touch of G23427: signal is true;
	signal G23428: std_logic; attribute dont_touch of G23428: signal is true;
	signal G23429: std_logic; attribute dont_touch of G23429: signal is true;
	signal G23432: std_logic; attribute dont_touch of G23432: signal is true;
	signal G23433: std_logic; attribute dont_touch of G23433: signal is true;
	signal G23434: std_logic; attribute dont_touch of G23434: signal is true;
	signal G23435: std_logic; attribute dont_touch of G23435: signal is true;
	signal G23438: std_logic; attribute dont_touch of G23438: signal is true;
	signal G23439: std_logic; attribute dont_touch of G23439: signal is true;
	signal G23440: std_logic; attribute dont_touch of G23440: signal is true;
	signal G23441: std_logic; attribute dont_touch of G23441: signal is true;
	signal G23444: std_logic; attribute dont_touch of G23444: signal is true;
	signal G23448: std_logic; attribute dont_touch of G23448: signal is true;
	signal G23451: std_logic; attribute dont_touch of G23451: signal is true;
	signal G23452: std_logic; attribute dont_touch of G23452: signal is true;
	signal G23453: std_logic; attribute dont_touch of G23453: signal is true;
	signal G23454: std_logic; attribute dont_touch of G23454: signal is true;
	signal G23455: std_logic; attribute dont_touch of G23455: signal is true;
	signal G23458: std_logic; attribute dont_touch of G23458: signal is true;
	signal G23459: std_logic; attribute dont_touch of G23459: signal is true;
	signal G23460: std_logic; attribute dont_touch of G23460: signal is true;
	signal G23461: std_logic; attribute dont_touch of G23461: signal is true;
	signal G23462: std_logic; attribute dont_touch of G23462: signal is true;
	signal G23463: std_logic; attribute dont_touch of G23463: signal is true;
	signal G23464: std_logic; attribute dont_touch of G23464: signal is true;
	signal G23467: std_logic; attribute dont_touch of G23467: signal is true;
	signal G23468: std_logic; attribute dont_touch of G23468: signal is true;
	signal G23469: std_logic; attribute dont_touch of G23469: signal is true;
	signal G23470: std_logic; attribute dont_touch of G23470: signal is true;
	signal G23471: std_logic; attribute dont_touch of G23471: signal is true;
	signal G23472: std_logic; attribute dont_touch of G23472: signal is true;
	signal G23473: std_logic; attribute dont_touch of G23473: signal is true;
	signal G23476: std_logic; attribute dont_touch of G23476: signal is true;
	signal G23477: std_logic; attribute dont_touch of G23477: signal is true;
	signal G23478: std_logic; attribute dont_touch of G23478: signal is true;
	signal G23481: std_logic; attribute dont_touch of G23481: signal is true;
	signal G23482: std_logic; attribute dont_touch of G23482: signal is true;
	signal G23483: std_logic; attribute dont_touch of G23483: signal is true;
	signal G23484: std_logic; attribute dont_touch of G23484: signal is true;
	signal G23485: std_logic; attribute dont_touch of G23485: signal is true;
	signal G23486: std_logic; attribute dont_touch of G23486: signal is true;
	signal G23489: std_logic; attribute dont_touch of G23489: signal is true;
	signal G23492: std_logic; attribute dont_touch of G23492: signal is true;
	signal G23493: std_logic; attribute dont_touch of G23493: signal is true;
	signal G23494: std_logic; attribute dont_touch of G23494: signal is true;
	signal G23495: std_logic; attribute dont_touch of G23495: signal is true;
	signal G23496: std_logic; attribute dont_touch of G23496: signal is true;
	signal G23497: std_logic; attribute dont_touch of G23497: signal is true;
	signal G23500: std_logic; attribute dont_touch of G23500: signal is true;
	signal G23501: std_logic; attribute dont_touch of G23501: signal is true;
	signal G23502: std_logic; attribute dont_touch of G23502: signal is true;
	signal G23505: std_logic; attribute dont_touch of G23505: signal is true;
	signal G23508: std_logic; attribute dont_touch of G23508: signal is true;
	signal G23509: std_logic; attribute dont_touch of G23509: signal is true;
	signal G23510: std_logic; attribute dont_touch of G23510: signal is true;
	signal G23511: std_logic; attribute dont_touch of G23511: signal is true;
	signal G23512: std_logic; attribute dont_touch of G23512: signal is true;
	signal G23513: std_logic; attribute dont_touch of G23513: signal is true;
	signal G23516: std_logic; attribute dont_touch of G23516: signal is true;
	signal G23517: std_logic; attribute dont_touch of G23517: signal is true;
	signal G23518: std_logic; attribute dont_touch of G23518: signal is true;
	signal G23521: std_logic; attribute dont_touch of G23521: signal is true;
	signal G23524: std_logic; attribute dont_touch of G23524: signal is true;
	signal G23525: std_logic; attribute dont_touch of G23525: signal is true;
	signal G23526: std_logic; attribute dont_touch of G23526: signal is true;
	signal G23527: std_logic; attribute dont_touch of G23527: signal is true;
	signal G23528: std_logic; attribute dont_touch of G23528: signal is true;
	signal G23531: std_logic; attribute dont_touch of G23531: signal is true;
	signal G23532: std_logic; attribute dont_touch of G23532: signal is true;
	signal G23533: std_logic; attribute dont_touch of G23533: signal is true;
	signal G23536: std_logic; attribute dont_touch of G23536: signal is true;
	signal G23537: std_logic; attribute dont_touch of G23537: signal is true;
	signal G23538: std_logic; attribute dont_touch of G23538: signal is true;
	signal G23539: std_logic; attribute dont_touch of G23539: signal is true;
	signal G23542: std_logic; attribute dont_touch of G23542: signal is true;
	signal G23543: std_logic; attribute dont_touch of G23543: signal is true;
	signal G23544: std_logic; attribute dont_touch of G23544: signal is true;
	signal G23545: std_logic; attribute dont_touch of G23545: signal is true;
	signal G23546: std_logic; attribute dont_touch of G23546: signal is true;
	signal G23547: std_logic; attribute dont_touch of G23547: signal is true;
	signal G23548: std_logic; attribute dont_touch of G23548: signal is true;
	signal G23549: std_logic; attribute dont_touch of G23549: signal is true;
	signal G23550: std_logic; attribute dont_touch of G23550: signal is true;
	signal G23551: std_logic; attribute dont_touch of G23551: signal is true;
	signal G23552: std_logic; attribute dont_touch of G23552: signal is true;
	signal G23553: std_logic; attribute dont_touch of G23553: signal is true;
	signal G23554: std_logic; attribute dont_touch of G23554: signal is true;
	signal G23555: std_logic; attribute dont_touch of G23555: signal is true;
	signal G23556: std_logic; attribute dont_touch of G23556: signal is true;
	signal G23557: std_logic; attribute dont_touch of G23557: signal is true;
	signal G23558: std_logic; attribute dont_touch of G23558: signal is true;
	signal G23559: std_logic; attribute dont_touch of G23559: signal is true;
	signal G23560: std_logic; attribute dont_touch of G23560: signal is true;
	signal G23561: std_logic; attribute dont_touch of G23561: signal is true;
	signal G23562: std_logic; attribute dont_touch of G23562: signal is true;
	signal G23563: std_logic; attribute dont_touch of G23563: signal is true;
	signal G23564: std_logic; attribute dont_touch of G23564: signal is true;
	signal G23565: std_logic; attribute dont_touch of G23565: signal is true;
	signal G23566: std_logic; attribute dont_touch of G23566: signal is true;
	signal G23567: std_logic; attribute dont_touch of G23567: signal is true;
	signal G23568: std_logic; attribute dont_touch of G23568: signal is true;
	signal G23569: std_logic; attribute dont_touch of G23569: signal is true;
	signal G23570: std_logic; attribute dont_touch of G23570: signal is true;
	signal G23571: std_logic; attribute dont_touch of G23571: signal is true;
	signal G23572: std_logic; attribute dont_touch of G23572: signal is true;
	signal G23573: std_logic; attribute dont_touch of G23573: signal is true;
	signal G23574: std_logic; attribute dont_touch of G23574: signal is true;
	signal G23575: std_logic; attribute dont_touch of G23575: signal is true;
	signal G23576: std_logic; attribute dont_touch of G23576: signal is true;
	signal G23577: std_logic; attribute dont_touch of G23577: signal is true;
	signal G23578: std_logic; attribute dont_touch of G23578: signal is true;
	signal G23579: std_logic; attribute dont_touch of G23579: signal is true;
	signal G23580: std_logic; attribute dont_touch of G23580: signal is true;
	signal G23581: std_logic; attribute dont_touch of G23581: signal is true;
	signal G23582: std_logic; attribute dont_touch of G23582: signal is true;
	signal G23583: std_logic; attribute dont_touch of G23583: signal is true;
	signal G23584: std_logic; attribute dont_touch of G23584: signal is true;
	signal G23585: std_logic; attribute dont_touch of G23585: signal is true;
	signal G23586: std_logic; attribute dont_touch of G23586: signal is true;
	signal G23587: std_logic; attribute dont_touch of G23587: signal is true;
	signal G23588: std_logic; attribute dont_touch of G23588: signal is true;
	signal G23589: std_logic; attribute dont_touch of G23589: signal is true;
	signal G23590: std_logic; attribute dont_touch of G23590: signal is true;
	signal G23591: std_logic; attribute dont_touch of G23591: signal is true;
	signal G23592: std_logic; attribute dont_touch of G23592: signal is true;
	signal G23593: std_logic; attribute dont_touch of G23593: signal is true;
	signal G23594: std_logic; attribute dont_touch of G23594: signal is true;
	signal G23595: std_logic; attribute dont_touch of G23595: signal is true;
	signal G23596: std_logic; attribute dont_touch of G23596: signal is true;
	signal G23597: std_logic; attribute dont_touch of G23597: signal is true;
	signal G23598: std_logic; attribute dont_touch of G23598: signal is true;
	signal G23599: std_logic; attribute dont_touch of G23599: signal is true;
	signal G23600: std_logic; attribute dont_touch of G23600: signal is true;
	signal G23601: std_logic; attribute dont_touch of G23601: signal is true;
	signal G23602: std_logic; attribute dont_touch of G23602: signal is true;
	signal G23603: std_logic; attribute dont_touch of G23603: signal is true;
	signal G23604: std_logic; attribute dont_touch of G23604: signal is true;
	signal G23605: std_logic; attribute dont_touch of G23605: signal is true;
	signal G23606: std_logic; attribute dont_touch of G23606: signal is true;
	signal G23607: std_logic; attribute dont_touch of G23607: signal is true;
	signal G23608: std_logic; attribute dont_touch of G23608: signal is true;
	signal G23609: std_logic; attribute dont_touch of G23609: signal is true;
	signal G23610: std_logic; attribute dont_touch of G23610: signal is true;
	signal G23611: std_logic; attribute dont_touch of G23611: signal is true;
	signal G23612: std_logic; attribute dont_touch of G23612: signal is true;
	signal G23613: std_logic; attribute dont_touch of G23613: signal is true;
	signal G23614: std_logic; attribute dont_touch of G23614: signal is true;
	signal G23615: std_logic; attribute dont_touch of G23615: signal is true;
	signal G23616: std_logic; attribute dont_touch of G23616: signal is true;
	signal G23617: std_logic; attribute dont_touch of G23617: signal is true;
	signal G23618: std_logic; attribute dont_touch of G23618: signal is true;
	signal G23619: std_logic; attribute dont_touch of G23619: signal is true;
	signal G23620: std_logic; attribute dont_touch of G23620: signal is true;
	signal G23621: std_logic; attribute dont_touch of G23621: signal is true;
	signal G23622: std_logic; attribute dont_touch of G23622: signal is true;
	signal G23623: std_logic; attribute dont_touch of G23623: signal is true;
	signal G23624: std_logic; attribute dont_touch of G23624: signal is true;
	signal G23625: std_logic; attribute dont_touch of G23625: signal is true;
	signal G23626: std_logic; attribute dont_touch of G23626: signal is true;
	signal G23627: std_logic; attribute dont_touch of G23627: signal is true;
	signal G23628: std_logic; attribute dont_touch of G23628: signal is true;
	signal G23629: std_logic; attribute dont_touch of G23629: signal is true;
	signal G23630: std_logic; attribute dont_touch of G23630: signal is true;
	signal G23631: std_logic; attribute dont_touch of G23631: signal is true;
	signal G23632: std_logic; attribute dont_touch of G23632: signal is true;
	signal G23633: std_logic; attribute dont_touch of G23633: signal is true;
	signal G23634: std_logic; attribute dont_touch of G23634: signal is true;
	signal G23635: std_logic; attribute dont_touch of G23635: signal is true;
	signal G23636: std_logic; attribute dont_touch of G23636: signal is true;
	signal G23637: std_logic; attribute dont_touch of G23637: signal is true;
	signal G23638: std_logic; attribute dont_touch of G23638: signal is true;
	signal G23639: std_logic; attribute dont_touch of G23639: signal is true;
	signal G23640: std_logic; attribute dont_touch of G23640: signal is true;
	signal G23641: std_logic; attribute dont_touch of G23641: signal is true;
	signal G23642: std_logic; attribute dont_touch of G23642: signal is true;
	signal G23643: std_logic; attribute dont_touch of G23643: signal is true;
	signal G23644: std_logic; attribute dont_touch of G23644: signal is true;
	signal G23659: std_logic; attribute dont_touch of G23659: signal is true;
	signal G23660: std_logic; attribute dont_touch of G23660: signal is true;
	signal G23661: std_logic; attribute dont_touch of G23661: signal is true;
	signal G23662: std_logic; attribute dont_touch of G23662: signal is true;
	signal G23663: std_logic; attribute dont_touch of G23663: signal is true;
	signal G23664: std_logic; attribute dont_touch of G23664: signal is true;
	signal G23665: std_logic; attribute dont_touch of G23665: signal is true;
	signal G23666: std_logic; attribute dont_touch of G23666: signal is true;
	signal G23667: std_logic; attribute dont_touch of G23667: signal is true;
	signal G23668: std_logic; attribute dont_touch of G23668: signal is true;
	signal G23669: std_logic; attribute dont_touch of G23669: signal is true;
	signal G23670: std_logic; attribute dont_touch of G23670: signal is true;
	signal G23671: std_logic; attribute dont_touch of G23671: signal is true;
	signal G23672: std_logic; attribute dont_touch of G23672: signal is true;
	signal G23673: std_logic; attribute dont_touch of G23673: signal is true;
	signal G23674: std_logic; attribute dont_touch of G23674: signal is true;
	signal G23675: std_logic; attribute dont_touch of G23675: signal is true;
	signal G23676: std_logic; attribute dont_touch of G23676: signal is true;
	signal G23677: std_logic; attribute dont_touch of G23677: signal is true;
	signal G23678: std_logic; attribute dont_touch of G23678: signal is true;
	signal G23679: std_logic; attribute dont_touch of G23679: signal is true;
	signal G23680: std_logic; attribute dont_touch of G23680: signal is true;
	signal G23681: std_logic; attribute dont_touch of G23681: signal is true;
	signal G23682: std_logic; attribute dont_touch of G23682: signal is true;
	signal G23683: std_logic; attribute dont_touch of G23683: signal is true;
	signal G23684: std_logic; attribute dont_touch of G23684: signal is true;
	signal G23685: std_logic; attribute dont_touch of G23685: signal is true;
	signal G23686: std_logic; attribute dont_touch of G23686: signal is true;
	signal G23687: std_logic; attribute dont_touch of G23687: signal is true;
	signal G23688: std_logic; attribute dont_touch of G23688: signal is true;
	signal G23689: std_logic; attribute dont_touch of G23689: signal is true;
	signal G23690: std_logic; attribute dont_touch of G23690: signal is true;
	signal G23691: std_logic; attribute dont_touch of G23691: signal is true;
	signal G23692: std_logic; attribute dont_touch of G23692: signal is true;
	signal G23693: std_logic; attribute dont_touch of G23693: signal is true;
	signal G23694: std_logic; attribute dont_touch of G23694: signal is true;
	signal G23709: std_logic; attribute dont_touch of G23709: signal is true;
	signal G23710: std_logic; attribute dont_touch of G23710: signal is true;
	signal G23711: std_logic; attribute dont_touch of G23711: signal is true;
	signal G23712: std_logic; attribute dont_touch of G23712: signal is true;
	signal G23713: std_logic; attribute dont_touch of G23713: signal is true;
	signal G23714: std_logic; attribute dont_touch of G23714: signal is true;
	signal G23715: std_logic; attribute dont_touch of G23715: signal is true;
	signal G23716: std_logic; attribute dont_touch of G23716: signal is true;
	signal G23717: std_logic; attribute dont_touch of G23717: signal is true;
	signal G23718: std_logic; attribute dont_touch of G23718: signal is true;
	signal G23719: std_logic; attribute dont_touch of G23719: signal is true;
	signal G23720: std_logic; attribute dont_touch of G23720: signal is true;
	signal G23721: std_logic; attribute dont_touch of G23721: signal is true;
	signal G23722: std_logic; attribute dont_touch of G23722: signal is true;
	signal G23723: std_logic; attribute dont_touch of G23723: signal is true;
	signal G23724: std_logic; attribute dont_touch of G23724: signal is true;
	signal G23725: std_logic; attribute dont_touch of G23725: signal is true;
	signal G23726: std_logic; attribute dont_touch of G23726: signal is true;
	signal G23727: std_logic; attribute dont_touch of G23727: signal is true;
	signal G23728: std_logic; attribute dont_touch of G23728: signal is true;
	signal G23729: std_logic; attribute dont_touch of G23729: signal is true;
	signal G23730: std_logic; attribute dont_touch of G23730: signal is true;
	signal G23731: std_logic; attribute dont_touch of G23731: signal is true;
	signal G23734: std_logic; attribute dont_touch of G23734: signal is true;
	signal G23735: std_logic; attribute dont_touch of G23735: signal is true;
	signal G23736: std_logic; attribute dont_touch of G23736: signal is true;
	signal G23737: std_logic; attribute dont_touch of G23737: signal is true;
	signal G23738: std_logic; attribute dont_touch of G23738: signal is true;
	signal G23739: std_logic; attribute dont_touch of G23739: signal is true;
	signal G23740: std_logic; attribute dont_touch of G23740: signal is true;
	signal G23741: std_logic; attribute dont_touch of G23741: signal is true;
	signal G23742: std_logic; attribute dont_touch of G23742: signal is true;
	signal G23743: std_logic; attribute dont_touch of G23743: signal is true;
	signal G23744: std_logic; attribute dont_touch of G23744: signal is true;
	signal G23745: std_logic; attribute dont_touch of G23745: signal is true;
	signal G23746: std_logic; attribute dont_touch of G23746: signal is true;
	signal G23747: std_logic; attribute dont_touch of G23747: signal is true;
	signal G23748: std_logic; attribute dont_touch of G23748: signal is true;
	signal G23763: std_logic; attribute dont_touch of G23763: signal is true;
	signal G23764: std_logic; attribute dont_touch of G23764: signal is true;
	signal G23765: std_logic; attribute dont_touch of G23765: signal is true;
	signal G23766: std_logic; attribute dont_touch of G23766: signal is true;
	signal G23767: std_logic; attribute dont_touch of G23767: signal is true;
	signal G23768: std_logic; attribute dont_touch of G23768: signal is true;
	signal G23769: std_logic; attribute dont_touch of G23769: signal is true;
	signal G23770: std_logic; attribute dont_touch of G23770: signal is true;
	signal G23771: std_logic; attribute dont_touch of G23771: signal is true;
	signal G23772: std_logic; attribute dont_touch of G23772: signal is true;
	signal G23773: std_logic; attribute dont_touch of G23773: signal is true;
	signal G23774: std_logic; attribute dont_touch of G23774: signal is true;
	signal G23775: std_logic; attribute dont_touch of G23775: signal is true;
	signal G23776: std_logic; attribute dont_touch of G23776: signal is true;
	signal G23777: std_logic; attribute dont_touch of G23777: signal is true;
	signal G23778: std_logic; attribute dont_touch of G23778: signal is true;
	signal G23779: std_logic; attribute dont_touch of G23779: signal is true;
	signal G23782: std_logic; attribute dont_touch of G23782: signal is true;
	signal G23783: std_logic; attribute dont_touch of G23783: signal is true;
	signal G23784: std_logic; attribute dont_touch of G23784: signal is true;
	signal G23785: std_logic; attribute dont_touch of G23785: signal is true;
	signal G23786: std_logic; attribute dont_touch of G23786: signal is true;
	signal G23789: std_logic; attribute dont_touch of G23789: signal is true;
	signal G23790: std_logic; attribute dont_touch of G23790: signal is true;
	signal G23791: std_logic; attribute dont_touch of G23791: signal is true;
	signal G23792: std_logic; attribute dont_touch of G23792: signal is true;
	signal G23793: std_logic; attribute dont_touch of G23793: signal is true;
	signal G23794: std_logic; attribute dont_touch of G23794: signal is true;
	signal G23795: std_logic; attribute dont_touch of G23795: signal is true;
	signal G23796: std_logic; attribute dont_touch of G23796: signal is true;
	signal G23797: std_logic; attribute dont_touch of G23797: signal is true;
	signal G23798: std_logic; attribute dont_touch of G23798: signal is true;
	signal G23799: std_logic; attribute dont_touch of G23799: signal is true;
	signal G23800: std_logic; attribute dont_touch of G23800: signal is true;
	signal G23801: std_logic; attribute dont_touch of G23801: signal is true;
	signal G23802: std_logic; attribute dont_touch of G23802: signal is true;
	signal G23803: std_logic; attribute dont_touch of G23803: signal is true;
	signal G23818: std_logic; attribute dont_touch of G23818: signal is true;
	signal G23819: std_logic; attribute dont_touch of G23819: signal is true;
	signal G23820: std_logic; attribute dont_touch of G23820: signal is true;
	signal G23821: std_logic; attribute dont_touch of G23821: signal is true;
	signal G23822: std_logic; attribute dont_touch of G23822: signal is true;
	signal G23823: std_logic; attribute dont_touch of G23823: signal is true;
	signal G23824: std_logic; attribute dont_touch of G23824: signal is true;
	signal G23825: std_logic; attribute dont_touch of G23825: signal is true;
	signal G23826: std_logic; attribute dont_touch of G23826: signal is true;
	signal G23827: std_logic; attribute dont_touch of G23827: signal is true;
	signal G23828: std_logic; attribute dont_touch of G23828: signal is true;
	signal G23829: std_logic; attribute dont_touch of G23829: signal is true;
	signal G23830: std_logic; attribute dont_touch of G23830: signal is true;
	signal G23831: std_logic; attribute dont_touch of G23831: signal is true;
	signal G23832: std_logic; attribute dont_touch of G23832: signal is true;
	signal G23835: std_logic; attribute dont_touch of G23835: signal is true;
	signal G23836: std_logic; attribute dont_touch of G23836: signal is true;
	signal G23837: std_logic; attribute dont_touch of G23837: signal is true;
	signal G23838: std_logic; attribute dont_touch of G23838: signal is true;
	signal G23839: std_logic; attribute dont_touch of G23839: signal is true;
	signal G23842: std_logic; attribute dont_touch of G23842: signal is true;
	signal G23843: std_logic; attribute dont_touch of G23843: signal is true;
	signal G23844: std_logic; attribute dont_touch of G23844: signal is true;
	signal G23845: std_logic; attribute dont_touch of G23845: signal is true;
	signal G23846: std_logic; attribute dont_touch of G23846: signal is true;
	signal G23847: std_logic; attribute dont_touch of G23847: signal is true;
	signal G23848: std_logic; attribute dont_touch of G23848: signal is true;
	signal G23849: std_logic; attribute dont_touch of G23849: signal is true;
	signal G23850: std_logic; attribute dont_touch of G23850: signal is true;
	signal G23851: std_logic; attribute dont_touch of G23851: signal is true;
	signal G23852: std_logic; attribute dont_touch of G23852: signal is true;
	signal G23853: std_logic; attribute dont_touch of G23853: signal is true;
	signal G23854: std_logic; attribute dont_touch of G23854: signal is true;
	signal G23855: std_logic; attribute dont_touch of G23855: signal is true;
	signal G23856: std_logic; attribute dont_touch of G23856: signal is true;
	signal G23857: std_logic; attribute dont_touch of G23857: signal is true;
	signal G23858: std_logic; attribute dont_touch of G23858: signal is true;
	signal G23859: std_logic; attribute dont_touch of G23859: signal is true;
	signal G23860: std_logic; attribute dont_touch of G23860: signal is true;
	signal G23861: std_logic; attribute dont_touch of G23861: signal is true;
	signal G23862: std_logic; attribute dont_touch of G23862: signal is true;
	signal G23863: std_logic; attribute dont_touch of G23863: signal is true;
	signal G23864: std_logic; attribute dont_touch of G23864: signal is true;
	signal G23865: std_logic; attribute dont_touch of G23865: signal is true;
	signal G23866: std_logic; attribute dont_touch of G23866: signal is true;
	signal G23867: std_logic; attribute dont_touch of G23867: signal is true;
	signal G23870: std_logic; attribute dont_touch of G23870: signal is true;
	signal G23871: std_logic; attribute dont_touch of G23871: signal is true;
	signal G23872: std_logic; attribute dont_touch of G23872: signal is true;
	signal G23873: std_logic; attribute dont_touch of G23873: signal is true;
	signal G23874: std_logic; attribute dont_touch of G23874: signal is true;
	signal G23877: std_logic; attribute dont_touch of G23877: signal is true;
	signal G23878: std_logic; attribute dont_touch of G23878: signal is true;
	signal G23879: std_logic; attribute dont_touch of G23879: signal is true;
	signal G23882: std_logic; attribute dont_touch of G23882: signal is true;
	signal G23885: std_logic; attribute dont_touch of G23885: signal is true;
	signal G23886: std_logic; attribute dont_touch of G23886: signal is true;
	signal G23887: std_logic; attribute dont_touch of G23887: signal is true;
	signal G23888: std_logic; attribute dont_touch of G23888: signal is true;
	signal G23889: std_logic; attribute dont_touch of G23889: signal is true;
	signal G23890: std_logic; attribute dont_touch of G23890: signal is true;
	signal G23891: std_logic; attribute dont_touch of G23891: signal is true;
	signal G23892: std_logic; attribute dont_touch of G23892: signal is true;
	signal G23893: std_logic; attribute dont_touch of G23893: signal is true;
	signal G23894: std_logic; attribute dont_touch of G23894: signal is true;
	signal G23895: std_logic; attribute dont_touch of G23895: signal is true;
	signal G23896: std_logic; attribute dont_touch of G23896: signal is true;
	signal G23897: std_logic; attribute dont_touch of G23897: signal is true;
	signal G23898: std_logic; attribute dont_touch of G23898: signal is true;
	signal G23899: std_logic; attribute dont_touch of G23899: signal is true;
	signal G23900: std_logic; attribute dont_touch of G23900: signal is true;
	signal G23901: std_logic; attribute dont_touch of G23901: signal is true;
	signal G23904: std_logic; attribute dont_touch of G23904: signal is true;
	signal G23905: std_logic; attribute dont_touch of G23905: signal is true;
	signal G23906: std_logic; attribute dont_touch of G23906: signal is true;
	signal G23907: std_logic; attribute dont_touch of G23907: signal is true;
	signal G23908: std_logic; attribute dont_touch of G23908: signal is true;
	signal G23909: std_logic; attribute dont_touch of G23909: signal is true;
	signal G23910: std_logic; attribute dont_touch of G23910: signal is true;
	signal G23911: std_logic; attribute dont_touch of G23911: signal is true;
	signal G23912: std_logic; attribute dont_touch of G23912: signal is true;
	signal G23913: std_logic; attribute dont_touch of G23913: signal is true;
	signal G23914: std_logic; attribute dont_touch of G23914: signal is true;
	signal G23915: std_logic; attribute dont_touch of G23915: signal is true;
	signal G23916: std_logic; attribute dont_touch of G23916: signal is true;
	signal G23917: std_logic; attribute dont_touch of G23917: signal is true;
	signal G23918: std_logic; attribute dont_touch of G23918: signal is true;
	signal G23919: std_logic; attribute dont_touch of G23919: signal is true;
	signal G23922: std_logic; attribute dont_touch of G23922: signal is true;
	signal G23923: std_logic; attribute dont_touch of G23923: signal is true;
	signal G23936: std_logic; attribute dont_touch of G23936: signal is true;
	signal G23937: std_logic; attribute dont_touch of G23937: signal is true;
	signal G23938: std_logic; attribute dont_touch of G23938: signal is true;
	signal G23939: std_logic; attribute dont_touch of G23939: signal is true;
	signal G23940: std_logic; attribute dont_touch of G23940: signal is true;
	signal G23941: std_logic; attribute dont_touch of G23941: signal is true;
	signal G23942: std_logic; attribute dont_touch of G23942: signal is true;
	signal G23943: std_logic; attribute dont_touch of G23943: signal is true;
	signal G23944: std_logic; attribute dont_touch of G23944: signal is true;
	signal G23945: std_logic; attribute dont_touch of G23945: signal is true;
	signal G23950: std_logic; attribute dont_touch of G23950: signal is true;
	signal G23953: std_logic; attribute dont_touch of G23953: signal is true;
	signal G23954: std_logic; attribute dont_touch of G23954: signal is true;
	signal G23955: std_logic; attribute dont_touch of G23955: signal is true;
	signal G23968: std_logic; attribute dont_touch of G23968: signal is true;
	signal G23969: std_logic; attribute dont_touch of G23969: signal is true;
	signal G23970: std_logic; attribute dont_touch of G23970: signal is true;
	signal G23971: std_logic; attribute dont_touch of G23971: signal is true;
	signal G23972: std_logic; attribute dont_touch of G23972: signal is true;
	signal G23973: std_logic; attribute dont_touch of G23973: signal is true;
	signal G23974: std_logic; attribute dont_touch of G23974: signal is true;
	signal G23979: std_logic; attribute dont_touch of G23979: signal is true;
	signal G23982: std_logic; attribute dont_touch of G23982: signal is true;
	signal G23983: std_logic; attribute dont_touch of G23983: signal is true;
	signal G23984: std_logic; attribute dont_touch of G23984: signal is true;
	signal G23997: std_logic; attribute dont_touch of G23997: signal is true;
	signal G23998: std_logic; attribute dont_touch of G23998: signal is true;
	signal G23999: std_logic; attribute dont_touch of G23999: signal is true;
	signal G24000: std_logic; attribute dont_touch of G24000: signal is true;
	signal G24001: std_logic; attribute dont_touch of G24001: signal is true;
	signal G24002: std_logic; attribute dont_touch of G24002: signal is true;
	signal G24003: std_logic; attribute dont_touch of G24003: signal is true;
	signal G24004: std_logic; attribute dont_touch of G24004: signal is true;
	signal G24009: std_logic; attribute dont_touch of G24009: signal is true;
	signal G24012: std_logic; attribute dont_touch of G24012: signal is true;
	signal G24013: std_logic; attribute dont_touch of G24013: signal is true;
	signal G24014: std_logic; attribute dont_touch of G24014: signal is true;
	signal G24027: std_logic; attribute dont_touch of G24027: signal is true;
	signal G24028: std_logic; attribute dont_touch of G24028: signal is true;
	signal G24029: std_logic; attribute dont_touch of G24029: signal is true;
	signal G24030: std_logic; attribute dont_touch of G24030: signal is true;
	signal G24033: std_logic; attribute dont_touch of G24033: signal is true;
	signal G24034: std_logic; attribute dont_touch of G24034: signal is true;
	signal G24035: std_logic; attribute dont_touch of G24035: signal is true;
	signal G24036: std_logic; attribute dont_touch of G24036: signal is true;
	signal G24037: std_logic; attribute dont_touch of G24037: signal is true;
	signal G24038: std_logic; attribute dont_touch of G24038: signal is true;
	signal G24043: std_logic; attribute dont_touch of G24043: signal is true;
	signal G24046: std_logic; attribute dont_touch of G24046: signal is true;
	signal G24047: std_logic; attribute dont_touch of G24047: signal is true;
	signal G24051: std_logic; attribute dont_touch of G24051: signal is true;
	signal G24052: std_logic; attribute dont_touch of G24052: signal is true;
	signal G24053: std_logic; attribute dont_touch of G24053: signal is true;
	signal G24054: std_logic; attribute dont_touch of G24054: signal is true;
	signal G24055: std_logic; attribute dont_touch of G24055: signal is true;
	signal G24056: std_logic; attribute dont_touch of G24056: signal is true;
	signal G24057: std_logic; attribute dont_touch of G24057: signal is true;
	signal G24058: std_logic; attribute dont_touch of G24058: signal is true;
	signal G24059: std_logic; attribute dont_touch of G24059: signal is true;
	signal G24060: std_logic; attribute dont_touch of G24060: signal is true;
	signal G24064: std_logic; attribute dont_touch of G24064: signal is true;
	signal G24065: std_logic; attribute dont_touch of G24065: signal is true;
	signal G24066: std_logic; attribute dont_touch of G24066: signal is true;
	signal G24067: std_logic; attribute dont_touch of G24067: signal is true;
	signal G24068: std_logic; attribute dont_touch of G24068: signal is true;
	signal G24069: std_logic; attribute dont_touch of G24069: signal is true;
	signal G24070: std_logic; attribute dont_touch of G24070: signal is true;
	signal G24071: std_logic; attribute dont_touch of G24071: signal is true;
	signal G24072: std_logic; attribute dont_touch of G24072: signal is true;
	signal G24073: std_logic; attribute dont_touch of G24073: signal is true;
	signal G24077: std_logic; attribute dont_touch of G24077: signal is true;
	signal G24078: std_logic; attribute dont_touch of G24078: signal is true;
	signal G24079: std_logic; attribute dont_touch of G24079: signal is true;
	signal G24080: std_logic; attribute dont_touch of G24080: signal is true;
	signal G24081: std_logic; attribute dont_touch of G24081: signal is true;
	signal G24082: std_logic; attribute dont_touch of G24082: signal is true;
	signal G24083: std_logic; attribute dont_touch of G24083: signal is true;
	signal G24084: std_logic; attribute dont_touch of G24084: signal is true;
	signal G24088: std_logic; attribute dont_touch of G24088: signal is true;
	signal G24089: std_logic; attribute dont_touch of G24089: signal is true;
	signal G24090: std_logic; attribute dont_touch of G24090: signal is true;
	signal G24091: std_logic; attribute dont_touch of G24091: signal is true;
	signal G24092: std_logic; attribute dont_touch of G24092: signal is true;
	signal G24093: std_logic; attribute dont_touch of G24093: signal is true;
	signal G24094: std_logic; attribute dont_touch of G24094: signal is true;
	signal G24095: std_logic; attribute dont_touch of G24095: signal is true;
	signal G24096: std_logic; attribute dont_touch of G24096: signal is true;
	signal G24097: std_logic; attribute dont_touch of G24097: signal is true;
	signal G24098: std_logic; attribute dont_touch of G24098: signal is true;
	signal G24099: std_logic; attribute dont_touch of G24099: signal is true;
	signal G24100: std_logic; attribute dont_touch of G24100: signal is true;
	signal G24101: std_logic; attribute dont_touch of G24101: signal is true;
	signal G24102: std_logic; attribute dont_touch of G24102: signal is true;
	signal G24103: std_logic; attribute dont_touch of G24103: signal is true;
	signal G24104: std_logic; attribute dont_touch of G24104: signal is true;
	signal G24105: std_logic; attribute dont_touch of G24105: signal is true;
	signal G24106: std_logic; attribute dont_touch of G24106: signal is true;
	signal G24107: std_logic; attribute dont_touch of G24107: signal is true;
	signal G24108: std_logic; attribute dont_touch of G24108: signal is true;
	signal G24109: std_logic; attribute dont_touch of G24109: signal is true;
	signal G24110: std_logic; attribute dont_touch of G24110: signal is true;
	signal G24111: std_logic; attribute dont_touch of G24111: signal is true;
	signal G24112: std_logic; attribute dont_touch of G24112: signal is true;
	signal G24113: std_logic; attribute dont_touch of G24113: signal is true;
	signal G24114: std_logic; attribute dont_touch of G24114: signal is true;
	signal G24115: std_logic; attribute dont_touch of G24115: signal is true;
	signal G24121: std_logic; attribute dont_touch of G24121: signal is true;
	signal G24122: std_logic; attribute dont_touch of G24122: signal is true;
	signal G24123: std_logic; attribute dont_touch of G24123: signal is true;
	signal G24124: std_logic; attribute dont_touch of G24124: signal is true;
	signal G24125: std_logic; attribute dont_touch of G24125: signal is true;
	signal G24126: std_logic; attribute dont_touch of G24126: signal is true;
	signal G24127: std_logic; attribute dont_touch of G24127: signal is true;
	signal G24128: std_logic; attribute dont_touch of G24128: signal is true;
	signal G24129: std_logic; attribute dont_touch of G24129: signal is true;
	signal G24130: std_logic; attribute dont_touch of G24130: signal is true;
	signal G24131: std_logic; attribute dont_touch of G24131: signal is true;
	signal G24132: std_logic; attribute dont_touch of G24132: signal is true;
	signal G24133: std_logic; attribute dont_touch of G24133: signal is true;
	signal G24134: std_logic; attribute dont_touch of G24134: signal is true;
	signal G24140: std_logic; attribute dont_touch of G24140: signal is true;
	signal G24141: std_logic; attribute dont_touch of G24141: signal is true;
	signal G24142: std_logic; attribute dont_touch of G24142: signal is true;
	signal G24143: std_logic; attribute dont_touch of G24143: signal is true;
	signal G24144: std_logic; attribute dont_touch of G24144: signal is true;
	signal G24145: std_logic; attribute dont_touch of G24145: signal is true;
	signal G24146: std_logic; attribute dont_touch of G24146: signal is true;
	signal G24147: std_logic; attribute dont_touch of G24147: signal is true;
	signal G24148: std_logic; attribute dont_touch of G24148: signal is true;
	signal G24149: std_logic; attribute dont_touch of G24149: signal is true;
	signal G24150: std_logic; attribute dont_touch of G24150: signal is true;
	signal G24151: std_logic; attribute dont_touch of G24151: signal is true;
	signal G24152: std_logic; attribute dont_touch of G24152: signal is true;
	signal G24153: std_logic; attribute dont_touch of G24153: signal is true;
	signal G24159: std_logic; attribute dont_touch of G24159: signal is true;
	signal G24160: std_logic; attribute dont_touch of G24160: signal is true;
	signal G24161: std_logic; attribute dont_touch of G24161: signal is true;
	signal G24162: std_logic; attribute dont_touch of G24162: signal is true;
	signal G24163: std_logic; attribute dont_touch of G24163: signal is true;
	signal G24164: std_logic; attribute dont_touch of G24164: signal is true;
	signal G24165: std_logic; attribute dont_touch of G24165: signal is true;
	signal G24166: std_logic; attribute dont_touch of G24166: signal is true;
	signal G24167: std_logic; attribute dont_touch of G24167: signal is true;
	signal G24168: std_logic; attribute dont_touch of G24168: signal is true;
	signal G24174: std_logic; attribute dont_touch of G24174: signal is true;
	signal G24175: std_logic; attribute dont_touch of G24175: signal is true;
	signal G24176: std_logic; attribute dont_touch of G24176: signal is true;
	signal G24177: std_logic; attribute dont_touch of G24177: signal is true;
	signal G24178: std_logic; attribute dont_touch of G24178: signal is true;
	signal G24179: std_logic; attribute dont_touch of G24179: signal is true;
	signal G24180: std_logic; attribute dont_touch of G24180: signal is true;
	signal G24181: std_logic; attribute dont_touch of G24181: signal is true;
	signal G24182: std_logic; attribute dont_touch of G24182: signal is true;
	signal G24183: std_logic; attribute dont_touch of G24183: signal is true;
	signal G24206: std_logic; attribute dont_touch of G24206: signal is true;
	signal G24207: std_logic; attribute dont_touch of G24207: signal is true;
	signal G24208: std_logic; attribute dont_touch of G24208: signal is true;
	signal G24209: std_logic; attribute dont_touch of G24209: signal is true;
	signal G24210: std_logic; attribute dont_touch of G24210: signal is true;
	signal G24211: std_logic; attribute dont_touch of G24211: signal is true;
	signal G24212: std_logic; attribute dont_touch of G24212: signal is true;
	signal G24213: std_logic; attribute dont_touch of G24213: signal is true;
	signal G24214: std_logic; attribute dont_touch of G24214: signal is true;
	signal G24215: std_logic; attribute dont_touch of G24215: signal is true;
	signal G24216: std_logic; attribute dont_touch of G24216: signal is true;
	signal G24217: std_logic; attribute dont_touch of G24217: signal is true;
	signal G24218: std_logic; attribute dont_touch of G24218: signal is true;
	signal G24219: std_logic; attribute dont_touch of G24219: signal is true;
	signal G24220: std_logic; attribute dont_touch of G24220: signal is true;
	signal G24221: std_logic; attribute dont_touch of G24221: signal is true;
	signal G24222: std_logic; attribute dont_touch of G24222: signal is true;
	signal G24223: std_logic; attribute dont_touch of G24223: signal is true;
	signal G24224: std_logic; attribute dont_touch of G24224: signal is true;
	signal G24225: std_logic; attribute dont_touch of G24225: signal is true;
	signal G24226: std_logic; attribute dont_touch of G24226: signal is true;
	signal G24227: std_logic; attribute dont_touch of G24227: signal is true;
	signal G24228: std_logic; attribute dont_touch of G24228: signal is true;
	signal G24229: std_logic; attribute dont_touch of G24229: signal is true;
	signal G24230: std_logic; attribute dont_touch of G24230: signal is true;
	signal G24231: std_logic; attribute dont_touch of G24231: signal is true;
	signal G24232: std_logic; attribute dont_touch of G24232: signal is true;
	signal G24233: std_logic; attribute dont_touch of G24233: signal is true;
	signal G24234: std_logic; attribute dont_touch of G24234: signal is true;
	signal G24235: std_logic; attribute dont_touch of G24235: signal is true;
	signal G24236: std_logic; attribute dont_touch of G24236: signal is true;
	signal G24237: std_logic; attribute dont_touch of G24237: signal is true;
	signal G24238: std_logic; attribute dont_touch of G24238: signal is true;
	signal G24239: std_logic; attribute dont_touch of G24239: signal is true;
	signal G24240: std_logic; attribute dont_touch of G24240: signal is true;
	signal G24241: std_logic; attribute dont_touch of G24241: signal is true;
	signal G24242: std_logic; attribute dont_touch of G24242: signal is true;
	signal G24243: std_logic; attribute dont_touch of G24243: signal is true;
	signal G24244: std_logic; attribute dont_touch of G24244: signal is true;
	signal G24245: std_logic; attribute dont_touch of G24245: signal is true;
	signal G24246: std_logic; attribute dont_touch of G24246: signal is true;
	signal G24247: std_logic; attribute dont_touch of G24247: signal is true;
	signal G24248: std_logic; attribute dont_touch of G24248: signal is true;
	signal G24249: std_logic; attribute dont_touch of G24249: signal is true;
	signal G24250: std_logic; attribute dont_touch of G24250: signal is true;
	signal G24251: std_logic; attribute dont_touch of G24251: signal is true;
	signal G24252: std_logic; attribute dont_touch of G24252: signal is true;
	signal G24253: std_logic; attribute dont_touch of G24253: signal is true;
	signal G24254: std_logic; attribute dont_touch of G24254: signal is true;
	signal G24255: std_logic; attribute dont_touch of G24255: signal is true;
	signal G24256: std_logic; attribute dont_touch of G24256: signal is true;
	signal G24257: std_logic; attribute dont_touch of G24257: signal is true;
	signal G24258: std_logic; attribute dont_touch of G24258: signal is true;
	signal G24259: std_logic; attribute dont_touch of G24259: signal is true;
	signal G24260: std_logic; attribute dont_touch of G24260: signal is true;
	signal G24261: std_logic; attribute dont_touch of G24261: signal is true;
	signal G24262: std_logic; attribute dont_touch of G24262: signal is true;
	signal G24263: std_logic; attribute dont_touch of G24263: signal is true;
	signal G24264: std_logic; attribute dont_touch of G24264: signal is true;
	signal G24265: std_logic; attribute dont_touch of G24265: signal is true;
	signal G24266: std_logic; attribute dont_touch of G24266: signal is true;
	signal G24267: std_logic; attribute dont_touch of G24267: signal is true;
	signal G24268: std_logic; attribute dont_touch of G24268: signal is true;
	signal G24269: std_logic; attribute dont_touch of G24269: signal is true;
	signal G24270: std_logic; attribute dont_touch of G24270: signal is true;
	signal G24271: std_logic; attribute dont_touch of G24271: signal is true;
	signal G24272: std_logic; attribute dont_touch of G24272: signal is true;
	signal G24273: std_logic; attribute dont_touch of G24273: signal is true;
	signal G24274: std_logic; attribute dont_touch of G24274: signal is true;
	signal G24275: std_logic; attribute dont_touch of G24275: signal is true;
	signal G24276: std_logic; attribute dont_touch of G24276: signal is true;
	signal G24277: std_logic; attribute dont_touch of G24277: signal is true;
	signal G24278: std_logic; attribute dont_touch of G24278: signal is true;
	signal G24279: std_logic; attribute dont_touch of G24279: signal is true;
	signal G24280: std_logic; attribute dont_touch of G24280: signal is true;
	signal G24281: std_logic; attribute dont_touch of G24281: signal is true;
	signal G24282: std_logic; attribute dont_touch of G24282: signal is true;
	signal G24283: std_logic; attribute dont_touch of G24283: signal is true;
	signal G24284: std_logic; attribute dont_touch of G24284: signal is true;
	signal G24285: std_logic; attribute dont_touch of G24285: signal is true;
	signal G24286: std_logic; attribute dont_touch of G24286: signal is true;
	signal G24287: std_logic; attribute dont_touch of G24287: signal is true;
	signal G24288: std_logic; attribute dont_touch of G24288: signal is true;
	signal G24289: std_logic; attribute dont_touch of G24289: signal is true;
	signal G24290: std_logic; attribute dont_touch of G24290: signal is true;
	signal G24291: std_logic; attribute dont_touch of G24291: signal is true;
	signal G24292: std_logic; attribute dont_touch of G24292: signal is true;
	signal G24293: std_logic; attribute dont_touch of G24293: signal is true;
	signal G24294: std_logic; attribute dont_touch of G24294: signal is true;
	signal G24295: std_logic; attribute dont_touch of G24295: signal is true;
	signal G24296: std_logic; attribute dont_touch of G24296: signal is true;
	signal G24297: std_logic; attribute dont_touch of G24297: signal is true;
	signal G24298: std_logic; attribute dont_touch of G24298: signal is true;
	signal G24299: std_logic; attribute dont_touch of G24299: signal is true;
	signal G24300: std_logic; attribute dont_touch of G24300: signal is true;
	signal G24301: std_logic; attribute dont_touch of G24301: signal is true;
	signal G24302: std_logic; attribute dont_touch of G24302: signal is true;
	signal G24303: std_logic; attribute dont_touch of G24303: signal is true;
	signal G24304: std_logic; attribute dont_touch of G24304: signal is true;
	signal G24305: std_logic; attribute dont_touch of G24305: signal is true;
	signal G24306: std_logic; attribute dont_touch of G24306: signal is true;
	signal G24307: std_logic; attribute dont_touch of G24307: signal is true;
	signal G24308: std_logic; attribute dont_touch of G24308: signal is true;
	signal G24309: std_logic; attribute dont_touch of G24309: signal is true;
	signal G24310: std_logic; attribute dont_touch of G24310: signal is true;
	signal G24311: std_logic; attribute dont_touch of G24311: signal is true;
	signal G24312: std_logic; attribute dont_touch of G24312: signal is true;
	signal G24313: std_logic; attribute dont_touch of G24313: signal is true;
	signal G24314: std_logic; attribute dont_touch of G24314: signal is true;
	signal G24315: std_logic; attribute dont_touch of G24315: signal is true;
	signal G24316: std_logic; attribute dont_touch of G24316: signal is true;
	signal G24317: std_logic; attribute dont_touch of G24317: signal is true;
	signal G24318: std_logic; attribute dont_touch of G24318: signal is true;
	signal G24319: std_logic; attribute dont_touch of G24319: signal is true;
	signal G24320: std_logic; attribute dont_touch of G24320: signal is true;
	signal G24321: std_logic; attribute dont_touch of G24321: signal is true;
	signal G24322: std_logic; attribute dont_touch of G24322: signal is true;
	signal G24323: std_logic; attribute dont_touch of G24323: signal is true;
	signal G24324: std_logic; attribute dont_touch of G24324: signal is true;
	signal G24325: std_logic; attribute dont_touch of G24325: signal is true;
	signal G24326: std_logic; attribute dont_touch of G24326: signal is true;
	signal G24327: std_logic; attribute dont_touch of G24327: signal is true;
	signal G24328: std_logic; attribute dont_touch of G24328: signal is true;
	signal G24329: std_logic; attribute dont_touch of G24329: signal is true;
	signal G24330: std_logic; attribute dont_touch of G24330: signal is true;
	signal G24331: std_logic; attribute dont_touch of G24331: signal is true;
	signal G24332: std_logic; attribute dont_touch of G24332: signal is true;
	signal G24333: std_logic; attribute dont_touch of G24333: signal is true;
	signal G24334: std_logic; attribute dont_touch of G24334: signal is true;
	signal G24335: std_logic; attribute dont_touch of G24335: signal is true;
	signal G24336: std_logic; attribute dont_touch of G24336: signal is true;
	signal G24337: std_logic; attribute dont_touch of G24337: signal is true;
	signal G24338: std_logic; attribute dont_touch of G24338: signal is true;
	signal G24339: std_logic; attribute dont_touch of G24339: signal is true;
	signal G24340: std_logic; attribute dont_touch of G24340: signal is true;
	signal G24341: std_logic; attribute dont_touch of G24341: signal is true;
	signal G24342: std_logic; attribute dont_touch of G24342: signal is true;
	signal G24343: std_logic; attribute dont_touch of G24343: signal is true;
	signal G24344: std_logic; attribute dont_touch of G24344: signal is true;
	signal G24345: std_logic; attribute dont_touch of G24345: signal is true;
	signal G24346: std_logic; attribute dont_touch of G24346: signal is true;
	signal G24347: std_logic; attribute dont_touch of G24347: signal is true;
	signal G24348: std_logic; attribute dont_touch of G24348: signal is true;
	signal G24349: std_logic; attribute dont_touch of G24349: signal is true;
	signal G24350: std_logic; attribute dont_touch of G24350: signal is true;
	signal G24351: std_logic; attribute dont_touch of G24351: signal is true;
	signal G24352: std_logic; attribute dont_touch of G24352: signal is true;
	signal G24353: std_logic; attribute dont_touch of G24353: signal is true;
	signal G24354: std_logic; attribute dont_touch of G24354: signal is true;
	signal G24355: std_logic; attribute dont_touch of G24355: signal is true;
	signal G24356: std_logic; attribute dont_touch of G24356: signal is true;
	signal G24357: std_logic; attribute dont_touch of G24357: signal is true;
	signal G24358: std_logic; attribute dont_touch of G24358: signal is true;
	signal G24359: std_logic; attribute dont_touch of G24359: signal is true;
	signal G24360: std_logic; attribute dont_touch of G24360: signal is true;
	signal G24361: std_logic; attribute dont_touch of G24361: signal is true;
	signal G24362: std_logic; attribute dont_touch of G24362: signal is true;
	signal G24363: std_logic; attribute dont_touch of G24363: signal is true;
	signal G24364: std_logic; attribute dont_touch of G24364: signal is true;
	signal G24365: std_logic; attribute dont_touch of G24365: signal is true;
	signal G24366: std_logic; attribute dont_touch of G24366: signal is true;
	signal G24367: std_logic; attribute dont_touch of G24367: signal is true;
	signal G24368: std_logic; attribute dont_touch of G24368: signal is true;
	signal G24369: std_logic; attribute dont_touch of G24369: signal is true;
	signal G24370: std_logic; attribute dont_touch of G24370: signal is true;
	signal G24371: std_logic; attribute dont_touch of G24371: signal is true;
	signal G24372: std_logic; attribute dont_touch of G24372: signal is true;
	signal G24373: std_logic; attribute dont_touch of G24373: signal is true;
	signal G24374: std_logic; attribute dont_touch of G24374: signal is true;
	signal G24375: std_logic; attribute dont_touch of G24375: signal is true;
	signal G24376: std_logic; attribute dont_touch of G24376: signal is true;
	signal G24377: std_logic; attribute dont_touch of G24377: signal is true;
	signal G24378: std_logic; attribute dont_touch of G24378: signal is true;
	signal G24379: std_logic; attribute dont_touch of G24379: signal is true;
	signal G24380: std_logic; attribute dont_touch of G24380: signal is true;
	signal G24381: std_logic; attribute dont_touch of G24381: signal is true;
	signal G24382: std_logic; attribute dont_touch of G24382: signal is true;
	signal G24383: std_logic; attribute dont_touch of G24383: signal is true;
	signal G24384: std_logic; attribute dont_touch of G24384: signal is true;
	signal G24385: std_logic; attribute dont_touch of G24385: signal is true;
	signal G24386: std_logic; attribute dont_touch of G24386: signal is true;
	signal G24387: std_logic; attribute dont_touch of G24387: signal is true;
	signal G24388: std_logic; attribute dont_touch of G24388: signal is true;
	signal G24389: std_logic; attribute dont_touch of G24389: signal is true;
	signal G24390: std_logic; attribute dont_touch of G24390: signal is true;
	signal G24391: std_logic; attribute dont_touch of G24391: signal is true;
	signal G24392: std_logic; attribute dont_touch of G24392: signal is true;
	signal G24393: std_logic; attribute dont_touch of G24393: signal is true;
	signal G24394: std_logic; attribute dont_touch of G24394: signal is true;
	signal G24395: std_logic; attribute dont_touch of G24395: signal is true;
	signal G24396: std_logic; attribute dont_touch of G24396: signal is true;
	signal G24397: std_logic; attribute dont_touch of G24397: signal is true;
	signal G24398: std_logic; attribute dont_touch of G24398: signal is true;
	signal G24399: std_logic; attribute dont_touch of G24399: signal is true;
	signal G24400: std_logic; attribute dont_touch of G24400: signal is true;
	signal G24401: std_logic; attribute dont_touch of G24401: signal is true;
	signal G24402: std_logic; attribute dont_touch of G24402: signal is true;
	signal G24403: std_logic; attribute dont_touch of G24403: signal is true;
	signal G24404: std_logic; attribute dont_touch of G24404: signal is true;
	signal G24405: std_logic; attribute dont_touch of G24405: signal is true;
	signal G24406: std_logic; attribute dont_touch of G24406: signal is true;
	signal G24407: std_logic; attribute dont_touch of G24407: signal is true;
	signal G24408: std_logic; attribute dont_touch of G24408: signal is true;
	signal G24409: std_logic; attribute dont_touch of G24409: signal is true;
	signal G24410: std_logic; attribute dont_touch of G24410: signal is true;
	signal G24411: std_logic; attribute dont_touch of G24411: signal is true;
	signal G24412: std_logic; attribute dont_touch of G24412: signal is true;
	signal G24413: std_logic; attribute dont_touch of G24413: signal is true;
	signal G24414: std_logic; attribute dont_touch of G24414: signal is true;
	signal G24415: std_logic; attribute dont_touch of G24415: signal is true;
	signal G24416: std_logic; attribute dont_touch of G24416: signal is true;
	signal G24417: std_logic; attribute dont_touch of G24417: signal is true;
	signal G24418: std_logic; attribute dont_touch of G24418: signal is true;
	signal G24419: std_logic; attribute dont_touch of G24419: signal is true;
	signal G24420: std_logic; attribute dont_touch of G24420: signal is true;
	signal G24421: std_logic; attribute dont_touch of G24421: signal is true;
	signal G24422: std_logic; attribute dont_touch of G24422: signal is true;
	signal G24423: std_logic; attribute dont_touch of G24423: signal is true;
	signal G24424: std_logic; attribute dont_touch of G24424: signal is true;
	signal G24425: std_logic; attribute dont_touch of G24425: signal is true;
	signal G24426: std_logic; attribute dont_touch of G24426: signal is true;
	signal G24427: std_logic; attribute dont_touch of G24427: signal is true;
	signal G24428: std_logic; attribute dont_touch of G24428: signal is true;
	signal G24429: std_logic; attribute dont_touch of G24429: signal is true;
	signal G24430: std_logic; attribute dont_touch of G24430: signal is true;
	signal G24431: std_logic; attribute dont_touch of G24431: signal is true;
	signal G24432: std_logic; attribute dont_touch of G24432: signal is true;
	signal G24433: std_logic; attribute dont_touch of G24433: signal is true;
	signal G24434: std_logic; attribute dont_touch of G24434: signal is true;
	signal G24435: std_logic; attribute dont_touch of G24435: signal is true;
	signal G24436: std_logic; attribute dont_touch of G24436: signal is true;
	signal G24437: std_logic; attribute dont_touch of G24437: signal is true;
	signal G24438: std_logic; attribute dont_touch of G24438: signal is true;
	signal G24439: std_logic; attribute dont_touch of G24439: signal is true;
	signal G24440: std_logic; attribute dont_touch of G24440: signal is true;
	signal G24441: std_logic; attribute dont_touch of G24441: signal is true;
	signal G24442: std_logic; attribute dont_touch of G24442: signal is true;
	signal G24443: std_logic; attribute dont_touch of G24443: signal is true;
	signal G24444: std_logic; attribute dont_touch of G24444: signal is true;
	signal G24445: std_logic; attribute dont_touch of G24445: signal is true;
	signal G24446: std_logic; attribute dont_touch of G24446: signal is true;
	signal G24447: std_logic; attribute dont_touch of G24447: signal is true;
	signal G24448: std_logic; attribute dont_touch of G24448: signal is true;
	signal G24449: std_logic; attribute dont_touch of G24449: signal is true;
	signal G24450: std_logic; attribute dont_touch of G24450: signal is true;
	signal G24451: std_logic; attribute dont_touch of G24451: signal is true;
	signal G24452: std_logic; attribute dont_touch of G24452: signal is true;
	signal G24453: std_logic; attribute dont_touch of G24453: signal is true;
	signal G24454: std_logic; attribute dont_touch of G24454: signal is true;
	signal G24455: std_logic; attribute dont_touch of G24455: signal is true;
	signal G24456: std_logic; attribute dont_touch of G24456: signal is true;
	signal G24457: std_logic; attribute dont_touch of G24457: signal is true;
	signal G24458: std_logic; attribute dont_touch of G24458: signal is true;
	signal G24459: std_logic; attribute dont_touch of G24459: signal is true;
	signal G24460: std_logic; attribute dont_touch of G24460: signal is true;
	signal G24461: std_logic; attribute dont_touch of G24461: signal is true;
	signal G24462: std_logic; attribute dont_touch of G24462: signal is true;
	signal G24463: std_logic; attribute dont_touch of G24463: signal is true;
	signal G24464: std_logic; attribute dont_touch of G24464: signal is true;
	signal G24465: std_logic; attribute dont_touch of G24465: signal is true;
	signal G24466: std_logic; attribute dont_touch of G24466: signal is true;
	signal G24467: std_logic; attribute dont_touch of G24467: signal is true;
	signal G24468: std_logic; attribute dont_touch of G24468: signal is true;
	signal G24469: std_logic; attribute dont_touch of G24469: signal is true;
	signal G24470: std_logic; attribute dont_touch of G24470: signal is true;
	signal G24471: std_logic; attribute dont_touch of G24471: signal is true;
	signal G24472: std_logic; attribute dont_touch of G24472: signal is true;
	signal G24473: std_logic; attribute dont_touch of G24473: signal is true;
	signal G24474: std_logic; attribute dont_touch of G24474: signal is true;
	signal G24475: std_logic; attribute dont_touch of G24475: signal is true;
	signal G24476: std_logic; attribute dont_touch of G24476: signal is true;
	signal G24477: std_logic; attribute dont_touch of G24477: signal is true;
	signal G24478: std_logic; attribute dont_touch of G24478: signal is true;
	signal G24479: std_logic; attribute dont_touch of G24479: signal is true;
	signal G24480: std_logic; attribute dont_touch of G24480: signal is true;
	signal G24481: std_logic; attribute dont_touch of G24481: signal is true;
	signal G24482: std_logic; attribute dont_touch of G24482: signal is true;
	signal G24485: std_logic; attribute dont_touch of G24485: signal is true;
	signal G24486: std_logic; attribute dont_touch of G24486: signal is true;
	signal G24487: std_logic; attribute dont_touch of G24487: signal is true;
	signal G24488: std_logic; attribute dont_touch of G24488: signal is true;
	signal G24489: std_logic; attribute dont_touch of G24489: signal is true;
	signal G24490: std_logic; attribute dont_touch of G24490: signal is true;
	signal G24491: std_logic; attribute dont_touch of G24491: signal is true;
	signal G24492: std_logic; attribute dont_touch of G24492: signal is true;
	signal G24493: std_logic; attribute dont_touch of G24493: signal is true;
	signal G24494: std_logic; attribute dont_touch of G24494: signal is true;
	signal G24495: std_logic; attribute dont_touch of G24495: signal is true;
	signal G24496: std_logic; attribute dont_touch of G24496: signal is true;
	signal G24497: std_logic; attribute dont_touch of G24497: signal is true;
	signal G24498: std_logic; attribute dont_touch of G24498: signal is true;
	signal G24499: std_logic; attribute dont_touch of G24499: signal is true;
	signal G24500: std_logic; attribute dont_touch of G24500: signal is true;
	signal G24501: std_logic; attribute dont_touch of G24501: signal is true;
	signal G24502: std_logic; attribute dont_touch of G24502: signal is true;
	signal G24503: std_logic; attribute dont_touch of G24503: signal is true;
	signal G24504: std_logic; attribute dont_touch of G24504: signal is true;
	signal G24505: std_logic; attribute dont_touch of G24505: signal is true;
	signal G24506: std_logic; attribute dont_touch of G24506: signal is true;
	signal G24507: std_logic; attribute dont_touch of G24507: signal is true;
	signal G24508: std_logic; attribute dont_touch of G24508: signal is true;
	signal G24509: std_logic; attribute dont_touch of G24509: signal is true;
	signal G24510: std_logic; attribute dont_touch of G24510: signal is true;
	signal G24511: std_logic; attribute dont_touch of G24511: signal is true;
	signal G24512: std_logic; attribute dont_touch of G24512: signal is true;
	signal G24513: std_logic; attribute dont_touch of G24513: signal is true;
	signal G24514: std_logic; attribute dont_touch of G24514: signal is true;
	signal G24515: std_logic; attribute dont_touch of G24515: signal is true;
	signal G24516: std_logic; attribute dont_touch of G24516: signal is true;
	signal G24517: std_logic; attribute dont_touch of G24517: signal is true;
	signal G24518: std_logic; attribute dont_touch of G24518: signal is true;
	signal G24519: std_logic; attribute dont_touch of G24519: signal is true;
	signal G24520: std_logic; attribute dont_touch of G24520: signal is true;
	signal G24521: std_logic; attribute dont_touch of G24521: signal is true;
	signal G24522: std_logic; attribute dont_touch of G24522: signal is true;
	signal G24523: std_logic; attribute dont_touch of G24523: signal is true;
	signal G24524: std_logic; attribute dont_touch of G24524: signal is true;
	signal G24525: std_logic; attribute dont_touch of G24525: signal is true;
	signal G24526: std_logic; attribute dont_touch of G24526: signal is true;
	signal G24527: std_logic; attribute dont_touch of G24527: signal is true;
	signal G24528: std_logic; attribute dont_touch of G24528: signal is true;
	signal G24529: std_logic; attribute dont_touch of G24529: signal is true;
	signal G24530: std_logic; attribute dont_touch of G24530: signal is true;
	signal G24531: std_logic; attribute dont_touch of G24531: signal is true;
	signal G24532: std_logic; attribute dont_touch of G24532: signal is true;
	signal G24533: std_logic; attribute dont_touch of G24533: signal is true;
	signal G24534: std_logic; attribute dont_touch of G24534: signal is true;
	signal G24535: std_logic; attribute dont_touch of G24535: signal is true;
	signal G24536: std_logic; attribute dont_touch of G24536: signal is true;
	signal G24537: std_logic; attribute dont_touch of G24537: signal is true;
	signal G24538: std_logic; attribute dont_touch of G24538: signal is true;
	signal G24539: std_logic; attribute dont_touch of G24539: signal is true;
	signal G24540: std_logic; attribute dont_touch of G24540: signal is true;
	signal G24541: std_logic; attribute dont_touch of G24541: signal is true;
	signal G24542: std_logic; attribute dont_touch of G24542: signal is true;
	signal G24543: std_logic; attribute dont_touch of G24543: signal is true;
	signal G24544: std_logic; attribute dont_touch of G24544: signal is true;
	signal G24545: std_logic; attribute dont_touch of G24545: signal is true;
	signal G24546: std_logic; attribute dont_touch of G24546: signal is true;
	signal G24547: std_logic; attribute dont_touch of G24547: signal is true;
	signal G24548: std_logic; attribute dont_touch of G24548: signal is true;
	signal G24549: std_logic; attribute dont_touch of G24549: signal is true;
	signal G24550: std_logic; attribute dont_touch of G24550: signal is true;
	signal G24551: std_logic; attribute dont_touch of G24551: signal is true;
	signal G24552: std_logic; attribute dont_touch of G24552: signal is true;
	signal G24553: std_logic; attribute dont_touch of G24553: signal is true;
	signal G24554: std_logic; attribute dont_touch of G24554: signal is true;
	signal G24555: std_logic; attribute dont_touch of G24555: signal is true;
	signal G24556: std_logic; attribute dont_touch of G24556: signal is true;
	signal G24557: std_logic; attribute dont_touch of G24557: signal is true;
	signal G24558: std_logic; attribute dont_touch of G24558: signal is true;
	signal G24559: std_logic; attribute dont_touch of G24559: signal is true;
	signal G24560: std_logic; attribute dont_touch of G24560: signal is true;
	signal G24561: std_logic; attribute dont_touch of G24561: signal is true;
	signal G24562: std_logic; attribute dont_touch of G24562: signal is true;
	signal G24563: std_logic; attribute dont_touch of G24563: signal is true;
	signal G24564: std_logic; attribute dont_touch of G24564: signal is true;
	signal G24565: std_logic; attribute dont_touch of G24565: signal is true;
	signal G24566: std_logic; attribute dont_touch of G24566: signal is true;
	signal G24567: std_logic; attribute dont_touch of G24567: signal is true;
	signal G24568: std_logic; attribute dont_touch of G24568: signal is true;
	signal G24569: std_logic; attribute dont_touch of G24569: signal is true;
	signal G24570: std_logic; attribute dont_touch of G24570: signal is true;
	signal G24571: std_logic; attribute dont_touch of G24571: signal is true;
	signal G24572: std_logic; attribute dont_touch of G24572: signal is true;
	signal G24573: std_logic; attribute dont_touch of G24573: signal is true;
	signal G24574: std_logic; attribute dont_touch of G24574: signal is true;
	signal G24575: std_logic; attribute dont_touch of G24575: signal is true;
	signal G24576: std_logic; attribute dont_touch of G24576: signal is true;
	signal G24577: std_logic; attribute dont_touch of G24577: signal is true;
	signal G24578: std_logic; attribute dont_touch of G24578: signal is true;
	signal G24579: std_logic; attribute dont_touch of G24579: signal is true;
	signal G24580: std_logic; attribute dont_touch of G24580: signal is true;
	signal G24581: std_logic; attribute dont_touch of G24581: signal is true;
	signal G24582: std_logic; attribute dont_touch of G24582: signal is true;
	signal G24583: std_logic; attribute dont_touch of G24583: signal is true;
	signal G24584: std_logic; attribute dont_touch of G24584: signal is true;
	signal G24585: std_logic; attribute dont_touch of G24585: signal is true;
	signal G24586: std_logic; attribute dont_touch of G24586: signal is true;
	signal G24587: std_logic; attribute dont_touch of G24587: signal is true;
	signal G24588: std_logic; attribute dont_touch of G24588: signal is true;
	signal G24589: std_logic; attribute dont_touch of G24589: signal is true;
	signal G24590: std_logic; attribute dont_touch of G24590: signal is true;
	signal G24591: std_logic; attribute dont_touch of G24591: signal is true;
	signal G24592: std_logic; attribute dont_touch of G24592: signal is true;
	signal G24593: std_logic; attribute dont_touch of G24593: signal is true;
	signal G24594: std_logic; attribute dont_touch of G24594: signal is true;
	signal G24595: std_logic; attribute dont_touch of G24595: signal is true;
	signal G24596: std_logic; attribute dont_touch of G24596: signal is true;
	signal G24597: std_logic; attribute dont_touch of G24597: signal is true;
	signal G24598: std_logic; attribute dont_touch of G24598: signal is true;
	signal G24599: std_logic; attribute dont_touch of G24599: signal is true;
	signal G24600: std_logic; attribute dont_touch of G24600: signal is true;
	signal G24603: std_logic; attribute dont_touch of G24603: signal is true;
	signal G24604: std_logic; attribute dont_touch of G24604: signal is true;
	signal G24605: std_logic; attribute dont_touch of G24605: signal is true;
	signal G24606: std_logic; attribute dont_touch of G24606: signal is true;
	signal G24607: std_logic; attribute dont_touch of G24607: signal is true;
	signal G24610: std_logic; attribute dont_touch of G24610: signal is true;
	signal G24611: std_logic; attribute dont_touch of G24611: signal is true;
	signal G24612: std_logic; attribute dont_touch of G24612: signal is true;
	signal G24613: std_logic; attribute dont_touch of G24613: signal is true;
	signal G24616: std_logic; attribute dont_touch of G24616: signal is true;
	signal G24619: std_logic; attribute dont_touch of G24619: signal is true;
	signal G24622: std_logic; attribute dont_touch of G24622: signal is true;
	signal G24623: std_logic; attribute dont_touch of G24623: signal is true;
	signal G24624: std_logic; attribute dont_touch of G24624: signal is true;
	signal G24627: std_logic; attribute dont_touch of G24627: signal is true;
	signal G24630: std_logic; attribute dont_touch of G24630: signal is true;
	signal G24633: std_logic; attribute dont_touch of G24633: signal is true;
	signal G24636: std_logic; attribute dont_touch of G24636: signal is true;
	signal G24637: std_logic; attribute dont_touch of G24637: signal is true;
	signal G24638: std_logic; attribute dont_touch of G24638: signal is true;
	signal G24641: std_logic; attribute dont_touch of G24641: signal is true;
	signal G24644: std_logic; attribute dont_touch of G24644: signal is true;
	signal G24648: std_logic; attribute dont_touch of G24648: signal is true;
	signal G24652: std_logic; attribute dont_touch of G24652: signal is true;
	signal G24653: std_logic; attribute dont_touch of G24653: signal is true;
	signal G24656: std_logic; attribute dont_touch of G24656: signal is true;
	signal G24657: std_logic; attribute dont_touch of G24657: signal is true;
	signal G24660: std_logic; attribute dont_touch of G24660: signal is true;
	signal G24663: std_logic; attribute dont_touch of G24663: signal is true;
	signal G24664: std_logic; attribute dont_touch of G24664: signal is true;
	signal G24668: std_logic; attribute dont_touch of G24668: signal is true;
	signal G24672: std_logic; attribute dont_touch of G24672: signal is true;
	signal G24675: std_logic; attribute dont_touch of G24675: signal is true;
	signal G24676: std_logic; attribute dont_touch of G24676: signal is true;
	signal G24681: std_logic; attribute dont_touch of G24681: signal is true;
	signal G24682: std_logic; attribute dont_touch of G24682: signal is true;
	signal G24683: std_logic; attribute dont_touch of G24683: signal is true;
	signal G24687: std_logic; attribute dont_touch of G24687: signal is true;
	signal G24691: std_logic; attribute dont_touch of G24691: signal is true;
	signal G24694: std_logic; attribute dont_touch of G24694: signal is true;
	signal G24695: std_logic; attribute dont_touch of G24695: signal is true;
	signal G24700: std_logic; attribute dont_touch of G24700: signal is true;
	signal G24704: std_logic; attribute dont_touch of G24704: signal is true;
	signal G24708: std_logic; attribute dont_touch of G24708: signal is true;
	signal G24711: std_logic; attribute dont_touch of G24711: signal is true;
	signal G24712: std_logic; attribute dont_touch of G24712: signal is true;
	signal G24717: std_logic; attribute dont_touch of G24717: signal is true;
	signal G24720: std_logic; attribute dont_touch of G24720: signal is true;
	signal G24723: std_logic; attribute dont_touch of G24723: signal is true;
	signal G24728: std_logic; attribute dont_touch of G24728: signal is true;
	signal G24731: std_logic; attribute dont_touch of G24731: signal is true;
	signal G24735: std_logic; attribute dont_touch of G24735: signal is true;
	signal G24736: std_logic; attribute dont_touch of G24736: signal is true;
	signal G24739: std_logic; attribute dont_touch of G24739: signal is true;
	signal G24742: std_logic; attribute dont_touch of G24742: signal is true;
	signal G24745: std_logic; attribute dont_touch of G24745: signal is true;
	signal G24746: std_logic; attribute dont_touch of G24746: signal is true;
	signal G24747: std_logic; attribute dont_touch of G24747: signal is true;
	signal G24748: std_logic; attribute dont_touch of G24748: signal is true;
	signal G24749: std_logic; attribute dont_touch of G24749: signal is true;
	signal G24750: std_logic; attribute dont_touch of G24750: signal is true;
	signal G24751: std_logic; attribute dont_touch of G24751: signal is true;
	signal G24752: std_logic; attribute dont_touch of G24752: signal is true;
	signal G24753: std_logic; attribute dont_touch of G24753: signal is true;
	signal G24754: std_logic; attribute dont_touch of G24754: signal is true;
	signal G24755: std_logic; attribute dont_touch of G24755: signal is true;
	signal G24756: std_logic; attribute dont_touch of G24756: signal is true;
	signal G24757: std_logic; attribute dont_touch of G24757: signal is true;
	signal G24758: std_logic; attribute dont_touch of G24758: signal is true;
	signal G24759: std_logic; attribute dont_touch of G24759: signal is true;
	signal G24760: std_logic; attribute dont_touch of G24760: signal is true;
	signal G24761: std_logic; attribute dont_touch of G24761: signal is true;
	signal G24762: std_logic; attribute dont_touch of G24762: signal is true;
	signal G24763: std_logic; attribute dont_touch of G24763: signal is true;
	signal G24766: std_logic; attribute dont_touch of G24766: signal is true;
	signal G24767: std_logic; attribute dont_touch of G24767: signal is true;
	signal G24768: std_logic; attribute dont_touch of G24768: signal is true;
	signal G24769: std_logic; attribute dont_touch of G24769: signal is true;
	signal G24770: std_logic; attribute dont_touch of G24770: signal is true;
	signal G24771: std_logic; attribute dont_touch of G24771: signal is true;
	signal G24772: std_logic; attribute dont_touch of G24772: signal is true;
	signal G24773: std_logic; attribute dont_touch of G24773: signal is true;
	signal G24774: std_logic; attribute dont_touch of G24774: signal is true;
	signal G24775: std_logic; attribute dont_touch of G24775: signal is true;
	signal G24776: std_logic; attribute dont_touch of G24776: signal is true;
	signal G24777: std_logic; attribute dont_touch of G24777: signal is true;
	signal G24778: std_logic; attribute dont_touch of G24778: signal is true;
	signal G24779: std_logic; attribute dont_touch of G24779: signal is true;
	signal G24780: std_logic; attribute dont_touch of G24780: signal is true;
	signal G24781: std_logic; attribute dont_touch of G24781: signal is true;
	signal G24782: std_logic; attribute dont_touch of G24782: signal is true;
	signal G24783: std_logic; attribute dont_touch of G24783: signal is true;
	signal G24784: std_logic; attribute dont_touch of G24784: signal is true;
	signal G24787: std_logic; attribute dont_touch of G24787: signal is true;
	signal G24788: std_logic; attribute dont_touch of G24788: signal is true;
	signal G24789: std_logic; attribute dont_touch of G24789: signal is true;
	signal G24790: std_logic; attribute dont_touch of G24790: signal is true;
	signal G24791: std_logic; attribute dont_touch of G24791: signal is true;
	signal G24792: std_logic; attribute dont_touch of G24792: signal is true;
	signal G24793: std_logic; attribute dont_touch of G24793: signal is true;
	signal G24794: std_logic; attribute dont_touch of G24794: signal is true;
	signal G24795: std_logic; attribute dont_touch of G24795: signal is true;
	signal G24796: std_logic; attribute dont_touch of G24796: signal is true;
	signal G24797: std_logic; attribute dont_touch of G24797: signal is true;
	signal G24798: std_logic; attribute dont_touch of G24798: signal is true;
	signal G24799: std_logic; attribute dont_touch of G24799: signal is true;
	signal G24800: std_logic; attribute dont_touch of G24800: signal is true;
	signal G24801: std_logic; attribute dont_touch of G24801: signal is true;
	signal G24802: std_logic; attribute dont_touch of G24802: signal is true;
	signal G24803: std_logic; attribute dont_touch of G24803: signal is true;
	signal G24804: std_logic; attribute dont_touch of G24804: signal is true;
	signal G24805: std_logic; attribute dont_touch of G24805: signal is true;
	signal G24808: std_logic; attribute dont_touch of G24808: signal is true;
	signal G24809: std_logic; attribute dont_touch of G24809: signal is true;
	signal G24810: std_logic; attribute dont_touch of G24810: signal is true;
	signal G24811: std_logic; attribute dont_touch of G24811: signal is true;
	signal G24812: std_logic; attribute dont_touch of G24812: signal is true;
	signal G24813: std_logic; attribute dont_touch of G24813: signal is true;
	signal G24814: std_logic; attribute dont_touch of G24814: signal is true;
	signal G24815: std_logic; attribute dont_touch of G24815: signal is true;
	signal G24816: std_logic; attribute dont_touch of G24816: signal is true;
	signal G24817: std_logic; attribute dont_touch of G24817: signal is true;
	signal G24818: std_logic; attribute dont_touch of G24818: signal is true;
	signal G24819: std_logic; attribute dont_touch of G24819: signal is true;
	signal G24820: std_logic; attribute dont_touch of G24820: signal is true;
	signal G24821: std_logic; attribute dont_touch of G24821: signal is true;
	signal G24822: std_logic; attribute dont_touch of G24822: signal is true;
	signal G24823: std_logic; attribute dont_touch of G24823: signal is true;
	signal G24824: std_logic; attribute dont_touch of G24824: signal is true;
	signal G24825: std_logic; attribute dont_touch of G24825: signal is true;
	signal G24826: std_logic; attribute dont_touch of G24826: signal is true;
	signal G24827: std_logic; attribute dont_touch of G24827: signal is true;
	signal G24830: std_logic; attribute dont_touch of G24830: signal is true;
	signal G24831: std_logic; attribute dont_touch of G24831: signal is true;
	signal G24832: std_logic; attribute dont_touch of G24832: signal is true;
	signal G24833: std_logic; attribute dont_touch of G24833: signal is true;
	signal G24834: std_logic; attribute dont_touch of G24834: signal is true;
	signal G24835: std_logic; attribute dont_touch of G24835: signal is true;
	signal G24836: std_logic; attribute dont_touch of G24836: signal is true;
	signal G24837: std_logic; attribute dont_touch of G24837: signal is true;
	signal G24838: std_logic; attribute dont_touch of G24838: signal is true;
	signal G24839: std_logic; attribute dont_touch of G24839: signal is true;
	signal G24840: std_logic; attribute dont_touch of G24840: signal is true;
	signal G24841: std_logic; attribute dont_touch of G24841: signal is true;
	signal G24842: std_logic; attribute dont_touch of G24842: signal is true;
	signal G24843: std_logic; attribute dont_touch of G24843: signal is true;
	signal G24844: std_logic; attribute dont_touch of G24844: signal is true;
	signal G24845: std_logic; attribute dont_touch of G24845: signal is true;
	signal G24846: std_logic; attribute dont_touch of G24846: signal is true;
	signal G24847: std_logic; attribute dont_touch of G24847: signal is true;
	signal G24848: std_logic; attribute dont_touch of G24848: signal is true;
	signal G24849: std_logic; attribute dont_touch of G24849: signal is true;
	signal G24850: std_logic; attribute dont_touch of G24850: signal is true;
	signal G24851: std_logic; attribute dont_touch of G24851: signal is true;
	signal G24852: std_logic; attribute dont_touch of G24852: signal is true;
	signal G24853: std_logic; attribute dont_touch of G24853: signal is true;
	signal G24854: std_logic; attribute dont_touch of G24854: signal is true;
	signal G24855: std_logic; attribute dont_touch of G24855: signal is true;
	signal G24856: std_logic; attribute dont_touch of G24856: signal is true;
	signal G24857: std_logic; attribute dont_touch of G24857: signal is true;
	signal G24858: std_logic; attribute dont_touch of G24858: signal is true;
	signal G24859: std_logic; attribute dont_touch of G24859: signal is true;
	signal G24860: std_logic; attribute dont_touch of G24860: signal is true;
	signal G24861: std_logic; attribute dont_touch of G24861: signal is true;
	signal G24862: std_logic; attribute dont_touch of G24862: signal is true;
	signal G24863: std_logic; attribute dont_touch of G24863: signal is true;
	signal G24864: std_logic; attribute dont_touch of G24864: signal is true;
	signal G24865: std_logic; attribute dont_touch of G24865: signal is true;
	signal G24866: std_logic; attribute dont_touch of G24866: signal is true;
	signal G24867: std_logic; attribute dont_touch of G24867: signal is true;
	signal G24868: std_logic; attribute dont_touch of G24868: signal is true;
	signal G24869: std_logic; attribute dont_touch of G24869: signal is true;
	signal G24870: std_logic; attribute dont_touch of G24870: signal is true;
	signal G24871: std_logic; attribute dont_touch of G24871: signal is true;
	signal G24872: std_logic; attribute dont_touch of G24872: signal is true;
	signal G24873: std_logic; attribute dont_touch of G24873: signal is true;
	signal G24874: std_logic; attribute dont_touch of G24874: signal is true;
	signal G24875: std_logic; attribute dont_touch of G24875: signal is true;
	signal G24876: std_logic; attribute dont_touch of G24876: signal is true;
	signal G24877: std_logic; attribute dont_touch of G24877: signal is true;
	signal G24878: std_logic; attribute dont_touch of G24878: signal is true;
	signal G24879: std_logic; attribute dont_touch of G24879: signal is true;
	signal G24880: std_logic; attribute dont_touch of G24880: signal is true;
	signal G24881: std_logic; attribute dont_touch of G24881: signal is true;
	signal G24882: std_logic; attribute dont_touch of G24882: signal is true;
	signal G24883: std_logic; attribute dont_touch of G24883: signal is true;
	signal G24884: std_logic; attribute dont_touch of G24884: signal is true;
	signal G24885: std_logic; attribute dont_touch of G24885: signal is true;
	signal G24886: std_logic; attribute dont_touch of G24886: signal is true;
	signal G24887: std_logic; attribute dont_touch of G24887: signal is true;
	signal G24888: std_logic; attribute dont_touch of G24888: signal is true;
	signal G24889: std_logic; attribute dont_touch of G24889: signal is true;
	signal G24890: std_logic; attribute dont_touch of G24890: signal is true;
	signal G24893: std_logic; attribute dont_touch of G24893: signal is true;
	signal G24897: std_logic; attribute dont_touch of G24897: signal is true;
	signal G24898: std_logic; attribute dont_touch of G24898: signal is true;
	signal G24899: std_logic; attribute dont_touch of G24899: signal is true;
	signal G24900: std_logic; attribute dont_touch of G24900: signal is true;
	signal G24901: std_logic; attribute dont_touch of G24901: signal is true;
	signal G24902: std_logic; attribute dont_touch of G24902: signal is true;
	signal G24903: std_logic; attribute dont_touch of G24903: signal is true;
	signal G24904: std_logic; attribute dont_touch of G24904: signal is true;
	signal G24905: std_logic; attribute dont_touch of G24905: signal is true;
	signal G24906: std_logic; attribute dont_touch of G24906: signal is true;
	signal G24907: std_logic; attribute dont_touch of G24907: signal is true;
	signal G24908: std_logic; attribute dont_touch of G24908: signal is true;
	signal G24909: std_logic; attribute dont_touch of G24909: signal is true;
	signal G24912: std_logic; attribute dont_touch of G24912: signal is true;
	signal G24916: std_logic; attribute dont_touch of G24916: signal is true;
	signal G24920: std_logic; attribute dont_touch of G24920: signal is true;
	signal G24921: std_logic; attribute dont_touch of G24921: signal is true;
	signal G24922: std_logic; attribute dont_touch of G24922: signal is true;
	signal G24923: std_logic; attribute dont_touch of G24923: signal is true;
	signal G24924: std_logic; attribute dont_touch of G24924: signal is true;
	signal G24925: std_logic; attribute dont_touch of G24925: signal is true;
	signal G24928: std_logic; attribute dont_touch of G24928: signal is true;
	signal G24929: std_logic; attribute dont_touch of G24929: signal is true;
	signal G24933: std_logic; attribute dont_touch of G24933: signal is true;
	signal G24937: std_logic; attribute dont_touch of G24937: signal is true;
	signal G24938: std_logic; attribute dont_touch of G24938: signal is true;
	signal G24939: std_logic; attribute dont_touch of G24939: signal is true;
	signal G24940: std_logic; attribute dont_touch of G24940: signal is true;
	signal G24941: std_logic; attribute dont_touch of G24941: signal is true;
	signal G24945: std_logic; attribute dont_touch of G24945: signal is true;
	signal G24949: std_logic; attribute dont_touch of G24949: signal is true;
	signal G24950: std_logic; attribute dont_touch of G24950: signal is true;
	signal G24951: std_logic; attribute dont_touch of G24951: signal is true;
	signal G24952: std_logic; attribute dont_touch of G24952: signal is true;
	signal G24956: std_logic; attribute dont_touch of G24956: signal is true;
	signal G24957: std_logic; attribute dont_touch of G24957: signal is true;
	signal G24958: std_logic; attribute dont_touch of G24958: signal is true;
	signal G24962: std_logic; attribute dont_touch of G24962: signal is true;
	signal G24963: std_logic; attribute dont_touch of G24963: signal is true;
	signal G24964: std_logic; attribute dont_touch of G24964: signal is true;
	signal G24965: std_logic; attribute dont_touch of G24965: signal is true;
	signal G24969: std_logic; attribute dont_touch of G24969: signal is true;
	signal G24973: std_logic; attribute dont_touch of G24973: signal is true;
	signal G24974: std_logic; attribute dont_touch of G24974: signal is true;
	signal G24975: std_logic; attribute dont_touch of G24975: signal is true;
	signal G24978: std_logic; attribute dont_touch of G24978: signal is true;
	signal G24982: std_logic; attribute dont_touch of G24982: signal is true;
	signal G24986: std_logic; attribute dont_touch of G24986: signal is true;
	signal G24989: std_logic; attribute dont_touch of G24989: signal is true;
	signal G24993: std_logic; attribute dont_touch of G24993: signal is true;
	signal G24997: std_logic; attribute dont_touch of G24997: signal is true;
	signal G25000: std_logic; attribute dont_touch of G25000: signal is true;
	signal G25004: std_logic; attribute dont_touch of G25004: signal is true;
	signal G25005: std_logic; attribute dont_touch of G25005: signal is true;
	signal G25008: std_logic; attribute dont_touch of G25008: signal is true;
	signal G25009: std_logic; attribute dont_touch of G25009: signal is true;
	signal G25010: std_logic; attribute dont_touch of G25010: signal is true;
	signal G25011: std_logic; attribute dont_touch of G25011: signal is true;
	signal G25012: std_logic; attribute dont_touch of G25012: signal is true;
	signal G25013: std_logic; attribute dont_touch of G25013: signal is true;
	signal G25014: std_logic; attribute dont_touch of G25014: signal is true;
	signal G25015: std_logic; attribute dont_touch of G25015: signal is true;
	signal G25016: std_logic; attribute dont_touch of G25016: signal is true;
	signal G25017: std_logic; attribute dont_touch of G25017: signal is true;
	signal G25018: std_logic; attribute dont_touch of G25018: signal is true;
	signal G25019: std_logic; attribute dont_touch of G25019: signal is true;
	signal G25020: std_logic; attribute dont_touch of G25020: signal is true;
	signal G25021: std_logic; attribute dont_touch of G25021: signal is true;
	signal G25022: std_logic; attribute dont_touch of G25022: signal is true;
	signal G25023: std_logic; attribute dont_touch of G25023: signal is true;
	signal G25024: std_logic; attribute dont_touch of G25024: signal is true;
	signal G25025: std_logic; attribute dont_touch of G25025: signal is true;
	signal G25026: std_logic; attribute dont_touch of G25026: signal is true;
	signal G25027: std_logic; attribute dont_touch of G25027: signal is true;
	signal G25028: std_logic; attribute dont_touch of G25028: signal is true;
	signal G25029: std_logic; attribute dont_touch of G25029: signal is true;
	signal G25030: std_logic; attribute dont_touch of G25030: signal is true;
	signal G25031: std_logic; attribute dont_touch of G25031: signal is true;
	signal G25032: std_logic; attribute dont_touch of G25032: signal is true;
	signal G25033: std_logic; attribute dont_touch of G25033: signal is true;
	signal G25034: std_logic; attribute dont_touch of G25034: signal is true;
	signal G25035: std_logic; attribute dont_touch of G25035: signal is true;
	signal G25036: std_logic; attribute dont_touch of G25036: signal is true;
	signal G25037: std_logic; attribute dont_touch of G25037: signal is true;
	signal G25038: std_logic; attribute dont_touch of G25038: signal is true;
	signal G25039: std_logic; attribute dont_touch of G25039: signal is true;
	signal G25040: std_logic; attribute dont_touch of G25040: signal is true;
	signal G25041: std_logic; attribute dont_touch of G25041: signal is true;
	signal G25042: std_logic; attribute dont_touch of G25042: signal is true;
	signal G25043: std_logic; attribute dont_touch of G25043: signal is true;
	signal G25044: std_logic; attribute dont_touch of G25044: signal is true;
	signal G25045: std_logic; attribute dont_touch of G25045: signal is true;
	signal G25046: std_logic; attribute dont_touch of G25046: signal is true;
	signal G25047: std_logic; attribute dont_touch of G25047: signal is true;
	signal G25048: std_logic; attribute dont_touch of G25048: signal is true;
	signal G25049: std_logic; attribute dont_touch of G25049: signal is true;
	signal G25050: std_logic; attribute dont_touch of G25050: signal is true;
	signal G25051: std_logic; attribute dont_touch of G25051: signal is true;
	signal G25052: std_logic; attribute dont_touch of G25052: signal is true;
	signal G25053: std_logic; attribute dont_touch of G25053: signal is true;
	signal G25054: std_logic; attribute dont_touch of G25054: signal is true;
	signal G25055: std_logic; attribute dont_touch of G25055: signal is true;
	signal G25056: std_logic; attribute dont_touch of G25056: signal is true;
	signal G25057: std_logic; attribute dont_touch of G25057: signal is true;
	signal G25058: std_logic; attribute dont_touch of G25058: signal is true;
	signal G25059: std_logic; attribute dont_touch of G25059: signal is true;
	signal G25060: std_logic; attribute dont_touch of G25060: signal is true;
	signal G25061: std_logic; attribute dont_touch of G25061: signal is true;
	signal G25062: std_logic; attribute dont_touch of G25062: signal is true;
	signal G25063: std_logic; attribute dont_touch of G25063: signal is true;
	signal G25064: std_logic; attribute dont_touch of G25064: signal is true;
	signal G25065: std_logic; attribute dont_touch of G25065: signal is true;
	signal G25066: std_logic; attribute dont_touch of G25066: signal is true;
	signal G25067: std_logic; attribute dont_touch of G25067: signal is true;
	signal G25068: std_logic; attribute dont_touch of G25068: signal is true;
	signal G25069: std_logic; attribute dont_touch of G25069: signal is true;
	signal G25070: std_logic; attribute dont_touch of G25070: signal is true;
	signal G25071: std_logic; attribute dont_touch of G25071: signal is true;
	signal G25072: std_logic; attribute dont_touch of G25072: signal is true;
	signal G25073: std_logic; attribute dont_touch of G25073: signal is true;
	signal G25074: std_logic; attribute dont_touch of G25074: signal is true;
	signal G25075: std_logic; attribute dont_touch of G25075: signal is true;
	signal G25076: std_logic; attribute dont_touch of G25076: signal is true;
	signal G25077: std_logic; attribute dont_touch of G25077: signal is true;
	signal G25078: std_logic; attribute dont_touch of G25078: signal is true;
	signal G25081: std_logic; attribute dont_touch of G25081: signal is true;
	signal G25082: std_logic; attribute dont_touch of G25082: signal is true;
	signal G25085: std_logic; attribute dont_touch of G25085: signal is true;
	signal G25086: std_logic; attribute dont_touch of G25086: signal is true;
	signal G25087: std_logic; attribute dont_touch of G25087: signal is true;
	signal G25088: std_logic; attribute dont_touch of G25088: signal is true;
	signal G25091: std_logic; attribute dont_touch of G25091: signal is true;
	signal G25094: std_logic; attribute dont_touch of G25094: signal is true;
	signal G25095: std_logic; attribute dont_touch of G25095: signal is true;
	signal G25096: std_logic; attribute dont_touch of G25096: signal is true;
	signal G25099: std_logic; attribute dont_touch of G25099: signal is true;
	signal G25102: std_logic; attribute dont_touch of G25102: signal is true;
	signal G25103: std_logic; attribute dont_touch of G25103: signal is true;
	signal G25104: std_logic; attribute dont_touch of G25104: signal is true;
	signal G25105: std_logic; attribute dont_touch of G25105: signal is true;
	signal G25106: std_logic; attribute dont_touch of G25106: signal is true;
	signal G25109: std_logic; attribute dont_touch of G25109: signal is true;
	signal G25110: std_logic; attribute dont_touch of G25110: signal is true;
	signal G25111: std_logic; attribute dont_touch of G25111: signal is true;
	signal G25112: std_logic; attribute dont_touch of G25112: signal is true;
	signal G25115: std_logic; attribute dont_touch of G25115: signal is true;
	signal G25116: std_logic; attribute dont_touch of G25116: signal is true;
	signal G25117: std_logic; attribute dont_touch of G25117: signal is true;
	signal G25118: std_logic; attribute dont_touch of G25118: signal is true;
	signal G25119: std_logic; attribute dont_touch of G25119: signal is true;
	signal G25120: std_logic; attribute dont_touch of G25120: signal is true;
	signal G25121: std_logic; attribute dont_touch of G25121: signal is true;
	signal G25122: std_logic; attribute dont_touch of G25122: signal is true;
	signal G25123: std_logic; attribute dont_touch of G25123: signal is true;
	signal G25124: std_logic; attribute dont_touch of G25124: signal is true;
	signal G25125: std_logic; attribute dont_touch of G25125: signal is true;
	signal G25126: std_logic; attribute dont_touch of G25126: signal is true;
	signal G25127: std_logic; attribute dont_touch of G25127: signal is true;
	signal G25128: std_logic; attribute dont_touch of G25128: signal is true;
	signal G25129: std_logic; attribute dont_touch of G25129: signal is true;
	signal G25130: std_logic; attribute dont_touch of G25130: signal is true;
	signal G25131: std_logic; attribute dont_touch of G25131: signal is true;
	signal G25132: std_logic; attribute dont_touch of G25132: signal is true;
	signal G25133: std_logic; attribute dont_touch of G25133: signal is true;
	signal G25134: std_logic; attribute dont_touch of G25134: signal is true;
	signal G25135: std_logic; attribute dont_touch of G25135: signal is true;
	signal G25136: std_logic; attribute dont_touch of G25136: signal is true;
	signal G25137: std_logic; attribute dont_touch of G25137: signal is true;
	signal G25138: std_logic; attribute dont_touch of G25138: signal is true;
	signal G25139: std_logic; attribute dont_touch of G25139: signal is true;
	signal G25140: std_logic; attribute dont_touch of G25140: signal is true;
	signal G25141: std_logic; attribute dont_touch of G25141: signal is true;
	signal G25142: std_logic; attribute dont_touch of G25142: signal is true;
	signal G25143: std_logic; attribute dont_touch of G25143: signal is true;
	signal G25144: std_logic; attribute dont_touch of G25144: signal is true;
	signal G25145: std_logic; attribute dont_touch of G25145: signal is true;
	signal G25146: std_logic; attribute dont_touch of G25146: signal is true;
	signal G25147: std_logic; attribute dont_touch of G25147: signal is true;
	signal G25148: std_logic; attribute dont_touch of G25148: signal is true;
	signal G25149: std_logic; attribute dont_touch of G25149: signal is true;
	signal G25150: std_logic; attribute dont_touch of G25150: signal is true;
	signal G25151: std_logic; attribute dont_touch of G25151: signal is true;
	signal G25152: std_logic; attribute dont_touch of G25152: signal is true;
	signal G25153: std_logic; attribute dont_touch of G25153: signal is true;
	signal G25154: std_logic; attribute dont_touch of G25154: signal is true;
	signal G25155: std_logic; attribute dont_touch of G25155: signal is true;
	signal G25156: std_logic; attribute dont_touch of G25156: signal is true;
	signal G25157: std_logic; attribute dont_touch of G25157: signal is true;
	signal G25158: std_logic; attribute dont_touch of G25158: signal is true;
	signal G25159: std_logic; attribute dont_touch of G25159: signal is true;
	signal G25160: std_logic; attribute dont_touch of G25160: signal is true;
	signal G25161: std_logic; attribute dont_touch of G25161: signal is true;
	signal G25162: std_logic; attribute dont_touch of G25162: signal is true;
	signal G25163: std_logic; attribute dont_touch of G25163: signal is true;
	signal G25164: std_logic; attribute dont_touch of G25164: signal is true;
	signal G25165: std_logic; attribute dont_touch of G25165: signal is true;
	signal G25166: std_logic; attribute dont_touch of G25166: signal is true;
	signal G25167: std_logic; attribute dont_touch of G25167: signal is true;
	signal G25168: std_logic; attribute dont_touch of G25168: signal is true;
	signal G25169: std_logic; attribute dont_touch of G25169: signal is true;
	signal G25170: std_logic; attribute dont_touch of G25170: signal is true;
	signal G25171: std_logic; attribute dont_touch of G25171: signal is true;
	signal G25172: std_logic; attribute dont_touch of G25172: signal is true;
	signal G25173: std_logic; attribute dont_touch of G25173: signal is true;
	signal G25174: std_logic; attribute dont_touch of G25174: signal is true;
	signal G25175: std_logic; attribute dont_touch of G25175: signal is true;
	signal G25176: std_logic; attribute dont_touch of G25176: signal is true;
	signal G25177: std_logic; attribute dont_touch of G25177: signal is true;
	signal G25178: std_logic; attribute dont_touch of G25178: signal is true;
	signal G25179: std_logic; attribute dont_touch of G25179: signal is true;
	signal G25180: std_logic; attribute dont_touch of G25180: signal is true;
	signal G25181: std_logic; attribute dont_touch of G25181: signal is true;
	signal G25182: std_logic; attribute dont_touch of G25182: signal is true;
	signal G25183: std_logic; attribute dont_touch of G25183: signal is true;
	signal G25184: std_logic; attribute dont_touch of G25184: signal is true;
	signal G25185: std_logic; attribute dont_touch of G25185: signal is true;
	signal G25186: std_logic; attribute dont_touch of G25186: signal is true;
	signal G25187: std_logic; attribute dont_touch of G25187: signal is true;
	signal G25188: std_logic; attribute dont_touch of G25188: signal is true;
	signal G25189: std_logic; attribute dont_touch of G25189: signal is true;
	signal G25190: std_logic; attribute dont_touch of G25190: signal is true;
	signal G25191: std_logic; attribute dont_touch of G25191: signal is true;
	signal G25192: std_logic; attribute dont_touch of G25192: signal is true;
	signal G25193: std_logic; attribute dont_touch of G25193: signal is true;
	signal G25194: std_logic; attribute dont_touch of G25194: signal is true;
	signal G25195: std_logic; attribute dont_touch of G25195: signal is true;
	signal G25196: std_logic; attribute dont_touch of G25196: signal is true;
	signal G25197: std_logic; attribute dont_touch of G25197: signal is true;
	signal G25198: std_logic; attribute dont_touch of G25198: signal is true;
	signal G25199: std_logic; attribute dont_touch of G25199: signal is true;
	signal G25200: std_logic; attribute dont_touch of G25200: signal is true;
	signal G25201: std_logic; attribute dont_touch of G25201: signal is true;
	signal G25202: std_logic; attribute dont_touch of G25202: signal is true;
	signal G25203: std_logic; attribute dont_touch of G25203: signal is true;
	signal G25204: std_logic; attribute dont_touch of G25204: signal is true;
	signal G25205: std_logic; attribute dont_touch of G25205: signal is true;
	signal G25206: std_logic; attribute dont_touch of G25206: signal is true;
	signal G25207: std_logic; attribute dont_touch of G25207: signal is true;
	signal G25208: std_logic; attribute dont_touch of G25208: signal is true;
	signal G25209: std_logic; attribute dont_touch of G25209: signal is true;
	signal G25210: std_logic; attribute dont_touch of G25210: signal is true;
	signal G25211: std_logic; attribute dont_touch of G25211: signal is true;
	signal G25212: std_logic; attribute dont_touch of G25212: signal is true;
	signal G25213: std_logic; attribute dont_touch of G25213: signal is true;
	signal G25214: std_logic; attribute dont_touch of G25214: signal is true;
	signal G25215: std_logic; attribute dont_touch of G25215: signal is true;
	signal G25216: std_logic; attribute dont_touch of G25216: signal is true;
	signal G25217: std_logic; attribute dont_touch of G25217: signal is true;
	signal G25218: std_logic; attribute dont_touch of G25218: signal is true;
	signal G25219: std_logic; attribute dont_touch of G25219: signal is true;
	signal G25220: std_logic; attribute dont_touch of G25220: signal is true;
	signal G25221: std_logic; attribute dont_touch of G25221: signal is true;
	signal G25222: std_logic; attribute dont_touch of G25222: signal is true;
	signal G25223: std_logic; attribute dont_touch of G25223: signal is true;
	signal G25224: std_logic; attribute dont_touch of G25224: signal is true;
	signal G25225: std_logic; attribute dont_touch of G25225: signal is true;
	signal G25226: std_logic; attribute dont_touch of G25226: signal is true;
	signal G25227: std_logic; attribute dont_touch of G25227: signal is true;
	signal G25228: std_logic; attribute dont_touch of G25228: signal is true;
	signal G25229: std_logic; attribute dont_touch of G25229: signal is true;
	signal G25230: std_logic; attribute dont_touch of G25230: signal is true;
	signal G25231: std_logic; attribute dont_touch of G25231: signal is true;
	signal G25232: std_logic; attribute dont_touch of G25232: signal is true;
	signal G25233: std_logic; attribute dont_touch of G25233: signal is true;
	signal G25234: std_logic; attribute dont_touch of G25234: signal is true;
	signal G25235: std_logic; attribute dont_touch of G25235: signal is true;
	signal G25236: std_logic; attribute dont_touch of G25236: signal is true;
	signal G25237: std_logic; attribute dont_touch of G25237: signal is true;
	signal G25238: std_logic; attribute dont_touch of G25238: signal is true;
	signal G25239: std_logic; attribute dont_touch of G25239: signal is true;
	signal G25240: std_logic; attribute dont_touch of G25240: signal is true;
	signal G25241: std_logic; attribute dont_touch of G25241: signal is true;
	signal G25242: std_logic; attribute dont_touch of G25242: signal is true;
	signal G25243: std_logic; attribute dont_touch of G25243: signal is true;
	signal G25244: std_logic; attribute dont_touch of G25244: signal is true;
	signal G25245: std_logic; attribute dont_touch of G25245: signal is true;
	signal G25246: std_logic; attribute dont_touch of G25246: signal is true;
	signal G25247: std_logic; attribute dont_touch of G25247: signal is true;
	signal G25248: std_logic; attribute dont_touch of G25248: signal is true;
	signal G25249: std_logic; attribute dont_touch of G25249: signal is true;
	signal G25250: std_logic; attribute dont_touch of G25250: signal is true;
	signal G25251: std_logic; attribute dont_touch of G25251: signal is true;
	signal G25252: std_logic; attribute dont_touch of G25252: signal is true;
	signal G25253: std_logic; attribute dont_touch of G25253: signal is true;
	signal G25254: std_logic; attribute dont_touch of G25254: signal is true;
	signal G25255: std_logic; attribute dont_touch of G25255: signal is true;
	signal G25256: std_logic; attribute dont_touch of G25256: signal is true;
	signal G25257: std_logic; attribute dont_touch of G25257: signal is true;
	signal G25258: std_logic; attribute dont_touch of G25258: signal is true;
	signal G25259: std_logic; attribute dont_touch of G25259: signal is true;
	signal G25260: std_logic; attribute dont_touch of G25260: signal is true;
	signal G25261: std_logic; attribute dont_touch of G25261: signal is true;
	signal G25262: std_logic; attribute dont_touch of G25262: signal is true;
	signal G25263: std_logic; attribute dont_touch of G25263: signal is true;
	signal G25264: std_logic; attribute dont_touch of G25264: signal is true;
	signal G25265: std_logic; attribute dont_touch of G25265: signal is true;
	signal G25266: std_logic; attribute dont_touch of G25266: signal is true;
	signal G25267: std_logic; attribute dont_touch of G25267: signal is true;
	signal G25268: std_logic; attribute dont_touch of G25268: signal is true;
	signal G25269: std_logic; attribute dont_touch of G25269: signal is true;
	signal G25270: std_logic; attribute dont_touch of G25270: signal is true;
	signal G25271: std_logic; attribute dont_touch of G25271: signal is true;
	signal G25272: std_logic; attribute dont_touch of G25272: signal is true;
	signal G25273: std_logic; attribute dont_touch of G25273: signal is true;
	signal G25274: std_logic; attribute dont_touch of G25274: signal is true;
	signal G25277: std_logic; attribute dont_touch of G25277: signal is true;
	signal G25278: std_logic; attribute dont_touch of G25278: signal is true;
	signal G25279: std_logic; attribute dont_touch of G25279: signal is true;
	signal G25280: std_logic; attribute dont_touch of G25280: signal is true;
	signal G25281: std_logic; attribute dont_touch of G25281: signal is true;
	signal G25282: std_logic; attribute dont_touch of G25282: signal is true;
	signal G25283: std_logic; attribute dont_touch of G25283: signal is true;
	signal G25286: std_logic; attribute dont_touch of G25286: signal is true;
	signal G25287: std_logic; attribute dont_touch of G25287: signal is true;
	signal G25288: std_logic; attribute dont_touch of G25288: signal is true;
	signal G25289: std_logic; attribute dont_touch of G25289: signal is true;
	signal G25290: std_logic; attribute dont_touch of G25290: signal is true;
	signal G25291: std_logic; attribute dont_touch of G25291: signal is true;
	signal G25294: std_logic; attribute dont_touch of G25294: signal is true;
	signal G25295: std_logic; attribute dont_touch of G25295: signal is true;
	signal G25296: std_logic; attribute dont_touch of G25296: signal is true;
	signal G25299: std_logic; attribute dont_touch of G25299: signal is true;
	signal G25300: std_logic; attribute dont_touch of G25300: signal is true;
	signal G25301: std_logic; attribute dont_touch of G25301: signal is true;
	signal G25304: std_logic; attribute dont_touch of G25304: signal is true;
	signal G25305: std_logic; attribute dont_touch of G25305: signal is true;
	signal G25306: std_logic; attribute dont_touch of G25306: signal is true;
	signal G25309: std_logic; attribute dont_touch of G25309: signal is true;
	signal G25310: std_logic; attribute dont_touch of G25310: signal is true;
	signal G25311: std_logic; attribute dont_touch of G25311: signal is true;
	signal G25312: std_logic; attribute dont_touch of G25312: signal is true;
	signal G25313: std_logic; attribute dont_touch of G25313: signal is true;
	signal G25314: std_logic; attribute dont_touch of G25314: signal is true;
	signal G25315: std_logic; attribute dont_touch of G25315: signal is true;
	signal G25318: std_logic; attribute dont_touch of G25318: signal is true;
	signal G25319: std_logic; attribute dont_touch of G25319: signal is true;
	signal G25320: std_logic; attribute dont_touch of G25320: signal is true;
	signal G25321: std_logic; attribute dont_touch of G25321: signal is true;
	signal G25322: std_logic; attribute dont_touch of G25322: signal is true;
	signal G25323: std_logic; attribute dont_touch of G25323: signal is true;
	signal G25324: std_logic; attribute dont_touch of G25324: signal is true;
	signal G25327: std_logic; attribute dont_touch of G25327: signal is true;
	signal G25328: std_logic; attribute dont_touch of G25328: signal is true;
	signal G25329: std_logic; attribute dont_touch of G25329: signal is true;
	signal G25330: std_logic; attribute dont_touch of G25330: signal is true;
	signal G25331: std_logic; attribute dont_touch of G25331: signal is true;
	signal G25332: std_logic; attribute dont_touch of G25332: signal is true;
	signal G25333: std_logic; attribute dont_touch of G25333: signal is true;
	signal G25334: std_logic; attribute dont_touch of G25334: signal is true;
	signal G25335: std_logic; attribute dont_touch of G25335: signal is true;
	signal G25336: std_logic; attribute dont_touch of G25336: signal is true;
	signal G25337: std_logic; attribute dont_touch of G25337: signal is true;
	signal G25338: std_logic; attribute dont_touch of G25338: signal is true;
	signal G25339: std_logic; attribute dont_touch of G25339: signal is true;
	signal G25340: std_logic; attribute dont_touch of G25340: signal is true;
	signal G25341: std_logic; attribute dont_touch of G25341: signal is true;
	signal G25342: std_logic; attribute dont_touch of G25342: signal is true;
	signal G25343: std_logic; attribute dont_touch of G25343: signal is true;
	signal G25346: std_logic; attribute dont_touch of G25346: signal is true;
	signal G25347: std_logic; attribute dont_touch of G25347: signal is true;
	signal G25348: std_logic; attribute dont_touch of G25348: signal is true;
	signal G25349: std_logic; attribute dont_touch of G25349: signal is true;
	signal G25350: std_logic; attribute dont_touch of G25350: signal is true;
	signal G25351: std_logic; attribute dont_touch of G25351: signal is true;
	signal G25352: std_logic; attribute dont_touch of G25352: signal is true;
	signal G25353: std_logic; attribute dont_touch of G25353: signal is true;
	signal G25354: std_logic; attribute dont_touch of G25354: signal is true;
	signal G25355: std_logic; attribute dont_touch of G25355: signal is true;
	signal G25356: std_logic; attribute dont_touch of G25356: signal is true;
	signal G25357: std_logic; attribute dont_touch of G25357: signal is true;
	signal G25360: std_logic; attribute dont_touch of G25360: signal is true;
	signal G25361: std_logic; attribute dont_touch of G25361: signal is true;
	signal G25362: std_logic; attribute dont_touch of G25362: signal is true;
	signal G25363: std_logic; attribute dont_touch of G25363: signal is true;
	signal G25364: std_logic; attribute dont_touch of G25364: signal is true;
	signal G25365: std_logic; attribute dont_touch of G25365: signal is true;
	signal G25366: std_logic; attribute dont_touch of G25366: signal is true;
	signal G25367: std_logic; attribute dont_touch of G25367: signal is true;
	signal G25368: std_logic; attribute dont_touch of G25368: signal is true;
	signal G25369: std_logic; attribute dont_touch of G25369: signal is true;
	signal G25370: std_logic; attribute dont_touch of G25370: signal is true;
	signal G25371: std_logic; attribute dont_touch of G25371: signal is true;
	signal G25372: std_logic; attribute dont_touch of G25372: signal is true;
	signal G25375: std_logic; attribute dont_touch of G25375: signal is true;
	signal G25376: std_logic; attribute dont_touch of G25376: signal is true;
	signal G25377: std_logic; attribute dont_touch of G25377: signal is true;
	signal G25378: std_logic; attribute dont_touch of G25378: signal is true;
	signal G25379: std_logic; attribute dont_touch of G25379: signal is true;
	signal G25383: std_logic; attribute dont_touch of G25383: signal is true;
	signal G25384: std_logic; attribute dont_touch of G25384: signal is true;
	signal G25385: std_logic; attribute dont_touch of G25385: signal is true;
	signal G25386: std_logic; attribute dont_touch of G25386: signal is true;
	signal G25387: std_logic; attribute dont_touch of G25387: signal is true;
	signal G25388: std_logic; attribute dont_touch of G25388: signal is true;
	signal G25389: std_logic; attribute dont_touch of G25389: signal is true;
	signal G25392: std_logic; attribute dont_touch of G25392: signal is true;
	signal G25393: std_logic; attribute dont_touch of G25393: signal is true;
	signal G25394: std_logic; attribute dont_touch of G25394: signal is true;
	signal G25395: std_logic; attribute dont_touch of G25395: signal is true;
	signal G25399: std_logic; attribute dont_touch of G25399: signal is true;
	signal G25400: std_logic; attribute dont_touch of G25400: signal is true;
	signal G25401: std_logic; attribute dont_touch of G25401: signal is true;
	signal G25402: std_logic; attribute dont_touch of G25402: signal is true;
	signal G25403: std_logic; attribute dont_touch of G25403: signal is true;
	signal G25404: std_logic; attribute dont_touch of G25404: signal is true;
	signal G25405: std_logic; attribute dont_touch of G25405: signal is true;
	signal G25409: std_logic; attribute dont_touch of G25409: signal is true;
	signal G25410: std_logic; attribute dont_touch of G25410: signal is true;
	signal G25411: std_logic; attribute dont_touch of G25411: signal is true;
	signal G25412: std_logic; attribute dont_touch of G25412: signal is true;
	signal G25413: std_logic; attribute dont_touch of G25413: signal is true;
	signal G25417: std_logic; attribute dont_touch of G25417: signal is true;
	signal G25418: std_logic; attribute dont_touch of G25418: signal is true;
	signal G25419: std_logic; attribute dont_touch of G25419: signal is true;
	signal G25421: std_logic; attribute dont_touch of G25421: signal is true;
	signal G25422: std_logic; attribute dont_touch of G25422: signal is true;
	signal G25426: std_logic; attribute dont_touch of G25426: signal is true;
	signal G25429: std_logic; attribute dont_touch of G25429: signal is true;
	signal G25430: std_logic; attribute dont_touch of G25430: signal is true;
	signal G25431: std_logic; attribute dont_touch of G25431: signal is true;
	signal G25436: std_logic; attribute dont_touch of G25436: signal is true;
	signal G25437: std_logic; attribute dont_touch of G25437: signal is true;
	signal G25438: std_logic; attribute dont_touch of G25438: signal is true;
	signal G25443: std_logic; attribute dont_touch of G25443: signal is true;
	signal G25444: std_logic; attribute dont_touch of G25444: signal is true;
	signal G25445: std_logic; attribute dont_touch of G25445: signal is true;
	signal G25449: std_logic; attribute dont_touch of G25449: signal is true;
	signal G25450: std_logic; attribute dont_touch of G25450: signal is true;
	signal G25451: std_logic; attribute dont_touch of G25451: signal is true;
	signal G25452: std_logic; attribute dont_touch of G25452: signal is true;
	signal G25453: std_logic; attribute dont_touch of G25453: signal is true;
	signal G25454: std_logic; attribute dont_touch of G25454: signal is true;
	signal G25457: std_logic; attribute dont_touch of G25457: signal is true;
	signal G25458: std_logic; attribute dont_touch of G25458: signal is true;
	signal G25461: std_logic; attribute dont_touch of G25461: signal is true;
	signal G25462: std_logic; attribute dont_touch of G25462: signal is true;
	signal G25463: std_logic; attribute dont_touch of G25463: signal is true;
	signal G25466: std_logic; attribute dont_touch of G25466: signal is true;
	signal G25467: std_logic; attribute dont_touch of G25467: signal is true;
	signal G25470: std_logic; attribute dont_touch of G25470: signal is true;
	signal G25471: std_logic; attribute dont_touch of G25471: signal is true;
	signal G25472: std_logic; attribute dont_touch of G25472: signal is true;
	signal G25475: std_logic; attribute dont_touch of G25475: signal is true;
	signal G25476: std_logic; attribute dont_touch of G25476: signal is true;
	signal G25479: std_logic; attribute dont_touch of G25479: signal is true;
	signal G25482: std_logic; attribute dont_touch of G25482: signal is true;
	signal G25483: std_logic; attribute dont_touch of G25483: signal is true;
	signal G25484: std_logic; attribute dont_touch of G25484: signal is true;
	signal G25487: std_logic; attribute dont_touch of G25487: signal is true;
	signal G25488: std_logic; attribute dont_touch of G25488: signal is true;
	signal G25490: std_logic; attribute dont_touch of G25490: signal is true;
	signal G25493: std_logic; attribute dont_touch of G25493: signal is true;
	signal G25496: std_logic; attribute dont_touch of G25496: signal is true;
	signal G25499: std_logic; attribute dont_touch of G25499: signal is true;
	signal G25502: std_logic; attribute dont_touch of G25502: signal is true;
	signal G25505: std_logic; attribute dont_touch of G25505: signal is true;
	signal G25506: std_logic; attribute dont_touch of G25506: signal is true;
	signal G25507: std_logic; attribute dont_touch of G25507: signal is true;
	signal G25510: std_logic; attribute dont_touch of G25510: signal is true;
	signal G25513: std_logic; attribute dont_touch of G25513: signal is true;
	signal G25514: std_logic; attribute dont_touch of G25514: signal is true;
	signal G25515: std_logic; attribute dont_touch of G25515: signal is true;
	signal G25518: std_logic; attribute dont_touch of G25518: signal is true;
	signal G25519: std_logic; attribute dont_touch of G25519: signal is true;
	signal G25520: std_logic; attribute dont_touch of G25520: signal is true;
	signal G25523: std_logic; attribute dont_touch of G25523: signal is true;
	signal G25524: std_logic; attribute dont_touch of G25524: signal is true;
	signal G25527: std_logic; attribute dont_touch of G25527: signal is true;
	signal G25530: std_logic; attribute dont_touch of G25530: signal is true;
	signal G25533: std_logic; attribute dont_touch of G25533: signal is true;
	signal G25536: std_logic; attribute dont_touch of G25536: signal is true;
	signal G25539: std_logic; attribute dont_touch of G25539: signal is true;
	signal G25540: std_logic; attribute dont_touch of G25540: signal is true;
	signal G25543: std_logic; attribute dont_touch of G25543: signal is true;
	signal G25546: std_logic; attribute dont_touch of G25546: signal is true;
	signal G25549: std_logic; attribute dont_touch of G25549: signal is true;
	signal G25552: std_logic; attribute dont_touch of G25552: signal is true;
	signal G25553: std_logic; attribute dont_touch of G25553: signal is true;
	signal G25554: std_logic; attribute dont_touch of G25554: signal is true;
	signal G25557: std_logic; attribute dont_touch of G25557: signal is true;
	signal G25560: std_logic; attribute dont_touch of G25560: signal is true;
	signal G25561: std_logic; attribute dont_touch of G25561: signal is true;
	signal G25562: std_logic; attribute dont_touch of G25562: signal is true;
	signal G25565: std_logic; attribute dont_touch of G25565: signal is true;
	signal G25566: std_logic; attribute dont_touch of G25566: signal is true;
	signal G25569: std_logic; attribute dont_touch of G25569: signal is true;
	signal G25573: std_logic; attribute dont_touch of G25573: signal is true;
	signal G25576: std_logic; attribute dont_touch of G25576: signal is true;
	signal G25579: std_logic; attribute dont_touch of G25579: signal is true;
	signal G25582: std_logic; attribute dont_touch of G25582: signal is true;
	signal G25585: std_logic; attribute dont_touch of G25585: signal is true;
	signal G25588: std_logic; attribute dont_touch of G25588: signal is true;
	signal G25589: std_logic; attribute dont_touch of G25589: signal is true;
	signal G25590: std_logic; attribute dont_touch of G25590: signal is true;
	signal G25593: std_logic; attribute dont_touch of G25593: signal is true;
	signal G25596: std_logic; attribute dont_touch of G25596: signal is true;
	signal G25599: std_logic; attribute dont_touch of G25599: signal is true;
	signal G25602: std_logic; attribute dont_touch of G25602: signal is true;
	signal G25605: std_logic; attribute dont_touch of G25605: signal is true;
	signal G25606: std_logic; attribute dont_touch of G25606: signal is true;
	signal G25609: std_logic; attribute dont_touch of G25609: signal is true;
	signal G25612: std_logic; attribute dont_touch of G25612: signal is true;
	signal G25615: std_logic; attribute dont_touch of G25615: signal is true;
	signal G25618: std_logic; attribute dont_touch of G25618: signal is true;
	signal G25619: std_logic; attribute dont_touch of G25619: signal is true;
	signal G25620: std_logic; attribute dont_touch of G25620: signal is true;
	signal G25623: std_logic; attribute dont_touch of G25623: signal is true;
	signal G25626: std_logic; attribute dont_touch of G25626: signal is true;
	signal G25627: std_logic; attribute dont_touch of G25627: signal is true;
	signal G25628: std_logic; attribute dont_touch of G25628: signal is true;
	signal G25629: std_logic; attribute dont_touch of G25629: signal is true;
	signal G25630: std_logic; attribute dont_touch of G25630: signal is true;
	signal G25631: std_logic; attribute dont_touch of G25631: signal is true;
	signal G25634: std_logic; attribute dont_touch of G25634: signal is true;
	signal G25637: std_logic; attribute dont_touch of G25637: signal is true;
	signal G25640: std_logic; attribute dont_touch of G25640: signal is true;
	signal G25643: std_logic; attribute dont_touch of G25643: signal is true;
	signal G25646: std_logic; attribute dont_touch of G25646: signal is true;
	signal G25647: std_logic; attribute dont_touch of G25647: signal is true;
	signal G25648: std_logic; attribute dont_touch of G25648: signal is true;
	signal G25652: std_logic; attribute dont_touch of G25652: signal is true;
	signal G25655: std_logic; attribute dont_touch of G25655: signal is true;
	signal G25658: std_logic; attribute dont_touch of G25658: signal is true;
	signal G25661: std_logic; attribute dont_touch of G25661: signal is true;
	signal G25664: std_logic; attribute dont_touch of G25664: signal is true;
	signal G25667: std_logic; attribute dont_touch of G25667: signal is true;
	signal G25668: std_logic; attribute dont_touch of G25668: signal is true;
	signal G25669: std_logic; attribute dont_touch of G25669: signal is true;
	signal G25672: std_logic; attribute dont_touch of G25672: signal is true;
	signal G25675: std_logic; attribute dont_touch of G25675: signal is true;
	signal G25678: std_logic; attribute dont_touch of G25678: signal is true;
	signal G25681: std_logic; attribute dont_touch of G25681: signal is true;
	signal G25684: std_logic; attribute dont_touch of G25684: signal is true;
	signal G25685: std_logic; attribute dont_touch of G25685: signal is true;
	signal G25688: std_logic; attribute dont_touch of G25688: signal is true;
	signal G25691: std_logic; attribute dont_touch of G25691: signal is true;
	signal G25694: std_logic; attribute dont_touch of G25694: signal is true;
	signal G25697: std_logic; attribute dont_touch of G25697: signal is true;
	signal G25698: std_logic; attribute dont_touch of G25698: signal is true;
	signal G25699: std_logic; attribute dont_touch of G25699: signal is true;
	signal G25700: std_logic; attribute dont_touch of G25700: signal is true;
	signal G25703: std_logic; attribute dont_touch of G25703: signal is true;
	signal G25706: std_logic; attribute dont_touch of G25706: signal is true;
	signal G25707: std_logic; attribute dont_touch of G25707: signal is true;
	signal G25708: std_logic; attribute dont_touch of G25708: signal is true;
	signal G25711: std_logic; attribute dont_touch of G25711: signal is true;
	signal G25714: std_logic; attribute dont_touch of G25714: signal is true;
	signal G25717: std_logic; attribute dont_touch of G25717: signal is true;
	signal G25720: std_logic; attribute dont_touch of G25720: signal is true;
	signal G25723: std_logic; attribute dont_touch of G25723: signal is true;
	signal G25724: std_logic; attribute dont_touch of G25724: signal is true;
	signal G25725: std_logic; attribute dont_touch of G25725: signal is true;
	signal G25729: std_logic; attribute dont_touch of G25729: signal is true;
	signal G25732: std_logic; attribute dont_touch of G25732: signal is true;
	signal G25735: std_logic; attribute dont_touch of G25735: signal is true;
	signal G25738: std_logic; attribute dont_touch of G25738: signal is true;
	signal G25741: std_logic; attribute dont_touch of G25741: signal is true;
	signal G25744: std_logic; attribute dont_touch of G25744: signal is true;
	signal G25745: std_logic; attribute dont_touch of G25745: signal is true;
	signal G25746: std_logic; attribute dont_touch of G25746: signal is true;
	signal G25749: std_logic; attribute dont_touch of G25749: signal is true;
	signal G25752: std_logic; attribute dont_touch of G25752: signal is true;
	signal G25755: std_logic; attribute dont_touch of G25755: signal is true;
	signal G25758: std_logic; attribute dont_touch of G25758: signal is true;
	signal G25761: std_logic; attribute dont_touch of G25761: signal is true;
	signal G25762: std_logic; attribute dont_touch of G25762: signal is true;
	signal G25763: std_logic; attribute dont_touch of G25763: signal is true;
	signal G25764: std_logic; attribute dont_touch of G25764: signal is true;
	signal G25767: std_logic; attribute dont_touch of G25767: signal is true;
	signal G25770: std_logic; attribute dont_touch of G25770: signal is true;
	signal G25771: std_logic; attribute dont_touch of G25771: signal is true;
	signal G25772: std_logic; attribute dont_touch of G25772: signal is true;
	signal G25773: std_logic; attribute dont_touch of G25773: signal is true;
	signal G25776: std_logic; attribute dont_touch of G25776: signal is true;
	signal G25779: std_logic; attribute dont_touch of G25779: signal is true;
	signal G25780: std_logic; attribute dont_touch of G25780: signal is true;
	signal G25781: std_logic; attribute dont_touch of G25781: signal is true;
	signal G25784: std_logic; attribute dont_touch of G25784: signal is true;
	signal G25787: std_logic; attribute dont_touch of G25787: signal is true;
	signal G25790: std_logic; attribute dont_touch of G25790: signal is true;
	signal G25793: std_logic; attribute dont_touch of G25793: signal is true;
	signal G25796: std_logic; attribute dont_touch of G25796: signal is true;
	signal G25797: std_logic; attribute dont_touch of G25797: signal is true;
	signal G25798: std_logic; attribute dont_touch of G25798: signal is true;
	signal G25802: std_logic; attribute dont_touch of G25802: signal is true;
	signal G25805: std_logic; attribute dont_touch of G25805: signal is true;
	signal G25808: std_logic; attribute dont_touch of G25808: signal is true;
	signal G25811: std_logic; attribute dont_touch of G25811: signal is true;
	signal G25814: std_logic; attribute dont_touch of G25814: signal is true;
	signal G25817: std_logic; attribute dont_touch of G25817: signal is true;
	signal G25818: std_logic; attribute dont_touch of G25818: signal is true;
	signal G25821: std_logic; attribute dont_touch of G25821: signal is true;
	signal G25824: std_logic; attribute dont_touch of G25824: signal is true;
	signal G25825: std_logic; attribute dont_touch of G25825: signal is true;
	signal G25826: std_logic; attribute dont_touch of G25826: signal is true;
	signal G25827: std_logic; attribute dont_touch of G25827: signal is true;
	signal G25830: std_logic; attribute dont_touch of G25830: signal is true;
	signal G25833: std_logic; attribute dont_touch of G25833: signal is true;
	signal G25834: std_logic; attribute dont_touch of G25834: signal is true;
	signal G25835: std_logic; attribute dont_touch of G25835: signal is true;
	signal G25838: std_logic; attribute dont_touch of G25838: signal is true;
	signal G25841: std_logic; attribute dont_touch of G25841: signal is true;
	signal G25844: std_logic; attribute dont_touch of G25844: signal is true;
	signal G25847: std_logic; attribute dont_touch of G25847: signal is true;
	signal G25850: std_logic; attribute dont_touch of G25850: signal is true;
	signal G25851: std_logic; attribute dont_touch of G25851: signal is true;
	signal G25852: std_logic; attribute dont_touch of G25852: signal is true;
	signal G25853: std_logic; attribute dont_touch of G25853: signal is true;
	signal G25856: std_logic; attribute dont_touch of G25856: signal is true;
	signal G25859: std_logic; attribute dont_touch of G25859: signal is true;
	signal G25860: std_logic; attribute dont_touch of G25860: signal is true;
	signal G25861: std_logic; attribute dont_touch of G25861: signal is true;
	signal G25862: std_logic; attribute dont_touch of G25862: signal is true;
	signal G25865: std_logic; attribute dont_touch of G25865: signal is true;
	signal G25868: std_logic; attribute dont_touch of G25868: signal is true;
	signal G25869: std_logic; attribute dont_touch of G25869: signal is true;
	signal G25870: std_logic; attribute dont_touch of G25870: signal is true;
	signal G25873: std_logic; attribute dont_touch of G25873: signal is true;
	signal G25874: std_logic; attribute dont_touch of G25874: signal is true;
	signal G25877: std_logic; attribute dont_touch of G25877: signal is true;
	signal G25880: std_logic; attribute dont_touch of G25880: signal is true;
	signal G25881: std_logic; attribute dont_touch of G25881: signal is true;
	signal G25882: std_logic; attribute dont_touch of G25882: signal is true;
	signal G25885: std_logic; attribute dont_touch of G25885: signal is true;
	signal G25886: std_logic; attribute dont_touch of G25886: signal is true;
	signal G25887: std_logic; attribute dont_touch of G25887: signal is true;
	signal G25890: std_logic; attribute dont_touch of G25890: signal is true;
	signal G25891: std_logic; attribute dont_touch of G25891: signal is true;
	signal G25892: std_logic; attribute dont_touch of G25892: signal is true;
	signal G25895: std_logic; attribute dont_touch of G25895: signal is true;
	signal G25899: std_logic; attribute dont_touch of G25899: signal is true;
	signal G25903: std_logic; attribute dont_touch of G25903: signal is true;
	signal G25907: std_logic; attribute dont_touch of G25907: signal is true;
	signal G25911: std_logic; attribute dont_touch of G25911: signal is true;
	signal G25915: std_logic; attribute dont_touch of G25915: signal is true;
	signal G25919: std_logic; attribute dont_touch of G25919: signal is true;
	signal G25923: std_logic; attribute dont_touch of G25923: signal is true;
	signal G25927: std_logic; attribute dont_touch of G25927: signal is true;
	signal G25928: std_logic; attribute dont_touch of G25928: signal is true;
	signal G25929: std_logic; attribute dont_touch of G25929: signal is true;
	signal G25930: std_logic; attribute dont_touch of G25930: signal is true;
	signal G25931: std_logic; attribute dont_touch of G25931: signal is true;
	signal G25932: std_logic; attribute dont_touch of G25932: signal is true;
	signal G25933: std_logic; attribute dont_touch of G25933: signal is true;
	signal G25934: std_logic; attribute dont_touch of G25934: signal is true;
	signal G25935: std_logic; attribute dont_touch of G25935: signal is true;
	signal G25936: std_logic; attribute dont_touch of G25936: signal is true;
	signal G25937: std_logic; attribute dont_touch of G25937: signal is true;
	signal G25938: std_logic; attribute dont_touch of G25938: signal is true;
	signal G25939: std_logic; attribute dont_touch of G25939: signal is true;
	signal G25940: std_logic; attribute dont_touch of G25940: signal is true;
	signal G25941: std_logic; attribute dont_touch of G25941: signal is true;
	signal G25942: std_logic; attribute dont_touch of G25942: signal is true;
	signal G25943: std_logic; attribute dont_touch of G25943: signal is true;
	signal G25944: std_logic; attribute dont_touch of G25944: signal is true;
	signal G25945: std_logic; attribute dont_touch of G25945: signal is true;
	signal G25946: std_logic; attribute dont_touch of G25946: signal is true;
	signal G25947: std_logic; attribute dont_touch of G25947: signal is true;
	signal G25948: std_logic; attribute dont_touch of G25948: signal is true;
	signal G25949: std_logic; attribute dont_touch of G25949: signal is true;
	signal G25950: std_logic; attribute dont_touch of G25950: signal is true;
	signal G25951: std_logic; attribute dont_touch of G25951: signal is true;
	signal G25952: std_logic; attribute dont_touch of G25952: signal is true;
	signal G25953: std_logic; attribute dont_touch of G25953: signal is true;
	signal G25954: std_logic; attribute dont_touch of G25954: signal is true;
	signal G25957: std_logic; attribute dont_touch of G25957: signal is true;
	signal G25958: std_logic; attribute dont_touch of G25958: signal is true;
	signal G25961: std_logic; attribute dont_touch of G25961: signal is true;
	signal G25962: std_logic; attribute dont_touch of G25962: signal is true;
	signal G25963: std_logic; attribute dont_touch of G25963: signal is true;
	signal G25964: std_logic; attribute dont_touch of G25964: signal is true;
	signal G25967: std_logic; attribute dont_touch of G25967: signal is true;
	signal G25968: std_logic; attribute dont_touch of G25968: signal is true;
	signal G25969: std_logic; attribute dont_touch of G25969: signal is true;
	signal G25972: std_logic; attribute dont_touch of G25972: signal is true;
	signal G25973: std_logic; attribute dont_touch of G25973: signal is true;
	signal G25974: std_logic; attribute dont_touch of G25974: signal is true;
	signal G25975: std_logic; attribute dont_touch of G25975: signal is true;
	signal G25976: std_logic; attribute dont_touch of G25976: signal is true;
	signal G25977: std_logic; attribute dont_touch of G25977: signal is true;
	signal G25978: std_logic; attribute dont_touch of G25978: signal is true;
	signal G25979: std_logic; attribute dont_touch of G25979: signal is true;
	signal G25980: std_logic; attribute dont_touch of G25980: signal is true;
	signal G25981: std_logic; attribute dont_touch of G25981: signal is true;
	signal G25982: std_logic; attribute dont_touch of G25982: signal is true;
	signal G25983: std_logic; attribute dont_touch of G25983: signal is true;
	signal G25984: std_logic; attribute dont_touch of G25984: signal is true;
	signal G25985: std_logic; attribute dont_touch of G25985: signal is true;
	signal G25986: std_logic; attribute dont_touch of G25986: signal is true;
	signal G25987: std_logic; attribute dont_touch of G25987: signal is true;
	signal G25988: std_logic; attribute dont_touch of G25988: signal is true;
	signal G25989: std_logic; attribute dont_touch of G25989: signal is true;
	signal G25990: std_logic; attribute dont_touch of G25990: signal is true;
	signal G25991: std_logic; attribute dont_touch of G25991: signal is true;
	signal G25992: std_logic; attribute dont_touch of G25992: signal is true;
	signal G25993: std_logic; attribute dont_touch of G25993: signal is true;
	signal G25994: std_logic; attribute dont_touch of G25994: signal is true;
	signal G25995: std_logic; attribute dont_touch of G25995: signal is true;
	signal G25996: std_logic; attribute dont_touch of G25996: signal is true;
	signal G25997: std_logic; attribute dont_touch of G25997: signal is true;
	signal G25998: std_logic; attribute dont_touch of G25998: signal is true;
	signal G25999: std_logic; attribute dont_touch of G25999: signal is true;
	signal G26000: std_logic; attribute dont_touch of G26000: signal is true;
	signal G26001: std_logic; attribute dont_touch of G26001: signal is true;
	signal G26002: std_logic; attribute dont_touch of G26002: signal is true;
	signal G26003: std_logic; attribute dont_touch of G26003: signal is true;
	signal G26004: std_logic; attribute dont_touch of G26004: signal is true;
	signal G26005: std_logic; attribute dont_touch of G26005: signal is true;
	signal G26006: std_logic; attribute dont_touch of G26006: signal is true;
	signal G26007: std_logic; attribute dont_touch of G26007: signal is true;
	signal G26008: std_logic; attribute dont_touch of G26008: signal is true;
	signal G26009: std_logic; attribute dont_touch of G26009: signal is true;
	signal G26010: std_logic; attribute dont_touch of G26010: signal is true;
	signal G26011: std_logic; attribute dont_touch of G26011: signal is true;
	signal G26012: std_logic; attribute dont_touch of G26012: signal is true;
	signal G26013: std_logic; attribute dont_touch of G26013: signal is true;
	signal G26014: std_logic; attribute dont_touch of G26014: signal is true;
	signal G26015: std_logic; attribute dont_touch of G26015: signal is true;
	signal G26016: std_logic; attribute dont_touch of G26016: signal is true;
	signal G26017: std_logic; attribute dont_touch of G26017: signal is true;
	signal G26018: std_logic; attribute dont_touch of G26018: signal is true;
	signal G26019: std_logic; attribute dont_touch of G26019: signal is true;
	signal G26020: std_logic; attribute dont_touch of G26020: signal is true;
	signal G26021: std_logic; attribute dont_touch of G26021: signal is true;
	signal G26022: std_logic; attribute dont_touch of G26022: signal is true;
	signal G26023: std_logic; attribute dont_touch of G26023: signal is true;
	signal G26024: std_logic; attribute dont_touch of G26024: signal is true;
	signal G26025: std_logic; attribute dont_touch of G26025: signal is true;
	signal G26026: std_logic; attribute dont_touch of G26026: signal is true;
	signal G26027: std_logic; attribute dont_touch of G26027: signal is true;
	signal G26028: std_logic; attribute dont_touch of G26028: signal is true;
	signal G26029: std_logic; attribute dont_touch of G26029: signal is true;
	signal G26030: std_logic; attribute dont_touch of G26030: signal is true;
	signal G26031: std_logic; attribute dont_touch of G26031: signal is true;
	signal G26032: std_logic; attribute dont_touch of G26032: signal is true;
	signal G26033: std_logic; attribute dont_touch of G26033: signal is true;
	signal G26034: std_logic; attribute dont_touch of G26034: signal is true;
	signal G26035: std_logic; attribute dont_touch of G26035: signal is true;
	signal G26036: std_logic; attribute dont_touch of G26036: signal is true;
	signal G26037: std_logic; attribute dont_touch of G26037: signal is true;
	signal G26038: std_logic; attribute dont_touch of G26038: signal is true;
	signal G26039: std_logic; attribute dont_touch of G26039: signal is true;
	signal G26040: std_logic; attribute dont_touch of G26040: signal is true;
	signal G26041: std_logic; attribute dont_touch of G26041: signal is true;
	signal G26042: std_logic; attribute dont_touch of G26042: signal is true;
	signal G26043: std_logic; attribute dont_touch of G26043: signal is true;
	signal G26044: std_logic; attribute dont_touch of G26044: signal is true;
	signal G26045: std_logic; attribute dont_touch of G26045: signal is true;
	signal G26046: std_logic; attribute dont_touch of G26046: signal is true;
	signal G26047: std_logic; attribute dont_touch of G26047: signal is true;
	signal G26048: std_logic; attribute dont_touch of G26048: signal is true;
	signal G26049: std_logic; attribute dont_touch of G26049: signal is true;
	signal G26050: std_logic; attribute dont_touch of G26050: signal is true;
	signal G26051: std_logic; attribute dont_touch of G26051: signal is true;
	signal G26052: std_logic; attribute dont_touch of G26052: signal is true;
	signal G26053: std_logic; attribute dont_touch of G26053: signal is true;
	signal G26054: std_logic; attribute dont_touch of G26054: signal is true;
	signal G26055: std_logic; attribute dont_touch of G26055: signal is true;
	signal G26056: std_logic; attribute dont_touch of G26056: signal is true;
	signal G26059: std_logic; attribute dont_touch of G26059: signal is true;
	signal G26060: std_logic; attribute dont_touch of G26060: signal is true;
	signal G26061: std_logic; attribute dont_touch of G26061: signal is true;
	signal G26062: std_logic; attribute dont_touch of G26062: signal is true;
	signal G26063: std_logic; attribute dont_touch of G26063: signal is true;
	signal G26066: std_logic; attribute dont_touch of G26066: signal is true;
	signal G26067: std_logic; attribute dont_touch of G26067: signal is true;
	signal G26068: std_logic; attribute dont_touch of G26068: signal is true;
	signal G26069: std_logic; attribute dont_touch of G26069: signal is true;
	signal G26070: std_logic; attribute dont_touch of G26070: signal is true;
	signal G26073: std_logic; attribute dont_touch of G26073: signal is true;
	signal G26074: std_logic; attribute dont_touch of G26074: signal is true;
	signal G26075: std_logic; attribute dont_touch of G26075: signal is true;
	signal G26076: std_logic; attribute dont_touch of G26076: signal is true;
	signal G26079: std_logic; attribute dont_touch of G26079: signal is true;
	signal G26080: std_logic; attribute dont_touch of G26080: signal is true;
	signal G26081: std_logic; attribute dont_touch of G26081: signal is true;
	signal G26082: std_logic; attribute dont_touch of G26082: signal is true;
	signal G26083: std_logic; attribute dont_touch of G26083: signal is true;
	signal G26084: std_logic; attribute dont_touch of G26084: signal is true;
	signal G26085: std_logic; attribute dont_touch of G26085: signal is true;
	signal G26086: std_logic; attribute dont_touch of G26086: signal is true;
	signal G26087: std_logic; attribute dont_touch of G26087: signal is true;
	signal G26090: std_logic; attribute dont_touch of G26090: signal is true;
	signal G26091: std_logic; attribute dont_touch of G26091: signal is true;
	signal G26092: std_logic; attribute dont_touch of G26092: signal is true;
	signal G26096: std_logic; attribute dont_touch of G26096: signal is true;
	signal G26099: std_logic; attribute dont_touch of G26099: signal is true;
	signal G26102: std_logic; attribute dont_touch of G26102: signal is true;
	signal G26103: std_logic; attribute dont_touch of G26103: signal is true;
	signal G26105: std_logic; attribute dont_touch of G26105: signal is true;
	signal G26106: std_logic; attribute dont_touch of G26106: signal is true;
	signal G26107: std_logic; attribute dont_touch of G26107: signal is true;
	signal G26110: std_logic; attribute dont_touch of G26110: signal is true;
	signal G26113: std_logic; attribute dont_touch of G26113: signal is true;
	signal G26114: std_logic; attribute dont_touch of G26114: signal is true;
	signal G26118: std_logic; attribute dont_touch of G26118: signal is true;
	signal G26119: std_logic; attribute dont_touch of G26119: signal is true;
	signal G26120: std_logic; attribute dont_touch of G26120: signal is true;
	signal G26121: std_logic; attribute dont_touch of G26121: signal is true;
	signal G26125: std_logic; attribute dont_touch of G26125: signal is true;
	signal G26126: std_logic; attribute dont_touch of G26126: signal is true;
	signal G26129: std_logic; attribute dont_touch of G26129: signal is true;
	signal G26130: std_logic; attribute dont_touch of G26130: signal is true;
	signal G26131: std_logic; attribute dont_touch of G26131: signal is true;
	signal G26136: std_logic; attribute dont_touch of G26136: signal is true;
	signal G26137: std_logic; attribute dont_touch of G26137: signal is true;
	signal G26140: std_logic; attribute dont_touch of G26140: signal is true;
	signal G26143: std_logic; attribute dont_touch of G26143: signal is true;
	signal G26144: std_logic; attribute dont_touch of G26144: signal is true;
	signal G26145: std_logic; attribute dont_touch of G26145: signal is true;
	signal G26148: std_logic; attribute dont_touch of G26148: signal is true;
	signal G26150: std_logic; attribute dont_touch of G26150: signal is true;
	signal G26151: std_logic; attribute dont_touch of G26151: signal is true;
	signal G26154: std_logic; attribute dont_touch of G26154: signal is true;
	signal G26157: std_logic; attribute dont_touch of G26157: signal is true;
	signal G26158: std_logic; attribute dont_touch of G26158: signal is true;
	signal G26159: std_logic; attribute dont_touch of G26159: signal is true;
	signal G26160: std_logic; attribute dont_touch of G26160: signal is true;
	signal G26163: std_logic; attribute dont_touch of G26163: signal is true;
	signal G26164: std_logic; attribute dont_touch of G26164: signal is true;
	signal G26165: std_logic; attribute dont_touch of G26165: signal is true;
	signal G26166: std_logic; attribute dont_touch of G26166: signal is true;
	signal G26167: std_logic; attribute dont_touch of G26167: signal is true;
	signal G26168: std_logic; attribute dont_touch of G26168: signal is true;
	signal G26171: std_logic; attribute dont_touch of G26171: signal is true;
	signal G26172: std_logic; attribute dont_touch of G26172: signal is true;
	signal G26173: std_logic; attribute dont_touch of G26173: signal is true;
	signal G26174: std_logic; attribute dont_touch of G26174: signal is true;
	signal G26175: std_logic; attribute dont_touch of G26175: signal is true;
	signal G26178: std_logic; attribute dont_touch of G26178: signal is true;
	signal G26181: std_logic; attribute dont_touch of G26181: signal is true;
	signal G26182: std_logic; attribute dont_touch of G26182: signal is true;
	signal G26183: std_logic; attribute dont_touch of G26183: signal is true;
	signal G26186: std_logic; attribute dont_touch of G26186: signal is true;
	signal G26187: std_logic; attribute dont_touch of G26187: signal is true;
	signal G26188: std_logic; attribute dont_touch of G26188: signal is true;
	signal G26189: std_logic; attribute dont_touch of G26189: signal is true;
	signal G26190: std_logic; attribute dont_touch of G26190: signal is true;
	signal G26191: std_logic; attribute dont_touch of G26191: signal is true;
	signal G26192: std_logic; attribute dont_touch of G26192: signal is true;
	signal G26193: std_logic; attribute dont_touch of G26193: signal is true;
	signal G26194: std_logic; attribute dont_touch of G26194: signal is true;
	signal G26195: std_logic; attribute dont_touch of G26195: signal is true;
	signal G26196: std_logic; attribute dont_touch of G26196: signal is true;
	signal G26199: std_logic; attribute dont_touch of G26199: signal is true;
	signal G26202: std_logic; attribute dont_touch of G26202: signal is true;
	signal G26205: std_logic; attribute dont_touch of G26205: signal is true;
	signal G26206: std_logic; attribute dont_touch of G26206: signal is true;
	signal G26207: std_logic; attribute dont_touch of G26207: signal is true;
	signal G26208: std_logic; attribute dont_touch of G26208: signal is true;
	signal G26209: std_logic; attribute dont_touch of G26209: signal is true;
	signal G26210: std_logic; attribute dont_touch of G26210: signal is true;
	signal G26211: std_logic; attribute dont_touch of G26211: signal is true;
	signal G26212: std_logic; attribute dont_touch of G26212: signal is true;
	signal G26213: std_logic; attribute dont_touch of G26213: signal is true;
	signal G26214: std_logic; attribute dont_touch of G26214: signal is true;
	signal G26215: std_logic; attribute dont_touch of G26215: signal is true;
	signal G26216: std_logic; attribute dont_touch of G26216: signal is true;
	signal G26217: std_logic; attribute dont_touch of G26217: signal is true;
	signal G26220: std_logic; attribute dont_touch of G26220: signal is true;
	signal G26221: std_logic; attribute dont_touch of G26221: signal is true;
	signal G26222: std_logic; attribute dont_touch of G26222: signal is true;
	signal G26223: std_logic; attribute dont_touch of G26223: signal is true;
	signal G26226: std_logic; attribute dont_touch of G26226: signal is true;
	signal G26229: std_logic; attribute dont_touch of G26229: signal is true;
	signal G26230: std_logic; attribute dont_touch of G26230: signal is true;
	signal G26231: std_logic; attribute dont_touch of G26231: signal is true;
	signal G26232: std_logic; attribute dont_touch of G26232: signal is true;
	signal G26233: std_logic; attribute dont_touch of G26233: signal is true;
	signal G26234: std_logic; attribute dont_touch of G26234: signal is true;
	signal G26235: std_logic; attribute dont_touch of G26235: signal is true;
	signal G26236: std_logic; attribute dont_touch of G26236: signal is true;
	signal G26237: std_logic; attribute dont_touch of G26237: signal is true;
	signal G26238: std_logic; attribute dont_touch of G26238: signal is true;
	signal G26239: std_logic; attribute dont_touch of G26239: signal is true;
	signal G26240: std_logic; attribute dont_touch of G26240: signal is true;
	signal G26243: std_logic; attribute dont_touch of G26243: signal is true;
	signal G26244: std_logic; attribute dont_touch of G26244: signal is true;
	signal G26245: std_logic; attribute dont_touch of G26245: signal is true;
	signal G26246: std_logic; attribute dont_touch of G26246: signal is true;
	signal G26247: std_logic; attribute dont_touch of G26247: signal is true;
	signal G26248: std_logic; attribute dont_touch of G26248: signal is true;
	signal G26249: std_logic; attribute dont_touch of G26249: signal is true;
	signal G26250: std_logic; attribute dont_touch of G26250: signal is true;
	signal G26251: std_logic; attribute dont_touch of G26251: signal is true;
	signal G26254: std_logic; attribute dont_touch of G26254: signal is true;
	signal G26257: std_logic; attribute dont_touch of G26257: signal is true;
	signal G26258: std_logic; attribute dont_touch of G26258: signal is true;
	signal G26259: std_logic; attribute dont_touch of G26259: signal is true;
	signal G26260: std_logic; attribute dont_touch of G26260: signal is true;
	signal G26261: std_logic; attribute dont_touch of G26261: signal is true;
	signal G26262: std_logic; attribute dont_touch of G26262: signal is true;
	signal G26263: std_logic; attribute dont_touch of G26263: signal is true;
	signal G26264: std_logic; attribute dont_touch of G26264: signal is true;
	signal G26265: std_logic; attribute dont_touch of G26265: signal is true;
	signal G26268: std_logic; attribute dont_touch of G26268: signal is true;
	signal G26269: std_logic; attribute dont_touch of G26269: signal is true;
	signal G26270: std_logic; attribute dont_touch of G26270: signal is true;
	signal G26271: std_logic; attribute dont_touch of G26271: signal is true;
	signal G26272: std_logic; attribute dont_touch of G26272: signal is true;
	signal G26275: std_logic; attribute dont_touch of G26275: signal is true;
	signal G26276: std_logic; attribute dont_touch of G26276: signal is true;
	signal G26277: std_logic; attribute dont_touch of G26277: signal is true;
	signal G26278: std_logic; attribute dont_touch of G26278: signal is true;
	signal G26279: std_logic; attribute dont_touch of G26279: signal is true;
	signal G26280: std_logic; attribute dont_touch of G26280: signal is true;
	signal G26281: std_logic; attribute dont_touch of G26281: signal is true;
	signal G26282: std_logic; attribute dont_touch of G26282: signal is true;
	signal G26283: std_logic; attribute dont_touch of G26283: signal is true;
	signal G26288: std_logic; attribute dont_touch of G26288: signal is true;
	signal G26289: std_logic; attribute dont_touch of G26289: signal is true;
	signal G26290: std_logic; attribute dont_touch of G26290: signal is true;
	signal G26291: std_logic; attribute dont_touch of G26291: signal is true;
	signal G26292: std_logic; attribute dont_touch of G26292: signal is true;
	signal G26293: std_logic; attribute dont_touch of G26293: signal is true;
	signal G26294: std_logic; attribute dont_touch of G26294: signal is true;
	signal G26295: std_logic; attribute dont_touch of G26295: signal is true;
	signal G26298: std_logic; attribute dont_touch of G26298: signal is true;
	signal G26299: std_logic; attribute dont_touch of G26299: signal is true;
	signal G26300: std_logic; attribute dont_touch of G26300: signal is true;
	signal G26301: std_logic; attribute dont_touch of G26301: signal is true;
	signal G26302: std_logic; attribute dont_touch of G26302: signal is true;
	signal G26303: std_logic; attribute dont_touch of G26303: signal is true;
	signal G26304: std_logic; attribute dont_touch of G26304: signal is true;
	signal G26307: std_logic; attribute dont_touch of G26307: signal is true;
	signal G26308: std_logic; attribute dont_touch of G26308: signal is true;
	signal G26309: std_logic; attribute dont_touch of G26309: signal is true;
	signal G26310: std_logic; attribute dont_touch of G26310: signal is true;
	signal G26311: std_logic; attribute dont_touch of G26311: signal is true;
	signal G26312: std_logic; attribute dont_touch of G26312: signal is true;
	signal G26313: std_logic; attribute dont_touch of G26313: signal is true;
	signal G26314: std_logic; attribute dont_touch of G26314: signal is true;
	signal G26315: std_logic; attribute dont_touch of G26315: signal is true;
	signal G26316: std_logic; attribute dont_touch of G26316: signal is true;
	signal G26317: std_logic; attribute dont_touch of G26317: signal is true;
	signal G26318: std_logic; attribute dont_touch of G26318: signal is true;
	signal G26319: std_logic; attribute dont_touch of G26319: signal is true;
	signal G26320: std_logic; attribute dont_touch of G26320: signal is true;
	signal G26324: std_logic; attribute dont_touch of G26324: signal is true;
	signal G26325: std_logic; attribute dont_touch of G26325: signal is true;
	signal G26326: std_logic; attribute dont_touch of G26326: signal is true;
	signal G26327: std_logic; attribute dont_touch of G26327: signal is true;
	signal G26332: std_logic; attribute dont_touch of G26332: signal is true;
	signal G26333: std_logic; attribute dont_touch of G26333: signal is true;
	signal G26334: std_logic; attribute dont_touch of G26334: signal is true;
	signal G26335: std_logic; attribute dont_touch of G26335: signal is true;
	signal G26336: std_logic; attribute dont_touch of G26336: signal is true;
	signal G26339: std_logic; attribute dont_touch of G26339: signal is true;
	signal G26340: std_logic; attribute dont_touch of G26340: signal is true;
	signal G26341: std_logic; attribute dont_touch of G26341: signal is true;
	signal G26342: std_logic; attribute dont_touch of G26342: signal is true;
	signal G26343: std_logic; attribute dont_touch of G26343: signal is true;
	signal G26344: std_logic; attribute dont_touch of G26344: signal is true;
	signal G26345: std_logic; attribute dont_touch of G26345: signal is true;
	signal G26346: std_logic; attribute dont_touch of G26346: signal is true;
	signal G26347: std_logic; attribute dont_touch of G26347: signal is true;
	signal G26348: std_logic; attribute dont_touch of G26348: signal is true;
	signal G26349: std_logic; attribute dont_touch of G26349: signal is true;
	signal G26350: std_logic; attribute dont_touch of G26350: signal is true;
	signal G26351: std_logic; attribute dont_touch of G26351: signal is true;
	signal G26352: std_logic; attribute dont_touch of G26352: signal is true;
	signal G26353: std_logic; attribute dont_touch of G26353: signal is true;
	signal G26354: std_logic; attribute dont_touch of G26354: signal is true;
	signal G26355: std_logic; attribute dont_touch of G26355: signal is true;
	signal G26356: std_logic; attribute dont_touch of G26356: signal is true;
	signal G26357: std_logic; attribute dont_touch of G26357: signal is true;
	signal G26358: std_logic; attribute dont_touch of G26358: signal is true;
	signal G26361: std_logic; attribute dont_touch of G26361: signal is true;
	signal G26362: std_logic; attribute dont_touch of G26362: signal is true;
	signal G26363: std_logic; attribute dont_touch of G26363: signal is true;
	signal G26364: std_logic; attribute dont_touch of G26364: signal is true;
	signal G26365: std_logic; attribute dont_touch of G26365: signal is true;
	signal G26366: std_logic; attribute dont_touch of G26366: signal is true;
	signal G26367: std_logic; attribute dont_touch of G26367: signal is true;
	signal G26371: std_logic; attribute dont_touch of G26371: signal is true;
	signal G26372: std_logic; attribute dont_touch of G26372: signal is true;
	signal G26373: std_logic; attribute dont_touch of G26373: signal is true;
	signal G26374: std_logic; attribute dont_touch of G26374: signal is true;
	signal G26379: std_logic; attribute dont_touch of G26379: signal is true;
	signal G26380: std_logic; attribute dont_touch of G26380: signal is true;
	signal G26381: std_logic; attribute dont_touch of G26381: signal is true;
	signal G26382: std_logic; attribute dont_touch of G26382: signal is true;
	signal G26383: std_logic; attribute dont_touch of G26383: signal is true;
	signal G26384: std_logic; attribute dont_touch of G26384: signal is true;
	signal G26385: std_logic; attribute dont_touch of G26385: signal is true;
	signal G26386: std_logic; attribute dont_touch of G26386: signal is true;
	signal G26387: std_logic; attribute dont_touch of G26387: signal is true;
	signal G26388: std_logic; attribute dont_touch of G26388: signal is true;
	signal G26389: std_logic; attribute dont_touch of G26389: signal is true;
	signal G26390: std_logic; attribute dont_touch of G26390: signal is true;
	signal G26391: std_logic; attribute dont_touch of G26391: signal is true;
	signal G26392: std_logic; attribute dont_touch of G26392: signal is true;
	signal G26393: std_logic; attribute dont_touch of G26393: signal is true;
	signal G26396: std_logic; attribute dont_touch of G26396: signal is true;
	signal G26397: std_logic; attribute dont_touch of G26397: signal is true;
	signal G26398: std_logic; attribute dont_touch of G26398: signal is true;
	signal G26399: std_logic; attribute dont_touch of G26399: signal is true;
	signal G26400: std_logic; attribute dont_touch of G26400: signal is true;
	signal G26401: std_logic; attribute dont_touch of G26401: signal is true;
	signal G26404: std_logic; attribute dont_touch of G26404: signal is true;
	signal G26405: std_logic; attribute dont_touch of G26405: signal is true;
	signal G26406: std_logic; attribute dont_touch of G26406: signal is true;
	signal G26407: std_logic; attribute dont_touch of G26407: signal is true;
	signal G26408: std_logic; attribute dont_touch of G26408: signal is true;
	signal G26409: std_logic; attribute dont_touch of G26409: signal is true;
	signal G26410: std_logic; attribute dont_touch of G26410: signal is true;
	signal G26414: std_logic; attribute dont_touch of G26414: signal is true;
	signal G26415: std_logic; attribute dont_touch of G26415: signal is true;
	signal G26416: std_logic; attribute dont_touch of G26416: signal is true;
	signal G26417: std_logic; attribute dont_touch of G26417: signal is true;
	signal G26422: std_logic; attribute dont_touch of G26422: signal is true;
	signal G26423: std_logic; attribute dont_touch of G26423: signal is true;
	signal G26424: std_logic; attribute dont_touch of G26424: signal is true;
	signal G26425: std_logic; attribute dont_touch of G26425: signal is true;
	signal G26426: std_logic; attribute dont_touch of G26426: signal is true;
	signal G26427: std_logic; attribute dont_touch of G26427: signal is true;
	signal G26428: std_logic; attribute dont_touch of G26428: signal is true;
	signal G26429: std_logic; attribute dont_touch of G26429: signal is true;
	signal G26432: std_logic; attribute dont_touch of G26432: signal is true;
	signal G26433: std_logic; attribute dont_touch of G26433: signal is true;
	signal G26434: std_logic; attribute dont_touch of G26434: signal is true;
	signal G26437: std_logic; attribute dont_touch of G26437: signal is true;
	signal G26438: std_logic; attribute dont_touch of G26438: signal is true;
	signal G26439: std_logic; attribute dont_touch of G26439: signal is true;
	signal G26440: std_logic; attribute dont_touch of G26440: signal is true;
	signal G26441: std_logic; attribute dont_touch of G26441: signal is true;
	signal G26442: std_logic; attribute dont_touch of G26442: signal is true;
	signal G26445: std_logic; attribute dont_touch of G26445: signal is true;
	signal G26446: std_logic; attribute dont_touch of G26446: signal is true;
	signal G26447: std_logic; attribute dont_touch of G26447: signal is true;
	signal G26448: std_logic; attribute dont_touch of G26448: signal is true;
	signal G26449: std_logic; attribute dont_touch of G26449: signal is true;
	signal G26450: std_logic; attribute dont_touch of G26450: signal is true;
	signal G26451: std_logic; attribute dont_touch of G26451: signal is true;
	signal G26455: std_logic; attribute dont_touch of G26455: signal is true;
	signal G26456: std_logic; attribute dont_touch of G26456: signal is true;
	signal G26457: std_logic; attribute dont_touch of G26457: signal is true;
	signal G26458: std_logic; attribute dont_touch of G26458: signal is true;
	signal G26461: std_logic; attribute dont_touch of G26461: signal is true;
	signal G26464: std_logic; attribute dont_touch of G26464: signal is true;
	signal G26465: std_logic; attribute dont_touch of G26465: signal is true;
	signal G26466: std_logic; attribute dont_touch of G26466: signal is true;
	signal G26469: std_logic; attribute dont_touch of G26469: signal is true;
	signal G26470: std_logic; attribute dont_touch of G26470: signal is true;
	signal G26471: std_logic; attribute dont_touch of G26471: signal is true;
	signal G26472: std_logic; attribute dont_touch of G26472: signal is true;
	signal G26473: std_logic; attribute dont_touch of G26473: signal is true;
	signal G26474: std_logic; attribute dont_touch of G26474: signal is true;
	signal G26477: std_logic; attribute dont_touch of G26477: signal is true;
	signal G26478: std_logic; attribute dont_touch of G26478: signal is true;
	signal G26479: std_logic; attribute dont_touch of G26479: signal is true;
	signal G26480: std_logic; attribute dont_touch of G26480: signal is true;
	signal G26481: std_logic; attribute dont_touch of G26481: signal is true;
	signal G26482: std_logic; attribute dont_touch of G26482: signal is true;
	signal G26485: std_logic; attribute dont_touch of G26485: signal is true;
	signal G26488: std_logic; attribute dont_touch of G26488: signal is true;
	signal G26489: std_logic; attribute dont_touch of G26489: signal is true;
	signal G26490: std_logic; attribute dont_touch of G26490: signal is true;
	signal G26493: std_logic; attribute dont_touch of G26493: signal is true;
	signal G26494: std_logic; attribute dont_touch of G26494: signal is true;
	signal G26495: std_logic; attribute dont_touch of G26495: signal is true;
	signal G26496: std_logic; attribute dont_touch of G26496: signal is true;
	signal G26497: std_logic; attribute dont_touch of G26497: signal is true;
	signal G26498: std_logic; attribute dont_touch of G26498: signal is true;
	signal G26501: std_logic; attribute dont_touch of G26501: signal is true;
	signal G26504: std_logic; attribute dont_touch of G26504: signal is true;
	signal G26505: std_logic; attribute dont_touch of G26505: signal is true;
	signal G26506: std_logic; attribute dont_touch of G26506: signal is true;
	signal G26507: std_logic; attribute dont_touch of G26507: signal is true;
	signal G26508: std_logic; attribute dont_touch of G26508: signal is true;
	signal G26512: std_logic; attribute dont_touch of G26512: signal is true;
	signal G26513: std_logic; attribute dont_touch of G26513: signal is true;
	signal G26516: std_logic; attribute dont_touch of G26516: signal is true;
	signal G26520: std_logic; attribute dont_touch of G26520: signal is true;
	signal G26521: std_logic; attribute dont_touch of G26521: signal is true;
	signal G26525: std_logic; attribute dont_touch of G26525: signal is true;
	signal G26529: std_logic; attribute dont_touch of G26529: signal is true;
	signal G26530: std_logic; attribute dont_touch of G26530: signal is true;
	signal G26531: std_logic; attribute dont_touch of G26531: signal is true;
	signal G26532: std_logic; attribute dont_touch of G26532: signal is true;
	signal G26533: std_logic; attribute dont_touch of G26533: signal is true;
	signal G26534: std_logic; attribute dont_touch of G26534: signal is true;
	signal G26538: std_logic; attribute dont_touch of G26538: signal is true;
	signal G26539: std_logic; attribute dont_touch of G26539: signal is true;
	signal G26540: std_logic; attribute dont_touch of G26540: signal is true;
	signal G26541: std_logic; attribute dont_touch of G26541: signal is true;
	signal G26542: std_logic; attribute dont_touch of G26542: signal is true;
	signal G26543: std_logic; attribute dont_touch of G26543: signal is true;
	signal G26544: std_logic; attribute dont_touch of G26544: signal is true;
	signal G26545: std_logic; attribute dont_touch of G26545: signal is true;
	signal G26546: std_logic; attribute dont_touch of G26546: signal is true;
	signal G26547: std_logic; attribute dont_touch of G26547: signal is true;
	signal G26548: std_logic; attribute dont_touch of G26548: signal is true;
	signal G26549: std_logic; attribute dont_touch of G26549: signal is true;
	signal G26550: std_logic; attribute dont_touch of G26550: signal is true;
	signal G26551: std_logic; attribute dont_touch of G26551: signal is true;
	signal G26552: std_logic; attribute dont_touch of G26552: signal is true;
	signal G26553: std_logic; attribute dont_touch of G26553: signal is true;
	signal G26554: std_logic; attribute dont_touch of G26554: signal is true;
	signal G26555: std_logic; attribute dont_touch of G26555: signal is true;
	signal G26556: std_logic; attribute dont_touch of G26556: signal is true;
	signal G26557: std_logic; attribute dont_touch of G26557: signal is true;
	signal G26558: std_logic; attribute dont_touch of G26558: signal is true;
	signal G26559: std_logic; attribute dont_touch of G26559: signal is true;
	signal G26560: std_logic; attribute dont_touch of G26560: signal is true;
	signal G26561: std_logic; attribute dont_touch of G26561: signal is true;
	signal G26562: std_logic; attribute dont_touch of G26562: signal is true;
	signal G26563: std_logic; attribute dont_touch of G26563: signal is true;
	signal G26564: std_logic; attribute dont_touch of G26564: signal is true;
	signal G26565: std_logic; attribute dont_touch of G26565: signal is true;
	signal G26566: std_logic; attribute dont_touch of G26566: signal is true;
	signal G26567: std_logic; attribute dont_touch of G26567: signal is true;
	signal G26568: std_logic; attribute dont_touch of G26568: signal is true;
	signal G26569: std_logic; attribute dont_touch of G26569: signal is true;
	signal G26570: std_logic; attribute dont_touch of G26570: signal is true;
	signal G26571: std_logic; attribute dont_touch of G26571: signal is true;
	signal G26572: std_logic; attribute dont_touch of G26572: signal is true;
	signal G26573: std_logic; attribute dont_touch of G26573: signal is true;
	signal G26574: std_logic; attribute dont_touch of G26574: signal is true;
	signal G26575: std_logic; attribute dont_touch of G26575: signal is true;
	signal G26576: std_logic; attribute dont_touch of G26576: signal is true;
	signal G26577: std_logic; attribute dont_touch of G26577: signal is true;
	signal G26578: std_logic; attribute dont_touch of G26578: signal is true;
	signal G26579: std_logic; attribute dont_touch of G26579: signal is true;
	signal G26580: std_logic; attribute dont_touch of G26580: signal is true;
	signal G26581: std_logic; attribute dont_touch of G26581: signal is true;
	signal G26582: std_logic; attribute dont_touch of G26582: signal is true;
	signal G26583: std_logic; attribute dont_touch of G26583: signal is true;
	signal G26584: std_logic; attribute dont_touch of G26584: signal is true;
	signal G26585: std_logic; attribute dont_touch of G26585: signal is true;
	signal G26586: std_logic; attribute dont_touch of G26586: signal is true;
	signal G26587: std_logic; attribute dont_touch of G26587: signal is true;
	signal G26588: std_logic; attribute dont_touch of G26588: signal is true;
	signal G26589: std_logic; attribute dont_touch of G26589: signal is true;
	signal G26590: std_logic; attribute dont_touch of G26590: signal is true;
	signal G26591: std_logic; attribute dont_touch of G26591: signal is true;
	signal G26592: std_logic; attribute dont_touch of G26592: signal is true;
	signal G26593: std_logic; attribute dont_touch of G26593: signal is true;
	signal G26594: std_logic; attribute dont_touch of G26594: signal is true;
	signal G26595: std_logic; attribute dont_touch of G26595: signal is true;
	signal G26596: std_logic; attribute dont_touch of G26596: signal is true;
	signal G26597: std_logic; attribute dont_touch of G26597: signal is true;
	signal G26598: std_logic; attribute dont_touch of G26598: signal is true;
	signal G26599: std_logic; attribute dont_touch of G26599: signal is true;
	signal G26600: std_logic; attribute dont_touch of G26600: signal is true;
	signal G26601: std_logic; attribute dont_touch of G26601: signal is true;
	signal G26602: std_logic; attribute dont_touch of G26602: signal is true;
	signal G26603: std_logic; attribute dont_touch of G26603: signal is true;
	signal G26604: std_logic; attribute dont_touch of G26604: signal is true;
	signal G26605: std_logic; attribute dont_touch of G26605: signal is true;
	signal G26606: std_logic; attribute dont_touch of G26606: signal is true;
	signal G26607: std_logic; attribute dont_touch of G26607: signal is true;
	signal G26608: std_logic; attribute dont_touch of G26608: signal is true;
	signal G26609: std_logic; attribute dont_touch of G26609: signal is true;
	signal G26610: std_logic; attribute dont_touch of G26610: signal is true;
	signal G26611: std_logic; attribute dont_touch of G26611: signal is true;
	signal G26612: std_logic; attribute dont_touch of G26612: signal is true;
	signal G26613: std_logic; attribute dont_touch of G26613: signal is true;
	signal G26614: std_logic; attribute dont_touch of G26614: signal is true;
	signal G26615: std_logic; attribute dont_touch of G26615: signal is true;
	signal G26616: std_logic; attribute dont_touch of G26616: signal is true;
	signal G26617: std_logic; attribute dont_touch of G26617: signal is true;
	signal G26618: std_logic; attribute dont_touch of G26618: signal is true;
	signal G26619: std_logic; attribute dont_touch of G26619: signal is true;
	signal G26620: std_logic; attribute dont_touch of G26620: signal is true;
	signal G26621: std_logic; attribute dont_touch of G26621: signal is true;
	signal G26622: std_logic; attribute dont_touch of G26622: signal is true;
	signal G26623: std_logic; attribute dont_touch of G26623: signal is true;
	signal G26624: std_logic; attribute dont_touch of G26624: signal is true;
	signal G26625: std_logic; attribute dont_touch of G26625: signal is true;
	signal G26626: std_logic; attribute dont_touch of G26626: signal is true;
	signal G26627: std_logic; attribute dont_touch of G26627: signal is true;
	signal G26628: std_logic; attribute dont_touch of G26628: signal is true;
	signal G26629: std_logic; attribute dont_touch of G26629: signal is true;
	signal G26630: std_logic; attribute dont_touch of G26630: signal is true;
	signal G26631: std_logic; attribute dont_touch of G26631: signal is true;
	signal G26632: std_logic; attribute dont_touch of G26632: signal is true;
	signal G26633: std_logic; attribute dont_touch of G26633: signal is true;
	signal G26634: std_logic; attribute dont_touch of G26634: signal is true;
	signal G26635: std_logic; attribute dont_touch of G26635: signal is true;
	signal G26636: std_logic; attribute dont_touch of G26636: signal is true;
	signal G26637: std_logic; attribute dont_touch of G26637: signal is true;
	signal G26638: std_logic; attribute dont_touch of G26638: signal is true;
	signal G26639: std_logic; attribute dont_touch of G26639: signal is true;
	signal G26640: std_logic; attribute dont_touch of G26640: signal is true;
	signal G26641: std_logic; attribute dont_touch of G26641: signal is true;
	signal G26642: std_logic; attribute dont_touch of G26642: signal is true;
	signal G26643: std_logic; attribute dont_touch of G26643: signal is true;
	signal G26644: std_logic; attribute dont_touch of G26644: signal is true;
	signal G26645: std_logic; attribute dont_touch of G26645: signal is true;
	signal G26646: std_logic; attribute dont_touch of G26646: signal is true;
	signal G26647: std_logic; attribute dont_touch of G26647: signal is true;
	signal G26648: std_logic; attribute dont_touch of G26648: signal is true;
	signal G26649: std_logic; attribute dont_touch of G26649: signal is true;
	signal G26650: std_logic; attribute dont_touch of G26650: signal is true;
	signal G26651: std_logic; attribute dont_touch of G26651: signal is true;
	signal G26652: std_logic; attribute dont_touch of G26652: signal is true;
	signal G26653: std_logic; attribute dont_touch of G26653: signal is true;
	signal G26654: std_logic; attribute dont_touch of G26654: signal is true;
	signal G26655: std_logic; attribute dont_touch of G26655: signal is true;
	signal G26656: std_logic; attribute dont_touch of G26656: signal is true;
	signal G26657: std_logic; attribute dont_touch of G26657: signal is true;
	signal G26658: std_logic; attribute dont_touch of G26658: signal is true;
	signal G26659: std_logic; attribute dont_touch of G26659: signal is true;
	signal G26660: std_logic; attribute dont_touch of G26660: signal is true;
	signal G26661: std_logic; attribute dont_touch of G26661: signal is true;
	signal G26662: std_logic; attribute dont_touch of G26662: signal is true;
	signal G26663: std_logic; attribute dont_touch of G26663: signal is true;
	signal G26664: std_logic; attribute dont_touch of G26664: signal is true;
	signal G26665: std_logic; attribute dont_touch of G26665: signal is true;
	signal G26666: std_logic; attribute dont_touch of G26666: signal is true;
	signal G26667: std_logic; attribute dont_touch of G26667: signal is true;
	signal G26668: std_logic; attribute dont_touch of G26668: signal is true;
	signal G26669: std_logic; attribute dont_touch of G26669: signal is true;
	signal G26670: std_logic; attribute dont_touch of G26670: signal is true;
	signal G26671: std_logic; attribute dont_touch of G26671: signal is true;
	signal G26672: std_logic; attribute dont_touch of G26672: signal is true;
	signal G26673: std_logic; attribute dont_touch of G26673: signal is true;
	signal G26674: std_logic; attribute dont_touch of G26674: signal is true;
	signal G26675: std_logic; attribute dont_touch of G26675: signal is true;
	signal G26676: std_logic; attribute dont_touch of G26676: signal is true;
	signal G26677: std_logic; attribute dont_touch of G26677: signal is true;
	signal G26678: std_logic; attribute dont_touch of G26678: signal is true;
	signal G26679: std_logic; attribute dont_touch of G26679: signal is true;
	signal G26680: std_logic; attribute dont_touch of G26680: signal is true;
	signal G26681: std_logic; attribute dont_touch of G26681: signal is true;
	signal G26682: std_logic; attribute dont_touch of G26682: signal is true;
	signal G26683: std_logic; attribute dont_touch of G26683: signal is true;
	signal G26684: std_logic; attribute dont_touch of G26684: signal is true;
	signal G26685: std_logic; attribute dont_touch of G26685: signal is true;
	signal G26686: std_logic; attribute dont_touch of G26686: signal is true;
	signal G26687: std_logic; attribute dont_touch of G26687: signal is true;
	signal G26688: std_logic; attribute dont_touch of G26688: signal is true;
	signal G26689: std_logic; attribute dont_touch of G26689: signal is true;
	signal G26690: std_logic; attribute dont_touch of G26690: signal is true;
	signal G26691: std_logic; attribute dont_touch of G26691: signal is true;
	signal G26692: std_logic; attribute dont_touch of G26692: signal is true;
	signal G26693: std_logic; attribute dont_touch of G26693: signal is true;
	signal G26694: std_logic; attribute dont_touch of G26694: signal is true;
	signal G26695: std_logic; attribute dont_touch of G26695: signal is true;
	signal G26696: std_logic; attribute dont_touch of G26696: signal is true;
	signal G26697: std_logic; attribute dont_touch of G26697: signal is true;
	signal G26698: std_logic; attribute dont_touch of G26698: signal is true;
	signal G26699: std_logic; attribute dont_touch of G26699: signal is true;
	signal G26700: std_logic; attribute dont_touch of G26700: signal is true;
	signal G26701: std_logic; attribute dont_touch of G26701: signal is true;
	signal G26702: std_logic; attribute dont_touch of G26702: signal is true;
	signal G26703: std_logic; attribute dont_touch of G26703: signal is true;
	signal G26704: std_logic; attribute dont_touch of G26704: signal is true;
	signal G26705: std_logic; attribute dont_touch of G26705: signal is true;
	signal G26706: std_logic; attribute dont_touch of G26706: signal is true;
	signal G26707: std_logic; attribute dont_touch of G26707: signal is true;
	signal G26708: std_logic; attribute dont_touch of G26708: signal is true;
	signal G26709: std_logic; attribute dont_touch of G26709: signal is true;
	signal G26710: std_logic; attribute dont_touch of G26710: signal is true;
	signal G26711: std_logic; attribute dont_touch of G26711: signal is true;
	signal G26712: std_logic; attribute dont_touch of G26712: signal is true;
	signal G26713: std_logic; attribute dont_touch of G26713: signal is true;
	signal G26714: std_logic; attribute dont_touch of G26714: signal is true;
	signal G26715: std_logic; attribute dont_touch of G26715: signal is true;
	signal G26716: std_logic; attribute dont_touch of G26716: signal is true;
	signal G26717: std_logic; attribute dont_touch of G26717: signal is true;
	signal G26718: std_logic; attribute dont_touch of G26718: signal is true;
	signal G26719: std_logic; attribute dont_touch of G26719: signal is true;
	signal G26720: std_logic; attribute dont_touch of G26720: signal is true;
	signal G26721: std_logic; attribute dont_touch of G26721: signal is true;
	signal G26722: std_logic; attribute dont_touch of G26722: signal is true;
	signal G26723: std_logic; attribute dont_touch of G26723: signal is true;
	signal G26724: std_logic; attribute dont_touch of G26724: signal is true;
	signal G26725: std_logic; attribute dont_touch of G26725: signal is true;
	signal G26726: std_logic; attribute dont_touch of G26726: signal is true;
	signal G26727: std_logic; attribute dont_touch of G26727: signal is true;
	signal G26728: std_logic; attribute dont_touch of G26728: signal is true;
	signal G26729: std_logic; attribute dont_touch of G26729: signal is true;
	signal G26730: std_logic; attribute dont_touch of G26730: signal is true;
	signal G26731: std_logic; attribute dont_touch of G26731: signal is true;
	signal G26732: std_logic; attribute dont_touch of G26732: signal is true;
	signal G26733: std_logic; attribute dont_touch of G26733: signal is true;
	signal G26734: std_logic; attribute dont_touch of G26734: signal is true;
	signal G26735: std_logic; attribute dont_touch of G26735: signal is true;
	signal G26736: std_logic; attribute dont_touch of G26736: signal is true;
	signal G26737: std_logic; attribute dont_touch of G26737: signal is true;
	signal G26738: std_logic; attribute dont_touch of G26738: signal is true;
	signal G26739: std_logic; attribute dont_touch of G26739: signal is true;
	signal G26740: std_logic; attribute dont_touch of G26740: signal is true;
	signal G26741: std_logic; attribute dont_touch of G26741: signal is true;
	signal G26742: std_logic; attribute dont_touch of G26742: signal is true;
	signal G26743: std_logic; attribute dont_touch of G26743: signal is true;
	signal G26744: std_logic; attribute dont_touch of G26744: signal is true;
	signal G26745: std_logic; attribute dont_touch of G26745: signal is true;
	signal G26746: std_logic; attribute dont_touch of G26746: signal is true;
	signal G26747: std_logic; attribute dont_touch of G26747: signal is true;
	signal G26748: std_logic; attribute dont_touch of G26748: signal is true;
	signal G26749: std_logic; attribute dont_touch of G26749: signal is true;
	signal G26750: std_logic; attribute dont_touch of G26750: signal is true;
	signal G26751: std_logic; attribute dont_touch of G26751: signal is true;
	signal G26752: std_logic; attribute dont_touch of G26752: signal is true;
	signal G26753: std_logic; attribute dont_touch of G26753: signal is true;
	signal G26754: std_logic; attribute dont_touch of G26754: signal is true;
	signal G26755: std_logic; attribute dont_touch of G26755: signal is true;
	signal G26756: std_logic; attribute dont_touch of G26756: signal is true;
	signal G26757: std_logic; attribute dont_touch of G26757: signal is true;
	signal G26758: std_logic; attribute dont_touch of G26758: signal is true;
	signal G26759: std_logic; attribute dont_touch of G26759: signal is true;
	signal G26760: std_logic; attribute dont_touch of G26760: signal is true;
	signal G26761: std_logic; attribute dont_touch of G26761: signal is true;
	signal G26762: std_logic; attribute dont_touch of G26762: signal is true;
	signal G26763: std_logic; attribute dont_touch of G26763: signal is true;
	signal G26764: std_logic; attribute dont_touch of G26764: signal is true;
	signal G26765: std_logic; attribute dont_touch of G26765: signal is true;
	signal G26766: std_logic; attribute dont_touch of G26766: signal is true;
	signal G26767: std_logic; attribute dont_touch of G26767: signal is true;
	signal G26768: std_logic; attribute dont_touch of G26768: signal is true;
	signal G26769: std_logic; attribute dont_touch of G26769: signal is true;
	signal G26770: std_logic; attribute dont_touch of G26770: signal is true;
	signal G26771: std_logic; attribute dont_touch of G26771: signal is true;
	signal G26772: std_logic; attribute dont_touch of G26772: signal is true;
	signal G26773: std_logic; attribute dont_touch of G26773: signal is true;
	signal G26774: std_logic; attribute dont_touch of G26774: signal is true;
	signal G26775: std_logic; attribute dont_touch of G26775: signal is true;
	signal G26776: std_logic; attribute dont_touch of G26776: signal is true;
	signal G26777: std_logic; attribute dont_touch of G26777: signal is true;
	signal G26778: std_logic; attribute dont_touch of G26778: signal is true;
	signal G26779: std_logic; attribute dont_touch of G26779: signal is true;
	signal G26780: std_logic; attribute dont_touch of G26780: signal is true;
	signal G26781: std_logic; attribute dont_touch of G26781: signal is true;
	signal G26782: std_logic; attribute dont_touch of G26782: signal is true;
	signal G26783: std_logic; attribute dont_touch of G26783: signal is true;
	signal G26784: std_logic; attribute dont_touch of G26784: signal is true;
	signal G26785: std_logic; attribute dont_touch of G26785: signal is true;
	signal G26786: std_logic; attribute dont_touch of G26786: signal is true;
	signal G26787: std_logic; attribute dont_touch of G26787: signal is true;
	signal G26788: std_logic; attribute dont_touch of G26788: signal is true;
	signal G26789: std_logic; attribute dont_touch of G26789: signal is true;
	signal G26790: std_logic; attribute dont_touch of G26790: signal is true;
	signal G26791: std_logic; attribute dont_touch of G26791: signal is true;
	signal G26792: std_logic; attribute dont_touch of G26792: signal is true;
	signal G26793: std_logic; attribute dont_touch of G26793: signal is true;
	signal G26794: std_logic; attribute dont_touch of G26794: signal is true;
	signal G26795: std_logic; attribute dont_touch of G26795: signal is true;
	signal G26796: std_logic; attribute dont_touch of G26796: signal is true;
	signal G26797: std_logic; attribute dont_touch of G26797: signal is true;
	signal G26798: std_logic; attribute dont_touch of G26798: signal is true;
	signal G26799: std_logic; attribute dont_touch of G26799: signal is true;
	signal G26800: std_logic; attribute dont_touch of G26800: signal is true;
	signal G26801: std_logic; attribute dont_touch of G26801: signal is true;
	signal G26802: std_logic; attribute dont_touch of G26802: signal is true;
	signal G26803: std_logic; attribute dont_touch of G26803: signal is true;
	signal G26804: std_logic; attribute dont_touch of G26804: signal is true;
	signal G26805: std_logic; attribute dont_touch of G26805: signal is true;
	signal G26806: std_logic; attribute dont_touch of G26806: signal is true;
	signal G26807: std_logic; attribute dont_touch of G26807: signal is true;
	signal G26808: std_logic; attribute dont_touch of G26808: signal is true;
	signal G26809: std_logic; attribute dont_touch of G26809: signal is true;
	signal G26810: std_logic; attribute dont_touch of G26810: signal is true;
	signal G26811: std_logic; attribute dont_touch of G26811: signal is true;
	signal G26812: std_logic; attribute dont_touch of G26812: signal is true;
	signal G26813: std_logic; attribute dont_touch of G26813: signal is true;
	signal G26814: std_logic; attribute dont_touch of G26814: signal is true;
	signal G26815: std_logic; attribute dont_touch of G26815: signal is true;
	signal G26816: std_logic; attribute dont_touch of G26816: signal is true;
	signal G26817: std_logic; attribute dont_touch of G26817: signal is true;
	signal G26818: std_logic; attribute dont_touch of G26818: signal is true;
	signal G26819: std_logic; attribute dont_touch of G26819: signal is true;
	signal G26820: std_logic; attribute dont_touch of G26820: signal is true;
	signal G26821: std_logic; attribute dont_touch of G26821: signal is true;
	signal G26822: std_logic; attribute dont_touch of G26822: signal is true;
	signal G26823: std_logic; attribute dont_touch of G26823: signal is true;
	signal G26824: std_logic; attribute dont_touch of G26824: signal is true;
	signal G26825: std_logic; attribute dont_touch of G26825: signal is true;
	signal G26826: std_logic; attribute dont_touch of G26826: signal is true;
	signal G26827: std_logic; attribute dont_touch of G26827: signal is true;
	signal G26828: std_logic; attribute dont_touch of G26828: signal is true;
	signal G26829: std_logic; attribute dont_touch of G26829: signal is true;
	signal G26830: std_logic; attribute dont_touch of G26830: signal is true;
	signal G26831: std_logic; attribute dont_touch of G26831: signal is true;
	signal G26832: std_logic; attribute dont_touch of G26832: signal is true;
	signal G26833: std_logic; attribute dont_touch of G26833: signal is true;
	signal G26834: std_logic; attribute dont_touch of G26834: signal is true;
	signal G26835: std_logic; attribute dont_touch of G26835: signal is true;
	signal G26836: std_logic; attribute dont_touch of G26836: signal is true;
	signal G26837: std_logic; attribute dont_touch of G26837: signal is true;
	signal G26840: std_logic; attribute dont_touch of G26840: signal is true;
	signal G26841: std_logic; attribute dont_touch of G26841: signal is true;
	signal G26842: std_logic; attribute dont_touch of G26842: signal is true;
	signal G26843: std_logic; attribute dont_touch of G26843: signal is true;
	signal G26844: std_logic; attribute dont_touch of G26844: signal is true;
	signal G26845: std_logic; attribute dont_touch of G26845: signal is true;
	signal G26846: std_logic; attribute dont_touch of G26846: signal is true;
	signal G26849: std_logic; attribute dont_touch of G26849: signal is true;
	signal G26850: std_logic; attribute dont_touch of G26850: signal is true;
	signal G26851: std_logic; attribute dont_touch of G26851: signal is true;
	signal G26852: std_logic; attribute dont_touch of G26852: signal is true;
	signal G26853: std_logic; attribute dont_touch of G26853: signal is true;
	signal G26854: std_logic; attribute dont_touch of G26854: signal is true;
	signal G26855: std_logic; attribute dont_touch of G26855: signal is true;
	signal G26858: std_logic; attribute dont_touch of G26858: signal is true;
	signal G26859: std_logic; attribute dont_touch of G26859: signal is true;
	signal G26860: std_logic; attribute dont_touch of G26860: signal is true;
	signal G26861: std_logic; attribute dont_touch of G26861: signal is true;
	signal G26864: std_logic; attribute dont_touch of G26864: signal is true;
	signal G26865: std_logic; attribute dont_touch of G26865: signal is true;
	signal G26866: std_logic; attribute dont_touch of G26866: signal is true;
	signal G26867: std_logic; attribute dont_touch of G26867: signal is true;
	signal G26868: std_logic; attribute dont_touch of G26868: signal is true;
	signal G26869: std_logic; attribute dont_touch of G26869: signal is true;
	signal G26872: std_logic; attribute dont_touch of G26872: signal is true;
	signal G26873: std_logic; attribute dont_touch of G26873: signal is true;
	signal G26874: std_logic; attribute dont_touch of G26874: signal is true;
	signal G26875: std_logic; attribute dont_touch of G26875: signal is true;
	signal G26876: std_logic; attribute dont_touch of G26876: signal is true;
	signal G26877: std_logic; attribute dont_touch of G26877: signal is true;
	signal G26878: std_logic; attribute dont_touch of G26878: signal is true;
	signal G26881: std_logic; attribute dont_touch of G26881: signal is true;
	signal G26882: std_logic; attribute dont_touch of G26882: signal is true;
	signal G26883: std_logic; attribute dont_touch of G26883: signal is true;
	signal G26884: std_logic; attribute dont_touch of G26884: signal is true;
	signal G26885: std_logic; attribute dont_touch of G26885: signal is true;
	signal G26886: std_logic; attribute dont_touch of G26886: signal is true;
	signal G26887: std_logic; attribute dont_touch of G26887: signal is true;
	signal G26890: std_logic; attribute dont_touch of G26890: signal is true;
	signal G26891: std_logic; attribute dont_touch of G26891: signal is true;
	signal G26892: std_logic; attribute dont_touch of G26892: signal is true;
	signal G26895: std_logic; attribute dont_touch of G26895: signal is true;
	signal G26896: std_logic; attribute dont_touch of G26896: signal is true;
	signal G26897: std_logic; attribute dont_touch of G26897: signal is true;
	signal G26900: std_logic; attribute dont_touch of G26900: signal is true;
	signal G26901: std_logic; attribute dont_touch of G26901: signal is true;
	signal G26902: std_logic; attribute dont_touch of G26902: signal is true;
	signal G26905: std_logic; attribute dont_touch of G26905: signal is true;
	signal G26906: std_logic; attribute dont_touch of G26906: signal is true;
	signal G26909: std_logic; attribute dont_touch of G26909: signal is true;
	signal G26910: std_logic; attribute dont_touch of G26910: signal is true;
	signal G26911: std_logic; attribute dont_touch of G26911: signal is true;
	signal G26914: std_logic; attribute dont_touch of G26914: signal is true;
	signal G26915: std_logic; attribute dont_touch of G26915: signal is true;
	signal G26918: std_logic; attribute dont_touch of G26918: signal is true;
	signal G26921: std_logic; attribute dont_touch of G26921: signal is true;
	signal G26922: std_logic; attribute dont_touch of G26922: signal is true;
	signal G26925: std_logic; attribute dont_touch of G26925: signal is true;
	signal G26928: std_logic; attribute dont_touch of G26928: signal is true;
	signal G26931: std_logic; attribute dont_touch of G26931: signal is true;
	signal G26934: std_logic; attribute dont_touch of G26934: signal is true;
	signal G26935: std_logic; attribute dont_touch of G26935: signal is true;
	signal G26938: std_logic; attribute dont_touch of G26938: signal is true;
	signal G26941: std_logic; attribute dont_touch of G26941: signal is true;
	signal G26944: std_logic; attribute dont_touch of G26944: signal is true;
	signal G26947: std_logic; attribute dont_touch of G26947: signal is true;
	signal G26950: std_logic; attribute dont_touch of G26950: signal is true;
	signal G26953: std_logic; attribute dont_touch of G26953: signal is true;
	signal G26954: std_logic; attribute dont_touch of G26954: signal is true;
	signal G26955: std_logic; attribute dont_touch of G26955: signal is true;
	signal G26956: std_logic; attribute dont_touch of G26956: signal is true;
	signal G26957: std_logic; attribute dont_touch of G26957: signal is true;
	signal G26958: std_logic; attribute dont_touch of G26958: signal is true;
	signal G26959: std_logic; attribute dont_touch of G26959: signal is true;
	signal G26960: std_logic; attribute dont_touch of G26960: signal is true;
	signal G26961: std_logic; attribute dont_touch of G26961: signal is true;
	signal G26962: std_logic; attribute dont_touch of G26962: signal is true;
	signal G26963: std_logic; attribute dont_touch of G26963: signal is true;
	signal G26964: std_logic; attribute dont_touch of G26964: signal is true;
	signal G26965: std_logic; attribute dont_touch of G26965: signal is true;
	signal G26966: std_logic; attribute dont_touch of G26966: signal is true;
	signal G26967: std_logic; attribute dont_touch of G26967: signal is true;
	signal G26968: std_logic; attribute dont_touch of G26968: signal is true;
	signal G26969: std_logic; attribute dont_touch of G26969: signal is true;
	signal G26970: std_logic; attribute dont_touch of G26970: signal is true;
	signal G26971: std_logic; attribute dont_touch of G26971: signal is true;
	signal G26972: std_logic; attribute dont_touch of G26972: signal is true;
	signal G26973: std_logic; attribute dont_touch of G26973: signal is true;
	signal G26974: std_logic; attribute dont_touch of G26974: signal is true;
	signal G26977: std_logic; attribute dont_touch of G26977: signal is true;
	signal G26978: std_logic; attribute dont_touch of G26978: signal is true;
	signal G26979: std_logic; attribute dont_touch of G26979: signal is true;
	signal G26980: std_logic; attribute dont_touch of G26980: signal is true;
	signal G26981: std_logic; attribute dont_touch of G26981: signal is true;
	signal G26982: std_logic; attribute dont_touch of G26982: signal is true;
	signal G26983: std_logic; attribute dont_touch of G26983: signal is true;
	signal G26984: std_logic; attribute dont_touch of G26984: signal is true;
	signal G26985: std_logic; attribute dont_touch of G26985: signal is true;
	signal G26986: std_logic; attribute dont_touch of G26986: signal is true;
	signal G26987: std_logic; attribute dont_touch of G26987: signal is true;
	signal G26988: std_logic; attribute dont_touch of G26988: signal is true;
	signal G26989: std_logic; attribute dont_touch of G26989: signal is true;
	signal G26993: std_logic; attribute dont_touch of G26993: signal is true;
	signal G26994: std_logic; attribute dont_touch of G26994: signal is true;
	signal G26995: std_logic; attribute dont_touch of G26995: signal is true;
	signal G26996: std_logic; attribute dont_touch of G26996: signal is true;
	signal G26997: std_logic; attribute dont_touch of G26997: signal is true;
	signal G26998: std_logic; attribute dont_touch of G26998: signal is true;
	signal G26999: std_logic; attribute dont_touch of G26999: signal is true;
	signal G27000: std_logic; attribute dont_touch of G27000: signal is true;
	signal G27001: std_logic; attribute dont_touch of G27001: signal is true;
	signal G27002: std_logic; attribute dont_touch of G27002: signal is true;
	signal G27003: std_logic; attribute dont_touch of G27003: signal is true;
	signal G27004: std_logic; attribute dont_touch of G27004: signal is true;
	signal G27005: std_logic; attribute dont_touch of G27005: signal is true;
	signal G27006: std_logic; attribute dont_touch of G27006: signal is true;
	signal G27007: std_logic; attribute dont_touch of G27007: signal is true;
	signal G27008: std_logic; attribute dont_touch of G27008: signal is true;
	signal G27009: std_logic; attribute dont_touch of G27009: signal is true;
	signal G27010: std_logic; attribute dont_touch of G27010: signal is true;
	signal G27011: std_logic; attribute dont_touch of G27011: signal is true;
	signal G27012: std_logic; attribute dont_touch of G27012: signal is true;
	signal G27016: std_logic; attribute dont_touch of G27016: signal is true;
	signal G27017: std_logic; attribute dont_touch of G27017: signal is true;
	signal G27018: std_logic; attribute dont_touch of G27018: signal is true;
	signal G27019: std_logic; attribute dont_touch of G27019: signal is true;
	signal G27020: std_logic; attribute dont_touch of G27020: signal is true;
	signal G27021: std_logic; attribute dont_touch of G27021: signal is true;
	signal G27022: std_logic; attribute dont_touch of G27022: signal is true;
	signal G27023: std_logic; attribute dont_touch of G27023: signal is true;
	signal G27024: std_logic; attribute dont_touch of G27024: signal is true;
	signal G27025: std_logic; attribute dont_touch of G27025: signal is true;
	signal G27026: std_logic; attribute dont_touch of G27026: signal is true;
	signal G27027: std_logic; attribute dont_touch of G27027: signal is true;
	signal G27028: std_logic; attribute dont_touch of G27028: signal is true;
	signal G27029: std_logic; attribute dont_touch of G27029: signal is true;
	signal G27030: std_logic; attribute dont_touch of G27030: signal is true;
	signal G27031: std_logic; attribute dont_touch of G27031: signal is true;
	signal G27032: std_logic; attribute dont_touch of G27032: signal is true;
	signal G27033: std_logic; attribute dont_touch of G27033: signal is true;
	signal G27034: std_logic; attribute dont_touch of G27034: signal is true;
	signal G27035: std_logic; attribute dont_touch of G27035: signal is true;
	signal G27036: std_logic; attribute dont_touch of G27036: signal is true;
	signal G27037: std_logic; attribute dont_touch of G27037: signal is true;
	signal G27038: std_logic; attribute dont_touch of G27038: signal is true;
	signal G27042: std_logic; attribute dont_touch of G27042: signal is true;
	signal G27043: std_logic; attribute dont_touch of G27043: signal is true;
	signal G27044: std_logic; attribute dont_touch of G27044: signal is true;
	signal G27045: std_logic; attribute dont_touch of G27045: signal is true;
	signal G27046: std_logic; attribute dont_touch of G27046: signal is true;
	signal G27047: std_logic; attribute dont_touch of G27047: signal is true;
	signal G27048: std_logic; attribute dont_touch of G27048: signal is true;
	signal G27049: std_logic; attribute dont_touch of G27049: signal is true;
	signal G27050: std_logic; attribute dont_touch of G27050: signal is true;
	signal G27051: std_logic; attribute dont_touch of G27051: signal is true;
	signal G27052: std_logic; attribute dont_touch of G27052: signal is true;
	signal G27053: std_logic; attribute dont_touch of G27053: signal is true;
	signal G27054: std_logic; attribute dont_touch of G27054: signal is true;
	signal G27055: std_logic; attribute dont_touch of G27055: signal is true;
	signal G27056: std_logic; attribute dont_touch of G27056: signal is true;
	signal G27057: std_logic; attribute dont_touch of G27057: signal is true;
	signal G27058: std_logic; attribute dont_touch of G27058: signal is true;
	signal G27059: std_logic; attribute dont_touch of G27059: signal is true;
	signal G27060: std_logic; attribute dont_touch of G27060: signal is true;
	signal G27061: std_logic; attribute dont_touch of G27061: signal is true;
	signal G27062: std_logic; attribute dont_touch of G27062: signal is true;
	signal G27063: std_logic; attribute dont_touch of G27063: signal is true;
	signal G27064: std_logic; attribute dont_touch of G27064: signal is true;
	signal G27065: std_logic; attribute dont_touch of G27065: signal is true;
	signal G27066: std_logic; attribute dont_touch of G27066: signal is true;
	signal G27070: std_logic; attribute dont_touch of G27070: signal is true;
	signal G27071: std_logic; attribute dont_touch of G27071: signal is true;
	signal G27072: std_logic; attribute dont_touch of G27072: signal is true;
	signal G27073: std_logic; attribute dont_touch of G27073: signal is true;
	signal G27074: std_logic; attribute dont_touch of G27074: signal is true;
	signal G27075: std_logic; attribute dont_touch of G27075: signal is true;
	signal G27076: std_logic; attribute dont_touch of G27076: signal is true;
	signal G27077: std_logic; attribute dont_touch of G27077: signal is true;
	signal G27078: std_logic; attribute dont_touch of G27078: signal is true;
	signal G27079: std_logic; attribute dont_touch of G27079: signal is true;
	signal G27080: std_logic; attribute dont_touch of G27080: signal is true;
	signal G27081: std_logic; attribute dont_touch of G27081: signal is true;
	signal G27082: std_logic; attribute dont_touch of G27082: signal is true;
	signal G27083: std_logic; attribute dont_touch of G27083: signal is true;
	signal G27084: std_logic; attribute dont_touch of G27084: signal is true;
	signal G27085: std_logic; attribute dont_touch of G27085: signal is true;
	signal G27086: std_logic; attribute dont_touch of G27086: signal is true;
	signal G27087: std_logic; attribute dont_touch of G27087: signal is true;
	signal G27088: std_logic; attribute dont_touch of G27088: signal is true;
	signal G27089: std_logic; attribute dont_touch of G27089: signal is true;
	signal G27090: std_logic; attribute dont_touch of G27090: signal is true;
	signal G27091: std_logic; attribute dont_touch of G27091: signal is true;
	signal G27092: std_logic; attribute dont_touch of G27092: signal is true;
	signal G27093: std_logic; attribute dont_touch of G27093: signal is true;
	signal G27094: std_logic; attribute dont_touch of G27094: signal is true;
	signal G27095: std_logic; attribute dont_touch of G27095: signal is true;
	signal G27096: std_logic; attribute dont_touch of G27096: signal is true;
	signal G27097: std_logic; attribute dont_touch of G27097: signal is true;
	signal G27098: std_logic; attribute dont_touch of G27098: signal is true;
	signal G27099: std_logic; attribute dont_touch of G27099: signal is true;
	signal G27100: std_logic; attribute dont_touch of G27100: signal is true;
	signal G27101: std_logic; attribute dont_touch of G27101: signal is true;
	signal G27102: std_logic; attribute dont_touch of G27102: signal is true;
	signal G27103: std_logic; attribute dont_touch of G27103: signal is true;
	signal G27104: std_logic; attribute dont_touch of G27104: signal is true;
	signal G27105: std_logic; attribute dont_touch of G27105: signal is true;
	signal G27106: std_logic; attribute dont_touch of G27106: signal is true;
	signal G27107: std_logic; attribute dont_touch of G27107: signal is true;
	signal G27108: std_logic; attribute dont_touch of G27108: signal is true;
	signal G27109: std_logic; attribute dont_touch of G27109: signal is true;
	signal G27110: std_logic; attribute dont_touch of G27110: signal is true;
	signal G27111: std_logic; attribute dont_touch of G27111: signal is true;
	signal G27112: std_logic; attribute dont_touch of G27112: signal is true;
	signal G27113: std_logic; attribute dont_touch of G27113: signal is true;
	signal G27114: std_logic; attribute dont_touch of G27114: signal is true;
	signal G27115: std_logic; attribute dont_touch of G27115: signal is true;
	signal G27116: std_logic; attribute dont_touch of G27116: signal is true;
	signal G27117: std_logic; attribute dont_touch of G27117: signal is true;
	signal G27118: std_logic; attribute dont_touch of G27118: signal is true;
	signal G27119: std_logic; attribute dont_touch of G27119: signal is true;
	signal G27120: std_logic; attribute dont_touch of G27120: signal is true;
	signal G27121: std_logic; attribute dont_touch of G27121: signal is true;
	signal G27122: std_logic; attribute dont_touch of G27122: signal is true;
	signal G27123: std_logic; attribute dont_touch of G27123: signal is true;
	signal G27124: std_logic; attribute dont_touch of G27124: signal is true;
	signal G27125: std_logic; attribute dont_touch of G27125: signal is true;
	signal G27126: std_logic; attribute dont_touch of G27126: signal is true;
	signal G27129: std_logic; attribute dont_touch of G27129: signal is true;
	signal G27130: std_logic; attribute dont_touch of G27130: signal is true;
	signal G27131: std_logic; attribute dont_touch of G27131: signal is true;
	signal G27132: std_logic; attribute dont_touch of G27132: signal is true;
	signal G27133: std_logic; attribute dont_touch of G27133: signal is true;
	signal G27134: std_logic; attribute dont_touch of G27134: signal is true;
	signal G27135: std_logic; attribute dont_touch of G27135: signal is true;
	signal G27136: std_logic; attribute dont_touch of G27136: signal is true;
	signal G27137: std_logic; attribute dont_touch of G27137: signal is true;
	signal G27138: std_logic; attribute dont_touch of G27138: signal is true;
	signal G27139: std_logic; attribute dont_touch of G27139: signal is true;
	signal G27140: std_logic; attribute dont_touch of G27140: signal is true;
	signal G27141: std_logic; attribute dont_touch of G27141: signal is true;
	signal G27142: std_logic; attribute dont_touch of G27142: signal is true;
	signal G27143: std_logic; attribute dont_touch of G27143: signal is true;
	signal G27144: std_logic; attribute dont_touch of G27144: signal is true;
	signal G27145: std_logic; attribute dont_touch of G27145: signal is true;
	signal G27146: std_logic; attribute dont_touch of G27146: signal is true;
	signal G27147: std_logic; attribute dont_touch of G27147: signal is true;
	signal G27148: std_logic; attribute dont_touch of G27148: signal is true;
	signal G27149: std_logic; attribute dont_touch of G27149: signal is true;
	signal G27150: std_logic; attribute dont_touch of G27150: signal is true;
	signal G27151: std_logic; attribute dont_touch of G27151: signal is true;
	signal G27152: std_logic; attribute dont_touch of G27152: signal is true;
	signal G27153: std_logic; attribute dont_touch of G27153: signal is true;
	signal G27154: std_logic; attribute dont_touch of G27154: signal is true;
	signal G27155: std_logic; attribute dont_touch of G27155: signal is true;
	signal G27156: std_logic; attribute dont_touch of G27156: signal is true;
	signal G27157: std_logic; attribute dont_touch of G27157: signal is true;
	signal G27158: std_logic; attribute dont_touch of G27158: signal is true;
	signal G27159: std_logic; attribute dont_touch of G27159: signal is true;
	signal G27160: std_logic; attribute dont_touch of G27160: signal is true;
	signal G27161: std_logic; attribute dont_touch of G27161: signal is true;
	signal G27162: std_logic; attribute dont_touch of G27162: signal is true;
	signal G27163: std_logic; attribute dont_touch of G27163: signal is true;
	signal G27164: std_logic; attribute dont_touch of G27164: signal is true;
	signal G27165: std_logic; attribute dont_touch of G27165: signal is true;
	signal G27166: std_logic; attribute dont_touch of G27166: signal is true;
	signal G27167: std_logic; attribute dont_touch of G27167: signal is true;
	signal G27168: std_logic; attribute dont_touch of G27168: signal is true;
	signal G27171: std_logic; attribute dont_touch of G27171: signal is true;
	signal G27172: std_logic; attribute dont_touch of G27172: signal is true;
	signal G27173: std_logic; attribute dont_touch of G27173: signal is true;
	signal G27174: std_logic; attribute dont_touch of G27174: signal is true;
	signal G27175: std_logic; attribute dont_touch of G27175: signal is true;
	signal G27176: std_logic; attribute dont_touch of G27176: signal is true;
	signal G27177: std_logic; attribute dont_touch of G27177: signal is true;
	signal G27178: std_logic; attribute dont_touch of G27178: signal is true;
	signal G27179: std_logic; attribute dont_touch of G27179: signal is true;
	signal G27180: std_logic; attribute dont_touch of G27180: signal is true;
	signal G27181: std_logic; attribute dont_touch of G27181: signal is true;
	signal G27182: std_logic; attribute dont_touch of G27182: signal is true;
	signal G27183: std_logic; attribute dont_touch of G27183: signal is true;
	signal G27184: std_logic; attribute dont_touch of G27184: signal is true;
	signal G27185: std_logic; attribute dont_touch of G27185: signal is true;
	signal G27186: std_logic; attribute dont_touch of G27186: signal is true;
	signal G27187: std_logic; attribute dont_touch of G27187: signal is true;
	signal G27188: std_logic; attribute dont_touch of G27188: signal is true;
	signal G27189: std_logic; attribute dont_touch of G27189: signal is true;
	signal G27190: std_logic; attribute dont_touch of G27190: signal is true;
	signal G27191: std_logic; attribute dont_touch of G27191: signal is true;
	signal G27192: std_logic; attribute dont_touch of G27192: signal is true;
	signal G27193: std_logic; attribute dont_touch of G27193: signal is true;
	signal G27194: std_logic; attribute dont_touch of G27194: signal is true;
	signal G27195: std_logic; attribute dont_touch of G27195: signal is true;
	signal G27196: std_logic; attribute dont_touch of G27196: signal is true;
	signal G27197: std_logic; attribute dont_touch of G27197: signal is true;
	signal G27198: std_logic; attribute dont_touch of G27198: signal is true;
	signal G27199: std_logic; attribute dont_touch of G27199: signal is true;
	signal G27200: std_logic; attribute dont_touch of G27200: signal is true;
	signal G27201: std_logic; attribute dont_touch of G27201: signal is true;
	signal G27202: std_logic; attribute dont_touch of G27202: signal is true;
	signal G27203: std_logic; attribute dont_touch of G27203: signal is true;
	signal G27204: std_logic; attribute dont_touch of G27204: signal is true;
	signal G27205: std_logic; attribute dont_touch of G27205: signal is true;
	signal G27206: std_logic; attribute dont_touch of G27206: signal is true;
	signal G27207: std_logic; attribute dont_touch of G27207: signal is true;
	signal G27208: std_logic; attribute dont_touch of G27208: signal is true;
	signal G27209: std_logic; attribute dont_touch of G27209: signal is true;
	signal G27210: std_logic; attribute dont_touch of G27210: signal is true;
	signal G27211: std_logic; attribute dont_touch of G27211: signal is true;
	signal G27212: std_logic; attribute dont_touch of G27212: signal is true;
	signal G27213: std_logic; attribute dont_touch of G27213: signal is true;
	signal G27214: std_logic; attribute dont_touch of G27214: signal is true;
	signal G27215: std_logic; attribute dont_touch of G27215: signal is true;
	signal G27216: std_logic; attribute dont_touch of G27216: signal is true;
	signal G27217: std_logic; attribute dont_touch of G27217: signal is true;
	signal G27218: std_logic; attribute dont_touch of G27218: signal is true;
	signal G27219: std_logic; attribute dont_touch of G27219: signal is true;
	signal G27220: std_logic; attribute dont_touch of G27220: signal is true;
	signal G27221: std_logic; attribute dont_touch of G27221: signal is true;
	signal G27222: std_logic; attribute dont_touch of G27222: signal is true;
	signal G27223: std_logic; attribute dont_touch of G27223: signal is true;
	signal G27224: std_logic; attribute dont_touch of G27224: signal is true;
	signal G27225: std_logic; attribute dont_touch of G27225: signal is true;
	signal G27226: std_logic; attribute dont_touch of G27226: signal is true;
	signal G27227: std_logic; attribute dont_touch of G27227: signal is true;
	signal G27228: std_logic; attribute dont_touch of G27228: signal is true;
	signal G27229: std_logic; attribute dont_touch of G27229: signal is true;
	signal G27230: std_logic; attribute dont_touch of G27230: signal is true;
	signal G27231: std_logic; attribute dont_touch of G27231: signal is true;
	signal G27232: std_logic; attribute dont_touch of G27232: signal is true;
	signal G27233: std_logic; attribute dont_touch of G27233: signal is true;
	signal G27234: std_logic; attribute dont_touch of G27234: signal is true;
	signal G27235: std_logic; attribute dont_touch of G27235: signal is true;
	signal G27236: std_logic; attribute dont_touch of G27236: signal is true;
	signal G27237: std_logic; attribute dont_touch of G27237: signal is true;
	signal G27238: std_logic; attribute dont_touch of G27238: signal is true;
	signal G27239: std_logic; attribute dont_touch of G27239: signal is true;
	signal G27240: std_logic; attribute dont_touch of G27240: signal is true;
	signal G27241: std_logic; attribute dont_touch of G27241: signal is true;
	signal G27242: std_logic; attribute dont_touch of G27242: signal is true;
	signal G27243: std_logic; attribute dont_touch of G27243: signal is true;
	signal G27244: std_logic; attribute dont_touch of G27244: signal is true;
	signal G27245: std_logic; attribute dont_touch of G27245: signal is true;
	signal G27246: std_logic; attribute dont_touch of G27246: signal is true;
	signal G27247: std_logic; attribute dont_touch of G27247: signal is true;
	signal G27248: std_logic; attribute dont_touch of G27248: signal is true;
	signal G27249: std_logic; attribute dont_touch of G27249: signal is true;
	signal G27250: std_logic; attribute dont_touch of G27250: signal is true;
	signal G27251: std_logic; attribute dont_touch of G27251: signal is true;
	signal G27252: std_logic; attribute dont_touch of G27252: signal is true;
	signal G27253: std_logic; attribute dont_touch of G27253: signal is true;
	signal G27254: std_logic; attribute dont_touch of G27254: signal is true;
	signal G27255: std_logic; attribute dont_touch of G27255: signal is true;
	signal G27256: std_logic; attribute dont_touch of G27256: signal is true;
	signal G27257: std_logic; attribute dont_touch of G27257: signal is true;
	signal G27258: std_logic; attribute dont_touch of G27258: signal is true;
	signal G27259: std_logic; attribute dont_touch of G27259: signal is true;
	signal G27260: std_logic; attribute dont_touch of G27260: signal is true;
	signal G27261: std_logic; attribute dont_touch of G27261: signal is true;
	signal G27262: std_logic; attribute dont_touch of G27262: signal is true;
	signal G27263: std_logic; attribute dont_touch of G27263: signal is true;
	signal G27264: std_logic; attribute dont_touch of G27264: signal is true;
	signal G27265: std_logic; attribute dont_touch of G27265: signal is true;
	signal G27266: std_logic; attribute dont_touch of G27266: signal is true;
	signal G27267: std_logic; attribute dont_touch of G27267: signal is true;
	signal G27268: std_logic; attribute dont_touch of G27268: signal is true;
	signal G27269: std_logic; attribute dont_touch of G27269: signal is true;
	signal G27270: std_logic; attribute dont_touch of G27270: signal is true;
	signal G27271: std_logic; attribute dont_touch of G27271: signal is true;
	signal G27272: std_logic; attribute dont_touch of G27272: signal is true;
	signal G27273: std_logic; attribute dont_touch of G27273: signal is true;
	signal G27274: std_logic; attribute dont_touch of G27274: signal is true;
	signal G27275: std_logic; attribute dont_touch of G27275: signal is true;
	signal G27276: std_logic; attribute dont_touch of G27276: signal is true;
	signal G27277: std_logic; attribute dont_touch of G27277: signal is true;
	signal G27278: std_logic; attribute dont_touch of G27278: signal is true;
	signal G27279: std_logic; attribute dont_touch of G27279: signal is true;
	signal G27280: std_logic; attribute dont_touch of G27280: signal is true;
	signal G27281: std_logic; attribute dont_touch of G27281: signal is true;
	signal G27282: std_logic; attribute dont_touch of G27282: signal is true;
	signal G27283: std_logic; attribute dont_touch of G27283: signal is true;
	signal G27284: std_logic; attribute dont_touch of G27284: signal is true;
	signal G27285: std_logic; attribute dont_touch of G27285: signal is true;
	signal G27286: std_logic; attribute dont_touch of G27286: signal is true;
	signal G27287: std_logic; attribute dont_touch of G27287: signal is true;
	signal G27288: std_logic; attribute dont_touch of G27288: signal is true;
	signal G27289: std_logic; attribute dont_touch of G27289: signal is true;
	signal G27290: std_logic; attribute dont_touch of G27290: signal is true;
	signal G27291: std_logic; attribute dont_touch of G27291: signal is true;
	signal G27292: std_logic; attribute dont_touch of G27292: signal is true;
	signal G27293: std_logic; attribute dont_touch of G27293: signal is true;
	signal G27294: std_logic; attribute dont_touch of G27294: signal is true;
	signal G27295: std_logic; attribute dont_touch of G27295: signal is true;
	signal G27296: std_logic; attribute dont_touch of G27296: signal is true;
	signal G27297: std_logic; attribute dont_touch of G27297: signal is true;
	signal G27298: std_logic; attribute dont_touch of G27298: signal is true;
	signal G27299: std_logic; attribute dont_touch of G27299: signal is true;
	signal G27300: std_logic; attribute dont_touch of G27300: signal is true;
	signal G27301: std_logic; attribute dont_touch of G27301: signal is true;
	signal G27302: std_logic; attribute dont_touch of G27302: signal is true;
	signal G27303: std_logic; attribute dont_touch of G27303: signal is true;
	signal G27304: std_logic; attribute dont_touch of G27304: signal is true;
	signal G27305: std_logic; attribute dont_touch of G27305: signal is true;
	signal G27306: std_logic; attribute dont_touch of G27306: signal is true;
	signal G27307: std_logic; attribute dont_touch of G27307: signal is true;
	signal G27308: std_logic; attribute dont_touch of G27308: signal is true;
	signal G27309: std_logic; attribute dont_touch of G27309: signal is true;
	signal G27310: std_logic; attribute dont_touch of G27310: signal is true;
	signal G27311: std_logic; attribute dont_touch of G27311: signal is true;
	signal G27312: std_logic; attribute dont_touch of G27312: signal is true;
	signal G27313: std_logic; attribute dont_touch of G27313: signal is true;
	signal G27314: std_logic; attribute dont_touch of G27314: signal is true;
	signal G27315: std_logic; attribute dont_touch of G27315: signal is true;
	signal G27316: std_logic; attribute dont_touch of G27316: signal is true;
	signal G27317: std_logic; attribute dont_touch of G27317: signal is true;
	signal G27318: std_logic; attribute dont_touch of G27318: signal is true;
	signal G27319: std_logic; attribute dont_touch of G27319: signal is true;
	signal G27320: std_logic; attribute dont_touch of G27320: signal is true;
	signal G27321: std_logic; attribute dont_touch of G27321: signal is true;
	signal G27322: std_logic; attribute dont_touch of G27322: signal is true;
	signal G27323: std_logic; attribute dont_touch of G27323: signal is true;
	signal G27324: std_logic; attribute dont_touch of G27324: signal is true;
	signal G27325: std_logic; attribute dont_touch of G27325: signal is true;
	signal G27326: std_logic; attribute dont_touch of G27326: signal is true;
	signal G27327: std_logic; attribute dont_touch of G27327: signal is true;
	signal G27328: std_logic; attribute dont_touch of G27328: signal is true;
	signal G27329: std_logic; attribute dont_touch of G27329: signal is true;
	signal G27330: std_logic; attribute dont_touch of G27330: signal is true;
	signal G27331: std_logic; attribute dont_touch of G27331: signal is true;
	signal G27332: std_logic; attribute dont_touch of G27332: signal is true;
	signal G27333: std_logic; attribute dont_touch of G27333: signal is true;
	signal G27334: std_logic; attribute dont_touch of G27334: signal is true;
	signal G27335: std_logic; attribute dont_touch of G27335: signal is true;
	signal G27336: std_logic; attribute dont_touch of G27336: signal is true;
	signal G27337: std_logic; attribute dont_touch of G27337: signal is true;
	signal G27338: std_logic; attribute dont_touch of G27338: signal is true;
	signal G27339: std_logic; attribute dont_touch of G27339: signal is true;
	signal G27340: std_logic; attribute dont_touch of G27340: signal is true;
	signal G27341: std_logic; attribute dont_touch of G27341: signal is true;
	signal G27342: std_logic; attribute dont_touch of G27342: signal is true;
	signal G27343: std_logic; attribute dont_touch of G27343: signal is true;
	signal G27344: std_logic; attribute dont_touch of G27344: signal is true;
	signal G27345: std_logic; attribute dont_touch of G27345: signal is true;
	signal G27346: std_logic; attribute dont_touch of G27346: signal is true;
	signal G27347: std_logic; attribute dont_touch of G27347: signal is true;
	signal G27348: std_logic; attribute dont_touch of G27348: signal is true;
	signal G27349: std_logic; attribute dont_touch of G27349: signal is true;
	signal G27353: std_logic; attribute dont_touch of G27353: signal is true;
	signal G27354: std_logic; attribute dont_touch of G27354: signal is true;
	signal G27355: std_logic; attribute dont_touch of G27355: signal is true;
	signal G27356: std_logic; attribute dont_touch of G27356: signal is true;
	signal G27357: std_logic; attribute dont_touch of G27357: signal is true;
	signal G27358: std_logic; attribute dont_touch of G27358: signal is true;
	signal G27359: std_logic; attribute dont_touch of G27359: signal is true;
	signal G27360: std_logic; attribute dont_touch of G27360: signal is true;
	signal G27361: std_logic; attribute dont_touch of G27361: signal is true;
	signal G27364: std_logic; attribute dont_touch of G27364: signal is true;
	signal G27365: std_logic; attribute dont_touch of G27365: signal is true;
	signal G27366: std_logic; attribute dont_touch of G27366: signal is true;
	signal G27367: std_logic; attribute dont_touch of G27367: signal is true;
	signal G27370: std_logic; attribute dont_touch of G27370: signal is true;
	signal G27371: std_logic; attribute dont_touch of G27371: signal is true;
	signal G27372: std_logic; attribute dont_touch of G27372: signal is true;
	signal G27373: std_logic; attribute dont_touch of G27373: signal is true;
	signal G27376: std_logic; attribute dont_touch of G27376: signal is true;
	signal G27379: std_logic; attribute dont_touch of G27379: signal is true;
	signal G27381: std_logic; attribute dont_touch of G27381: signal is true;
	signal G27382: std_logic; attribute dont_touch of G27382: signal is true;
	signal G27383: std_logic; attribute dont_touch of G27383: signal is true;
	signal G27384: std_logic; attribute dont_touch of G27384: signal is true;
	signal G27385: std_logic; attribute dont_touch of G27385: signal is true;
	signal G27386: std_logic; attribute dont_touch of G27386: signal is true;
	signal G27387: std_logic; attribute dont_touch of G27387: signal is true;
	signal G27390: std_logic; attribute dont_touch of G27390: signal is true;
	signal G27391: std_logic; attribute dont_touch of G27391: signal is true;
	signal G27394: std_logic; attribute dont_touch of G27394: signal is true;
	signal G27395: std_logic; attribute dont_touch of G27395: signal is true;
	signal G27396: std_logic; attribute dont_touch of G27396: signal is true;
	signal G27397: std_logic; attribute dont_touch of G27397: signal is true;
	signal G27400: std_logic; attribute dont_touch of G27400: signal is true;
	signal G27401: std_logic; attribute dont_touch of G27401: signal is true;
	signal G27404: std_logic; attribute dont_touch of G27404: signal is true;
	signal G27407: std_logic; attribute dont_touch of G27407: signal is true;
	signal G27408: std_logic; attribute dont_touch of G27408: signal is true;
	signal G27409: std_logic; attribute dont_touch of G27409: signal is true;
	signal G27410: std_logic; attribute dont_touch of G27410: signal is true;
	signal G27413: std_logic; attribute dont_touch of G27413: signal is true;
	signal G27414: std_logic; attribute dont_touch of G27414: signal is true;
	signal G27415: std_logic; attribute dont_touch of G27415: signal is true;
	signal G27416: std_logic; attribute dont_touch of G27416: signal is true;
	signal G27419: std_logic; attribute dont_touch of G27419: signal is true;
	signal G27422: std_logic; attribute dont_touch of G27422: signal is true;
	signal G27425: std_logic; attribute dont_touch of G27425: signal is true;
	signal G27426: std_logic; attribute dont_touch of G27426: signal is true;
	signal G27427: std_logic; attribute dont_touch of G27427: signal is true;
	signal G27428: std_logic; attribute dont_touch of G27428: signal is true;
	signal G27431: std_logic; attribute dont_touch of G27431: signal is true;
	signal G27432: std_logic; attribute dont_touch of G27432: signal is true;
	signal G27435: std_logic; attribute dont_touch of G27435: signal is true;
	signal G27436: std_logic; attribute dont_touch of G27436: signal is true;
	signal G27437: std_logic; attribute dont_touch of G27437: signal is true;
	signal G27440: std_logic; attribute dont_touch of G27440: signal is true;
	signal G27443: std_logic; attribute dont_touch of G27443: signal is true;
	signal G27446: std_logic; attribute dont_touch of G27446: signal is true;
	signal G27447: std_logic; attribute dont_touch of G27447: signal is true;
	signal G27448: std_logic; attribute dont_touch of G27448: signal is true;
	signal G27449: std_logic; attribute dont_touch of G27449: signal is true;
	signal G27450: std_logic; attribute dont_touch of G27450: signal is true;
	signal G27451: std_logic; attribute dont_touch of G27451: signal is true;
	signal G27454: std_logic; attribute dont_touch of G27454: signal is true;
	signal G27455: std_logic; attribute dont_touch of G27455: signal is true;
	signal G27456: std_logic; attribute dont_touch of G27456: signal is true;
	signal G27459: std_logic; attribute dont_touch of G27459: signal is true;
	signal G27462: std_logic; attribute dont_touch of G27462: signal is true;
	signal G27463: std_logic; attribute dont_touch of G27463: signal is true;
	signal G27464: std_logic; attribute dont_touch of G27464: signal is true;
	signal G27465: std_logic; attribute dont_touch of G27465: signal is true;
	signal G27466: std_logic; attribute dont_touch of G27466: signal is true;
	signal G27467: std_logic; attribute dont_touch of G27467: signal is true;
	signal G27470: std_logic; attribute dont_touch of G27470: signal is true;
	signal G27471: std_logic; attribute dont_touch of G27471: signal is true;
	signal G27472: std_logic; attribute dont_touch of G27472: signal is true;
	signal G27475: std_logic; attribute dont_touch of G27475: signal is true;
	signal G27478: std_logic; attribute dont_touch of G27478: signal is true;
	signal G27479: std_logic; attribute dont_touch of G27479: signal is true;
	signal G27480: std_logic; attribute dont_touch of G27480: signal is true;
	signal G27481: std_logic; attribute dont_touch of G27481: signal is true;
	signal G27482: std_logic; attribute dont_touch of G27482: signal is true;
	signal G27483: std_logic; attribute dont_touch of G27483: signal is true;
	signal G27484: std_logic; attribute dont_touch of G27484: signal is true;
	signal G27485: std_logic; attribute dont_touch of G27485: signal is true;
	signal G27486: std_logic; attribute dont_touch of G27486: signal is true;
	signal G27489: std_logic; attribute dont_touch of G27489: signal is true;
	signal G27492: std_logic; attribute dont_touch of G27492: signal is true;
	signal G27493: std_logic; attribute dont_touch of G27493: signal is true;
	signal G27494: std_logic; attribute dont_touch of G27494: signal is true;
	signal G27495: std_logic; attribute dont_touch of G27495: signal is true;
	signal G27496: std_logic; attribute dont_touch of G27496: signal is true;
	signal G27497: std_logic; attribute dont_touch of G27497: signal is true;
	signal G27498: std_logic; attribute dont_touch of G27498: signal is true;
	signal G27501: std_logic; attribute dont_touch of G27501: signal is true;
	signal G27502: std_logic; attribute dont_touch of G27502: signal is true;
	signal G27503: std_logic; attribute dont_touch of G27503: signal is true;
	signal G27504: std_logic; attribute dont_touch of G27504: signal is true;
	signal G27505: std_logic; attribute dont_touch of G27505: signal is true;
	signal G27506: std_logic; attribute dont_touch of G27506: signal is true;
	signal G27507: std_logic; attribute dont_touch of G27507: signal is true;
	signal G27508: std_logic; attribute dont_touch of G27508: signal is true;
	signal G27509: std_logic; attribute dont_touch of G27509: signal is true;
	signal G27510: std_logic; attribute dont_touch of G27510: signal is true;
	signal G27513: std_logic; attribute dont_touch of G27513: signal is true;
	signal G27514: std_logic; attribute dont_touch of G27514: signal is true;
	signal G27515: std_logic; attribute dont_touch of G27515: signal is true;
	signal G27516: std_logic; attribute dont_touch of G27516: signal is true;
	signal G27517: std_logic; attribute dont_touch of G27517: signal is true;
	signal G27518: std_logic; attribute dont_touch of G27518: signal is true;
	signal G27521: std_logic; attribute dont_touch of G27521: signal is true;
	signal G27522: std_logic; attribute dont_touch of G27522: signal is true;
	signal G27523: std_logic; attribute dont_touch of G27523: signal is true;
	signal G27524: std_logic; attribute dont_touch of G27524: signal is true;
	signal G27525: std_logic; attribute dont_touch of G27525: signal is true;
	signal G27526: std_logic; attribute dont_touch of G27526: signal is true;
	signal G27527: std_logic; attribute dont_touch of G27527: signal is true;
	signal G27528: std_logic; attribute dont_touch of G27528: signal is true;
	signal G27529: std_logic; attribute dont_touch of G27529: signal is true;
	signal G27530: std_logic; attribute dont_touch of G27530: signal is true;
	signal G27531: std_logic; attribute dont_touch of G27531: signal is true;
	signal G27532: std_logic; attribute dont_touch of G27532: signal is true;
	signal G27533: std_logic; attribute dont_touch of G27533: signal is true;
	signal G27534: std_logic; attribute dont_touch of G27534: signal is true;
	signal G27535: std_logic; attribute dont_touch of G27535: signal is true;
	signal G27538: std_logic; attribute dont_touch of G27538: signal is true;
	signal G27539: std_logic; attribute dont_touch of G27539: signal is true;
	signal G27540: std_logic; attribute dont_touch of G27540: signal is true;
	signal G27541: std_logic; attribute dont_touch of G27541: signal is true;
	signal G27542: std_logic; attribute dont_touch of G27542: signal is true;
	signal G27543: std_logic; attribute dont_touch of G27543: signal is true;
	signal G27546: std_logic; attribute dont_touch of G27546: signal is true;
	signal G27547: std_logic; attribute dont_touch of G27547: signal is true;
	signal G27548: std_logic; attribute dont_touch of G27548: signal is true;
	signal G27549: std_logic; attribute dont_touch of G27549: signal is true;
	signal G27550: std_logic; attribute dont_touch of G27550: signal is true;
	signal G27551: std_logic; attribute dont_touch of G27551: signal is true;
	signal G27552: std_logic; attribute dont_touch of G27552: signal is true;
	signal G27553: std_logic; attribute dont_touch of G27553: signal is true;
	signal G27554: std_logic; attribute dont_touch of G27554: signal is true;
	signal G27555: std_logic; attribute dont_touch of G27555: signal is true;
	signal G27558: std_logic; attribute dont_touch of G27558: signal is true;
	signal G27559: std_logic; attribute dont_touch of G27559: signal is true;
	signal G27560: std_logic; attribute dont_touch of G27560: signal is true;
	signal G27561: std_logic; attribute dont_touch of G27561: signal is true;
	signal G27562: std_logic; attribute dont_touch of G27562: signal is true;
	signal G27563: std_logic; attribute dont_touch of G27563: signal is true;
	signal G27564: std_logic; attribute dont_touch of G27564: signal is true;
	signal G27565: std_logic; attribute dont_touch of G27565: signal is true;
	signal G27566: std_logic; attribute dont_touch of G27566: signal is true;
	signal G27567: std_logic; attribute dont_touch of G27567: signal is true;
	signal G27568: std_logic; attribute dont_touch of G27568: signal is true;
	signal G27569: std_logic; attribute dont_touch of G27569: signal is true;
	signal G27570: std_logic; attribute dont_touch of G27570: signal is true;
	signal G27571: std_logic; attribute dont_touch of G27571: signal is true;
	signal G27572: std_logic; attribute dont_touch of G27572: signal is true;
	signal G27573: std_logic; attribute dont_touch of G27573: signal is true;
	signal G27574: std_logic; attribute dont_touch of G27574: signal is true;
	signal G27575: std_logic; attribute dont_touch of G27575: signal is true;
	signal G27576: std_logic; attribute dont_touch of G27576: signal is true;
	signal G27577: std_logic; attribute dont_touch of G27577: signal is true;
	signal G27578: std_logic; attribute dont_touch of G27578: signal is true;
	signal G27579: std_logic; attribute dont_touch of G27579: signal is true;
	signal G27580: std_logic; attribute dont_touch of G27580: signal is true;
	signal G27581: std_logic; attribute dont_touch of G27581: signal is true;
	signal G27582: std_logic; attribute dont_touch of G27582: signal is true;
	signal G27583: std_logic; attribute dont_touch of G27583: signal is true;
	signal G27584: std_logic; attribute dont_touch of G27584: signal is true;
	signal G27585: std_logic; attribute dont_touch of G27585: signal is true;
	signal G27586: std_logic; attribute dont_touch of G27586: signal is true;
	signal G27587: std_logic; attribute dont_touch of G27587: signal is true;
	signal G27588: std_logic; attribute dont_touch of G27588: signal is true;
	signal G27589: std_logic; attribute dont_touch of G27589: signal is true;
	signal G27590: std_logic; attribute dont_touch of G27590: signal is true;
	signal G27594: std_logic; attribute dont_touch of G27594: signal is true;
	signal G27595: std_logic; attribute dont_touch of G27595: signal is true;
	signal G27599: std_logic; attribute dont_touch of G27599: signal is true;
	signal G27603: std_logic; attribute dont_touch of G27603: signal is true;
	signal G27604: std_logic; attribute dont_touch of G27604: signal is true;
	signal G27608: std_logic; attribute dont_touch of G27608: signal is true;
	signal G27612: std_logic; attribute dont_touch of G27612: signal is true;
	signal G27613: std_logic; attribute dont_touch of G27613: signal is true;
	signal G27617: std_logic; attribute dont_touch of G27617: signal is true;
	signal G27621: std_logic; attribute dont_touch of G27621: signal is true;
	signal G27622: std_logic; attribute dont_touch of G27622: signal is true;
	signal G27626: std_logic; attribute dont_touch of G27626: signal is true;
	signal G27627: std_logic; attribute dont_touch of G27627: signal is true;
	signal G27628: std_logic; attribute dont_touch of G27628: signal is true;
	signal G27629: std_logic; attribute dont_touch of G27629: signal is true;
	signal G27630: std_logic; attribute dont_touch of G27630: signal is true;
	signal G27631: std_logic; attribute dont_touch of G27631: signal is true;
	signal G27632: std_logic; attribute dont_touch of G27632: signal is true;
	signal G27655: std_logic; attribute dont_touch of G27655: signal is true;
	signal G27656: std_logic; attribute dont_touch of G27656: signal is true;
	signal G27657: std_logic; attribute dont_touch of G27657: signal is true;
	signal G27658: std_logic; attribute dont_touch of G27658: signal is true;
	signal G27659: std_logic; attribute dont_touch of G27659: signal is true;
	signal G27660: std_logic; attribute dont_touch of G27660: signal is true;
	signal G27661: std_logic; attribute dont_touch of G27661: signal is true;
	signal G27662: std_logic; attribute dont_touch of G27662: signal is true;
	signal G27666: std_logic; attribute dont_touch of G27666: signal is true;
	signal G27667: std_logic; attribute dont_touch of G27667: signal is true;
	signal G27671: std_logic; attribute dont_touch of G27671: signal is true;
	signal G27672: std_logic; attribute dont_touch of G27672: signal is true;
	signal G27673: std_logic; attribute dont_touch of G27673: signal is true;
	signal G27674: std_logic; attribute dont_touch of G27674: signal is true;
	signal G27678: std_logic; attribute dont_touch of G27678: signal is true;
	signal G27679: std_logic; attribute dont_touch of G27679: signal is true;
	signal G27680: std_logic; attribute dont_touch of G27680: signal is true;
	signal G27681: std_logic; attribute dont_touch of G27681: signal is true;
	signal G27682: std_logic; attribute dont_touch of G27682: signal is true;
	signal G27683: std_logic; attribute dont_touch of G27683: signal is true;
	signal G27684: std_logic; attribute dont_touch of G27684: signal is true;
	signal G27685: std_logic; attribute dont_touch of G27685: signal is true;
	signal G27686: std_logic; attribute dont_touch of G27686: signal is true;
	signal G27687: std_logic; attribute dont_touch of G27687: signal is true;
	signal G27688: std_logic; attribute dont_touch of G27688: signal is true;
	signal G27689: std_logic; attribute dont_touch of G27689: signal is true;
	signal G27690: std_logic; attribute dont_touch of G27690: signal is true;
	signal G27691: std_logic; attribute dont_touch of G27691: signal is true;
	signal G27692: std_logic; attribute dont_touch of G27692: signal is true;
	signal G27693: std_logic; attribute dont_touch of G27693: signal is true;
	signal G27694: std_logic; attribute dont_touch of G27694: signal is true;
	signal G27695: std_logic; attribute dont_touch of G27695: signal is true;
	signal G27696: std_logic; attribute dont_touch of G27696: signal is true;
	signal G27697: std_logic; attribute dont_touch of G27697: signal is true;
	signal G27698: std_logic; attribute dont_touch of G27698: signal is true;
	signal G27699: std_logic; attribute dont_touch of G27699: signal is true;
	signal G27700: std_logic; attribute dont_touch of G27700: signal is true;
	signal G27701: std_logic; attribute dont_touch of G27701: signal is true;
	signal G27702: std_logic; attribute dont_touch of G27702: signal is true;
	signal G27703: std_logic; attribute dont_touch of G27703: signal is true;
	signal G27704: std_logic; attribute dont_touch of G27704: signal is true;
	signal G27705: std_logic; attribute dont_touch of G27705: signal is true;
	signal G27706: std_logic; attribute dont_touch of G27706: signal is true;
	signal G27707: std_logic; attribute dont_touch of G27707: signal is true;
	signal G27708: std_logic; attribute dont_touch of G27708: signal is true;
	signal G27709: std_logic; attribute dont_touch of G27709: signal is true;
	signal G27710: std_logic; attribute dont_touch of G27710: signal is true;
	signal G27711: std_logic; attribute dont_touch of G27711: signal is true;
	signal G27712: std_logic; attribute dont_touch of G27712: signal is true;
	signal G27713: std_logic; attribute dont_touch of G27713: signal is true;
	signal G27714: std_logic; attribute dont_touch of G27714: signal is true;
	signal G27715: std_logic; attribute dont_touch of G27715: signal is true;
	signal G27716: std_logic; attribute dont_touch of G27716: signal is true;
	signal G27717: std_logic; attribute dont_touch of G27717: signal is true;
	signal G27718: std_logic; attribute dont_touch of G27718: signal is true;
	signal G27719: std_logic; attribute dont_touch of G27719: signal is true;
	signal G27720: std_logic; attribute dont_touch of G27720: signal is true;
	signal G27721: std_logic; attribute dont_touch of G27721: signal is true;
	signal G27722: std_logic; attribute dont_touch of G27722: signal is true;
	signal G27723: std_logic; attribute dont_touch of G27723: signal is true;
	signal G27724: std_logic; attribute dont_touch of G27724: signal is true;
	signal G27725: std_logic; attribute dont_touch of G27725: signal is true;
	signal G27726: std_logic; attribute dont_touch of G27726: signal is true;
	signal G27727: std_logic; attribute dont_touch of G27727: signal is true;
	signal G27728: std_logic; attribute dont_touch of G27728: signal is true;
	signal G27729: std_logic; attribute dont_touch of G27729: signal is true;
	signal G27730: std_logic; attribute dont_touch of G27730: signal is true;
	signal G27731: std_logic; attribute dont_touch of G27731: signal is true;
	signal G27732: std_logic; attribute dont_touch of G27732: signal is true;
	signal G27733: std_logic; attribute dont_touch of G27733: signal is true;
	signal G27734: std_logic; attribute dont_touch of G27734: signal is true;
	signal G27735: std_logic; attribute dont_touch of G27735: signal is true;
	signal G27736: std_logic; attribute dont_touch of G27736: signal is true;
	signal G27737: std_logic; attribute dont_touch of G27737: signal is true;
	signal G27738: std_logic; attribute dont_touch of G27738: signal is true;
	signal G27741: std_logic; attribute dont_touch of G27741: signal is true;
	signal G27742: std_logic; attribute dont_touch of G27742: signal is true;
	signal G27743: std_logic; attribute dont_touch of G27743: signal is true;
	signal G27746: std_logic; attribute dont_touch of G27746: signal is true;
	signal G27747: std_logic; attribute dont_touch of G27747: signal is true;
	signal G27748: std_logic; attribute dont_touch of G27748: signal is true;
	signal G27751: std_logic; attribute dont_touch of G27751: signal is true;
	signal G27754: std_logic; attribute dont_touch of G27754: signal is true;
	signal G27755: std_logic; attribute dont_touch of G27755: signal is true;
	signal G27756: std_logic; attribute dont_touch of G27756: signal is true;
	signal G27759: std_logic; attribute dont_touch of G27759: signal is true;
	signal G27760: std_logic; attribute dont_touch of G27760: signal is true;
	signal G27761: std_logic; attribute dont_touch of G27761: signal is true;
	signal G27762: std_logic; attribute dont_touch of G27762: signal is true;
	signal G27763: std_logic; attribute dont_touch of G27763: signal is true;
	signal G27764: std_logic; attribute dont_touch of G27764: signal is true;
	signal G27765: std_logic; attribute dont_touch of G27765: signal is true;
	signal G27766: std_logic; attribute dont_touch of G27766: signal is true;
	signal G27767: std_logic; attribute dont_touch of G27767: signal is true;
	signal G27768: std_logic; attribute dont_touch of G27768: signal is true;
	signal G27769: std_logic; attribute dont_touch of G27769: signal is true;
	signal G27770: std_logic; attribute dont_touch of G27770: signal is true;
	signal G27771: std_logic; attribute dont_touch of G27771: signal is true;
	signal G27772: std_logic; attribute dont_touch of G27772: signal is true;
	signal G27773: std_logic; attribute dont_touch of G27773: signal is true;
	signal G27774: std_logic; attribute dont_touch of G27774: signal is true;
	signal G27775: std_logic; attribute dont_touch of G27775: signal is true;
	signal G27776: std_logic; attribute dont_touch of G27776: signal is true;
	signal G27779: std_logic; attribute dont_touch of G27779: signal is true;
	signal G27780: std_logic; attribute dont_touch of G27780: signal is true;
	signal G27783: std_logic; attribute dont_touch of G27783: signal is true;
	signal G27784: std_logic; attribute dont_touch of G27784: signal is true;
	signal G27785: std_logic; attribute dont_touch of G27785: signal is true;
	signal G27786: std_logic; attribute dont_touch of G27786: signal is true;
	signal G27787: std_logic; attribute dont_touch of G27787: signal is true;
	signal G27790: std_logic; attribute dont_touch of G27790: signal is true;
	signal G27791: std_logic; attribute dont_touch of G27791: signal is true;
	signal G27792: std_logic; attribute dont_touch of G27792: signal is true;
	signal G27793: std_logic; attribute dont_touch of G27793: signal is true;
	signal G27794: std_logic; attribute dont_touch of G27794: signal is true;
	signal G27797: std_logic; attribute dont_touch of G27797: signal is true;
	signal G27798: std_logic; attribute dont_touch of G27798: signal is true;
	signal G27799: std_logic; attribute dont_touch of G27799: signal is true;
	signal G27800: std_logic; attribute dont_touch of G27800: signal is true;
	signal G27801: std_logic; attribute dont_touch of G27801: signal is true;
	signal G27802: std_logic; attribute dont_touch of G27802: signal is true;
	signal G27805: std_logic; attribute dont_touch of G27805: signal is true;
	signal G27806: std_logic; attribute dont_touch of G27806: signal is true;
	signal G27809: std_logic; attribute dont_touch of G27809: signal is true;
	signal G27810: std_logic; attribute dont_touch of G27810: signal is true;
	signal G27811: std_logic; attribute dont_touch of G27811: signal is true;
	signal G27814: std_logic; attribute dont_touch of G27814: signal is true;
	signal G27817: std_logic; attribute dont_touch of G27817: signal is true;
	signal G27820: std_logic; attribute dont_touch of G27820: signal is true;
	signal G27823: std_logic; attribute dont_touch of G27823: signal is true;
	signal G27824: std_logic; attribute dont_touch of G27824: signal is true;
	signal G27827: std_logic; attribute dont_touch of G27827: signal is true;
	signal G27830: std_logic; attribute dont_touch of G27830: signal is true;
	signal G27831: std_logic; attribute dont_touch of G27831: signal is true;
	signal G27834: std_logic; attribute dont_touch of G27834: signal is true;
	signal G27838: std_logic; attribute dont_touch of G27838: signal is true;
	signal G27839: std_logic; attribute dont_touch of G27839: signal is true;
	signal G27842: std_logic; attribute dont_touch of G27842: signal is true;
	signal G27843: std_logic; attribute dont_touch of G27843: signal is true;
	signal G27846: std_logic; attribute dont_touch of G27846: signal is true;
	signal G27847: std_logic; attribute dont_touch of G27847: signal is true;
	signal G27850: std_logic; attribute dont_touch of G27850: signal is true;
	signal G27854: std_logic; attribute dont_touch of G27854: signal is true;
	signal G27855: std_logic; attribute dont_touch of G27855: signal is true;
	signal G27858: std_logic; attribute dont_touch of G27858: signal is true;
	signal G27861: std_logic; attribute dont_touch of G27861: signal is true;
	signal G27864: std_logic; attribute dont_touch of G27864: signal is true;
	signal G27865: std_logic; attribute dont_touch of G27865: signal is true;
	signal G27868: std_logic; attribute dont_touch of G27868: signal is true;
	signal G27869: std_logic; attribute dont_touch of G27869: signal is true;
	signal G27872: std_logic; attribute dont_touch of G27872: signal is true;
	signal G27875: std_logic; attribute dont_touch of G27875: signal is true;
	signal G27879: std_logic; attribute dont_touch of G27879: signal is true;
	signal G27882: std_logic; attribute dont_touch of G27882: signal is true;
	signal G27883: std_logic; attribute dont_touch of G27883: signal is true;
	signal G27886: std_logic; attribute dont_touch of G27886: signal is true;
	signal G27889: std_logic; attribute dont_touch of G27889: signal is true;
	signal G27892: std_logic; attribute dont_touch of G27892: signal is true;
	signal G27896: std_logic; attribute dont_touch of G27896: signal is true;
	signal G27897: std_logic; attribute dont_touch of G27897: signal is true;
	signal G27900: std_logic; attribute dont_touch of G27900: signal is true;
	signal G27903: std_logic; attribute dont_touch of G27903: signal is true;
	signal G27904: std_logic; attribute dont_touch of G27904: signal is true;
	signal G27905: std_logic; attribute dont_touch of G27905: signal is true;
	signal G27906: std_logic; attribute dont_touch of G27906: signal is true;
	signal G27907: std_logic; attribute dont_touch of G27907: signal is true;
	signal G27908: std_logic; attribute dont_touch of G27908: signal is true;
	signal G27909: std_logic; attribute dont_touch of G27909: signal is true;
	signal G27910: std_logic; attribute dont_touch of G27910: signal is true;
	signal G27911: std_logic; attribute dont_touch of G27911: signal is true;
	signal G27912: std_logic; attribute dont_touch of G27912: signal is true;
	signal G27913: std_logic; attribute dont_touch of G27913: signal is true;
	signal G27914: std_logic; attribute dont_touch of G27914: signal is true;
	signal G27915: std_logic; attribute dont_touch of G27915: signal is true;
	signal G27916: std_logic; attribute dont_touch of G27916: signal is true;
	signal G27917: std_logic; attribute dont_touch of G27917: signal is true;
	signal G27918: std_logic; attribute dont_touch of G27918: signal is true;
	signal G27919: std_logic; attribute dont_touch of G27919: signal is true;
	signal G27922: std_logic; attribute dont_touch of G27922: signal is true;
	signal G27923: std_logic; attribute dont_touch of G27923: signal is true;
	signal G27924: std_logic; attribute dont_touch of G27924: signal is true;
	signal G27925: std_logic; attribute dont_touch of G27925: signal is true;
	signal G27926: std_logic; attribute dont_touch of G27926: signal is true;
	signal G27927: std_logic; attribute dont_touch of G27927: signal is true;
	signal G27928: std_logic; attribute dont_touch of G27928: signal is true;
	signal G27931: std_logic; attribute dont_touch of G27931: signal is true;
	signal G27932: std_logic; attribute dont_touch of G27932: signal is true;
	signal G27935: std_logic; attribute dont_touch of G27935: signal is true;
	signal G27936: std_logic; attribute dont_touch of G27936: signal is true;
	signal G27937: std_logic; attribute dont_touch of G27937: signal is true;
	signal G27938: std_logic; attribute dont_touch of G27938: signal is true;
	signal G27939: std_logic; attribute dont_touch of G27939: signal is true;
	signal G27942: std_logic; attribute dont_touch of G27942: signal is true;
	signal G27945: std_logic; attribute dont_touch of G27945: signal is true;
	signal G27946: std_logic; attribute dont_touch of G27946: signal is true;
	signal G27949: std_logic; attribute dont_touch of G27949: signal is true;
	signal G27950: std_logic; attribute dont_touch of G27950: signal is true;
	signal G27951: std_logic; attribute dont_touch of G27951: signal is true;
	signal G27952: std_logic; attribute dont_touch of G27952: signal is true;
	signal G27955: std_logic; attribute dont_touch of G27955: signal is true;
	signal G27956: std_logic; attribute dont_touch of G27956: signal is true;
	signal G27959: std_logic; attribute dont_touch of G27959: signal is true;
	signal G27962: std_logic; attribute dont_touch of G27962: signal is true;
	signal G27963: std_logic; attribute dont_touch of G27963: signal is true;
	signal G27964: std_logic; attribute dont_touch of G27964: signal is true;
	signal G27965: std_logic; attribute dont_touch of G27965: signal is true;
	signal G27968: std_logic; attribute dont_touch of G27968: signal is true;
	signal G27969: std_logic; attribute dont_touch of G27969: signal is true;
	signal G27970: std_logic; attribute dont_touch of G27970: signal is true;
	signal G27971: std_logic; attribute dont_touch of G27971: signal is true;
	signal G27972: std_logic; attribute dont_touch of G27972: signal is true;
	signal G27973: std_logic; attribute dont_touch of G27973: signal is true;
	signal G27976: std_logic; attribute dont_touch of G27976: signal is true;
	signal G27977: std_logic; attribute dont_touch of G27977: signal is true;
	signal G27980: std_logic; attribute dont_touch of G27980: signal is true;
	signal G27981: std_logic; attribute dont_touch of G27981: signal is true;
	signal G27984: std_logic; attribute dont_touch of G27984: signal is true;
	signal G27985: std_logic; attribute dont_touch of G27985: signal is true;
	signal G27986: std_logic; attribute dont_touch of G27986: signal is true;
	signal G27987: std_logic; attribute dont_touch of G27987: signal is true;
	signal G27988: std_logic; attribute dont_touch of G27988: signal is true;
	signal G27989: std_logic; attribute dont_touch of G27989: signal is true;
	signal G27990: std_logic; attribute dont_touch of G27990: signal is true;
	signal G27991: std_logic; attribute dont_touch of G27991: signal is true;
	signal G27992: std_logic; attribute dont_touch of G27992: signal is true;
	signal G27993: std_logic; attribute dont_touch of G27993: signal is true;
	signal G27994: std_logic; attribute dont_touch of G27994: signal is true;
	signal G27997: std_logic; attribute dont_touch of G27997: signal is true;
	signal G27998: std_logic; attribute dont_touch of G27998: signal is true;
	signal G27999: std_logic; attribute dont_touch of G27999: signal is true;
	signal G28002: std_logic; attribute dont_touch of G28002: signal is true;
	signal G28003: std_logic; attribute dont_touch of G28003: signal is true;
	signal G28004: std_logic; attribute dont_touch of G28004: signal is true;
	signal G28005: std_logic; attribute dont_touch of G28005: signal is true;
	signal G28006: std_logic; attribute dont_touch of G28006: signal is true;
	signal G28007: std_logic; attribute dont_touch of G28007: signal is true;
	signal G28008: std_logic; attribute dont_touch of G28008: signal is true;
	signal G28009: std_logic; attribute dont_touch of G28009: signal is true;
	signal G28010: std_logic; attribute dont_touch of G28010: signal is true;
	signal G28011: std_logic; attribute dont_touch of G28011: signal is true;
	signal G28012: std_logic; attribute dont_touch of G28012: signal is true;
	signal G28013: std_logic; attribute dont_touch of G28013: signal is true;
	signal G28014: std_logic; attribute dont_touch of G28014: signal is true;
	signal G28015: std_logic; attribute dont_touch of G28015: signal is true;
	signal G28016: std_logic; attribute dont_touch of G28016: signal is true;
	signal G28017: std_logic; attribute dont_touch of G28017: signal is true;
	signal G28018: std_logic; attribute dont_touch of G28018: signal is true;
	signal G28021: std_logic; attribute dont_touch of G28021: signal is true;
	signal G28022: std_logic; attribute dont_touch of G28022: signal is true;
	signal G28023: std_logic; attribute dont_touch of G28023: signal is true;
	signal G28024: std_logic; attribute dont_touch of G28024: signal is true;
	signal G28025: std_logic; attribute dont_touch of G28025: signal is true;
	signal G28026: std_logic; attribute dont_touch of G28026: signal is true;
	signal G28027: std_logic; attribute dont_touch of G28027: signal is true;
	signal G28028: std_logic; attribute dont_touch of G28028: signal is true;
	signal G28029: std_logic; attribute dont_touch of G28029: signal is true;
	signal G28030: std_logic; attribute dont_touch of G28030: signal is true;
	signal G28031: std_logic; attribute dont_touch of G28031: signal is true;
	signal G28032: std_logic; attribute dont_touch of G28032: signal is true;
	signal G28033: std_logic; attribute dont_touch of G28033: signal is true;
	signal G28034: std_logic; attribute dont_touch of G28034: signal is true;
	signal G28035: std_logic; attribute dont_touch of G28035: signal is true;
	signal G28036: std_logic; attribute dont_touch of G28036: signal is true;
	signal G28037: std_logic; attribute dont_touch of G28037: signal is true;
	signal G28038: std_logic; attribute dont_touch of G28038: signal is true;
	signal G28039: std_logic; attribute dont_touch of G28039: signal is true;
	signal G28040: std_logic; attribute dont_touch of G28040: signal is true;
	signal G28041: std_logic; attribute dont_touch of G28041: signal is true;
	signal G28042: std_logic; attribute dont_touch of G28042: signal is true;
	signal G28043: std_logic; attribute dont_touch of G28043: signal is true;
	signal G28044: std_logic; attribute dont_touch of G28044: signal is true;
	signal G28045: std_logic; attribute dont_touch of G28045: signal is true;
	signal G28046: std_logic; attribute dont_touch of G28046: signal is true;
	signal G28047: std_logic; attribute dont_touch of G28047: signal is true;
	signal G28048: std_logic; attribute dont_touch of G28048: signal is true;
	signal G28049: std_logic; attribute dont_touch of G28049: signal is true;
	signal G28050: std_logic; attribute dont_touch of G28050: signal is true;
	signal G28051: std_logic; attribute dont_touch of G28051: signal is true;
	signal G28052: std_logic; attribute dont_touch of G28052: signal is true;
	signal G28053: std_logic; attribute dont_touch of G28053: signal is true;
	signal G28054: std_logic; attribute dont_touch of G28054: signal is true;
	signal G28055: std_logic; attribute dont_touch of G28055: signal is true;
	signal G28056: std_logic; attribute dont_touch of G28056: signal is true;
	signal G28057: std_logic; attribute dont_touch of G28057: signal is true;
	signal G28058: std_logic; attribute dont_touch of G28058: signal is true;
	signal G28059: std_logic; attribute dont_touch of G28059: signal is true;
	signal G28060: std_logic; attribute dont_touch of G28060: signal is true;
	signal G28061: std_logic; attribute dont_touch of G28061: signal is true;
	signal G28062: std_logic; attribute dont_touch of G28062: signal is true;
	signal G28063: std_logic; attribute dont_touch of G28063: signal is true;
	signal G28064: std_logic; attribute dont_touch of G28064: signal is true;
	signal G28065: std_logic; attribute dont_touch of G28065: signal is true;
	signal G28066: std_logic; attribute dont_touch of G28066: signal is true;
	signal G28067: std_logic; attribute dont_touch of G28067: signal is true;
	signal G28068: std_logic; attribute dont_touch of G28068: signal is true;
	signal G28069: std_logic; attribute dont_touch of G28069: signal is true;
	signal G28070: std_logic; attribute dont_touch of G28070: signal is true;
	signal G28071: std_logic; attribute dont_touch of G28071: signal is true;
	signal G28072: std_logic; attribute dont_touch of G28072: signal is true;
	signal G28073: std_logic; attribute dont_touch of G28073: signal is true;
	signal G28074: std_logic; attribute dont_touch of G28074: signal is true;
	signal G28075: std_logic; attribute dont_touch of G28075: signal is true;
	signal G28076: std_logic; attribute dont_touch of G28076: signal is true;
	signal G28077: std_logic; attribute dont_touch of G28077: signal is true;
	signal G28078: std_logic; attribute dont_touch of G28078: signal is true;
	signal G28079: std_logic; attribute dont_touch of G28079: signal is true;
	signal G28080: std_logic; attribute dont_touch of G28080: signal is true;
	signal G28081: std_logic; attribute dont_touch of G28081: signal is true;
	signal G28082: std_logic; attribute dont_touch of G28082: signal is true;
	signal G28083: std_logic; attribute dont_touch of G28083: signal is true;
	signal G28084: std_logic; attribute dont_touch of G28084: signal is true;
	signal G28085: std_logic; attribute dont_touch of G28085: signal is true;
	signal G28086: std_logic; attribute dont_touch of G28086: signal is true;
	signal G28087: std_logic; attribute dont_touch of G28087: signal is true;
	signal G28088: std_logic; attribute dont_touch of G28088: signal is true;
	signal G28089: std_logic; attribute dont_touch of G28089: signal is true;
	signal G28090: std_logic; attribute dont_touch of G28090: signal is true;
	signal G28091: std_logic; attribute dont_touch of G28091: signal is true;
	signal G28092: std_logic; attribute dont_touch of G28092: signal is true;
	signal G28093: std_logic; attribute dont_touch of G28093: signal is true;
	signal G28094: std_logic; attribute dont_touch of G28094: signal is true;
	signal G28095: std_logic; attribute dont_touch of G28095: signal is true;
	signal G28096: std_logic; attribute dont_touch of G28096: signal is true;
	signal G28097: std_logic; attribute dont_touch of G28097: signal is true;
	signal G28098: std_logic; attribute dont_touch of G28098: signal is true;
	signal G28099: std_logic; attribute dont_touch of G28099: signal is true;
	signal G28100: std_logic; attribute dont_touch of G28100: signal is true;
	signal G28101: std_logic; attribute dont_touch of G28101: signal is true;
	signal G28102: std_logic; attribute dont_touch of G28102: signal is true;
	signal G28103: std_logic; attribute dont_touch of G28103: signal is true;
	signal G28104: std_logic; attribute dont_touch of G28104: signal is true;
	signal G28105: std_logic; attribute dont_touch of G28105: signal is true;
	signal G28106: std_logic; attribute dont_touch of G28106: signal is true;
	signal G28107: std_logic; attribute dont_touch of G28107: signal is true;
	signal G28108: std_logic; attribute dont_touch of G28108: signal is true;
	signal G28109: std_logic; attribute dont_touch of G28109: signal is true;
	signal G28110: std_logic; attribute dont_touch of G28110: signal is true;
	signal G28111: std_logic; attribute dont_touch of G28111: signal is true;
	signal G28112: std_logic; attribute dont_touch of G28112: signal is true;
	signal G28113: std_logic; attribute dont_touch of G28113: signal is true;
	signal G28114: std_logic; attribute dont_touch of G28114: signal is true;
	signal G28115: std_logic; attribute dont_touch of G28115: signal is true;
	signal G28116: std_logic; attribute dont_touch of G28116: signal is true;
	signal G28117: std_logic; attribute dont_touch of G28117: signal is true;
	signal G28118: std_logic; attribute dont_touch of G28118: signal is true;
	signal G28119: std_logic; attribute dont_touch of G28119: signal is true;
	signal G28120: std_logic; attribute dont_touch of G28120: signal is true;
	signal G28121: std_logic; attribute dont_touch of G28121: signal is true;
	signal G28122: std_logic; attribute dont_touch of G28122: signal is true;
	signal G28123: std_logic; attribute dont_touch of G28123: signal is true;
	signal G28124: std_logic; attribute dont_touch of G28124: signal is true;
	signal G28125: std_logic; attribute dont_touch of G28125: signal is true;
	signal G28126: std_logic; attribute dont_touch of G28126: signal is true;
	signal G28127: std_logic; attribute dont_touch of G28127: signal is true;
	signal G28128: std_logic; attribute dont_touch of G28128: signal is true;
	signal G28132: std_logic; attribute dont_touch of G28132: signal is true;
	signal G28133: std_logic; attribute dont_touch of G28133: signal is true;
	signal G28137: std_logic; attribute dont_touch of G28137: signal is true;
	signal G28141: std_logic; attribute dont_touch of G28141: signal is true;
	signal G28145: std_logic; attribute dont_touch of G28145: signal is true;
	signal G28146: std_logic; attribute dont_touch of G28146: signal is true;
	signal G28147: std_logic; attribute dont_touch of G28147: signal is true;
	signal G28148: std_logic; attribute dont_touch of G28148: signal is true;
	signal G28149: std_logic; attribute dont_touch of G28149: signal is true;
	signal G28150: std_logic; attribute dont_touch of G28150: signal is true;
	signal G28151: std_logic; attribute dont_touch of G28151: signal is true;
	signal G28152: std_logic; attribute dont_touch of G28152: signal is true;
	signal G28153: std_logic; attribute dont_touch of G28153: signal is true;
	signal G28154: std_logic; attribute dont_touch of G28154: signal is true;
	signal G28155: std_logic; attribute dont_touch of G28155: signal is true;
	signal G28156: std_logic; attribute dont_touch of G28156: signal is true;
	signal G28157: std_logic; attribute dont_touch of G28157: signal is true;
	signal G28158: std_logic; attribute dont_touch of G28158: signal is true;
	signal G28159: std_logic; attribute dont_touch of G28159: signal is true;
	signal G28160: std_logic; attribute dont_touch of G28160: signal is true;
	signal G28161: std_logic; attribute dont_touch of G28161: signal is true;
	signal G28162: std_logic; attribute dont_touch of G28162: signal is true;
	signal G28163: std_logic; attribute dont_touch of G28163: signal is true;
	signal G28164: std_logic; attribute dont_touch of G28164: signal is true;
	signal G28165: std_logic; attribute dont_touch of G28165: signal is true;
	signal G28166: std_logic; attribute dont_touch of G28166: signal is true;
	signal G28167: std_logic; attribute dont_touch of G28167: signal is true;
	signal G28168: std_logic; attribute dont_touch of G28168: signal is true;
	signal G28169: std_logic; attribute dont_touch of G28169: signal is true;
	signal G28170: std_logic; attribute dont_touch of G28170: signal is true;
	signal G28171: std_logic; attribute dont_touch of G28171: signal is true;
	signal G28172: std_logic; attribute dont_touch of G28172: signal is true;
	signal G28173: std_logic; attribute dont_touch of G28173: signal is true;
	signal G28174: std_logic; attribute dont_touch of G28174: signal is true;
	signal G28175: std_logic; attribute dont_touch of G28175: signal is true;
	signal G28176: std_logic; attribute dont_touch of G28176: signal is true;
	signal G28177: std_logic; attribute dont_touch of G28177: signal is true;
	signal G28178: std_logic; attribute dont_touch of G28178: signal is true;
	signal G28179: std_logic; attribute dont_touch of G28179: signal is true;
	signal G28185: std_logic; attribute dont_touch of G28185: signal is true;
	signal G28186: std_logic; attribute dont_touch of G28186: signal is true;
	signal G28187: std_logic; attribute dont_touch of G28187: signal is true;
	signal G28188: std_logic; attribute dont_touch of G28188: signal is true;
	signal G28189: std_logic; attribute dont_touch of G28189: signal is true;
	signal G28190: std_logic; attribute dont_touch of G28190: signal is true;
	signal G28191: std_logic; attribute dont_touch of G28191: signal is true;
	signal G28192: std_logic; attribute dont_touch of G28192: signal is true;
	signal G28193: std_logic; attribute dont_touch of G28193: signal is true;
	signal G28194: std_logic; attribute dont_touch of G28194: signal is true;
	signal G28199: std_logic; attribute dont_touch of G28199: signal is true;
	signal G28200: std_logic; attribute dont_touch of G28200: signal is true;
	signal G28206: std_logic; attribute dont_touch of G28206: signal is true;
	signal G28207: std_logic; attribute dont_touch of G28207: signal is true;
	signal G28208: std_logic; attribute dont_touch of G28208: signal is true;
	signal G28209: std_logic; attribute dont_touch of G28209: signal is true;
	signal G28210: std_logic; attribute dont_touch of G28210: signal is true;
	signal G28211: std_logic; attribute dont_touch of G28211: signal is true;
	signal G28212: std_logic; attribute dont_touch of G28212: signal is true;
	signal G28213: std_logic; attribute dont_touch of G28213: signal is true;
	signal G28214: std_logic; attribute dont_touch of G28214: signal is true;
	signal G28215: std_logic; attribute dont_touch of G28215: signal is true;
	signal G28216: std_logic; attribute dont_touch of G28216: signal is true;
	signal G28217: std_logic; attribute dont_touch of G28217: signal is true;
	signal G28218: std_logic; attribute dont_touch of G28218: signal is true;
	signal G28219: std_logic; attribute dont_touch of G28219: signal is true;
	signal G28220: std_logic; attribute dont_touch of G28220: signal is true;
	signal G28221: std_logic; attribute dont_touch of G28221: signal is true;
	signal G28222: std_logic; attribute dont_touch of G28222: signal is true;
	signal G28223: std_logic; attribute dont_touch of G28223: signal is true;
	signal G28224: std_logic; attribute dont_touch of G28224: signal is true;
	signal G28225: std_logic; attribute dont_touch of G28225: signal is true;
	signal G28226: std_logic; attribute dont_touch of G28226: signal is true;
	signal G28227: std_logic; attribute dont_touch of G28227: signal is true;
	signal G28228: std_logic; attribute dont_touch of G28228: signal is true;
	signal G28229: std_logic; attribute dont_touch of G28229: signal is true;
	signal G28230: std_logic; attribute dont_touch of G28230: signal is true;
	signal G28231: std_logic; attribute dont_touch of G28231: signal is true;
	signal G28232: std_logic; attribute dont_touch of G28232: signal is true;
	signal G28233: std_logic; attribute dont_touch of G28233: signal is true;
	signal G28234: std_logic; attribute dont_touch of G28234: signal is true;
	signal G28235: std_logic; attribute dont_touch of G28235: signal is true;
	signal G28236: std_logic; attribute dont_touch of G28236: signal is true;
	signal G28237: std_logic; attribute dont_touch of G28237: signal is true;
	signal G28238: std_logic; attribute dont_touch of G28238: signal is true;
	signal G28239: std_logic; attribute dont_touch of G28239: signal is true;
	signal G28240: std_logic; attribute dont_touch of G28240: signal is true;
	signal G28241: std_logic; attribute dont_touch of G28241: signal is true;
	signal G28242: std_logic; attribute dont_touch of G28242: signal is true;
	signal G28243: std_logic; attribute dont_touch of G28243: signal is true;
	signal G28244: std_logic; attribute dont_touch of G28244: signal is true;
	signal G28245: std_logic; attribute dont_touch of G28245: signal is true;
	signal G28246: std_logic; attribute dont_touch of G28246: signal is true;
	signal G28247: std_logic; attribute dont_touch of G28247: signal is true;
	signal G28248: std_logic; attribute dont_touch of G28248: signal is true;
	signal G28249: std_logic; attribute dont_touch of G28249: signal is true;
	signal G28250: std_logic; attribute dont_touch of G28250: signal is true;
	signal G28251: std_logic; attribute dont_touch of G28251: signal is true;
	signal G28252: std_logic; attribute dont_touch of G28252: signal is true;
	signal G28253: std_logic; attribute dont_touch of G28253: signal is true;
	signal G28254: std_logic; attribute dont_touch of G28254: signal is true;
	signal G28255: std_logic; attribute dont_touch of G28255: signal is true;
	signal G28256: std_logic; attribute dont_touch of G28256: signal is true;
	signal G28257: std_logic; attribute dont_touch of G28257: signal is true;
	signal G28258: std_logic; attribute dont_touch of G28258: signal is true;
	signal G28259: std_logic; attribute dont_touch of G28259: signal is true;
	signal G28260: std_logic; attribute dont_touch of G28260: signal is true;
	signal G28261: std_logic; attribute dont_touch of G28261: signal is true;
	signal G28262: std_logic; attribute dont_touch of G28262: signal is true;
	signal G28263: std_logic; attribute dont_touch of G28263: signal is true;
	signal G28264: std_logic; attribute dont_touch of G28264: signal is true;
	signal G28265: std_logic; attribute dont_touch of G28265: signal is true;
	signal G28266: std_logic; attribute dont_touch of G28266: signal is true;
	signal G28267: std_logic; attribute dont_touch of G28267: signal is true;
	signal G28268: std_logic; attribute dont_touch of G28268: signal is true;
	signal G28269: std_logic; attribute dont_touch of G28269: signal is true;
	signal G28270: std_logic; attribute dont_touch of G28270: signal is true;
	signal G28271: std_logic; attribute dont_touch of G28271: signal is true;
	signal G28272: std_logic; attribute dont_touch of G28272: signal is true;
	signal G28273: std_logic; attribute dont_touch of G28273: signal is true;
	signal G28274: std_logic; attribute dont_touch of G28274: signal is true;
	signal G28275: std_logic; attribute dont_touch of G28275: signal is true;
	signal G28276: std_logic; attribute dont_touch of G28276: signal is true;
	signal G28277: std_logic; attribute dont_touch of G28277: signal is true;
	signal G28278: std_logic; attribute dont_touch of G28278: signal is true;
	signal G28279: std_logic; attribute dont_touch of G28279: signal is true;
	signal G28280: std_logic; attribute dont_touch of G28280: signal is true;
	signal G28281: std_logic; attribute dont_touch of G28281: signal is true;
	signal G28282: std_logic; attribute dont_touch of G28282: signal is true;
	signal G28283: std_logic; attribute dont_touch of G28283: signal is true;
	signal G28284: std_logic; attribute dont_touch of G28284: signal is true;
	signal G28285: std_logic; attribute dont_touch of G28285: signal is true;
	signal G28286: std_logic; attribute dont_touch of G28286: signal is true;
	signal G28287: std_logic; attribute dont_touch of G28287: signal is true;
	signal G28288: std_logic; attribute dont_touch of G28288: signal is true;
	signal G28289: std_logic; attribute dont_touch of G28289: signal is true;
	signal G28290: std_logic; attribute dont_touch of G28290: signal is true;
	signal G28291: std_logic; attribute dont_touch of G28291: signal is true;
	signal G28292: std_logic; attribute dont_touch of G28292: signal is true;
	signal G28293: std_logic; attribute dont_touch of G28293: signal is true;
	signal G28294: std_logic; attribute dont_touch of G28294: signal is true;
	signal G28295: std_logic; attribute dont_touch of G28295: signal is true;
	signal G28296: std_logic; attribute dont_touch of G28296: signal is true;
	signal G28297: std_logic; attribute dont_touch of G28297: signal is true;
	signal G28298: std_logic; attribute dont_touch of G28298: signal is true;
	signal G28299: std_logic; attribute dont_touch of G28299: signal is true;
	signal G28300: std_logic; attribute dont_touch of G28300: signal is true;
	signal G28301: std_logic; attribute dont_touch of G28301: signal is true;
	signal G28302: std_logic; attribute dont_touch of G28302: signal is true;
	signal G28303: std_logic; attribute dont_touch of G28303: signal is true;
	signal G28304: std_logic; attribute dont_touch of G28304: signal is true;
	signal G28305: std_logic; attribute dont_touch of G28305: signal is true;
	signal G28306: std_logic; attribute dont_touch of G28306: signal is true;
	signal G28307: std_logic; attribute dont_touch of G28307: signal is true;
	signal G28308: std_logic; attribute dont_touch of G28308: signal is true;
	signal G28309: std_logic; attribute dont_touch of G28309: signal is true;
	signal G28310: std_logic; attribute dont_touch of G28310: signal is true;
	signal G28311: std_logic; attribute dont_touch of G28311: signal is true;
	signal G28312: std_logic; attribute dont_touch of G28312: signal is true;
	signal G28313: std_logic; attribute dont_touch of G28313: signal is true;
	signal G28314: std_logic; attribute dont_touch of G28314: signal is true;
	signal G28315: std_logic; attribute dont_touch of G28315: signal is true;
	signal G28316: std_logic; attribute dont_touch of G28316: signal is true;
	signal G28317: std_logic; attribute dont_touch of G28317: signal is true;
	signal G28318: std_logic; attribute dont_touch of G28318: signal is true;
	signal G28319: std_logic; attribute dont_touch of G28319: signal is true;
	signal G28320: std_logic; attribute dont_touch of G28320: signal is true;
	signal G28321: std_logic; attribute dont_touch of G28321: signal is true;
	signal G28322: std_logic; attribute dont_touch of G28322: signal is true;
	signal G28323: std_logic; attribute dont_touch of G28323: signal is true;
	signal G28324: std_logic; attribute dont_touch of G28324: signal is true;
	signal G28325: std_logic; attribute dont_touch of G28325: signal is true;
	signal G28326: std_logic; attribute dont_touch of G28326: signal is true;
	signal G28327: std_logic; attribute dont_touch of G28327: signal is true;
	signal G28328: std_logic; attribute dont_touch of G28328: signal is true;
	signal G28329: std_logic; attribute dont_touch of G28329: signal is true;
	signal G28330: std_logic; attribute dont_touch of G28330: signal is true;
	signal G28331: std_logic; attribute dont_touch of G28331: signal is true;
	signal G28332: std_logic; attribute dont_touch of G28332: signal is true;
	signal G28333: std_logic; attribute dont_touch of G28333: signal is true;
	signal G28334: std_logic; attribute dont_touch of G28334: signal is true;
	signal G28335: std_logic; attribute dont_touch of G28335: signal is true;
	signal G28336: std_logic; attribute dont_touch of G28336: signal is true;
	signal G28337: std_logic; attribute dont_touch of G28337: signal is true;
	signal G28338: std_logic; attribute dont_touch of G28338: signal is true;
	signal G28339: std_logic; attribute dont_touch of G28339: signal is true;
	signal G28340: std_logic; attribute dont_touch of G28340: signal is true;
	signal G28341: std_logic; attribute dont_touch of G28341: signal is true;
	signal G28342: std_logic; attribute dont_touch of G28342: signal is true;
	signal G28343: std_logic; attribute dont_touch of G28343: signal is true;
	signal G28344: std_logic; attribute dont_touch of G28344: signal is true;
	signal G28345: std_logic; attribute dont_touch of G28345: signal is true;
	signal G28346: std_logic; attribute dont_touch of G28346: signal is true;
	signal G28347: std_logic; attribute dont_touch of G28347: signal is true;
	signal G28348: std_logic; attribute dont_touch of G28348: signal is true;
	signal G28349: std_logic; attribute dont_touch of G28349: signal is true;
	signal G28350: std_logic; attribute dont_touch of G28350: signal is true;
	signal G28351: std_logic; attribute dont_touch of G28351: signal is true;
	signal G28352: std_logic; attribute dont_touch of G28352: signal is true;
	signal G28353: std_logic; attribute dont_touch of G28353: signal is true;
	signal G28354: std_logic; attribute dont_touch of G28354: signal is true;
	signal G28355: std_logic; attribute dont_touch of G28355: signal is true;
	signal G28356: std_logic; attribute dont_touch of G28356: signal is true;
	signal G28357: std_logic; attribute dont_touch of G28357: signal is true;
	signal G28358: std_logic; attribute dont_touch of G28358: signal is true;
	signal G28359: std_logic; attribute dont_touch of G28359: signal is true;
	signal G28360: std_logic; attribute dont_touch of G28360: signal is true;
	signal G28361: std_logic; attribute dont_touch of G28361: signal is true;
	signal G28362: std_logic; attribute dont_touch of G28362: signal is true;
	signal G28363: std_logic; attribute dont_touch of G28363: signal is true;
	signal G28364: std_logic; attribute dont_touch of G28364: signal is true;
	signal G28365: std_logic; attribute dont_touch of G28365: signal is true;
	signal G28366: std_logic; attribute dont_touch of G28366: signal is true;
	signal G28367: std_logic; attribute dont_touch of G28367: signal is true;
	signal G28368: std_logic; attribute dont_touch of G28368: signal is true;
	signal G28369: std_logic; attribute dont_touch of G28369: signal is true;
	signal G28370: std_logic; attribute dont_touch of G28370: signal is true;
	signal G28371: std_logic; attribute dont_touch of G28371: signal is true;
	signal G28372: std_logic; attribute dont_touch of G28372: signal is true;
	signal G28373: std_logic; attribute dont_touch of G28373: signal is true;
	signal G28374: std_logic; attribute dont_touch of G28374: signal is true;
	signal G28375: std_logic; attribute dont_touch of G28375: signal is true;
	signal G28376: std_logic; attribute dont_touch of G28376: signal is true;
	signal G28377: std_logic; attribute dont_touch of G28377: signal is true;
	signal G28378: std_logic; attribute dont_touch of G28378: signal is true;
	signal G28379: std_logic; attribute dont_touch of G28379: signal is true;
	signal G28380: std_logic; attribute dont_touch of G28380: signal is true;
	signal G28381: std_logic; attribute dont_touch of G28381: signal is true;
	signal G28382: std_logic; attribute dont_touch of G28382: signal is true;
	signal G28383: std_logic; attribute dont_touch of G28383: signal is true;
	signal G28384: std_logic; attribute dont_touch of G28384: signal is true;
	signal G28385: std_logic; attribute dont_touch of G28385: signal is true;
	signal G28386: std_logic; attribute dont_touch of G28386: signal is true;
	signal G28387: std_logic; attribute dont_touch of G28387: signal is true;
	signal G28388: std_logic; attribute dont_touch of G28388: signal is true;
	signal G28389: std_logic; attribute dont_touch of G28389: signal is true;
	signal G28390: std_logic; attribute dont_touch of G28390: signal is true;
	signal G28391: std_logic; attribute dont_touch of G28391: signal is true;
	signal G28392: std_logic; attribute dont_touch of G28392: signal is true;
	signal G28393: std_logic; attribute dont_touch of G28393: signal is true;
	signal G28394: std_logic; attribute dont_touch of G28394: signal is true;
	signal G28395: std_logic; attribute dont_touch of G28395: signal is true;
	signal G28396: std_logic; attribute dont_touch of G28396: signal is true;
	signal G28397: std_logic; attribute dont_touch of G28397: signal is true;
	signal G28398: std_logic; attribute dont_touch of G28398: signal is true;
	signal G28399: std_logic; attribute dont_touch of G28399: signal is true;
	signal G28400: std_logic; attribute dont_touch of G28400: signal is true;
	signal G28401: std_logic; attribute dont_touch of G28401: signal is true;
	signal G28402: std_logic; attribute dont_touch of G28402: signal is true;
	signal G28403: std_logic; attribute dont_touch of G28403: signal is true;
	signal G28404: std_logic; attribute dont_touch of G28404: signal is true;
	signal G28405: std_logic; attribute dont_touch of G28405: signal is true;
	signal G28406: std_logic; attribute dont_touch of G28406: signal is true;
	signal G28407: std_logic; attribute dont_touch of G28407: signal is true;
	signal G28408: std_logic; attribute dont_touch of G28408: signal is true;
	signal G28409: std_logic; attribute dont_touch of G28409: signal is true;
	signal G28410: std_logic; attribute dont_touch of G28410: signal is true;
	signal G28411: std_logic; attribute dont_touch of G28411: signal is true;
	signal G28412: std_logic; attribute dont_touch of G28412: signal is true;
	signal G28413: std_logic; attribute dont_touch of G28413: signal is true;
	signal G28414: std_logic; attribute dont_touch of G28414: signal is true;
	signal G28415: std_logic; attribute dont_touch of G28415: signal is true;
	signal G28416: std_logic; attribute dont_touch of G28416: signal is true;
	signal G28417: std_logic; attribute dont_touch of G28417: signal is true;
	signal G28418: std_logic; attribute dont_touch of G28418: signal is true;
	signal G28419: std_logic; attribute dont_touch of G28419: signal is true;
	signal G28420: std_logic; attribute dont_touch of G28420: signal is true;
	signal G28421: std_logic; attribute dont_touch of G28421: signal is true;
	signal G28422: std_logic; attribute dont_touch of G28422: signal is true;
	signal G28423: std_logic; attribute dont_touch of G28423: signal is true;
	signal G28424: std_logic; attribute dont_touch of G28424: signal is true;
	signal G28425: std_logic; attribute dont_touch of G28425: signal is true;
	signal G28426: std_logic; attribute dont_touch of G28426: signal is true;
	signal G28427: std_logic; attribute dont_touch of G28427: signal is true;
	signal G28428: std_logic; attribute dont_touch of G28428: signal is true;
	signal G28429: std_logic; attribute dont_touch of G28429: signal is true;
	signal G28430: std_logic; attribute dont_touch of G28430: signal is true;
	signal G28431: std_logic; attribute dont_touch of G28431: signal is true;
	signal G28432: std_logic; attribute dont_touch of G28432: signal is true;
	signal G28433: std_logic; attribute dont_touch of G28433: signal is true;
	signal G28434: std_logic; attribute dont_touch of G28434: signal is true;
	signal G28435: std_logic; attribute dont_touch of G28435: signal is true;
	signal G28436: std_logic; attribute dont_touch of G28436: signal is true;
	signal G28437: std_logic; attribute dont_touch of G28437: signal is true;
	signal G28438: std_logic; attribute dont_touch of G28438: signal is true;
	signal G28439: std_logic; attribute dont_touch of G28439: signal is true;
	signal G28440: std_logic; attribute dont_touch of G28440: signal is true;
	signal G28441: std_logic; attribute dont_touch of G28441: signal is true;
	signal G28442: std_logic; attribute dont_touch of G28442: signal is true;
	signal G28443: std_logic; attribute dont_touch of G28443: signal is true;
	signal G28444: std_logic; attribute dont_touch of G28444: signal is true;
	signal G28445: std_logic; attribute dont_touch of G28445: signal is true;
	signal G28446: std_logic; attribute dont_touch of G28446: signal is true;
	signal G28447: std_logic; attribute dont_touch of G28447: signal is true;
	signal G28448: std_logic; attribute dont_touch of G28448: signal is true;
	signal G28449: std_logic; attribute dont_touch of G28449: signal is true;
	signal G28450: std_logic; attribute dont_touch of G28450: signal is true;
	signal G28451: std_logic; attribute dont_touch of G28451: signal is true;
	signal G28452: std_logic; attribute dont_touch of G28452: signal is true;
	signal G28453: std_logic; attribute dont_touch of G28453: signal is true;
	signal G28454: std_logic; attribute dont_touch of G28454: signal is true;
	signal G28455: std_logic; attribute dont_touch of G28455: signal is true;
	signal G28456: std_logic; attribute dont_touch of G28456: signal is true;
	signal G28457: std_logic; attribute dont_touch of G28457: signal is true;
	signal G28458: std_logic; attribute dont_touch of G28458: signal is true;
	signal G28459: std_logic; attribute dont_touch of G28459: signal is true;
	signal G28460: std_logic; attribute dont_touch of G28460: signal is true;
	signal G28461: std_logic; attribute dont_touch of G28461: signal is true;
	signal G28462: std_logic; attribute dont_touch of G28462: signal is true;
	signal G28463: std_logic; attribute dont_touch of G28463: signal is true;
	signal G28464: std_logic; attribute dont_touch of G28464: signal is true;
	signal G28465: std_logic; attribute dont_touch of G28465: signal is true;
	signal G28466: std_logic; attribute dont_touch of G28466: signal is true;
	signal G28467: std_logic; attribute dont_touch of G28467: signal is true;
	signal G28468: std_logic; attribute dont_touch of G28468: signal is true;
	signal G28469: std_logic; attribute dont_touch of G28469: signal is true;
	signal G28470: std_logic; attribute dont_touch of G28470: signal is true;
	signal G28471: std_logic; attribute dont_touch of G28471: signal is true;
	signal G28472: std_logic; attribute dont_touch of G28472: signal is true;
	signal G28473: std_logic; attribute dont_touch of G28473: signal is true;
	signal G28474: std_logic; attribute dont_touch of G28474: signal is true;
	signal G28475: std_logic; attribute dont_touch of G28475: signal is true;
	signal G28476: std_logic; attribute dont_touch of G28476: signal is true;
	signal G28477: std_logic; attribute dont_touch of G28477: signal is true;
	signal G28478: std_logic; attribute dont_touch of G28478: signal is true;
	signal G28479: std_logic; attribute dont_touch of G28479: signal is true;
	signal G28480: std_logic; attribute dont_touch of G28480: signal is true;
	signal G28481: std_logic; attribute dont_touch of G28481: signal is true;
	signal G28482: std_logic; attribute dont_touch of G28482: signal is true;
	signal G28483: std_logic; attribute dont_touch of G28483: signal is true;
	signal G28484: std_logic; attribute dont_touch of G28484: signal is true;
	signal G28485: std_logic; attribute dont_touch of G28485: signal is true;
	signal G28486: std_logic; attribute dont_touch of G28486: signal is true;
	signal G28487: std_logic; attribute dont_touch of G28487: signal is true;
	signal G28488: std_logic; attribute dont_touch of G28488: signal is true;
	signal G28489: std_logic; attribute dont_touch of G28489: signal is true;
	signal G28490: std_logic; attribute dont_touch of G28490: signal is true;
	signal G28491: std_logic; attribute dont_touch of G28491: signal is true;
	signal G28492: std_logic; attribute dont_touch of G28492: signal is true;
	signal G28493: std_logic; attribute dont_touch of G28493: signal is true;
	signal G28494: std_logic; attribute dont_touch of G28494: signal is true;
	signal G28495: std_logic; attribute dont_touch of G28495: signal is true;
	signal G28496: std_logic; attribute dont_touch of G28496: signal is true;
	signal G28497: std_logic; attribute dont_touch of G28497: signal is true;
	signal G28498: std_logic; attribute dont_touch of G28498: signal is true;
	signal G28499: std_logic; attribute dont_touch of G28499: signal is true;
	signal G28500: std_logic; attribute dont_touch of G28500: signal is true;
	signal G28501: std_logic; attribute dont_touch of G28501: signal is true;
	signal G28512: std_logic; attribute dont_touch of G28512: signal is true;
	signal G28523: std_logic; attribute dont_touch of G28523: signal is true;
	signal G28524: std_logic; attribute dont_touch of G28524: signal is true;
	signal G28525: std_logic; attribute dont_touch of G28525: signal is true;
	signal G28526: std_logic; attribute dont_touch of G28526: signal is true;
	signal G28527: std_logic; attribute dont_touch of G28527: signal is true;
	signal G28528: std_logic; attribute dont_touch of G28528: signal is true;
	signal G28529: std_logic; attribute dont_touch of G28529: signal is true;
	signal G28540: std_logic; attribute dont_touch of G28540: signal is true;
	signal G28551: std_logic; attribute dont_touch of G28551: signal is true;
	signal G28552: std_logic; attribute dont_touch of G28552: signal is true;
	signal G28553: std_logic; attribute dont_touch of G28553: signal is true;
	signal G28554: std_logic; attribute dont_touch of G28554: signal is true;
	signal G28555: std_logic; attribute dont_touch of G28555: signal is true;
	signal G28556: std_logic; attribute dont_touch of G28556: signal is true;
	signal G28567: std_logic; attribute dont_touch of G28567: signal is true;
	signal G28578: std_logic; attribute dont_touch of G28578: signal is true;
	signal G28579: std_logic; attribute dont_touch of G28579: signal is true;
	signal G28580: std_logic; attribute dont_touch of G28580: signal is true;
	signal G28581: std_logic; attribute dont_touch of G28581: signal is true;
	signal G28582: std_logic; attribute dont_touch of G28582: signal is true;
	signal G28583: std_logic; attribute dont_touch of G28583: signal is true;
	signal G28584: std_logic; attribute dont_touch of G28584: signal is true;
	signal G28595: std_logic; attribute dont_touch of G28595: signal is true;
	signal G28606: std_logic; attribute dont_touch of G28606: signal is true;
	signal G28607: std_logic; attribute dont_touch of G28607: signal is true;
	signal G28608: std_logic; attribute dont_touch of G28608: signal is true;
	signal G28609: std_logic; attribute dont_touch of G28609: signal is true;
	signal G28610: std_logic; attribute dont_touch of G28610: signal is true;
	signal G28611: std_logic; attribute dont_touch of G28611: signal is true;
	signal G28612: std_logic; attribute dont_touch of G28612: signal is true;
	signal G28616: std_logic; attribute dont_touch of G28616: signal is true;
	signal G28617: std_logic; attribute dont_touch of G28617: signal is true;
	signal G28618: std_logic; attribute dont_touch of G28618: signal is true;
	signal G28619: std_logic; attribute dont_touch of G28619: signal is true;
	signal G28623: std_logic; attribute dont_touch of G28623: signal is true;
	signal G28624: std_logic; attribute dont_touch of G28624: signal is true;
	signal G28625: std_logic; attribute dont_touch of G28625: signal is true;
	signal G28629: std_logic; attribute dont_touch of G28629: signal is true;
	signal G28630: std_logic; attribute dont_touch of G28630: signal is true;
	signal G28634: std_logic; attribute dont_touch of G28634: signal is true;
	signal G28635: std_logic; attribute dont_touch of G28635: signal is true;
	signal G28636: std_logic; attribute dont_touch of G28636: signal is true;
	signal G28637: std_logic; attribute dont_touch of G28637: signal is true;
	signal G28638: std_logic; attribute dont_touch of G28638: signal is true;
	signal G28639: std_logic; attribute dont_touch of G28639: signal is true;
	signal G28640: std_logic; attribute dont_touch of G28640: signal is true;
	signal G28641: std_logic; attribute dont_touch of G28641: signal is true;
	signal G28642: std_logic; attribute dont_touch of G28642: signal is true;
	signal G28643: std_logic; attribute dont_touch of G28643: signal is true;
	signal G28644: std_logic; attribute dont_touch of G28644: signal is true;
	signal G28645: std_logic; attribute dont_touch of G28645: signal is true;
	signal G28646: std_logic; attribute dont_touch of G28646: signal is true;
	signal G28647: std_logic; attribute dont_touch of G28647: signal is true;
	signal G28648: std_logic; attribute dont_touch of G28648: signal is true;
	signal G28649: std_logic; attribute dont_touch of G28649: signal is true;
	signal G28650: std_logic; attribute dont_touch of G28650: signal is true;
	signal G28651: std_logic; attribute dont_touch of G28651: signal is true;
	signal G28652: std_logic; attribute dont_touch of G28652: signal is true;
	signal G28653: std_logic; attribute dont_touch of G28653: signal is true;
	signal G28654: std_logic; attribute dont_touch of G28654: signal is true;
	signal G28655: std_logic; attribute dont_touch of G28655: signal is true;
	signal G28656: std_logic; attribute dont_touch of G28656: signal is true;
	signal G28657: std_logic; attribute dont_touch of G28657: signal is true;
	signal G28658: std_logic; attribute dont_touch of G28658: signal is true;
	signal G28659: std_logic; attribute dont_touch of G28659: signal is true;
	signal G28660: std_logic; attribute dont_touch of G28660: signal is true;
	signal G28661: std_logic; attribute dont_touch of G28661: signal is true;
	signal G28662: std_logic; attribute dont_touch of G28662: signal is true;
	signal G28663: std_logic; attribute dont_touch of G28663: signal is true;
	signal G28664: std_logic; attribute dont_touch of G28664: signal is true;
	signal G28665: std_logic; attribute dont_touch of G28665: signal is true;
	signal G28666: std_logic; attribute dont_touch of G28666: signal is true;
	signal G28667: std_logic; attribute dont_touch of G28667: signal is true;
	signal G28668: std_logic; attribute dont_touch of G28668: signal is true;
	signal G28669: std_logic; attribute dont_touch of G28669: signal is true;
	signal G28670: std_logic; attribute dont_touch of G28670: signal is true;
	signal G28671: std_logic; attribute dont_touch of G28671: signal is true;
	signal G28672: std_logic; attribute dont_touch of G28672: signal is true;
	signal G28673: std_logic; attribute dont_touch of G28673: signal is true;
	signal G28674: std_logic; attribute dont_touch of G28674: signal is true;
	signal G28675: std_logic; attribute dont_touch of G28675: signal is true;
	signal G28676: std_logic; attribute dont_touch of G28676: signal is true;
	signal G28677: std_logic; attribute dont_touch of G28677: signal is true;
	signal G28678: std_logic; attribute dont_touch of G28678: signal is true;
	signal G28679: std_logic; attribute dont_touch of G28679: signal is true;
	signal G28680: std_logic; attribute dont_touch of G28680: signal is true;
	signal G28681: std_logic; attribute dont_touch of G28681: signal is true;
	signal G28682: std_logic; attribute dont_touch of G28682: signal is true;
	signal G28683: std_logic; attribute dont_touch of G28683: signal is true;
	signal G28684: std_logic; attribute dont_touch of G28684: signal is true;
	signal G28685: std_logic; attribute dont_touch of G28685: signal is true;
	signal G28686: std_logic; attribute dont_touch of G28686: signal is true;
	signal G28687: std_logic; attribute dont_touch of G28687: signal is true;
	signal G28688: std_logic; attribute dont_touch of G28688: signal is true;
	signal G28689: std_logic; attribute dont_touch of G28689: signal is true;
	signal G28690: std_logic; attribute dont_touch of G28690: signal is true;
	signal G28691: std_logic; attribute dont_touch of G28691: signal is true;
	signal G28692: std_logic; attribute dont_touch of G28692: signal is true;
	signal G28693: std_logic; attribute dont_touch of G28693: signal is true;
	signal G28694: std_logic; attribute dont_touch of G28694: signal is true;
	signal G28695: std_logic; attribute dont_touch of G28695: signal is true;
	signal G28696: std_logic; attribute dont_touch of G28696: signal is true;
	signal G28697: std_logic; attribute dont_touch of G28697: signal is true;
	signal G28698: std_logic; attribute dont_touch of G28698: signal is true;
	signal G28699: std_logic; attribute dont_touch of G28699: signal is true;
	signal G28700: std_logic; attribute dont_touch of G28700: signal is true;
	signal G28701: std_logic; attribute dont_touch of G28701: signal is true;
	signal G28702: std_logic; attribute dont_touch of G28702: signal is true;
	signal G28703: std_logic; attribute dont_touch of G28703: signal is true;
	signal G28704: std_logic; attribute dont_touch of G28704: signal is true;
	signal G28705: std_logic; attribute dont_touch of G28705: signal is true;
	signal G28706: std_logic; attribute dont_touch of G28706: signal is true;
	signal G28707: std_logic; attribute dont_touch of G28707: signal is true;
	signal G28708: std_logic; attribute dont_touch of G28708: signal is true;
	signal G28709: std_logic; attribute dont_touch of G28709: signal is true;
	signal G28710: std_logic; attribute dont_touch of G28710: signal is true;
	signal G28711: std_logic; attribute dont_touch of G28711: signal is true;
	signal G28712: std_logic; attribute dont_touch of G28712: signal is true;
	signal G28713: std_logic; attribute dont_touch of G28713: signal is true;
	signal G28714: std_logic; attribute dont_touch of G28714: signal is true;
	signal G28715: std_logic; attribute dont_touch of G28715: signal is true;
	signal G28716: std_logic; attribute dont_touch of G28716: signal is true;
	signal G28717: std_logic; attribute dont_touch of G28717: signal is true;
	signal G28718: std_logic; attribute dont_touch of G28718: signal is true;
	signal G28719: std_logic; attribute dont_touch of G28719: signal is true;
	signal G28720: std_logic; attribute dont_touch of G28720: signal is true;
	signal G28721: std_logic; attribute dont_touch of G28721: signal is true;
	signal G28722: std_logic; attribute dont_touch of G28722: signal is true;
	signal G28723: std_logic; attribute dont_touch of G28723: signal is true;
	signal G28724: std_logic; attribute dont_touch of G28724: signal is true;
	signal G28725: std_logic; attribute dont_touch of G28725: signal is true;
	signal G28726: std_logic; attribute dont_touch of G28726: signal is true;
	signal G28727: std_logic; attribute dont_touch of G28727: signal is true;
	signal G28728: std_logic; attribute dont_touch of G28728: signal is true;
	signal G28729: std_logic; attribute dont_touch of G28729: signal is true;
	signal G28730: std_logic; attribute dont_touch of G28730: signal is true;
	signal G28731: std_logic; attribute dont_touch of G28731: signal is true;
	signal G28732: std_logic; attribute dont_touch of G28732: signal is true;
	signal G28733: std_logic; attribute dont_touch of G28733: signal is true;
	signal G28734: std_logic; attribute dont_touch of G28734: signal is true;
	signal G28735: std_logic; attribute dont_touch of G28735: signal is true;
	signal G28736: std_logic; attribute dont_touch of G28736: signal is true;
	signal G28737: std_logic; attribute dont_touch of G28737: signal is true;
	signal G28738: std_logic; attribute dont_touch of G28738: signal is true;
	signal G28739: std_logic; attribute dont_touch of G28739: signal is true;
	signal G28740: std_logic; attribute dont_touch of G28740: signal is true;
	signal G28741: std_logic; attribute dont_touch of G28741: signal is true;
	signal G28744: std_logic; attribute dont_touch of G28744: signal is true;
	signal G28745: std_logic; attribute dont_touch of G28745: signal is true;
	signal G28746: std_logic; attribute dont_touch of G28746: signal is true;
	signal G28747: std_logic; attribute dont_touch of G28747: signal is true;
	signal G28748: std_logic; attribute dont_touch of G28748: signal is true;
	signal G28749: std_logic; attribute dont_touch of G28749: signal is true;
	signal G28750: std_logic; attribute dont_touch of G28750: signal is true;
	signal G28751: std_logic; attribute dont_touch of G28751: signal is true;
	signal G28754: std_logic; attribute dont_touch of G28754: signal is true;
	signal G28755: std_logic; attribute dont_touch of G28755: signal is true;
	signal G28758: std_logic; attribute dont_touch of G28758: signal is true;
	signal G28759: std_logic; attribute dont_touch of G28759: signal is true;
	signal G28760: std_logic; attribute dont_touch of G28760: signal is true;
	signal G28761: std_logic; attribute dont_touch of G28761: signal is true;
	signal G28762: std_logic; attribute dont_touch of G28762: signal is true;
	signal G28763: std_logic; attribute dont_touch of G28763: signal is true;
	signal G28764: std_logic; attribute dont_touch of G28764: signal is true;
	signal G28767: std_logic; attribute dont_touch of G28767: signal is true;
	signal G28768: std_logic; attribute dont_touch of G28768: signal is true;
	signal G28771: std_logic; attribute dont_touch of G28771: signal is true;
	signal G28772: std_logic; attribute dont_touch of G28772: signal is true;
	signal G28773: std_logic; attribute dont_touch of G28773: signal is true;
	signal G28774: std_logic; attribute dont_touch of G28774: signal is true;
	signal G28775: std_logic; attribute dont_touch of G28775: signal is true;
	signal G28778: std_logic; attribute dont_touch of G28778: signal is true;
	signal G28779: std_logic; attribute dont_touch of G28779: signal is true;
	signal G28782: std_logic; attribute dont_touch of G28782: signal is true;
	signal G28783: std_logic; attribute dont_touch of G28783: signal is true;
	signal G28784: std_logic; attribute dont_touch of G28784: signal is true;
	signal G28785: std_logic; attribute dont_touch of G28785: signal is true;
	signal G28788: std_logic; attribute dont_touch of G28788: signal is true;
	signal G28789: std_logic; attribute dont_touch of G28789: signal is true;
	signal G28790: std_logic; attribute dont_touch of G28790: signal is true;
	signal G28791: std_logic; attribute dont_touch of G28791: signal is true;
	signal G28794: std_logic; attribute dont_touch of G28794: signal is true;
	signal G28795: std_logic; attribute dont_touch of G28795: signal is true;
	signal G28796: std_logic; attribute dont_touch of G28796: signal is true;
	signal G28799: std_logic; attribute dont_touch of G28799: signal is true;
	signal G28802: std_logic; attribute dont_touch of G28802: signal is true;
	signal G28803: std_logic; attribute dont_touch of G28803: signal is true;
	signal G28804: std_logic; attribute dont_touch of G28804: signal is true;
	signal G28807: std_logic; attribute dont_touch of G28807: signal is true;
	signal G28810: std_logic; attribute dont_touch of G28810: signal is true;
	signal G28813: std_logic; attribute dont_touch of G28813: signal is true;
	signal G28814: std_logic; attribute dont_touch of G28814: signal is true;
	signal G28817: std_logic; attribute dont_touch of G28817: signal is true;
	signal G28820: std_logic; attribute dont_touch of G28820: signal is true;
	signal G28823: std_logic; attribute dont_touch of G28823: signal is true;
	signal G28826: std_logic; attribute dont_touch of G28826: signal is true;
	signal G28829: std_logic; attribute dont_touch of G28829: signal is true;
	signal G28832: std_logic; attribute dont_touch of G28832: signal is true;
	signal G28833: std_logic; attribute dont_touch of G28833: signal is true;
	signal G28834: std_logic; attribute dont_touch of G28834: signal is true;
	signal G28835: std_logic; attribute dont_touch of G28835: signal is true;
	signal G28836: std_logic; attribute dont_touch of G28836: signal is true;
	signal G28837: std_logic; attribute dont_touch of G28837: signal is true;
	signal G28838: std_logic; attribute dont_touch of G28838: signal is true;
	signal G28839: std_logic; attribute dont_touch of G28839: signal is true;
	signal G28840: std_logic; attribute dont_touch of G28840: signal is true;
	signal G28841: std_logic; attribute dont_touch of G28841: signal is true;
	signal G28842: std_logic; attribute dont_touch of G28842: signal is true;
	signal G28843: std_logic; attribute dont_touch of G28843: signal is true;
	signal G28844: std_logic; attribute dont_touch of G28844: signal is true;
	signal G28845: std_logic; attribute dont_touch of G28845: signal is true;
	signal G28846: std_logic; attribute dont_touch of G28846: signal is true;
	signal G28847: std_logic; attribute dont_touch of G28847: signal is true;
	signal G28848: std_logic; attribute dont_touch of G28848: signal is true;
	signal G28849: std_logic; attribute dont_touch of G28849: signal is true;
	signal G28850: std_logic; attribute dont_touch of G28850: signal is true;
	signal G28851: std_logic; attribute dont_touch of G28851: signal is true;
	signal G28852: std_logic; attribute dont_touch of G28852: signal is true;
	signal G28853: std_logic; attribute dont_touch of G28853: signal is true;
	signal G28854: std_logic; attribute dont_touch of G28854: signal is true;
	signal G28855: std_logic; attribute dont_touch of G28855: signal is true;
	signal G28859: std_logic; attribute dont_touch of G28859: signal is true;
	signal G28863: std_logic; attribute dont_touch of G28863: signal is true;
	signal G28867: std_logic; attribute dont_touch of G28867: signal is true;
	signal G28871: std_logic; attribute dont_touch of G28871: signal is true;
	signal G28874: std_logic; attribute dont_touch of G28874: signal is true;
	signal G28877: std_logic; attribute dont_touch of G28877: signal is true;
	signal G28880: std_logic; attribute dont_touch of G28880: signal is true;
	signal G28881: std_logic; attribute dont_touch of G28881: signal is true;
	signal G28882: std_logic; attribute dont_touch of G28882: signal is true;
	signal G28883: std_logic; attribute dont_touch of G28883: signal is true;
	signal G28886: std_logic; attribute dont_touch of G28886: signal is true;
	signal G28889: std_logic; attribute dont_touch of G28889: signal is true;
	signal G28892: std_logic; attribute dont_touch of G28892: signal is true;
	signal G28893: std_logic; attribute dont_touch of G28893: signal is true;
	signal G28894: std_logic; attribute dont_touch of G28894: signal is true;
	signal G28897: std_logic; attribute dont_touch of G28897: signal is true;
	signal G28898: std_logic; attribute dont_touch of G28898: signal is true;
	signal G28899: std_logic; attribute dont_touch of G28899: signal is true;
	signal G28900: std_logic; attribute dont_touch of G28900: signal is true;
	signal G28903: std_logic; attribute dont_touch of G28903: signal is true;
	signal G28906: std_logic; attribute dont_touch of G28906: signal is true;
	signal G28909: std_logic; attribute dont_touch of G28909: signal is true;
	signal G28910: std_logic; attribute dont_touch of G28910: signal is true;
	signal G28911: std_logic; attribute dont_touch of G28911: signal is true;
	signal G28914: std_logic; attribute dont_touch of G28914: signal is true;
	signal G28915: std_logic; attribute dont_touch of G28915: signal is true;
	signal G28916: std_logic; attribute dont_touch of G28916: signal is true;
	signal G28919: std_logic; attribute dont_touch of G28919: signal is true;
	signal G28920: std_logic; attribute dont_touch of G28920: signal is true;
	signal G28923: std_logic; attribute dont_touch of G28923: signal is true;
	signal G28924: std_logic; attribute dont_touch of G28924: signal is true;
	signal G28925: std_logic; attribute dont_touch of G28925: signal is true;
	signal G28928: std_logic; attribute dont_touch of G28928: signal is true;
	signal G28931: std_logic; attribute dont_touch of G28931: signal is true;
	signal G28932: std_logic; attribute dont_touch of G28932: signal is true;
	signal G28935: std_logic; attribute dont_touch of G28935: signal is true;
	signal G28936: std_logic; attribute dont_touch of G28936: signal is true;
	signal G28937: std_logic; attribute dont_touch of G28937: signal is true;
	signal G28940: std_logic; attribute dont_touch of G28940: signal is true;
	signal G28941: std_logic; attribute dont_touch of G28941: signal is true;
	signal G28944: std_logic; attribute dont_touch of G28944: signal is true;
	signal G28945: std_logic; attribute dont_touch of G28945: signal is true;
	signal G28948: std_logic; attribute dont_touch of G28948: signal is true;
	signal G28949: std_logic; attribute dont_touch of G28949: signal is true;
	signal G28950: std_logic; attribute dont_touch of G28950: signal is true;
	signal G28951: std_logic; attribute dont_touch of G28951: signal is true;
	signal G28954: std_logic; attribute dont_touch of G28954: signal is true;
	signal G28955: std_logic; attribute dont_touch of G28955: signal is true;
	signal G28958: std_logic; attribute dont_touch of G28958: signal is true;
	signal G28959: std_logic; attribute dont_touch of G28959: signal is true;
	signal G28962: std_logic; attribute dont_touch of G28962: signal is true;
	signal G28963: std_logic; attribute dont_touch of G28963: signal is true;
	signal G28966: std_logic; attribute dont_touch of G28966: signal is true;
	signal G28967: std_logic; attribute dont_touch of G28967: signal is true;
	signal G28970: std_logic; attribute dont_touch of G28970: signal is true;
	signal G28971: std_logic; attribute dont_touch of G28971: signal is true;
	signal G28972: std_logic; attribute dont_touch of G28972: signal is true;
	signal G28975: std_logic; attribute dont_touch of G28975: signal is true;
	signal G28978: std_logic; attribute dont_touch of G28978: signal is true;
	signal G28979: std_logic; attribute dont_touch of G28979: signal is true;
	signal G28982: std_logic; attribute dont_touch of G28982: signal is true;
	signal G28983: std_logic; attribute dont_touch of G28983: signal is true;
	signal G28986: std_logic; attribute dont_touch of G28986: signal is true;
	signal G28987: std_logic; attribute dont_touch of G28987: signal is true;
	signal G28990: std_logic; attribute dont_touch of G28990: signal is true;
	signal G28993: std_logic; attribute dont_touch of G28993: signal is true;
	signal G28996: std_logic; attribute dont_touch of G28996: signal is true;
	signal G28997: std_logic; attribute dont_touch of G28997: signal is true;
	signal G28998: std_logic; attribute dont_touch of G28998: signal is true;
	signal G29001: std_logic; attribute dont_touch of G29001: signal is true;
	signal G29002: std_logic; attribute dont_touch of G29002: signal is true;
	signal G29005: std_logic; attribute dont_touch of G29005: signal is true;
	signal G29008: std_logic; attribute dont_touch of G29008: signal is true;
	signal G29009: std_logic; attribute dont_touch of G29009: signal is true;
	signal G29010: std_logic; attribute dont_touch of G29010: signal is true;
	signal G29013: std_logic; attribute dont_touch of G29013: signal is true;
	signal G29016: std_logic; attribute dont_touch of G29016: signal is true;
	signal G29019: std_logic; attribute dont_touch of G29019: signal is true;
	signal G29022: std_logic; attribute dont_touch of G29022: signal is true;
	signal G29023: std_logic; attribute dont_touch of G29023: signal is true;
	signal G29026: std_logic; attribute dont_touch of G29026: signal is true;
	signal G29027: std_logic; attribute dont_touch of G29027: signal is true;
	signal G29030: std_logic; attribute dont_touch of G29030: signal is true;
	signal G29031: std_logic; attribute dont_touch of G29031: signal is true;
	signal G29032: std_logic; attribute dont_touch of G29032: signal is true;
	signal G29035: std_logic; attribute dont_touch of G29035: signal is true;
	signal G29038: std_logic; attribute dont_touch of G29038: signal is true;
	signal G29039: std_logic; attribute dont_touch of G29039: signal is true;
	signal G29042: std_logic; attribute dont_touch of G29042: signal is true;
	signal G29045: std_logic; attribute dont_touch of G29045: signal is true;
	signal G29046: std_logic; attribute dont_touch of G29046: signal is true;
	signal G29049: std_logic; attribute dont_touch of G29049: signal is true;
	signal G29050: std_logic; attribute dont_touch of G29050: signal is true;
	signal G29053: std_logic; attribute dont_touch of G29053: signal is true;
	signal G29054: std_logic; attribute dont_touch of G29054: signal is true;
	signal G29057: std_logic; attribute dont_touch of G29057: signal is true;
	signal G29060: std_logic; attribute dont_touch of G29060: signal is true;
	signal G29061: std_logic; attribute dont_touch of G29061: signal is true;
	signal G29062: std_logic; attribute dont_touch of G29062: signal is true;
	signal G29063: std_logic; attribute dont_touch of G29063: signal is true;
	signal G29064: std_logic; attribute dont_touch of G29064: signal is true;
	signal G29065: std_logic; attribute dont_touch of G29065: signal is true;
	signal G29068: std_logic; attribute dont_touch of G29068: signal is true;
	signal G29069: std_logic; attribute dont_touch of G29069: signal is true;
	signal G29072: std_logic; attribute dont_touch of G29072: signal is true;
	signal G29073: std_logic; attribute dont_touch of G29073: signal is true;
	signal G29074: std_logic; attribute dont_touch of G29074: signal is true;
	signal G29075: std_logic; attribute dont_touch of G29075: signal is true;
	signal G29076: std_logic; attribute dont_touch of G29076: signal is true;
	signal G29077: std_logic; attribute dont_touch of G29077: signal is true;
	signal G29080: std_logic; attribute dont_touch of G29080: signal is true;
	signal G29081: std_logic; attribute dont_touch of G29081: signal is true;
	signal G29082: std_logic; attribute dont_touch of G29082: signal is true;
	signal G29083: std_logic; attribute dont_touch of G29083: signal is true;
	signal G29084: std_logic; attribute dont_touch of G29084: signal is true;
	signal G29085: std_logic; attribute dont_touch of G29085: signal is true;
	signal G29086: std_logic; attribute dont_touch of G29086: signal is true;
	signal G29087: std_logic; attribute dont_touch of G29087: signal is true;
	signal G29088: std_logic; attribute dont_touch of G29088: signal is true;
	signal G29089: std_logic; attribute dont_touch of G29089: signal is true;
	signal G29090: std_logic; attribute dont_touch of G29090: signal is true;
	signal G29091: std_logic; attribute dont_touch of G29091: signal is true;
	signal G29092: std_logic; attribute dont_touch of G29092: signal is true;
	signal G29093: std_logic; attribute dont_touch of G29093: signal is true;
	signal G29094: std_logic; attribute dont_touch of G29094: signal is true;
	signal G29095: std_logic; attribute dont_touch of G29095: signal is true;
	signal G29096: std_logic; attribute dont_touch of G29096: signal is true;
	signal G29097: std_logic; attribute dont_touch of G29097: signal is true;
	signal G29098: std_logic; attribute dont_touch of G29098: signal is true;
	signal G29099: std_logic; attribute dont_touch of G29099: signal is true;
	signal G29100: std_logic; attribute dont_touch of G29100: signal is true;
	signal G29101: std_logic; attribute dont_touch of G29101: signal is true;
	signal G29102: std_logic; attribute dont_touch of G29102: signal is true;
	signal G29103: std_logic; attribute dont_touch of G29103: signal is true;
	signal G29104: std_logic; attribute dont_touch of G29104: signal is true;
	signal G29105: std_logic; attribute dont_touch of G29105: signal is true;
	signal G29106: std_logic; attribute dont_touch of G29106: signal is true;
	signal G29107: std_logic; attribute dont_touch of G29107: signal is true;
	signal G29108: std_logic; attribute dont_touch of G29108: signal is true;
	signal G29109: std_logic; attribute dont_touch of G29109: signal is true;
	signal G29110: std_logic; attribute dont_touch of G29110: signal is true;
	signal G29111: std_logic; attribute dont_touch of G29111: signal is true;
	signal G29112: std_logic; attribute dont_touch of G29112: signal is true;
	signal G29113: std_logic; attribute dont_touch of G29113: signal is true;
	signal G29117: std_logic; attribute dont_touch of G29117: signal is true;
	signal G29118: std_logic; attribute dont_touch of G29118: signal is true;
	signal G29119: std_logic; attribute dont_touch of G29119: signal is true;
	signal G29120: std_logic; attribute dont_touch of G29120: signal is true;
	signal G29126: std_logic; attribute dont_touch of G29126: signal is true;
	signal G29127: std_logic; attribute dont_touch of G29127: signal is true;
	signal G29128: std_logic; attribute dont_touch of G29128: signal is true;
	signal G29129: std_logic; attribute dont_touch of G29129: signal is true;
	signal G29130: std_logic; attribute dont_touch of G29130: signal is true;
	signal G29131: std_logic; attribute dont_touch of G29131: signal is true;
	signal G29132: std_logic; attribute dont_touch of G29132: signal is true;
	signal G29133: std_logic; attribute dont_touch of G29133: signal is true;
	signal G29134: std_logic; attribute dont_touch of G29134: signal is true;
	signal G29135: std_logic; attribute dont_touch of G29135: signal is true;
	signal G29136: std_logic; attribute dont_touch of G29136: signal is true;
	signal G29137: std_logic; attribute dont_touch of G29137: signal is true;
	signal G29138: std_logic; attribute dont_touch of G29138: signal is true;
	signal G29139: std_logic; attribute dont_touch of G29139: signal is true;
	signal G29140: std_logic; attribute dont_touch of G29140: signal is true;
	signal G29141: std_logic; attribute dont_touch of G29141: signal is true;
	signal G29142: std_logic; attribute dont_touch of G29142: signal is true;
	signal G29143: std_logic; attribute dont_touch of G29143: signal is true;
	signal G29144: std_logic; attribute dont_touch of G29144: signal is true;
	signal G29145: std_logic; attribute dont_touch of G29145: signal is true;
	signal G29146: std_logic; attribute dont_touch of G29146: signal is true;
	signal G29147: std_logic; attribute dont_touch of G29147: signal is true;
	signal G29148: std_logic; attribute dont_touch of G29148: signal is true;
	signal G29149: std_logic; attribute dont_touch of G29149: signal is true;
	signal G29150: std_logic; attribute dont_touch of G29150: signal is true;
	signal G29151: std_logic; attribute dont_touch of G29151: signal is true;
	signal G29152: std_logic; attribute dont_touch of G29152: signal is true;
	signal G29153: std_logic; attribute dont_touch of G29153: signal is true;
	signal G29154: std_logic; attribute dont_touch of G29154: signal is true;
	signal G29155: std_logic; attribute dont_touch of G29155: signal is true;
	signal G29156: std_logic; attribute dont_touch of G29156: signal is true;
	signal G29157: std_logic; attribute dont_touch of G29157: signal is true;
	signal G29158: std_logic; attribute dont_touch of G29158: signal is true;
	signal G29159: std_logic; attribute dont_touch of G29159: signal is true;
	signal G29160: std_logic; attribute dont_touch of G29160: signal is true;
	signal G29161: std_logic; attribute dont_touch of G29161: signal is true;
	signal G29162: std_logic; attribute dont_touch of G29162: signal is true;
	signal G29163: std_logic; attribute dont_touch of G29163: signal is true;
	signal G29164: std_logic; attribute dont_touch of G29164: signal is true;
	signal G29165: std_logic; attribute dont_touch of G29165: signal is true;
	signal G29166: std_logic; attribute dont_touch of G29166: signal is true;
	signal G29167: std_logic; attribute dont_touch of G29167: signal is true;
	signal G29168: std_logic; attribute dont_touch of G29168: signal is true;
	signal G29169: std_logic; attribute dont_touch of G29169: signal is true;
	signal G29170: std_logic; attribute dont_touch of G29170: signal is true;
	signal G29171: std_logic; attribute dont_touch of G29171: signal is true;
	signal G29172: std_logic; attribute dont_touch of G29172: signal is true;
	signal G29173: std_logic; attribute dont_touch of G29173: signal is true;
	signal G29174: std_logic; attribute dont_touch of G29174: signal is true;
	signal G29175: std_logic; attribute dont_touch of G29175: signal is true;
	signal G29176: std_logic; attribute dont_touch of G29176: signal is true;
	signal G29177: std_logic; attribute dont_touch of G29177: signal is true;
	signal G29178: std_logic; attribute dont_touch of G29178: signal is true;
	signal G29179: std_logic; attribute dont_touch of G29179: signal is true;
	signal G29180: std_logic; attribute dont_touch of G29180: signal is true;
	signal G29181: std_logic; attribute dont_touch of G29181: signal is true;
	signal G29182: std_logic; attribute dont_touch of G29182: signal is true;
	signal G29183: std_logic; attribute dont_touch of G29183: signal is true;
	signal G29184: std_logic; attribute dont_touch of G29184: signal is true;
	signal G29185: std_logic; attribute dont_touch of G29185: signal is true;
	signal G29186: std_logic; attribute dont_touch of G29186: signal is true;
	signal G29187: std_logic; attribute dont_touch of G29187: signal is true;
	signal G29188: std_logic; attribute dont_touch of G29188: signal is true;
	signal G29189: std_logic; attribute dont_touch of G29189: signal is true;
	signal G29190: std_logic; attribute dont_touch of G29190: signal is true;
	signal G29191: std_logic; attribute dont_touch of G29191: signal is true;
	signal G29192: std_logic; attribute dont_touch of G29192: signal is true;
	signal G29193: std_logic; attribute dont_touch of G29193: signal is true;
	signal G29194: std_logic; attribute dont_touch of G29194: signal is true;
	signal G29195: std_logic; attribute dont_touch of G29195: signal is true;
	signal G29196: std_logic; attribute dont_touch of G29196: signal is true;
	signal G29197: std_logic; attribute dont_touch of G29197: signal is true;
	signal G29198: std_logic; attribute dont_touch of G29198: signal is true;
	signal G29199: std_logic; attribute dont_touch of G29199: signal is true;
	signal G29200: std_logic; attribute dont_touch of G29200: signal is true;
	signal G29201: std_logic; attribute dont_touch of G29201: signal is true;
	signal G29202: std_logic; attribute dont_touch of G29202: signal is true;
	signal G29203: std_logic; attribute dont_touch of G29203: signal is true;
	signal G29204: std_logic; attribute dont_touch of G29204: signal is true;
	signal G29205: std_logic; attribute dont_touch of G29205: signal is true;
	signal G29206: std_logic; attribute dont_touch of G29206: signal is true;
	signal G29207: std_logic; attribute dont_touch of G29207: signal is true;
	signal G29208: std_logic; attribute dont_touch of G29208: signal is true;
	signal G29209: std_logic; attribute dont_touch of G29209: signal is true;
	signal G29210: std_logic; attribute dont_touch of G29210: signal is true;
	signal G29211: std_logic; attribute dont_touch of G29211: signal is true;
	signal G29212: std_logic; attribute dont_touch of G29212: signal is true;
	signal G29213: std_logic; attribute dont_touch of G29213: signal is true;
	signal G29214: std_logic; attribute dont_touch of G29214: signal is true;
	signal G29215: std_logic; attribute dont_touch of G29215: signal is true;
	signal G29216: std_logic; attribute dont_touch of G29216: signal is true;
	signal G29217: std_logic; attribute dont_touch of G29217: signal is true;
	signal G29218: std_logic; attribute dont_touch of G29218: signal is true;
	signal G29219: std_logic; attribute dont_touch of G29219: signal is true;
	signal G29220: std_logic; attribute dont_touch of G29220: signal is true;
	signal G29221: std_logic; attribute dont_touch of G29221: signal is true;
	signal G29222: std_logic; attribute dont_touch of G29222: signal is true;
	signal G29223: std_logic; attribute dont_touch of G29223: signal is true;
	signal G29224: std_logic; attribute dont_touch of G29224: signal is true;
	signal G29225: std_logic; attribute dont_touch of G29225: signal is true;
	signal G29226: std_logic; attribute dont_touch of G29226: signal is true;
	signal G29227: std_logic; attribute dont_touch of G29227: signal is true;
	signal G29228: std_logic; attribute dont_touch of G29228: signal is true;
	signal G29229: std_logic; attribute dont_touch of G29229: signal is true;
	signal G29230: std_logic; attribute dont_touch of G29230: signal is true;
	signal G29231: std_logic; attribute dont_touch of G29231: signal is true;
	signal G29232: std_logic; attribute dont_touch of G29232: signal is true;
	signal G29233: std_logic; attribute dont_touch of G29233: signal is true;
	signal G29234: std_logic; attribute dont_touch of G29234: signal is true;
	signal G29235: std_logic; attribute dont_touch of G29235: signal is true;
	signal G29236: std_logic; attribute dont_touch of G29236: signal is true;
	signal G29237: std_logic; attribute dont_touch of G29237: signal is true;
	signal G29238: std_logic; attribute dont_touch of G29238: signal is true;
	signal G29239: std_logic; attribute dont_touch of G29239: signal is true;
	signal G29240: std_logic; attribute dont_touch of G29240: signal is true;
	signal G29241: std_logic; attribute dont_touch of G29241: signal is true;
	signal G29242: std_logic; attribute dont_touch of G29242: signal is true;
	signal G29243: std_logic; attribute dont_touch of G29243: signal is true;
	signal G29244: std_logic; attribute dont_touch of G29244: signal is true;
	signal G29245: std_logic; attribute dont_touch of G29245: signal is true;
	signal G29246: std_logic; attribute dont_touch of G29246: signal is true;
	signal G29247: std_logic; attribute dont_touch of G29247: signal is true;
	signal G29248: std_logic; attribute dont_touch of G29248: signal is true;
	signal G29249: std_logic; attribute dont_touch of G29249: signal is true;
	signal G29250: std_logic; attribute dont_touch of G29250: signal is true;
	signal G29251: std_logic; attribute dont_touch of G29251: signal is true;
	signal G29252: std_logic; attribute dont_touch of G29252: signal is true;
	signal G29253: std_logic; attribute dont_touch of G29253: signal is true;
	signal G29254: std_logic; attribute dont_touch of G29254: signal is true;
	signal G29255: std_logic; attribute dont_touch of G29255: signal is true;
	signal G29256: std_logic; attribute dont_touch of G29256: signal is true;
	signal G29257: std_logic; attribute dont_touch of G29257: signal is true;
	signal G29258: std_logic; attribute dont_touch of G29258: signal is true;
	signal G29259: std_logic; attribute dont_touch of G29259: signal is true;
	signal G29260: std_logic; attribute dont_touch of G29260: signal is true;
	signal G29261: std_logic; attribute dont_touch of G29261: signal is true;
	signal G29262: std_logic; attribute dont_touch of G29262: signal is true;
	signal G29263: std_logic; attribute dont_touch of G29263: signal is true;
	signal G29264: std_logic; attribute dont_touch of G29264: signal is true;
	signal G29265: std_logic; attribute dont_touch of G29265: signal is true;
	signal G29266: std_logic; attribute dont_touch of G29266: signal is true;
	signal G29267: std_logic; attribute dont_touch of G29267: signal is true;
	signal G29268: std_logic; attribute dont_touch of G29268: signal is true;
	signal G29269: std_logic; attribute dont_touch of G29269: signal is true;
	signal G29270: std_logic; attribute dont_touch of G29270: signal is true;
	signal G29271: std_logic; attribute dont_touch of G29271: signal is true;
	signal G29272: std_logic; attribute dont_touch of G29272: signal is true;
	signal G29273: std_logic; attribute dont_touch of G29273: signal is true;
	signal G29274: std_logic; attribute dont_touch of G29274: signal is true;
	signal G29275: std_logic; attribute dont_touch of G29275: signal is true;
	signal G29276: std_logic; attribute dont_touch of G29276: signal is true;
	signal G29277: std_logic; attribute dont_touch of G29277: signal is true;
	signal G29278: std_logic; attribute dont_touch of G29278: signal is true;
	signal G29279: std_logic; attribute dont_touch of G29279: signal is true;
	signal G29280: std_logic; attribute dont_touch of G29280: signal is true;
	signal G29281: std_logic; attribute dont_touch of G29281: signal is true;
	signal G29282: std_logic; attribute dont_touch of G29282: signal is true;
	signal G29283: std_logic; attribute dont_touch of G29283: signal is true;
	signal G29284: std_logic; attribute dont_touch of G29284: signal is true;
	signal G29285: std_logic; attribute dont_touch of G29285: signal is true;
	signal G29286: std_logic; attribute dont_touch of G29286: signal is true;
	signal G29287: std_logic; attribute dont_touch of G29287: signal is true;
	signal G29288: std_logic; attribute dont_touch of G29288: signal is true;
	signal G29289: std_logic; attribute dont_touch of G29289: signal is true;
	signal G29290: std_logic; attribute dont_touch of G29290: signal is true;
	signal G29291: std_logic; attribute dont_touch of G29291: signal is true;
	signal G29292: std_logic; attribute dont_touch of G29292: signal is true;
	signal G29293: std_logic; attribute dont_touch of G29293: signal is true;
	signal G29294: std_logic; attribute dont_touch of G29294: signal is true;
	signal G29295: std_logic; attribute dont_touch of G29295: signal is true;
	signal G29296: std_logic; attribute dont_touch of G29296: signal is true;
	signal G29297: std_logic; attribute dont_touch of G29297: signal is true;
	signal G29298: std_logic; attribute dont_touch of G29298: signal is true;
	signal G29299: std_logic; attribute dont_touch of G29299: signal is true;
	signal G29300: std_logic; attribute dont_touch of G29300: signal is true;
	signal G29301: std_logic; attribute dont_touch of G29301: signal is true;
	signal G29302: std_logic; attribute dont_touch of G29302: signal is true;
	signal G29303: std_logic; attribute dont_touch of G29303: signal is true;
	signal G29304: std_logic; attribute dont_touch of G29304: signal is true;
	signal G29305: std_logic; attribute dont_touch of G29305: signal is true;
	signal G29306: std_logic; attribute dont_touch of G29306: signal is true;
	signal G29307: std_logic; attribute dont_touch of G29307: signal is true;
	signal G29308: std_logic; attribute dont_touch of G29308: signal is true;
	signal G29309: std_logic; attribute dont_touch of G29309: signal is true;
	signal G29310: std_logic; attribute dont_touch of G29310: signal is true;
	signal G29311: std_logic; attribute dont_touch of G29311: signal is true;
	signal G29312: std_logic; attribute dont_touch of G29312: signal is true;
	signal G29313: std_logic; attribute dont_touch of G29313: signal is true;
	signal G29314: std_logic; attribute dont_touch of G29314: signal is true;
	signal G29315: std_logic; attribute dont_touch of G29315: signal is true;
	signal G29316: std_logic; attribute dont_touch of G29316: signal is true;
	signal G29317: std_logic; attribute dont_touch of G29317: signal is true;
	signal G29318: std_logic; attribute dont_touch of G29318: signal is true;
	signal G29319: std_logic; attribute dont_touch of G29319: signal is true;
	signal G29320: std_logic; attribute dont_touch of G29320: signal is true;
	signal G29321: std_logic; attribute dont_touch of G29321: signal is true;
	signal G29322: std_logic; attribute dont_touch of G29322: signal is true;
	signal G29323: std_logic; attribute dont_touch of G29323: signal is true;
	signal G29324: std_logic; attribute dont_touch of G29324: signal is true;
	signal G29325: std_logic; attribute dont_touch of G29325: signal is true;
	signal G29326: std_logic; attribute dont_touch of G29326: signal is true;
	signal G29327: std_logic; attribute dont_touch of G29327: signal is true;
	signal G29328: std_logic; attribute dont_touch of G29328: signal is true;
	signal G29329: std_logic; attribute dont_touch of G29329: signal is true;
	signal G29330: std_logic; attribute dont_touch of G29330: signal is true;
	signal G29331: std_logic; attribute dont_touch of G29331: signal is true;
	signal G29332: std_logic; attribute dont_touch of G29332: signal is true;
	signal G29333: std_logic; attribute dont_touch of G29333: signal is true;
	signal G29334: std_logic; attribute dont_touch of G29334: signal is true;
	signal G29335: std_logic; attribute dont_touch of G29335: signal is true;
	signal G29336: std_logic; attribute dont_touch of G29336: signal is true;
	signal G29337: std_logic; attribute dont_touch of G29337: signal is true;
	signal G29338: std_logic; attribute dont_touch of G29338: signal is true;
	signal G29339: std_logic; attribute dont_touch of G29339: signal is true;
	signal G29340: std_logic; attribute dont_touch of G29340: signal is true;
	signal G29341: std_logic; attribute dont_touch of G29341: signal is true;
	signal G29342: std_logic; attribute dont_touch of G29342: signal is true;
	signal G29343: std_logic; attribute dont_touch of G29343: signal is true;
	signal G29344: std_logic; attribute dont_touch of G29344: signal is true;
	signal G29345: std_logic; attribute dont_touch of G29345: signal is true;
	signal G29346: std_logic; attribute dont_touch of G29346: signal is true;
	signal G29347: std_logic; attribute dont_touch of G29347: signal is true;
	signal G29348: std_logic; attribute dont_touch of G29348: signal is true;
	signal G29349: std_logic; attribute dont_touch of G29349: signal is true;
	signal G29350: std_logic; attribute dont_touch of G29350: signal is true;
	signal G29353: std_logic; attribute dont_touch of G29353: signal is true;
	signal G29354: std_logic; attribute dont_touch of G29354: signal is true;
	signal G29355: std_logic; attribute dont_touch of G29355: signal is true;
	signal G29356: std_logic; attribute dont_touch of G29356: signal is true;
	signal G29357: std_logic; attribute dont_touch of G29357: signal is true;
	signal G29358: std_logic; attribute dont_touch of G29358: signal is true;
	signal G29359: std_logic; attribute dont_touch of G29359: signal is true;
	signal G29360: std_logic; attribute dont_touch of G29360: signal is true;
	signal G29361: std_logic; attribute dont_touch of G29361: signal is true;
	signal G29362: std_logic; attribute dont_touch of G29362: signal is true;
	signal G29363: std_logic; attribute dont_touch of G29363: signal is true;
	signal G29364: std_logic; attribute dont_touch of G29364: signal is true;
	signal G29365: std_logic; attribute dont_touch of G29365: signal is true;
	signal G29366: std_logic; attribute dont_touch of G29366: signal is true;
	signal G29367: std_logic; attribute dont_touch of G29367: signal is true;
	signal G29368: std_logic; attribute dont_touch of G29368: signal is true;
	signal G29369: std_logic; attribute dont_touch of G29369: signal is true;
	signal G29370: std_logic; attribute dont_touch of G29370: signal is true;
	signal G29371: std_logic; attribute dont_touch of G29371: signal is true;
	signal G29372: std_logic; attribute dont_touch of G29372: signal is true;
	signal G29373: std_logic; attribute dont_touch of G29373: signal is true;
	signal G29374: std_logic; attribute dont_touch of G29374: signal is true;
	signal G29375: std_logic; attribute dont_touch of G29375: signal is true;
	signal G29376: std_logic; attribute dont_touch of G29376: signal is true;
	signal G29377: std_logic; attribute dont_touch of G29377: signal is true;
	signal G29378: std_logic; attribute dont_touch of G29378: signal is true;
	signal G29379: std_logic; attribute dont_touch of G29379: signal is true;
	signal G29380: std_logic; attribute dont_touch of G29380: signal is true;
	signal G29381: std_logic; attribute dont_touch of G29381: signal is true;
	signal G29382: std_logic; attribute dont_touch of G29382: signal is true;
	signal G29383: std_logic; attribute dont_touch of G29383: signal is true;
	signal G29384: std_logic; attribute dont_touch of G29384: signal is true;
	signal G29385: std_logic; attribute dont_touch of G29385: signal is true;
	signal G29386: std_logic; attribute dont_touch of G29386: signal is true;
	signal G29387: std_logic; attribute dont_touch of G29387: signal is true;
	signal G29388: std_logic; attribute dont_touch of G29388: signal is true;
	signal G29389: std_logic; attribute dont_touch of G29389: signal is true;
	signal G29390: std_logic; attribute dont_touch of G29390: signal is true;
	signal G29391: std_logic; attribute dont_touch of G29391: signal is true;
	signal G29392: std_logic; attribute dont_touch of G29392: signal is true;
	signal G29393: std_logic; attribute dont_touch of G29393: signal is true;
	signal G29394: std_logic; attribute dont_touch of G29394: signal is true;
	signal G29395: std_logic; attribute dont_touch of G29395: signal is true;
	signal G29396: std_logic; attribute dont_touch of G29396: signal is true;
	signal G29397: std_logic; attribute dont_touch of G29397: signal is true;
	signal G29398: std_logic; attribute dont_touch of G29398: signal is true;
	signal G29399: std_logic; attribute dont_touch of G29399: signal is true;
	signal G29400: std_logic; attribute dont_touch of G29400: signal is true;
	signal G29401: std_logic; attribute dont_touch of G29401: signal is true;
	signal G29402: std_logic; attribute dont_touch of G29402: signal is true;
	signal G29403: std_logic; attribute dont_touch of G29403: signal is true;
	signal G29404: std_logic; attribute dont_touch of G29404: signal is true;
	signal G29405: std_logic; attribute dont_touch of G29405: signal is true;
	signal G29406: std_logic; attribute dont_touch of G29406: signal is true;
	signal G29407: std_logic; attribute dont_touch of G29407: signal is true;
	signal G29408: std_logic; attribute dont_touch of G29408: signal is true;
	signal G29409: std_logic; attribute dont_touch of G29409: signal is true;
	signal G29410: std_logic; attribute dont_touch of G29410: signal is true;
	signal G29411: std_logic; attribute dont_touch of G29411: signal is true;
	signal G29412: std_logic; attribute dont_touch of G29412: signal is true;
	signal G29413: std_logic; attribute dont_touch of G29413: signal is true;
	signal G29414: std_logic; attribute dont_touch of G29414: signal is true;
	signal G29415: std_logic; attribute dont_touch of G29415: signal is true;
	signal G29416: std_logic; attribute dont_touch of G29416: signal is true;
	signal G29417: std_logic; attribute dont_touch of G29417: signal is true;
	signal G29418: std_logic; attribute dont_touch of G29418: signal is true;
	signal G29419: std_logic; attribute dont_touch of G29419: signal is true;
	signal G29420: std_logic; attribute dont_touch of G29420: signal is true;
	signal G29421: std_logic; attribute dont_touch of G29421: signal is true;
	signal G29422: std_logic; attribute dont_touch of G29422: signal is true;
	signal G29423: std_logic; attribute dont_touch of G29423: signal is true;
	signal G29424: std_logic; attribute dont_touch of G29424: signal is true;
	signal G29425: std_logic; attribute dont_touch of G29425: signal is true;
	signal G29426: std_logic; attribute dont_touch of G29426: signal is true;
	signal G29427: std_logic; attribute dont_touch of G29427: signal is true;
	signal G29428: std_logic; attribute dont_touch of G29428: signal is true;
	signal G29429: std_logic; attribute dont_touch of G29429: signal is true;
	signal G29430: std_logic; attribute dont_touch of G29430: signal is true;
	signal G29431: std_logic; attribute dont_touch of G29431: signal is true;
	signal G29432: std_logic; attribute dont_touch of G29432: signal is true;
	signal G29433: std_logic; attribute dont_touch of G29433: signal is true;
	signal G29434: std_logic; attribute dont_touch of G29434: signal is true;
	signal G29435: std_logic; attribute dont_touch of G29435: signal is true;
	signal G29436: std_logic; attribute dont_touch of G29436: signal is true;
	signal G29437: std_logic; attribute dont_touch of G29437: signal is true;
	signal G29438: std_logic; attribute dont_touch of G29438: signal is true;
	signal G29439: std_logic; attribute dont_touch of G29439: signal is true;
	signal G29440: std_logic; attribute dont_touch of G29440: signal is true;
	signal G29441: std_logic; attribute dont_touch of G29441: signal is true;
	signal G29442: std_logic; attribute dont_touch of G29442: signal is true;
	signal G29443: std_logic; attribute dont_touch of G29443: signal is true;
	signal G29444: std_logic; attribute dont_touch of G29444: signal is true;
	signal G29445: std_logic; attribute dont_touch of G29445: signal is true;
	signal G29446: std_logic; attribute dont_touch of G29446: signal is true;
	signal G29447: std_logic; attribute dont_touch of G29447: signal is true;
	signal G29448: std_logic; attribute dont_touch of G29448: signal is true;
	signal G29449: std_logic; attribute dont_touch of G29449: signal is true;
	signal G29450: std_logic; attribute dont_touch of G29450: signal is true;
	signal G29451: std_logic; attribute dont_touch of G29451: signal is true;
	signal G29452: std_logic; attribute dont_touch of G29452: signal is true;
	signal G29453: std_logic; attribute dont_touch of G29453: signal is true;
	signal G29454: std_logic; attribute dont_touch of G29454: signal is true;
	signal G29455: std_logic; attribute dont_touch of G29455: signal is true;
	signal G29456: std_logic; attribute dont_touch of G29456: signal is true;
	signal G29457: std_logic; attribute dont_touch of G29457: signal is true;
	signal G29458: std_logic; attribute dont_touch of G29458: signal is true;
	signal G29459: std_logic; attribute dont_touch of G29459: signal is true;
	signal G29460: std_logic; attribute dont_touch of G29460: signal is true;
	signal G29461: std_logic; attribute dont_touch of G29461: signal is true;
	signal G29462: std_logic; attribute dont_touch of G29462: signal is true;
	signal G29463: std_logic; attribute dont_touch of G29463: signal is true;
	signal G29464: std_logic; attribute dont_touch of G29464: signal is true;
	signal G29465: std_logic; attribute dont_touch of G29465: signal is true;
	signal G29466: std_logic; attribute dont_touch of G29466: signal is true;
	signal G29467: std_logic; attribute dont_touch of G29467: signal is true;
	signal G29468: std_logic; attribute dont_touch of G29468: signal is true;
	signal G29469: std_logic; attribute dont_touch of G29469: signal is true;
	signal G29470: std_logic; attribute dont_touch of G29470: signal is true;
	signal G29471: std_logic; attribute dont_touch of G29471: signal is true;
	signal G29472: std_logic; attribute dont_touch of G29472: signal is true;
	signal G29473: std_logic; attribute dont_touch of G29473: signal is true;
	signal G29474: std_logic; attribute dont_touch of G29474: signal is true;
	signal G29475: std_logic; attribute dont_touch of G29475: signal is true;
	signal G29476: std_logic; attribute dont_touch of G29476: signal is true;
	signal G29477: std_logic; attribute dont_touch of G29477: signal is true;
	signal G29478: std_logic; attribute dont_touch of G29478: signal is true;
	signal G29479: std_logic; attribute dont_touch of G29479: signal is true;
	signal G29480: std_logic; attribute dont_touch of G29480: signal is true;
	signal G29481: std_logic; attribute dont_touch of G29481: signal is true;
	signal G29482: std_logic; attribute dont_touch of G29482: signal is true;
	signal G29483: std_logic; attribute dont_touch of G29483: signal is true;
	signal G29484: std_logic; attribute dont_touch of G29484: signal is true;
	signal G29485: std_logic; attribute dont_touch of G29485: signal is true;
	signal G29486: std_logic; attribute dont_touch of G29486: signal is true;
	signal G29487: std_logic; attribute dont_touch of G29487: signal is true;
	signal G29488: std_logic; attribute dont_touch of G29488: signal is true;
	signal G29489: std_logic; attribute dont_touch of G29489: signal is true;
	signal G29490: std_logic; attribute dont_touch of G29490: signal is true;
	signal G29491: std_logic; attribute dont_touch of G29491: signal is true;
	signal G29495: std_logic; attribute dont_touch of G29495: signal is true;
	signal G29496: std_logic; attribute dont_touch of G29496: signal is true;
	signal G29497: std_logic; attribute dont_touch of G29497: signal is true;
	signal G29498: std_logic; attribute dont_touch of G29498: signal is true;
	signal G29499: std_logic; attribute dont_touch of G29499: signal is true;
	signal G29500: std_logic; attribute dont_touch of G29500: signal is true;
	signal G29501: std_logic; attribute dont_touch of G29501: signal is true;
	signal G29502: std_logic; attribute dont_touch of G29502: signal is true;
	signal G29503: std_logic; attribute dont_touch of G29503: signal is true;
	signal G29504: std_logic; attribute dont_touch of G29504: signal is true;
	signal G29505: std_logic; attribute dont_touch of G29505: signal is true;
	signal G29506: std_logic; attribute dont_touch of G29506: signal is true;
	signal G29507: std_logic; attribute dont_touch of G29507: signal is true;
	signal G29508: std_logic; attribute dont_touch of G29508: signal is true;
	signal G29509: std_logic; attribute dont_touch of G29509: signal is true;
	signal G29510: std_logic; attribute dont_touch of G29510: signal is true;
	signal G29511: std_logic; attribute dont_touch of G29511: signal is true;
	signal G29512: std_logic; attribute dont_touch of G29512: signal is true;
	signal G29513: std_logic; attribute dont_touch of G29513: signal is true;
	signal G29514: std_logic; attribute dont_touch of G29514: signal is true;
	signal G29515: std_logic; attribute dont_touch of G29515: signal is true;
	signal G29516: std_logic; attribute dont_touch of G29516: signal is true;
	signal G29517: std_logic; attribute dont_touch of G29517: signal is true;
	signal G29518: std_logic; attribute dont_touch of G29518: signal is true;
	signal G29519: std_logic; attribute dont_touch of G29519: signal is true;
	signal G29520: std_logic; attribute dont_touch of G29520: signal is true;
	signal G29521: std_logic; attribute dont_touch of G29521: signal is true;
	signal G29522: std_logic; attribute dont_touch of G29522: signal is true;
	signal G29523: std_logic; attribute dont_touch of G29523: signal is true;
	signal G29524: std_logic; attribute dont_touch of G29524: signal is true;
	signal G29525: std_logic; attribute dont_touch of G29525: signal is true;
	signal G29526: std_logic; attribute dont_touch of G29526: signal is true;
	signal G29527: std_logic; attribute dont_touch of G29527: signal is true;
	signal G29528: std_logic; attribute dont_touch of G29528: signal is true;
	signal G29529: std_logic; attribute dont_touch of G29529: signal is true;
	signal G29530: std_logic; attribute dont_touch of G29530: signal is true;
	signal G29531: std_logic; attribute dont_touch of G29531: signal is true;
	signal G29532: std_logic; attribute dont_touch of G29532: signal is true;
	signal G29533: std_logic; attribute dont_touch of G29533: signal is true;
	signal G29534: std_logic; attribute dont_touch of G29534: signal is true;
	signal G29535: std_logic; attribute dont_touch of G29535: signal is true;
	signal G29536: std_logic; attribute dont_touch of G29536: signal is true;
	signal G29537: std_logic; attribute dont_touch of G29537: signal is true;
	signal G29538: std_logic; attribute dont_touch of G29538: signal is true;
	signal G29539: std_logic; attribute dont_touch of G29539: signal is true;
	signal G29540: std_logic; attribute dont_touch of G29540: signal is true;
	signal G29541: std_logic; attribute dont_touch of G29541: signal is true;
	signal G29542: std_logic; attribute dont_touch of G29542: signal is true;
	signal G29543: std_logic; attribute dont_touch of G29543: signal is true;
	signal G29544: std_logic; attribute dont_touch of G29544: signal is true;
	signal G29545: std_logic; attribute dont_touch of G29545: signal is true;
	signal G29546: std_logic; attribute dont_touch of G29546: signal is true;
	signal G29547: std_logic; attribute dont_touch of G29547: signal is true;
	signal G29548: std_logic; attribute dont_touch of G29548: signal is true;
	signal G29549: std_logic; attribute dont_touch of G29549: signal is true;
	signal G29550: std_logic; attribute dont_touch of G29550: signal is true;
	signal G29551: std_logic; attribute dont_touch of G29551: signal is true;
	signal G29552: std_logic; attribute dont_touch of G29552: signal is true;
	signal G29553: std_logic; attribute dont_touch of G29553: signal is true;
	signal G29554: std_logic; attribute dont_touch of G29554: signal is true;
	signal G29555: std_logic; attribute dont_touch of G29555: signal is true;
	signal G29556: std_logic; attribute dont_touch of G29556: signal is true;
	signal G29557: std_logic; attribute dont_touch of G29557: signal is true;
	signal G29558: std_logic; attribute dont_touch of G29558: signal is true;
	signal G29559: std_logic; attribute dont_touch of G29559: signal is true;
	signal G29560: std_logic; attribute dont_touch of G29560: signal is true;
	signal G29561: std_logic; attribute dont_touch of G29561: signal is true;
	signal G29562: std_logic; attribute dont_touch of G29562: signal is true;
	signal G29563: std_logic; attribute dont_touch of G29563: signal is true;
	signal G29564: std_logic; attribute dont_touch of G29564: signal is true;
	signal G29565: std_logic; attribute dont_touch of G29565: signal is true;
	signal G29566: std_logic; attribute dont_touch of G29566: signal is true;
	signal G29567: std_logic; attribute dont_touch of G29567: signal is true;
	signal G29568: std_logic; attribute dont_touch of G29568: signal is true;
	signal G29569: std_logic; attribute dont_touch of G29569: signal is true;
	signal G29570: std_logic; attribute dont_touch of G29570: signal is true;
	signal G29571: std_logic; attribute dont_touch of G29571: signal is true;
	signal G29572: std_logic; attribute dont_touch of G29572: signal is true;
	signal G29573: std_logic; attribute dont_touch of G29573: signal is true;
	signal G29574: std_logic; attribute dont_touch of G29574: signal is true;
	signal G29575: std_logic; attribute dont_touch of G29575: signal is true;
	signal G29576: std_logic; attribute dont_touch of G29576: signal is true;
	signal G29577: std_logic; attribute dont_touch of G29577: signal is true;
	signal G29578: std_logic; attribute dont_touch of G29578: signal is true;
	signal G29579: std_logic; attribute dont_touch of G29579: signal is true;
	signal G29580: std_logic; attribute dont_touch of G29580: signal is true;
	signal G29581: std_logic; attribute dont_touch of G29581: signal is true;
	signal G29582: std_logic; attribute dont_touch of G29582: signal is true;
	signal G29583: std_logic; attribute dont_touch of G29583: signal is true;
	signal G29606: std_logic; attribute dont_touch of G29606: signal is true;
	signal G29607: std_logic; attribute dont_touch of G29607: signal is true;
	signal G29608: std_logic; attribute dont_touch of G29608: signal is true;
	signal G29609: std_logic; attribute dont_touch of G29609: signal is true;
	signal G29610: std_logic; attribute dont_touch of G29610: signal is true;
	signal G29611: std_logic; attribute dont_touch of G29611: signal is true;
	signal G29612: std_logic; attribute dont_touch of G29612: signal is true;
	signal G29613: std_logic; attribute dont_touch of G29613: signal is true;
	signal G29614: std_logic; attribute dont_touch of G29614: signal is true;
	signal G29615: std_logic; attribute dont_touch of G29615: signal is true;
	signal G29616: std_logic; attribute dont_touch of G29616: signal is true;
	signal G29617: std_logic; attribute dont_touch of G29617: signal is true;
	signal G29618: std_logic; attribute dont_touch of G29618: signal is true;
	signal G29619: std_logic; attribute dont_touch of G29619: signal is true;
	signal G29620: std_logic; attribute dont_touch of G29620: signal is true;
	signal G29621: std_logic; attribute dont_touch of G29621: signal is true;
	signal G29622: std_logic; attribute dont_touch of G29622: signal is true;
	signal G29623: std_logic; attribute dont_touch of G29623: signal is true;
	signal G29624: std_logic; attribute dont_touch of G29624: signal is true;
	signal G29625: std_logic; attribute dont_touch of G29625: signal is true;
	signal G29626: std_logic; attribute dont_touch of G29626: signal is true;
	signal G29627: std_logic; attribute dont_touch of G29627: signal is true;
	signal G29628: std_logic; attribute dont_touch of G29628: signal is true;
	signal G29629: std_logic; attribute dont_touch of G29629: signal is true;
	signal G29630: std_logic; attribute dont_touch of G29630: signal is true;
	signal G29631: std_logic; attribute dont_touch of G29631: signal is true;
	signal G29632: std_logic; attribute dont_touch of G29632: signal is true;
	signal G29633: std_logic; attribute dont_touch of G29633: signal is true;
	signal G29634: std_logic; attribute dont_touch of G29634: signal is true;
	signal G29635: std_logic; attribute dont_touch of G29635: signal is true;
	signal G29636: std_logic; attribute dont_touch of G29636: signal is true;
	signal G29637: std_logic; attribute dont_touch of G29637: signal is true;
	signal G29638: std_logic; attribute dont_touch of G29638: signal is true;
	signal G29639: std_logic; attribute dont_touch of G29639: signal is true;
	signal G29640: std_logic; attribute dont_touch of G29640: signal is true;
	signal G29641: std_logic; attribute dont_touch of G29641: signal is true;
	signal G29642: std_logic; attribute dont_touch of G29642: signal is true;
	signal G29643: std_logic; attribute dont_touch of G29643: signal is true;
	signal G29644: std_logic; attribute dont_touch of G29644: signal is true;
	signal G29645: std_logic; attribute dont_touch of G29645: signal is true;
	signal G29646: std_logic; attribute dont_touch of G29646: signal is true;
	signal G29647: std_logic; attribute dont_touch of G29647: signal is true;
	signal G29648: std_logic; attribute dont_touch of G29648: signal is true;
	signal G29649: std_logic; attribute dont_touch of G29649: signal is true;
	signal G29650: std_logic; attribute dont_touch of G29650: signal is true;
	signal G29651: std_logic; attribute dont_touch of G29651: signal is true;
	signal G29652: std_logic; attribute dont_touch of G29652: signal is true;
	signal G29653: std_logic; attribute dont_touch of G29653: signal is true;
	signal G29654: std_logic; attribute dont_touch of G29654: signal is true;
	signal G29655: std_logic; attribute dont_touch of G29655: signal is true;
	signal G29656: std_logic; attribute dont_touch of G29656: signal is true;
	signal G29657: std_logic; attribute dont_touch of G29657: signal is true;
	signal G29658: std_logic; attribute dont_touch of G29658: signal is true;
	signal G29659: std_logic; attribute dont_touch of G29659: signal is true;
	signal G29660: std_logic; attribute dont_touch of G29660: signal is true;
	signal G29661: std_logic; attribute dont_touch of G29661: signal is true;
	signal G29662: std_logic; attribute dont_touch of G29662: signal is true;
	signal G29663: std_logic; attribute dont_touch of G29663: signal is true;
	signal G29664: std_logic; attribute dont_touch of G29664: signal is true;
	signal G29665: std_logic; attribute dont_touch of G29665: signal is true;
	signal G29666: std_logic; attribute dont_touch of G29666: signal is true;
	signal G29667: std_logic; attribute dont_touch of G29667: signal is true;
	signal G29668: std_logic; attribute dont_touch of G29668: signal is true;
	signal G29669: std_logic; attribute dont_touch of G29669: signal is true;
	signal G29670: std_logic; attribute dont_touch of G29670: signal is true;
	signal G29671: std_logic; attribute dont_touch of G29671: signal is true;
	signal G29672: std_logic; attribute dont_touch of G29672: signal is true;
	signal G29673: std_logic; attribute dont_touch of G29673: signal is true;
	signal G29676: std_logic; attribute dont_touch of G29676: signal is true;
	signal G29677: std_logic; attribute dont_touch of G29677: signal is true;
	signal G29678: std_logic; attribute dont_touch of G29678: signal is true;
	signal G29679: std_logic; attribute dont_touch of G29679: signal is true;
	signal G29680: std_logic; attribute dont_touch of G29680: signal is true;
	signal G29681: std_logic; attribute dont_touch of G29681: signal is true;
	signal G29682: std_logic; attribute dont_touch of G29682: signal is true;
	signal G29683: std_logic; attribute dont_touch of G29683: signal is true;
	signal G29684: std_logic; attribute dont_touch of G29684: signal is true;
	signal G29685: std_logic; attribute dont_touch of G29685: signal is true;
	signal G29686: std_logic; attribute dont_touch of G29686: signal is true;
	signal G29687: std_logic; attribute dont_touch of G29687: signal is true;
	signal G29688: std_logic; attribute dont_touch of G29688: signal is true;
	signal G29689: std_logic; attribute dont_touch of G29689: signal is true;
	signal G29690: std_logic; attribute dont_touch of G29690: signal is true;
	signal G29691: std_logic; attribute dont_touch of G29691: signal is true;
	signal G29692: std_logic; attribute dont_touch of G29692: signal is true;
	signal G29693: std_logic; attribute dont_touch of G29693: signal is true;
	signal G29694: std_logic; attribute dont_touch of G29694: signal is true;
	signal G29695: std_logic; attribute dont_touch of G29695: signal is true;
	signal G29696: std_logic; attribute dont_touch of G29696: signal is true;
	signal G29697: std_logic; attribute dont_touch of G29697: signal is true;
	signal G29698: std_logic; attribute dont_touch of G29698: signal is true;
	signal G29699: std_logic; attribute dont_touch of G29699: signal is true;
	signal G29700: std_logic; attribute dont_touch of G29700: signal is true;
	signal G29701: std_logic; attribute dont_touch of G29701: signal is true;
	signal G29702: std_logic; attribute dont_touch of G29702: signal is true;
	signal G29703: std_logic; attribute dont_touch of G29703: signal is true;
	signal G29704: std_logic; attribute dont_touch of G29704: signal is true;
	signal G29705: std_logic; attribute dont_touch of G29705: signal is true;
	signal G29708: std_logic; attribute dont_touch of G29708: signal is true;
	signal G29709: std_logic; attribute dont_touch of G29709: signal is true;
	signal G29710: std_logic; attribute dont_touch of G29710: signal is true;
	signal G29713: std_logic; attribute dont_touch of G29713: signal is true;
	signal G29716: std_logic; attribute dont_touch of G29716: signal is true;
	signal G29717: std_logic; attribute dont_touch of G29717: signal is true;
	signal G29718: std_logic; attribute dont_touch of G29718: signal is true;
	signal G29721: std_logic; attribute dont_touch of G29721: signal is true;
	signal G29724: std_logic; attribute dont_touch of G29724: signal is true;
	signal G29725: std_logic; attribute dont_touch of G29725: signal is true;
	signal G29726: std_logic; attribute dont_touch of G29726: signal is true;
	signal G29727: std_logic; attribute dont_touch of G29727: signal is true;
	signal G29728: std_logic; attribute dont_touch of G29728: signal is true;
	signal G29731: std_logic; attribute dont_touch of G29731: signal is true;
	signal G29732: std_logic; attribute dont_touch of G29732: signal is true;
	signal G29735: std_logic; attribute dont_touch of G29735: signal is true;
	signal G29736: std_logic; attribute dont_touch of G29736: signal is true;
	signal G29739: std_logic; attribute dont_touch of G29739: signal is true;
	signal G29740: std_logic; attribute dont_touch of G29740: signal is true;
	signal G29741: std_logic; attribute dont_touch of G29741: signal is true;
	signal G29744: std_logic; attribute dont_touch of G29744: signal is true;
	signal G29747: std_logic; attribute dont_touch of G29747: signal is true;
	signal G29748: std_logic; attribute dont_touch of G29748: signal is true;
	signal G29751: std_logic; attribute dont_touch of G29751: signal is true;
	signal G29754: std_logic; attribute dont_touch of G29754: signal is true;
	signal G29755: std_logic; attribute dont_touch of G29755: signal is true;
	signal G29756: std_logic; attribute dont_touch of G29756: signal is true;
	signal G29757: std_logic; attribute dont_touch of G29757: signal is true;
	signal G29758: std_logic; attribute dont_touch of G29758: signal is true;
	signal G29759: std_logic; attribute dont_touch of G29759: signal is true;
	signal G29760: std_logic; attribute dont_touch of G29760: signal is true;
	signal G29761: std_logic; attribute dont_touch of G29761: signal is true;
	signal G29762: std_logic; attribute dont_touch of G29762: signal is true;
	signal G29763: std_logic; attribute dont_touch of G29763: signal is true;
	signal G29764: std_logic; attribute dont_touch of G29764: signal is true;
	signal G29765: std_logic; attribute dont_touch of G29765: signal is true;
	signal G29766: std_logic; attribute dont_touch of G29766: signal is true;
	signal G29767: std_logic; attribute dont_touch of G29767: signal is true;
	signal G29768: std_logic; attribute dont_touch of G29768: signal is true;
	signal G29769: std_logic; attribute dont_touch of G29769: signal is true;
	signal G29770: std_logic; attribute dont_touch of G29770: signal is true;
	signal G29771: std_logic; attribute dont_touch of G29771: signal is true;
	signal G29772: std_logic; attribute dont_touch of G29772: signal is true;
	signal G29773: std_logic; attribute dont_touch of G29773: signal is true;
	signal G29774: std_logic; attribute dont_touch of G29774: signal is true;
	signal G29775: std_logic; attribute dont_touch of G29775: signal is true;
	signal G29776: std_logic; attribute dont_touch of G29776: signal is true;
	signal G29777: std_logic; attribute dont_touch of G29777: signal is true;
	signal G29778: std_logic; attribute dont_touch of G29778: signal is true;
	signal G29779: std_logic; attribute dont_touch of G29779: signal is true;
	signal G29780: std_logic; attribute dont_touch of G29780: signal is true;
	signal G29781: std_logic; attribute dont_touch of G29781: signal is true;
	signal G29782: std_logic; attribute dont_touch of G29782: signal is true;
	signal G29783: std_logic; attribute dont_touch of G29783: signal is true;
	signal G29784: std_logic; attribute dont_touch of G29784: signal is true;
	signal G29785: std_logic; attribute dont_touch of G29785: signal is true;
	signal G29786: std_logic; attribute dont_touch of G29786: signal is true;
	signal G29787: std_logic; attribute dont_touch of G29787: signal is true;
	signal G29788: std_logic; attribute dont_touch of G29788: signal is true;
	signal G29789: std_logic; attribute dont_touch of G29789: signal is true;
	signal G29790: std_logic; attribute dont_touch of G29790: signal is true;
	signal G29791: std_logic; attribute dont_touch of G29791: signal is true;
	signal G29792: std_logic; attribute dont_touch of G29792: signal is true;
	signal G29793: std_logic; attribute dont_touch of G29793: signal is true;
	signal G29794: std_logic; attribute dont_touch of G29794: signal is true;
	signal G29795: std_logic; attribute dont_touch of G29795: signal is true;
	signal G29796: std_logic; attribute dont_touch of G29796: signal is true;
	signal G29797: std_logic; attribute dont_touch of G29797: signal is true;
	signal G29798: std_logic; attribute dont_touch of G29798: signal is true;
	signal G29799: std_logic; attribute dont_touch of G29799: signal is true;
	signal G29800: std_logic; attribute dont_touch of G29800: signal is true;
	signal G29801: std_logic; attribute dont_touch of G29801: signal is true;
	signal G29802: std_logic; attribute dont_touch of G29802: signal is true;
	signal G29803: std_logic; attribute dont_touch of G29803: signal is true;
	signal G29804: std_logic; attribute dont_touch of G29804: signal is true;
	signal G29805: std_logic; attribute dont_touch of G29805: signal is true;
	signal G29806: std_logic; attribute dont_touch of G29806: signal is true;
	signal G29807: std_logic; attribute dont_touch of G29807: signal is true;
	signal G29808: std_logic; attribute dont_touch of G29808: signal is true;
	signal G29809: std_logic; attribute dont_touch of G29809: signal is true;
	signal G29810: std_logic; attribute dont_touch of G29810: signal is true;
	signal G29811: std_logic; attribute dont_touch of G29811: signal is true;
	signal G29812: std_logic; attribute dont_touch of G29812: signal is true;
	signal G29813: std_logic; attribute dont_touch of G29813: signal is true;
	signal G29814: std_logic; attribute dont_touch of G29814: signal is true;
	signal G29815: std_logic; attribute dont_touch of G29815: signal is true;
	signal G29816: std_logic; attribute dont_touch of G29816: signal is true;
	signal G29817: std_logic; attribute dont_touch of G29817: signal is true;
	signal G29818: std_logic; attribute dont_touch of G29818: signal is true;
	signal G29819: std_logic; attribute dont_touch of G29819: signal is true;
	signal G29820: std_logic; attribute dont_touch of G29820: signal is true;
	signal G29821: std_logic; attribute dont_touch of G29821: signal is true;
	signal G29822: std_logic; attribute dont_touch of G29822: signal is true;
	signal G29823: std_logic; attribute dont_touch of G29823: signal is true;
	signal G29827: std_logic; attribute dont_touch of G29827: signal is true;
	signal G29828: std_logic; attribute dont_touch of G29828: signal is true;
	signal G29829: std_logic; attribute dont_touch of G29829: signal is true;
	signal G29833: std_logic; attribute dont_touch of G29833: signal is true;
	signal G29834: std_logic; attribute dont_touch of G29834: signal is true;
	signal G29835: std_logic; attribute dont_touch of G29835: signal is true;
	signal G29839: std_logic; attribute dont_touch of G29839: signal is true;
	signal G29840: std_logic; attribute dont_touch of G29840: signal is true;
	signal G29844: std_logic; attribute dont_touch of G29844: signal is true;
	signal G29848: std_logic; attribute dont_touch of G29848: signal is true;
	signal G29849: std_logic; attribute dont_touch of G29849: signal is true;
	signal G29853: std_logic; attribute dont_touch of G29853: signal is true;
	signal G29857: std_logic; attribute dont_touch of G29857: signal is true;
	signal G29861: std_logic; attribute dont_touch of G29861: signal is true;
	signal G29865: std_logic; attribute dont_touch of G29865: signal is true;
	signal G29869: std_logic; attribute dont_touch of G29869: signal is true;
	signal G29873: std_logic; attribute dont_touch of G29873: signal is true;
	signal G29877: std_logic; attribute dont_touch of G29877: signal is true;
	signal G29881: std_logic; attribute dont_touch of G29881: signal is true;
	signal G29885: std_logic; attribute dont_touch of G29885: signal is true;
	signal G29889: std_logic; attribute dont_touch of G29889: signal is true;
	signal G29893: std_logic; attribute dont_touch of G29893: signal is true;
	signal G29897: std_logic; attribute dont_touch of G29897: signal is true;
	signal G29901: std_logic; attribute dont_touch of G29901: signal is true;
	signal G29905: std_logic; attribute dont_touch of G29905: signal is true;
	signal G29909: std_logic; attribute dont_touch of G29909: signal is true;
	signal G29910: std_logic; attribute dont_touch of G29910: signal is true;
	signal G29911: std_logic; attribute dont_touch of G29911: signal is true;
	signal G29912: std_logic; attribute dont_touch of G29912: signal is true;
	signal G29913: std_logic; attribute dont_touch of G29913: signal is true;
	signal G29914: std_logic; attribute dont_touch of G29914: signal is true;
	signal G29915: std_logic; attribute dont_touch of G29915: signal is true;
	signal G29916: std_logic; attribute dont_touch of G29916: signal is true;
	signal G29917: std_logic; attribute dont_touch of G29917: signal is true;
	signal G29918: std_logic; attribute dont_touch of G29918: signal is true;
	signal G29919: std_logic; attribute dont_touch of G29919: signal is true;
	signal G29920: std_logic; attribute dont_touch of G29920: signal is true;
	signal G29921: std_logic; attribute dont_touch of G29921: signal is true;
	signal G29922: std_logic; attribute dont_touch of G29922: signal is true;
	signal G29923: std_logic; attribute dont_touch of G29923: signal is true;
	signal G29924: std_logic; attribute dont_touch of G29924: signal is true;
	signal G29925: std_logic; attribute dont_touch of G29925: signal is true;
	signal G29926: std_logic; attribute dont_touch of G29926: signal is true;
	signal G29927: std_logic; attribute dont_touch of G29927: signal is true;
	signal G29928: std_logic; attribute dont_touch of G29928: signal is true;
	signal G29929: std_logic; attribute dont_touch of G29929: signal is true;
	signal G29930: std_logic; attribute dont_touch of G29930: signal is true;
	signal G29931: std_logic; attribute dont_touch of G29931: signal is true;
	signal G29932: std_logic; attribute dont_touch of G29932: signal is true;
	signal G29933: std_logic; attribute dont_touch of G29933: signal is true;
	signal G29934: std_logic; attribute dont_touch of G29934: signal is true;
	signal G29935: std_logic; attribute dont_touch of G29935: signal is true;
	signal G29936: std_logic; attribute dont_touch of G29936: signal is true;
	signal G29937: std_logic; attribute dont_touch of G29937: signal is true;
	signal G29938: std_logic; attribute dont_touch of G29938: signal is true;
	signal G29939: std_logic; attribute dont_touch of G29939: signal is true;
	signal G29940: std_logic; attribute dont_touch of G29940: signal is true;
	signal G29941: std_logic; attribute dont_touch of G29941: signal is true;
	signal G29942: std_logic; attribute dont_touch of G29942: signal is true;
	signal G29943: std_logic; attribute dont_touch of G29943: signal is true;
	signal G29944: std_logic; attribute dont_touch of G29944: signal is true;
	signal G29945: std_logic; attribute dont_touch of G29945: signal is true;
	signal G29946: std_logic; attribute dont_touch of G29946: signal is true;
	signal G29947: std_logic; attribute dont_touch of G29947: signal is true;
	signal G29948: std_logic; attribute dont_touch of G29948: signal is true;
	signal G29949: std_logic; attribute dont_touch of G29949: signal is true;
	signal G29950: std_logic; attribute dont_touch of G29950: signal is true;
	signal G29951: std_logic; attribute dont_touch of G29951: signal is true;
	signal G29952: std_logic; attribute dont_touch of G29952: signal is true;
	signal G29953: std_logic; attribute dont_touch of G29953: signal is true;
	signal G29954: std_logic; attribute dont_touch of G29954: signal is true;
	signal G29955: std_logic; attribute dont_touch of G29955: signal is true;
	signal G29956: std_logic; attribute dont_touch of G29956: signal is true;
	signal G29957: std_logic; attribute dont_touch of G29957: signal is true;
	signal G29958: std_logic; attribute dont_touch of G29958: signal is true;
	signal G29959: std_logic; attribute dont_touch of G29959: signal is true;
	signal G29960: std_logic; attribute dont_touch of G29960: signal is true;
	signal G29961: std_logic; attribute dont_touch of G29961: signal is true;
	signal G29962: std_logic; attribute dont_touch of G29962: signal is true;
	signal G29963: std_logic; attribute dont_touch of G29963: signal is true;
	signal G29964: std_logic; attribute dont_touch of G29964: signal is true;
	signal G29965: std_logic; attribute dont_touch of G29965: signal is true;
	signal G29966: std_logic; attribute dont_touch of G29966: signal is true;
	signal G29967: std_logic; attribute dont_touch of G29967: signal is true;
	signal G29968: std_logic; attribute dont_touch of G29968: signal is true;
	signal G29969: std_logic; attribute dont_touch of G29969: signal is true;
	signal G29970: std_logic; attribute dont_touch of G29970: signal is true;
	signal G29971: std_logic; attribute dont_touch of G29971: signal is true;
	signal G29972: std_logic; attribute dont_touch of G29972: signal is true;
	signal G29973: std_logic; attribute dont_touch of G29973: signal is true;
	signal G29974: std_logic; attribute dont_touch of G29974: signal is true;
	signal G29975: std_logic; attribute dont_touch of G29975: signal is true;
	signal G29976: std_logic; attribute dont_touch of G29976: signal is true;
	signal G29977: std_logic; attribute dont_touch of G29977: signal is true;
	signal G29978: std_logic; attribute dont_touch of G29978: signal is true;
	signal G29979: std_logic; attribute dont_touch of G29979: signal is true;
	signal G29980: std_logic; attribute dont_touch of G29980: signal is true;
	signal G29981: std_logic; attribute dont_touch of G29981: signal is true;
	signal G29982: std_logic; attribute dont_touch of G29982: signal is true;
	signal G29983: std_logic; attribute dont_touch of G29983: signal is true;
	signal G29984: std_logic; attribute dont_touch of G29984: signal is true;
	signal G29985: std_logic; attribute dont_touch of G29985: signal is true;
	signal G29986: std_logic; attribute dont_touch of G29986: signal is true;
	signal G29987: std_logic; attribute dont_touch of G29987: signal is true;
	signal G29988: std_logic; attribute dont_touch of G29988: signal is true;
	signal G29989: std_logic; attribute dont_touch of G29989: signal is true;
	signal G29990: std_logic; attribute dont_touch of G29990: signal is true;
	signal G29991: std_logic; attribute dont_touch of G29991: signal is true;
	signal G29992: std_logic; attribute dont_touch of G29992: signal is true;
	signal G29993: std_logic; attribute dont_touch of G29993: signal is true;
	signal G29994: std_logic; attribute dont_touch of G29994: signal is true;
	signal G29995: std_logic; attribute dont_touch of G29995: signal is true;
	signal G29996: std_logic; attribute dont_touch of G29996: signal is true;
	signal G29997: std_logic; attribute dont_touch of G29997: signal is true;
	signal G29998: std_logic; attribute dont_touch of G29998: signal is true;
	signal G29999: std_logic; attribute dont_touch of G29999: signal is true;
	signal G30000: std_logic; attribute dont_touch of G30000: signal is true;
	signal G30001: std_logic; attribute dont_touch of G30001: signal is true;
	signal G30002: std_logic; attribute dont_touch of G30002: signal is true;
	signal G30003: std_logic; attribute dont_touch of G30003: signal is true;
	signal G30004: std_logic; attribute dont_touch of G30004: signal is true;
	signal G30005: std_logic; attribute dont_touch of G30005: signal is true;
	signal G30006: std_logic; attribute dont_touch of G30006: signal is true;
	signal G30007: std_logic; attribute dont_touch of G30007: signal is true;
	signal G30008: std_logic; attribute dont_touch of G30008: signal is true;
	signal G30009: std_logic; attribute dont_touch of G30009: signal is true;
	signal G30010: std_logic; attribute dont_touch of G30010: signal is true;
	signal G30011: std_logic; attribute dont_touch of G30011: signal is true;
	signal G30012: std_logic; attribute dont_touch of G30012: signal is true;
	signal G30013: std_logic; attribute dont_touch of G30013: signal is true;
	signal G30014: std_logic; attribute dont_touch of G30014: signal is true;
	signal G30015: std_logic; attribute dont_touch of G30015: signal is true;
	signal G30016: std_logic; attribute dont_touch of G30016: signal is true;
	signal G30017: std_logic; attribute dont_touch of G30017: signal is true;
	signal G30018: std_logic; attribute dont_touch of G30018: signal is true;
	signal G30019: std_logic; attribute dont_touch of G30019: signal is true;
	signal G30020: std_logic; attribute dont_touch of G30020: signal is true;
	signal G30021: std_logic; attribute dont_touch of G30021: signal is true;
	signal G30022: std_logic; attribute dont_touch of G30022: signal is true;
	signal G30023: std_logic; attribute dont_touch of G30023: signal is true;
	signal G30024: std_logic; attribute dont_touch of G30024: signal is true;
	signal G30025: std_logic; attribute dont_touch of G30025: signal is true;
	signal G30026: std_logic; attribute dont_touch of G30026: signal is true;
	signal G30027: std_logic; attribute dont_touch of G30027: signal is true;
	signal G30028: std_logic; attribute dont_touch of G30028: signal is true;
	signal G30029: std_logic; attribute dont_touch of G30029: signal is true;
	signal G30030: std_logic; attribute dont_touch of G30030: signal is true;
	signal G30031: std_logic; attribute dont_touch of G30031: signal is true;
	signal G30032: std_logic; attribute dont_touch of G30032: signal is true;
	signal G30033: std_logic; attribute dont_touch of G30033: signal is true;
	signal G30034: std_logic; attribute dont_touch of G30034: signal is true;
	signal G30035: std_logic; attribute dont_touch of G30035: signal is true;
	signal G30036: std_logic; attribute dont_touch of G30036: signal is true;
	signal G30040: std_logic; attribute dont_touch of G30040: signal is true;
	signal G30044: std_logic; attribute dont_touch of G30044: signal is true;
	signal G30048: std_logic; attribute dont_touch of G30048: signal is true;
	signal G30052: std_logic; attribute dont_touch of G30052: signal is true;
	signal G30053: std_logic; attribute dont_touch of G30053: signal is true;
	signal G30054: std_logic; attribute dont_touch of G30054: signal is true;
	signal G30055: std_logic; attribute dont_touch of G30055: signal is true;
	signal G30056: std_logic; attribute dont_touch of G30056: signal is true;
	signal G30057: std_logic; attribute dont_touch of G30057: signal is true;
	signal G30058: std_logic; attribute dont_touch of G30058: signal is true;
	signal G30059: std_logic; attribute dont_touch of G30059: signal is true;
	signal G30060: std_logic; attribute dont_touch of G30060: signal is true;
	signal G30061: std_logic; attribute dont_touch of G30061: signal is true;
	signal G30062: std_logic; attribute dont_touch of G30062: signal is true;
	signal G30063: std_logic; attribute dont_touch of G30063: signal is true;
	signal G30064: std_logic; attribute dont_touch of G30064: signal is true;
	signal G30065: std_logic; attribute dont_touch of G30065: signal is true;
	signal G30066: std_logic; attribute dont_touch of G30066: signal is true;
	signal G30067: std_logic; attribute dont_touch of G30067: signal is true;
	signal G30068: std_logic; attribute dont_touch of G30068: signal is true;
	signal G30069: std_logic; attribute dont_touch of G30069: signal is true;
	signal G30070: std_logic; attribute dont_touch of G30070: signal is true;
	signal G30071: std_logic; attribute dont_touch of G30071: signal is true;
	signal G30072: std_logic; attribute dont_touch of G30072: signal is true;
	signal G30076: std_logic; attribute dont_touch of G30076: signal is true;
	signal G30077: std_logic; attribute dont_touch of G30077: signal is true;
	signal G30078: std_logic; attribute dont_touch of G30078: signal is true;
	signal G30079: std_logic; attribute dont_touch of G30079: signal is true;
	signal G30080: std_logic; attribute dont_touch of G30080: signal is true;
	signal G30081: std_logic; attribute dont_touch of G30081: signal is true;
	signal G30082: std_logic; attribute dont_touch of G30082: signal is true;
	signal G30083: std_logic; attribute dont_touch of G30083: signal is true;
	signal G30084: std_logic; attribute dont_touch of G30084: signal is true;
	signal G30085: std_logic; attribute dont_touch of G30085: signal is true;
	signal G30086: std_logic; attribute dont_touch of G30086: signal is true;
	signal G30087: std_logic; attribute dont_touch of G30087: signal is true;
	signal G30088: std_logic; attribute dont_touch of G30088: signal is true;
	signal G30089: std_logic; attribute dont_touch of G30089: signal is true;
	signal G30090: std_logic; attribute dont_touch of G30090: signal is true;
	signal G30091: std_logic; attribute dont_touch of G30091: signal is true;
	signal G30092: std_logic; attribute dont_touch of G30092: signal is true;
	signal G30093: std_logic; attribute dont_touch of G30093: signal is true;
	signal G30094: std_logic; attribute dont_touch of G30094: signal is true;
	signal G30095: std_logic; attribute dont_touch of G30095: signal is true;
	signal G30096: std_logic; attribute dont_touch of G30096: signal is true;
	signal G30097: std_logic; attribute dont_touch of G30097: signal is true;
	signal G30098: std_logic; attribute dont_touch of G30098: signal is true;
	signal G30099: std_logic; attribute dont_touch of G30099: signal is true;
	signal G30100: std_logic; attribute dont_touch of G30100: signal is true;
	signal G30101: std_logic; attribute dont_touch of G30101: signal is true;
	signal G30102: std_logic; attribute dont_touch of G30102: signal is true;
	signal G30103: std_logic; attribute dont_touch of G30103: signal is true;
	signal G30104: std_logic; attribute dont_touch of G30104: signal is true;
	signal G30105: std_logic; attribute dont_touch of G30105: signal is true;
	signal G30106: std_logic; attribute dont_touch of G30106: signal is true;
	signal G30107: std_logic; attribute dont_touch of G30107: signal is true;
	signal G30108: std_logic; attribute dont_touch of G30108: signal is true;
	signal G30109: std_logic; attribute dont_touch of G30109: signal is true;
	signal G30110: std_logic; attribute dont_touch of G30110: signal is true;
	signal G30111: std_logic; attribute dont_touch of G30111: signal is true;
	signal G30112: std_logic; attribute dont_touch of G30112: signal is true;
	signal G30113: std_logic; attribute dont_touch of G30113: signal is true;
	signal G30114: std_logic; attribute dont_touch of G30114: signal is true;
	signal G30115: std_logic; attribute dont_touch of G30115: signal is true;
	signal G30116: std_logic; attribute dont_touch of G30116: signal is true;
	signal G30117: std_logic; attribute dont_touch of G30117: signal is true;
	signal G30118: std_logic; attribute dont_touch of G30118: signal is true;
	signal G30119: std_logic; attribute dont_touch of G30119: signal is true;
	signal G30120: std_logic; attribute dont_touch of G30120: signal is true;
	signal G30121: std_logic; attribute dont_touch of G30121: signal is true;
	signal G30122: std_logic; attribute dont_touch of G30122: signal is true;
	signal G30123: std_logic; attribute dont_touch of G30123: signal is true;
	signal G30124: std_logic; attribute dont_touch of G30124: signal is true;
	signal G30125: std_logic; attribute dont_touch of G30125: signal is true;
	signal G30126: std_logic; attribute dont_touch of G30126: signal is true;
	signal G30127: std_logic; attribute dont_touch of G30127: signal is true;
	signal G30128: std_logic; attribute dont_touch of G30128: signal is true;
	signal G30129: std_logic; attribute dont_touch of G30129: signal is true;
	signal G30130: std_logic; attribute dont_touch of G30130: signal is true;
	signal G30131: std_logic; attribute dont_touch of G30131: signal is true;
	signal G30132: std_logic; attribute dont_touch of G30132: signal is true;
	signal G30133: std_logic; attribute dont_touch of G30133: signal is true;
	signal G30134: std_logic; attribute dont_touch of G30134: signal is true;
	signal G30138: std_logic; attribute dont_touch of G30138: signal is true;
	signal G30139: std_logic; attribute dont_touch of G30139: signal is true;
	signal G30143: std_logic; attribute dont_touch of G30143: signal is true;
	signal G30147: std_logic; attribute dont_touch of G30147: signal is true;
	signal G30151: std_logic; attribute dont_touch of G30151: signal is true;
	signal G30155: std_logic; attribute dont_touch of G30155: signal is true;
	signal G30159: std_logic; attribute dont_touch of G30159: signal is true;
	signal G30163: std_logic; attribute dont_touch of G30163: signal is true;
	signal G30167: std_logic; attribute dont_touch of G30167: signal is true;
	signal G30171: std_logic; attribute dont_touch of G30171: signal is true;
	signal G30175: std_logic; attribute dont_touch of G30175: signal is true;
	signal G30179: std_logic; attribute dont_touch of G30179: signal is true;
	signal G30183: std_logic; attribute dont_touch of G30183: signal is true;
	signal G30187: std_logic; attribute dont_touch of G30187: signal is true;
	signal G30191: std_logic; attribute dont_touch of G30191: signal is true;
	signal G30195: std_logic; attribute dont_touch of G30195: signal is true;
	signal G30199: std_logic; attribute dont_touch of G30199: signal is true;
	signal G30203: std_logic; attribute dont_touch of G30203: signal is true;
	signal G30207: std_logic; attribute dont_touch of G30207: signal is true;
	signal G30211: std_logic; attribute dont_touch of G30211: signal is true;
	signal G30215: std_logic; attribute dont_touch of G30215: signal is true;
	signal G30216: std_logic; attribute dont_touch of G30216: signal is true;
	signal G30217: std_logic; attribute dont_touch of G30217: signal is true;
	signal G30218: std_logic; attribute dont_touch of G30218: signal is true;
	signal G30219: std_logic; attribute dont_touch of G30219: signal is true;
	signal G30220: std_logic; attribute dont_touch of G30220: signal is true;
	signal G30221: std_logic; attribute dont_touch of G30221: signal is true;
	signal G30222: std_logic; attribute dont_touch of G30222: signal is true;
	signal G30223: std_logic; attribute dont_touch of G30223: signal is true;
	signal G30224: std_logic; attribute dont_touch of G30224: signal is true;
	signal G30225: std_logic; attribute dont_touch of G30225: signal is true;
	signal G30226: std_logic; attribute dont_touch of G30226: signal is true;
	signal G30227: std_logic; attribute dont_touch of G30227: signal is true;
	signal G30228: std_logic; attribute dont_touch of G30228: signal is true;
	signal G30229: std_logic; attribute dont_touch of G30229: signal is true;
	signal G30233: std_logic; attribute dont_touch of G30233: signal is true;
	signal G30237: std_logic; attribute dont_touch of G30237: signal is true;
	signal G30241: std_logic; attribute dont_touch of G30241: signal is true;
	signal G30245: std_logic; attribute dont_touch of G30245: signal is true;
	signal G30246: std_logic; attribute dont_touch of G30246: signal is true;
	signal G30247: std_logic; attribute dont_touch of G30247: signal is true;
	signal G30248: std_logic; attribute dont_touch of G30248: signal is true;
	signal G30249: std_logic; attribute dont_touch of G30249: signal is true;
	signal G30250: std_logic; attribute dont_touch of G30250: signal is true;
	signal G30251: std_logic; attribute dont_touch of G30251: signal is true;
	signal G30252: std_logic; attribute dont_touch of G30252: signal is true;
	signal G30253: std_logic; attribute dont_touch of G30253: signal is true;
	signal G30254: std_logic; attribute dont_touch of G30254: signal is true;
	signal G30255: std_logic; attribute dont_touch of G30255: signal is true;
	signal G30256: std_logic; attribute dont_touch of G30256: signal is true;
	signal G30257: std_logic; attribute dont_touch of G30257: signal is true;
	signal G30258: std_logic; attribute dont_touch of G30258: signal is true;
	signal G30259: std_logic; attribute dont_touch of G30259: signal is true;
	signal G30260: std_logic; attribute dont_touch of G30260: signal is true;
	signal G30261: std_logic; attribute dont_touch of G30261: signal is true;
	signal G30262: std_logic; attribute dont_touch of G30262: signal is true;
	signal G30263: std_logic; attribute dont_touch of G30263: signal is true;
	signal G30264: std_logic; attribute dont_touch of G30264: signal is true;
	signal G30265: std_logic; attribute dont_touch of G30265: signal is true;
	signal G30266: std_logic; attribute dont_touch of G30266: signal is true;
	signal G30267: std_logic; attribute dont_touch of G30267: signal is true;
	signal G30268: std_logic; attribute dont_touch of G30268: signal is true;
	signal G30269: std_logic; attribute dont_touch of G30269: signal is true;
	signal G30270: std_logic; attribute dont_touch of G30270: signal is true;
	signal G30271: std_logic; attribute dont_touch of G30271: signal is true;
	signal G30272: std_logic; attribute dont_touch of G30272: signal is true;
	signal G30273: std_logic; attribute dont_touch of G30273: signal is true;
	signal G30274: std_logic; attribute dont_touch of G30274: signal is true;
	signal G30275: std_logic; attribute dont_touch of G30275: signal is true;
	signal G30276: std_logic; attribute dont_touch of G30276: signal is true;
	signal G30277: std_logic; attribute dont_touch of G30277: signal is true;
	signal G30278: std_logic; attribute dont_touch of G30278: signal is true;
	signal G30279: std_logic; attribute dont_touch of G30279: signal is true;
	signal G30280: std_logic; attribute dont_touch of G30280: signal is true;
	signal G30281: std_logic; attribute dont_touch of G30281: signal is true;
	signal G30282: std_logic; attribute dont_touch of G30282: signal is true;
	signal G30283: std_logic; attribute dont_touch of G30283: signal is true;
	signal G30284: std_logic; attribute dont_touch of G30284: signal is true;
	signal G30285: std_logic; attribute dont_touch of G30285: signal is true;
	signal G30286: std_logic; attribute dont_touch of G30286: signal is true;
	signal G30287: std_logic; attribute dont_touch of G30287: signal is true;
	signal G30288: std_logic; attribute dont_touch of G30288: signal is true;
	signal G30289: std_logic; attribute dont_touch of G30289: signal is true;
	signal G30290: std_logic; attribute dont_touch of G30290: signal is true;
	signal G30291: std_logic; attribute dont_touch of G30291: signal is true;
	signal G30292: std_logic; attribute dont_touch of G30292: signal is true;
	signal G30293: std_logic; attribute dont_touch of G30293: signal is true;
	signal G30294: std_logic; attribute dont_touch of G30294: signal is true;
	signal G30295: std_logic; attribute dont_touch of G30295: signal is true;
	signal G30296: std_logic; attribute dont_touch of G30296: signal is true;
	signal G30297: std_logic; attribute dont_touch of G30297: signal is true;
	signal G30298: std_logic; attribute dont_touch of G30298: signal is true;
	signal G30299: std_logic; attribute dont_touch of G30299: signal is true;
	signal G30300: std_logic; attribute dont_touch of G30300: signal is true;
	signal G30301: std_logic; attribute dont_touch of G30301: signal is true;
	signal G30302: std_logic; attribute dont_touch of G30302: signal is true;
	signal G30303: std_logic; attribute dont_touch of G30303: signal is true;
	signal G30304: std_logic; attribute dont_touch of G30304: signal is true;
	signal G30305: std_logic; attribute dont_touch of G30305: signal is true;
	signal G30306: std_logic; attribute dont_touch of G30306: signal is true;
	signal G30307: std_logic; attribute dont_touch of G30307: signal is true;
	signal G30308: std_logic; attribute dont_touch of G30308: signal is true;
	signal G30309: std_logic; attribute dont_touch of G30309: signal is true;
	signal G30310: std_logic; attribute dont_touch of G30310: signal is true;
	signal G30311: std_logic; attribute dont_touch of G30311: signal is true;
	signal G30312: std_logic; attribute dont_touch of G30312: signal is true;
	signal G30313: std_logic; attribute dont_touch of G30313: signal is true;
	signal G30314: std_logic; attribute dont_touch of G30314: signal is true;
	signal G30315: std_logic; attribute dont_touch of G30315: signal is true;
	signal G30316: std_logic; attribute dont_touch of G30316: signal is true;
	signal G30317: std_logic; attribute dont_touch of G30317: signal is true;
	signal G30318: std_logic; attribute dont_touch of G30318: signal is true;
	signal G30319: std_logic; attribute dont_touch of G30319: signal is true;
	signal G30320: std_logic; attribute dont_touch of G30320: signal is true;
	signal G30321: std_logic; attribute dont_touch of G30321: signal is true;
	signal G30322: std_logic; attribute dont_touch of G30322: signal is true;
	signal G30323: std_logic; attribute dont_touch of G30323: signal is true;
	signal G30324: std_logic; attribute dont_touch of G30324: signal is true;
	signal G30325: std_logic; attribute dont_touch of G30325: signal is true;
	signal G30326: std_logic; attribute dont_touch of G30326: signal is true;
	signal G30327: std_logic; attribute dont_touch of G30327: signal is true;
	signal G30328: std_logic; attribute dont_touch of G30328: signal is true;
	signal G30329: std_logic; attribute dont_touch of G30329: signal is true;
	signal G30330: std_logic; attribute dont_touch of G30330: signal is true;
	signal G30331: std_logic; attribute dont_touch of G30331: signal is true;
	signal G30332: std_logic; attribute dont_touch of G30332: signal is true;
	signal G30333: std_logic; attribute dont_touch of G30333: signal is true;
	signal G30334: std_logic; attribute dont_touch of G30334: signal is true;
	signal G30335: std_logic; attribute dont_touch of G30335: signal is true;
	signal G30336: std_logic; attribute dont_touch of G30336: signal is true;
	signal G30337: std_logic; attribute dont_touch of G30337: signal is true;
	signal G30338: std_logic; attribute dont_touch of G30338: signal is true;
	signal G30339: std_logic; attribute dont_touch of G30339: signal is true;
	signal G30340: std_logic; attribute dont_touch of G30340: signal is true;
	signal G30341: std_logic; attribute dont_touch of G30341: signal is true;
	signal G30342: std_logic; attribute dont_touch of G30342: signal is true;
	signal G30343: std_logic; attribute dont_touch of G30343: signal is true;
	signal G30344: std_logic; attribute dont_touch of G30344: signal is true;
	signal G30345: std_logic; attribute dont_touch of G30345: signal is true;
	signal G30346: std_logic; attribute dont_touch of G30346: signal is true;
	signal G30347: std_logic; attribute dont_touch of G30347: signal is true;
	signal G30348: std_logic; attribute dont_touch of G30348: signal is true;
	signal G30349: std_logic; attribute dont_touch of G30349: signal is true;
	signal G30350: std_logic; attribute dont_touch of G30350: signal is true;
	signal G30351: std_logic; attribute dont_touch of G30351: signal is true;
	signal G30352: std_logic; attribute dont_touch of G30352: signal is true;
	signal G30353: std_logic; attribute dont_touch of G30353: signal is true;
	signal G30354: std_logic; attribute dont_touch of G30354: signal is true;
	signal G30355: std_logic; attribute dont_touch of G30355: signal is true;
	signal G30356: std_logic; attribute dont_touch of G30356: signal is true;
	signal G30357: std_logic; attribute dont_touch of G30357: signal is true;
	signal G30358: std_logic; attribute dont_touch of G30358: signal is true;
	signal G30359: std_logic; attribute dont_touch of G30359: signal is true;
	signal G30360: std_logic; attribute dont_touch of G30360: signal is true;
	signal G30361: std_logic; attribute dont_touch of G30361: signal is true;
	signal G30362: std_logic; attribute dont_touch of G30362: signal is true;
	signal G30363: std_logic; attribute dont_touch of G30363: signal is true;
	signal G30364: std_logic; attribute dont_touch of G30364: signal is true;
	signal G30365: std_logic; attribute dont_touch of G30365: signal is true;
	signal G30366: std_logic; attribute dont_touch of G30366: signal is true;
	signal G30367: std_logic; attribute dont_touch of G30367: signal is true;
	signal G30368: std_logic; attribute dont_touch of G30368: signal is true;
	signal G30369: std_logic; attribute dont_touch of G30369: signal is true;
	signal G30370: std_logic; attribute dont_touch of G30370: signal is true;
	signal G30371: std_logic; attribute dont_touch of G30371: signal is true;
	signal G30372: std_logic; attribute dont_touch of G30372: signal is true;
	signal G30373: std_logic; attribute dont_touch of G30373: signal is true;
	signal G30374: std_logic; attribute dont_touch of G30374: signal is true;
	signal G30375: std_logic; attribute dont_touch of G30375: signal is true;
	signal G30376: std_logic; attribute dont_touch of G30376: signal is true;
	signal G30377: std_logic; attribute dont_touch of G30377: signal is true;
	signal G30378: std_logic; attribute dont_touch of G30378: signal is true;
	signal G30379: std_logic; attribute dont_touch of G30379: signal is true;
	signal G30380: std_logic; attribute dont_touch of G30380: signal is true;
	signal G30381: std_logic; attribute dont_touch of G30381: signal is true;
	signal G30382: std_logic; attribute dont_touch of G30382: signal is true;
	signal G30383: std_logic; attribute dont_touch of G30383: signal is true;
	signal G30387: std_logic; attribute dont_touch of G30387: signal is true;
	signal G30388: std_logic; attribute dont_touch of G30388: signal is true;
	signal G30389: std_logic; attribute dont_touch of G30389: signal is true;
	signal G30390: std_logic; attribute dont_touch of G30390: signal is true;
	signal G30391: std_logic; attribute dont_touch of G30391: signal is true;
	signal G30392: std_logic; attribute dont_touch of G30392: signal is true;
	signal G30393: std_logic; attribute dont_touch of G30393: signal is true;
	signal G30394: std_logic; attribute dont_touch of G30394: signal is true;
	signal G30395: std_logic; attribute dont_touch of G30395: signal is true;
	signal G30396: std_logic; attribute dont_touch of G30396: signal is true;
	signal G30397: std_logic; attribute dont_touch of G30397: signal is true;
	signal G30398: std_logic; attribute dont_touch of G30398: signal is true;
	signal G30399: std_logic; attribute dont_touch of G30399: signal is true;
	signal G30400: std_logic; attribute dont_touch of G30400: signal is true;
	signal G30401: std_logic; attribute dont_touch of G30401: signal is true;
	signal G30402: std_logic; attribute dont_touch of G30402: signal is true;
	signal G30403: std_logic; attribute dont_touch of G30403: signal is true;
	signal G30404: std_logic; attribute dont_touch of G30404: signal is true;
	signal G30405: std_logic; attribute dont_touch of G30405: signal is true;
	signal G30406: std_logic; attribute dont_touch of G30406: signal is true;
	signal G30407: std_logic; attribute dont_touch of G30407: signal is true;
	signal G30408: std_logic; attribute dont_touch of G30408: signal is true;
	signal G30409: std_logic; attribute dont_touch of G30409: signal is true;
	signal G30410: std_logic; attribute dont_touch of G30410: signal is true;
	signal G30411: std_logic; attribute dont_touch of G30411: signal is true;
	signal G30412: std_logic; attribute dont_touch of G30412: signal is true;
	signal G30435: std_logic; attribute dont_touch of G30435: signal is true;
	signal G30436: std_logic; attribute dont_touch of G30436: signal is true;
	signal G30437: std_logic; attribute dont_touch of G30437: signal is true;
	signal G30438: std_logic; attribute dont_touch of G30438: signal is true;
	signal G30439: std_logic; attribute dont_touch of G30439: signal is true;
	signal G30440: std_logic; attribute dont_touch of G30440: signal is true;
	signal G30441: std_logic; attribute dont_touch of G30441: signal is true;
	signal G30442: std_logic; attribute dont_touch of G30442: signal is true;
	signal G30443: std_logic; attribute dont_touch of G30443: signal is true;
	signal G30444: std_logic; attribute dont_touch of G30444: signal is true;
	signal G30445: std_logic; attribute dont_touch of G30445: signal is true;
	signal G30446: std_logic; attribute dont_touch of G30446: signal is true;
	signal G30447: std_logic; attribute dont_touch of G30447: signal is true;
	signal G30448: std_logic; attribute dont_touch of G30448: signal is true;
	signal G30449: std_logic; attribute dont_touch of G30449: signal is true;
	signal G30450: std_logic; attribute dont_touch of G30450: signal is true;
	signal G30451: std_logic; attribute dont_touch of G30451: signal is true;
	signal G30452: std_logic; attribute dont_touch of G30452: signal is true;
	signal G30453: std_logic; attribute dont_touch of G30453: signal is true;
	signal G30454: std_logic; attribute dont_touch of G30454: signal is true;
	signal G30455: std_logic; attribute dont_touch of G30455: signal is true;
	signal G30456: std_logic; attribute dont_touch of G30456: signal is true;
	signal G30457: std_logic; attribute dont_touch of G30457: signal is true;
	signal G30458: std_logic; attribute dont_touch of G30458: signal is true;
	signal G30459: std_logic; attribute dont_touch of G30459: signal is true;
	signal G30460: std_logic; attribute dont_touch of G30460: signal is true;
	signal G30461: std_logic; attribute dont_touch of G30461: signal is true;
	signal G30462: std_logic; attribute dont_touch of G30462: signal is true;
	signal G30463: std_logic; attribute dont_touch of G30463: signal is true;
	signal G30464: std_logic; attribute dont_touch of G30464: signal is true;
	signal G30465: std_logic; attribute dont_touch of G30465: signal is true;
	signal G30466: std_logic; attribute dont_touch of G30466: signal is true;
	signal G30467: std_logic; attribute dont_touch of G30467: signal is true;
	signal G30468: std_logic; attribute dont_touch of G30468: signal is true;
	signal G30469: std_logic; attribute dont_touch of G30469: signal is true;
	signal G30470: std_logic; attribute dont_touch of G30470: signal is true;
	signal G30471: std_logic; attribute dont_touch of G30471: signal is true;
	signal G30472: std_logic; attribute dont_touch of G30472: signal is true;
	signal G30473: std_logic; attribute dont_touch of G30473: signal is true;
	signal G30474: std_logic; attribute dont_touch of G30474: signal is true;
	signal G30475: std_logic; attribute dont_touch of G30475: signal is true;
	signal G30476: std_logic; attribute dont_touch of G30476: signal is true;
	signal G30477: std_logic; attribute dont_touch of G30477: signal is true;
	signal G30478: std_logic; attribute dont_touch of G30478: signal is true;
	signal G30479: std_logic; attribute dont_touch of G30479: signal is true;
	signal G30480: std_logic; attribute dont_touch of G30480: signal is true;
	signal G30481: std_logic; attribute dont_touch of G30481: signal is true;
	signal G30482: std_logic; attribute dont_touch of G30482: signal is true;
	signal G30483: std_logic; attribute dont_touch of G30483: signal is true;
	signal G30484: std_logic; attribute dont_touch of G30484: signal is true;
	signal G30485: std_logic; attribute dont_touch of G30485: signal is true;
	signal G30486: std_logic; attribute dont_touch of G30486: signal is true;
	signal G30487: std_logic; attribute dont_touch of G30487: signal is true;
	signal G30488: std_logic; attribute dont_touch of G30488: signal is true;
	signal G30489: std_logic; attribute dont_touch of G30489: signal is true;
	signal G30490: std_logic; attribute dont_touch of G30490: signal is true;
	signal G30491: std_logic; attribute dont_touch of G30491: signal is true;
	signal G30492: std_logic; attribute dont_touch of G30492: signal is true;
	signal G30493: std_logic; attribute dont_touch of G30493: signal is true;
	signal G30494: std_logic; attribute dont_touch of G30494: signal is true;
	signal G30495: std_logic; attribute dont_touch of G30495: signal is true;
	signal G30496: std_logic; attribute dont_touch of G30496: signal is true;
	signal G30497: std_logic; attribute dont_touch of G30497: signal is true;
	signal G30498: std_logic; attribute dont_touch of G30498: signal is true;
	signal G30499: std_logic; attribute dont_touch of G30499: signal is true;
	signal G30500: std_logic; attribute dont_touch of G30500: signal is true;
	signal G30501: std_logic; attribute dont_touch of G30501: signal is true;
	signal G30502: std_logic; attribute dont_touch of G30502: signal is true;
	signal G30503: std_logic; attribute dont_touch of G30503: signal is true;
	signal G30504: std_logic; attribute dont_touch of G30504: signal is true;
	signal G30505: std_logic; attribute dont_touch of G30505: signal is true;
	signal G30506: std_logic; attribute dont_touch of G30506: signal is true;
	signal G30507: std_logic; attribute dont_touch of G30507: signal is true;
	signal G30508: std_logic; attribute dont_touch of G30508: signal is true;
	signal G30509: std_logic; attribute dont_touch of G30509: signal is true;
	signal G30510: std_logic; attribute dont_touch of G30510: signal is true;
	signal G30511: std_logic; attribute dont_touch of G30511: signal is true;
	signal G30512: std_logic; attribute dont_touch of G30512: signal is true;
	signal G30513: std_logic; attribute dont_touch of G30513: signal is true;
	signal G30514: std_logic; attribute dont_touch of G30514: signal is true;
	signal G30515: std_logic; attribute dont_touch of G30515: signal is true;
	signal G30516: std_logic; attribute dont_touch of G30516: signal is true;
	signal G30517: std_logic; attribute dont_touch of G30517: signal is true;
	signal G30518: std_logic; attribute dont_touch of G30518: signal is true;
	signal G30519: std_logic; attribute dont_touch of G30519: signal is true;
	signal G30520: std_logic; attribute dont_touch of G30520: signal is true;
	signal G30521: std_logic; attribute dont_touch of G30521: signal is true;
	signal G30522: std_logic; attribute dont_touch of G30522: signal is true;
	signal G30523: std_logic; attribute dont_touch of G30523: signal is true;
	signal G30524: std_logic; attribute dont_touch of G30524: signal is true;
	signal G30525: std_logic; attribute dont_touch of G30525: signal is true;
	signal G30526: std_logic; attribute dont_touch of G30526: signal is true;
	signal G30527: std_logic; attribute dont_touch of G30527: signal is true;
	signal G30528: std_logic; attribute dont_touch of G30528: signal is true;
	signal G30529: std_logic; attribute dont_touch of G30529: signal is true;
	signal G30530: std_logic; attribute dont_touch of G30530: signal is true;
	signal G30531: std_logic; attribute dont_touch of G30531: signal is true;
	signal G30532: std_logic; attribute dont_touch of G30532: signal is true;
	signal G30533: std_logic; attribute dont_touch of G30533: signal is true;
	signal G30534: std_logic; attribute dont_touch of G30534: signal is true;
	signal G30535: std_logic; attribute dont_touch of G30535: signal is true;
	signal G30536: std_logic; attribute dont_touch of G30536: signal is true;
	signal G30537: std_logic; attribute dont_touch of G30537: signal is true;
	signal G30538: std_logic; attribute dont_touch of G30538: signal is true;
	signal G30539: std_logic; attribute dont_touch of G30539: signal is true;
	signal G30540: std_logic; attribute dont_touch of G30540: signal is true;
	signal G30541: std_logic; attribute dont_touch of G30541: signal is true;
	signal G30542: std_logic; attribute dont_touch of G30542: signal is true;
	signal G30543: std_logic; attribute dont_touch of G30543: signal is true;
	signal G30544: std_logic; attribute dont_touch of G30544: signal is true;
	signal G30545: std_logic; attribute dont_touch of G30545: signal is true;
	signal G30546: std_logic; attribute dont_touch of G30546: signal is true;
	signal G30547: std_logic; attribute dont_touch of G30547: signal is true;
	signal G30548: std_logic; attribute dont_touch of G30548: signal is true;
	signal G30549: std_logic; attribute dont_touch of G30549: signal is true;
	signal G30550: std_logic; attribute dont_touch of G30550: signal is true;
	signal G30551: std_logic; attribute dont_touch of G30551: signal is true;
	signal G30552: std_logic; attribute dont_touch of G30552: signal is true;
	signal G30553: std_logic; attribute dont_touch of G30553: signal is true;
	signal G30554: std_logic; attribute dont_touch of G30554: signal is true;
	signal G30555: std_logic; attribute dont_touch of G30555: signal is true;
	signal G30556: std_logic; attribute dont_touch of G30556: signal is true;
	signal G30557: std_logic; attribute dont_touch of G30557: signal is true;
	signal G30558: std_logic; attribute dont_touch of G30558: signal is true;
	signal G30559: std_logic; attribute dont_touch of G30559: signal is true;
	signal G30560: std_logic; attribute dont_touch of G30560: signal is true;
	signal G30561: std_logic; attribute dont_touch of G30561: signal is true;
	signal G30562: std_logic; attribute dont_touch of G30562: signal is true;
	signal G30563: std_logic; attribute dont_touch of G30563: signal is true;
	signal G30564: std_logic; attribute dont_touch of G30564: signal is true;
	signal G30565: std_logic; attribute dont_touch of G30565: signal is true;
	signal G30566: std_logic; attribute dont_touch of G30566: signal is true;
	signal G30567: std_logic; attribute dont_touch of G30567: signal is true;
	signal G30568: std_logic; attribute dont_touch of G30568: signal is true;
	signal G30569: std_logic; attribute dont_touch of G30569: signal is true;
	signal G30570: std_logic; attribute dont_touch of G30570: signal is true;
	signal G30571: std_logic; attribute dont_touch of G30571: signal is true;
	signal G30572: std_logic; attribute dont_touch of G30572: signal is true;
	signal G30573: std_logic; attribute dont_touch of G30573: signal is true;
	signal G30574: std_logic; attribute dont_touch of G30574: signal is true;
	signal G30575: std_logic; attribute dont_touch of G30575: signal is true;
	signal G30578: std_logic; attribute dont_touch of G30578: signal is true;
	signal G30579: std_logic; attribute dont_touch of G30579: signal is true;
	signal G30580: std_logic; attribute dont_touch of G30580: signal is true;
	signal G30581: std_logic; attribute dont_touch of G30581: signal is true;
	signal G30582: std_logic; attribute dont_touch of G30582: signal is true;
	signal G30583: std_logic; attribute dont_touch of G30583: signal is true;
	signal G30584: std_logic; attribute dont_touch of G30584: signal is true;
	signal G30585: std_logic; attribute dont_touch of G30585: signal is true;
	signal G30586: std_logic; attribute dont_touch of G30586: signal is true;
	signal G30587: std_logic; attribute dont_touch of G30587: signal is true;
	signal G30588: std_logic; attribute dont_touch of G30588: signal is true;
	signal G30591: std_logic; attribute dont_touch of G30591: signal is true;
	signal G30592: std_logic; attribute dont_touch of G30592: signal is true;
	signal G30593: std_logic; attribute dont_touch of G30593: signal is true;
	signal G30594: std_logic; attribute dont_touch of G30594: signal is true;
	signal G30597: std_logic; attribute dont_touch of G30597: signal is true;
	signal G30600: std_logic; attribute dont_touch of G30600: signal is true;
	signal G30601: std_logic; attribute dont_touch of G30601: signal is true;
	signal G30602: std_logic; attribute dont_touch of G30602: signal is true;
	signal G30605: std_logic; attribute dont_touch of G30605: signal is true;
	signal G30608: std_logic; attribute dont_touch of G30608: signal is true;
	signal G30609: std_logic; attribute dont_touch of G30609: signal is true;
	signal G30610: std_logic; attribute dont_touch of G30610: signal is true;
	signal G30613: std_logic; attribute dont_touch of G30613: signal is true;
	signal G30614: std_logic; attribute dont_touch of G30614: signal is true;
	signal G30617: std_logic; attribute dont_touch of G30617: signal is true;
	signal G30618: std_logic; attribute dont_touch of G30618: signal is true;
	signal G30621: std_logic; attribute dont_touch of G30621: signal is true;
	signal G30622: std_logic; attribute dont_touch of G30622: signal is true;
	signal G30625: std_logic; attribute dont_touch of G30625: signal is true;
	signal G30628: std_logic; attribute dont_touch of G30628: signal is true;
	signal G30629: std_logic; attribute dont_touch of G30629: signal is true;
	signal G30632: std_logic; attribute dont_touch of G30632: signal is true;
	signal G30635: std_logic; attribute dont_touch of G30635: signal is true;
	signal G30636: std_logic; attribute dont_touch of G30636: signal is true;
	signal G30637: std_logic; attribute dont_touch of G30637: signal is true;
	signal G30638: std_logic; attribute dont_touch of G30638: signal is true;
	signal G30639: std_logic; attribute dont_touch of G30639: signal is true;
	signal G30640: std_logic; attribute dont_touch of G30640: signal is true;
	signal G30641: std_logic; attribute dont_touch of G30641: signal is true;
	signal G30642: std_logic; attribute dont_touch of G30642: signal is true;
	signal G30643: std_logic; attribute dont_touch of G30643: signal is true;
	signal G30644: std_logic; attribute dont_touch of G30644: signal is true;
	signal G30645: std_logic; attribute dont_touch of G30645: signal is true;
	signal G30646: std_logic; attribute dont_touch of G30646: signal is true;
	signal G30647: std_logic; attribute dont_touch of G30647: signal is true;
	signal G30648: std_logic; attribute dont_touch of G30648: signal is true;
	signal G30649: std_logic; attribute dont_touch of G30649: signal is true;
	signal G30650: std_logic; attribute dont_touch of G30650: signal is true;
	signal G30651: std_logic; attribute dont_touch of G30651: signal is true;
	signal G30652: std_logic; attribute dont_touch of G30652: signal is true;
	signal G30653: std_logic; attribute dont_touch of G30653: signal is true;
	signal G30654: std_logic; attribute dont_touch of G30654: signal is true;
	signal G30655: std_logic; attribute dont_touch of G30655: signal is true;
	signal G30656: std_logic; attribute dont_touch of G30656: signal is true;
	signal G30657: std_logic; attribute dont_touch of G30657: signal is true;
	signal G30658: std_logic; attribute dont_touch of G30658: signal is true;
	signal G30659: std_logic; attribute dont_touch of G30659: signal is true;
	signal G30660: std_logic; attribute dont_touch of G30660: signal is true;
	signal G30661: std_logic; attribute dont_touch of G30661: signal is true;
	signal G30662: std_logic; attribute dont_touch of G30662: signal is true;
	signal G30663: std_logic; attribute dont_touch of G30663: signal is true;
	signal G30664: std_logic; attribute dont_touch of G30664: signal is true;
	signal G30665: std_logic; attribute dont_touch of G30665: signal is true;
	signal G30666: std_logic; attribute dont_touch of G30666: signal is true;
	signal G30667: std_logic; attribute dont_touch of G30667: signal is true;
	signal G30668: std_logic; attribute dont_touch of G30668: signal is true;
	signal G30669: std_logic; attribute dont_touch of G30669: signal is true;
	signal G30670: std_logic; attribute dont_touch of G30670: signal is true;
	signal G30671: std_logic; attribute dont_touch of G30671: signal is true;
	signal G30672: std_logic; attribute dont_touch of G30672: signal is true;
	signal G30673: std_logic; attribute dont_touch of G30673: signal is true;
	signal G30674: std_logic; attribute dont_touch of G30674: signal is true;
	signal G30675: std_logic; attribute dont_touch of G30675: signal is true;
	signal G30676: std_logic; attribute dont_touch of G30676: signal is true;
	signal G30677: std_logic; attribute dont_touch of G30677: signal is true;
	signal G30678: std_logic; attribute dont_touch of G30678: signal is true;
	signal G30679: std_logic; attribute dont_touch of G30679: signal is true;
	signal G30680: std_logic; attribute dont_touch of G30680: signal is true;
	signal G30681: std_logic; attribute dont_touch of G30681: signal is true;
	signal G30682: std_logic; attribute dont_touch of G30682: signal is true;
	signal G30683: std_logic; attribute dont_touch of G30683: signal is true;
	signal G30684: std_logic; attribute dont_touch of G30684: signal is true;
	signal G30685: std_logic; attribute dont_touch of G30685: signal is true;
	signal G30686: std_logic; attribute dont_touch of G30686: signal is true;
	signal G30687: std_logic; attribute dont_touch of G30687: signal is true;
	signal G30688: std_logic; attribute dont_touch of G30688: signal is true;
	signal G30689: std_logic; attribute dont_touch of G30689: signal is true;
	signal G30690: std_logic; attribute dont_touch of G30690: signal is true;
	signal G30691: std_logic; attribute dont_touch of G30691: signal is true;
	signal G30692: std_logic; attribute dont_touch of G30692: signal is true;
	signal G30693: std_logic; attribute dont_touch of G30693: signal is true;
	signal G30694: std_logic; attribute dont_touch of G30694: signal is true;
	signal G30695: std_logic; attribute dont_touch of G30695: signal is true;
	signal G30696: std_logic; attribute dont_touch of G30696: signal is true;
	signal G30697: std_logic; attribute dont_touch of G30697: signal is true;
	signal G30698: std_logic; attribute dont_touch of G30698: signal is true;
	signal G30699: std_logic; attribute dont_touch of G30699: signal is true;
	signal G30700: std_logic; attribute dont_touch of G30700: signal is true;
	signal G30701: std_logic; attribute dont_touch of G30701: signal is true;
	signal G30702: std_logic; attribute dont_touch of G30702: signal is true;
	signal G30703: std_logic; attribute dont_touch of G30703: signal is true;
	signal G30704: std_logic; attribute dont_touch of G30704: signal is true;
	signal G30705: std_logic; attribute dont_touch of G30705: signal is true;
	signal G30706: std_logic; attribute dont_touch of G30706: signal is true;
	signal G30707: std_logic; attribute dont_touch of G30707: signal is true;
	signal G30708: std_logic; attribute dont_touch of G30708: signal is true;
	signal G30709: std_logic; attribute dont_touch of G30709: signal is true;
	signal G30710: std_logic; attribute dont_touch of G30710: signal is true;
	signal G30711: std_logic; attribute dont_touch of G30711: signal is true;
	signal G30712: std_logic; attribute dont_touch of G30712: signal is true;
	signal G30713: std_logic; attribute dont_touch of G30713: signal is true;
	signal G30714: std_logic; attribute dont_touch of G30714: signal is true;
	signal G30715: std_logic; attribute dont_touch of G30715: signal is true;
	signal G30716: std_logic; attribute dont_touch of G30716: signal is true;
	signal G30717: std_logic; attribute dont_touch of G30717: signal is true;
	signal G30718: std_logic; attribute dont_touch of G30718: signal is true;
	signal G30719: std_logic; attribute dont_touch of G30719: signal is true;
	signal G30720: std_logic; attribute dont_touch of G30720: signal is true;
	signal G30721: std_logic; attribute dont_touch of G30721: signal is true;
	signal G30722: std_logic; attribute dont_touch of G30722: signal is true;
	signal G30723: std_logic; attribute dont_touch of G30723: signal is true;
	signal G30724: std_logic; attribute dont_touch of G30724: signal is true;
	signal G30725: std_logic; attribute dont_touch of G30725: signal is true;
	signal G30726: std_logic; attribute dont_touch of G30726: signal is true;
	signal G30727: std_logic; attribute dont_touch of G30727: signal is true;
	signal G30728: std_logic; attribute dont_touch of G30728: signal is true;
	signal G30729: std_logic; attribute dont_touch of G30729: signal is true;
	signal G30730: std_logic; attribute dont_touch of G30730: signal is true;
	signal G30731: std_logic; attribute dont_touch of G30731: signal is true;
	signal G30732: std_logic; attribute dont_touch of G30732: signal is true;
	signal G30733: std_logic; attribute dont_touch of G30733: signal is true;
	signal G30734: std_logic; attribute dont_touch of G30734: signal is true;
	signal G30735: std_logic; attribute dont_touch of G30735: signal is true;
	signal G30736: std_logic; attribute dont_touch of G30736: signal is true;
	signal G30737: std_logic; attribute dont_touch of G30737: signal is true;
	signal G30738: std_logic; attribute dont_touch of G30738: signal is true;
	signal G30739: std_logic; attribute dont_touch of G30739: signal is true;
	signal G30740: std_logic; attribute dont_touch of G30740: signal is true;
	signal G30741: std_logic; attribute dont_touch of G30741: signal is true;
	signal G30742: std_logic; attribute dont_touch of G30742: signal is true;
	signal G30743: std_logic; attribute dont_touch of G30743: signal is true;
	signal G30744: std_logic; attribute dont_touch of G30744: signal is true;
	signal G30745: std_logic; attribute dont_touch of G30745: signal is true;
	signal G30746: std_logic; attribute dont_touch of G30746: signal is true;
	signal G30747: std_logic; attribute dont_touch of G30747: signal is true;
	signal G30748: std_logic; attribute dont_touch of G30748: signal is true;
	signal G30749: std_logic; attribute dont_touch of G30749: signal is true;
	signal G30750: std_logic; attribute dont_touch of G30750: signal is true;
	signal G30751: std_logic; attribute dont_touch of G30751: signal is true;
	signal G30752: std_logic; attribute dont_touch of G30752: signal is true;
	signal G30753: std_logic; attribute dont_touch of G30753: signal is true;
	signal G30754: std_logic; attribute dont_touch of G30754: signal is true;
	signal G30755: std_logic; attribute dont_touch of G30755: signal is true;
	signal G30756: std_logic; attribute dont_touch of G30756: signal is true;
	signal G30757: std_logic; attribute dont_touch of G30757: signal is true;
	signal G30758: std_logic; attribute dont_touch of G30758: signal is true;
	signal G30759: std_logic; attribute dont_touch of G30759: signal is true;
	signal G30760: std_logic; attribute dont_touch of G30760: signal is true;
	signal G30761: std_logic; attribute dont_touch of G30761: signal is true;
	signal G30762: std_logic; attribute dont_touch of G30762: signal is true;
	signal G30763: std_logic; attribute dont_touch of G30763: signal is true;
	signal G30764: std_logic; attribute dont_touch of G30764: signal is true;
	signal G30765: std_logic; attribute dont_touch of G30765: signal is true;
	signal G30766: std_logic; attribute dont_touch of G30766: signal is true;
	signal G30767: std_logic; attribute dont_touch of G30767: signal is true;
	signal G30768: std_logic; attribute dont_touch of G30768: signal is true;
	signal G30769: std_logic; attribute dont_touch of G30769: signal is true;
	signal G30770: std_logic; attribute dont_touch of G30770: signal is true;
	signal G30771: std_logic; attribute dont_touch of G30771: signal is true;
	signal G30772: std_logic; attribute dont_touch of G30772: signal is true;
	signal G30773: std_logic; attribute dont_touch of G30773: signal is true;
	signal G30774: std_logic; attribute dont_touch of G30774: signal is true;
	signal G30775: std_logic; attribute dont_touch of G30775: signal is true;
	signal G30776: std_logic; attribute dont_touch of G30776: signal is true;
	signal G30777: std_logic; attribute dont_touch of G30777: signal is true;
	signal G30778: std_logic; attribute dont_touch of G30778: signal is true;
	signal G30779: std_logic; attribute dont_touch of G30779: signal is true;
	signal G30780: std_logic; attribute dont_touch of G30780: signal is true;
	signal G30781: std_logic; attribute dont_touch of G30781: signal is true;
	signal G30782: std_logic; attribute dont_touch of G30782: signal is true;
	signal G30783: std_logic; attribute dont_touch of G30783: signal is true;
	signal G30784: std_logic; attribute dont_touch of G30784: signal is true;
	signal G30785: std_logic; attribute dont_touch of G30785: signal is true;
	signal G30786: std_logic; attribute dont_touch of G30786: signal is true;
	signal G30787: std_logic; attribute dont_touch of G30787: signal is true;
	signal G30788: std_logic; attribute dont_touch of G30788: signal is true;
	signal G30789: std_logic; attribute dont_touch of G30789: signal is true;
	signal G30790: std_logic; attribute dont_touch of G30790: signal is true;
	signal G30791: std_logic; attribute dont_touch of G30791: signal is true;
	signal G30792: std_logic; attribute dont_touch of G30792: signal is true;
	signal G30793: std_logic; attribute dont_touch of G30793: signal is true;
	signal G30794: std_logic; attribute dont_touch of G30794: signal is true;
	signal G30795: std_logic; attribute dont_touch of G30795: signal is true;
	signal G30796: std_logic; attribute dont_touch of G30796: signal is true;
	signal G30797: std_logic; attribute dont_touch of G30797: signal is true;
	signal G30798: std_logic; attribute dont_touch of G30798: signal is true;
	signal G30799: std_logic; attribute dont_touch of G30799: signal is true;
	signal G30800: std_logic; attribute dont_touch of G30800: signal is true;
	signal G30801: std_logic; attribute dont_touch of G30801: signal is true;
	signal G30802: std_logic; attribute dont_touch of G30802: signal is true;
	signal G30803: std_logic; attribute dont_touch of G30803: signal is true;
	signal G30804: std_logic; attribute dont_touch of G30804: signal is true;
	signal G30805: std_logic; attribute dont_touch of G30805: signal is true;
	signal G30806: std_logic; attribute dont_touch of G30806: signal is true;
	signal G30807: std_logic; attribute dont_touch of G30807: signal is true;
	signal G30808: std_logic; attribute dont_touch of G30808: signal is true;
	signal G30809: std_logic; attribute dont_touch of G30809: signal is true;
	signal G30810: std_logic; attribute dont_touch of G30810: signal is true;
	signal G30811: std_logic; attribute dont_touch of G30811: signal is true;
	signal G30812: std_logic; attribute dont_touch of G30812: signal is true;
	signal G30813: std_logic; attribute dont_touch of G30813: signal is true;
	signal G30814: std_logic; attribute dont_touch of G30814: signal is true;
	signal G30815: std_logic; attribute dont_touch of G30815: signal is true;
	signal G30816: std_logic; attribute dont_touch of G30816: signal is true;
	signal G30817: std_logic; attribute dont_touch of G30817: signal is true;
	signal G30818: std_logic; attribute dont_touch of G30818: signal is true;
	signal G30819: std_logic; attribute dont_touch of G30819: signal is true;
	signal G30820: std_logic; attribute dont_touch of G30820: signal is true;
	signal G30821: std_logic; attribute dont_touch of G30821: signal is true;
	signal G30822: std_logic; attribute dont_touch of G30822: signal is true;
	signal G30823: std_logic; attribute dont_touch of G30823: signal is true;
	signal G30824: std_logic; attribute dont_touch of G30824: signal is true;
	signal G30825: std_logic; attribute dont_touch of G30825: signal is true;
	signal G30826: std_logic; attribute dont_touch of G30826: signal is true;
	signal G30827: std_logic; attribute dont_touch of G30827: signal is true;
	signal G30828: std_logic; attribute dont_touch of G30828: signal is true;
	signal G30829: std_logic; attribute dont_touch of G30829: signal is true;
	signal G30830: std_logic; attribute dont_touch of G30830: signal is true;
	signal G30831: std_logic; attribute dont_touch of G30831: signal is true;
	signal G30832: std_logic; attribute dont_touch of G30832: signal is true;
	signal G30833: std_logic; attribute dont_touch of G30833: signal is true;
	signal G30834: std_logic; attribute dont_touch of G30834: signal is true;
	signal G30835: std_logic; attribute dont_touch of G30835: signal is true;
	signal G30836: std_logic; attribute dont_touch of G30836: signal is true;
	signal G30837: std_logic; attribute dont_touch of G30837: signal is true;
	signal G30838: std_logic; attribute dont_touch of G30838: signal is true;
	signal G30839: std_logic; attribute dont_touch of G30839: signal is true;
	signal G30840: std_logic; attribute dont_touch of G30840: signal is true;
	signal G30841: std_logic; attribute dont_touch of G30841: signal is true;
	signal G30842: std_logic; attribute dont_touch of G30842: signal is true;
	signal G30843: std_logic; attribute dont_touch of G30843: signal is true;
	signal G30844: std_logic; attribute dont_touch of G30844: signal is true;
	signal G30845: std_logic; attribute dont_touch of G30845: signal is true;
	signal G30846: std_logic; attribute dont_touch of G30846: signal is true;
	signal G30847: std_logic; attribute dont_touch of G30847: signal is true;
	signal G30848: std_logic; attribute dont_touch of G30848: signal is true;
	signal G30849: std_logic; attribute dont_touch of G30849: signal is true;
	signal G30850: std_logic; attribute dont_touch of G30850: signal is true;
	signal G30851: std_logic; attribute dont_touch of G30851: signal is true;
	signal G30852: std_logic; attribute dont_touch of G30852: signal is true;
	signal G30853: std_logic; attribute dont_touch of G30853: signal is true;
	signal G30854: std_logic; attribute dont_touch of G30854: signal is true;
	signal G30855: std_logic; attribute dont_touch of G30855: signal is true;
	signal G30856: std_logic; attribute dont_touch of G30856: signal is true;
	signal G30857: std_logic; attribute dont_touch of G30857: signal is true;
	signal G30858: std_logic; attribute dont_touch of G30858: signal is true;
	signal G30859: std_logic; attribute dont_touch of G30859: signal is true;
	signal G30860: std_logic; attribute dont_touch of G30860: signal is true;
	signal G30861: std_logic; attribute dont_touch of G30861: signal is true;
	signal G30862: std_logic; attribute dont_touch of G30862: signal is true;
	signal G30863: std_logic; attribute dont_touch of G30863: signal is true;
	signal G30864: std_logic; attribute dont_touch of G30864: signal is true;
	signal G30865: std_logic; attribute dont_touch of G30865: signal is true;
	signal G30866: std_logic; attribute dont_touch of G30866: signal is true;
	signal G30867: std_logic; attribute dont_touch of G30867: signal is true;
	signal G30868: std_logic; attribute dont_touch of G30868: signal is true;
	signal G30869: std_logic; attribute dont_touch of G30869: signal is true;
	signal G30870: std_logic; attribute dont_touch of G30870: signal is true;
	signal G30871: std_logic; attribute dont_touch of G30871: signal is true;
	signal G30872: std_logic; attribute dont_touch of G30872: signal is true;
	signal G30873: std_logic; attribute dont_touch of G30873: signal is true;
	signal G30874: std_logic; attribute dont_touch of G30874: signal is true;
	signal G30875: std_logic; attribute dont_touch of G30875: signal is true;
	signal G30876: std_logic; attribute dont_touch of G30876: signal is true;
	signal G30877: std_logic; attribute dont_touch of G30877: signal is true;
	signal G30878: std_logic; attribute dont_touch of G30878: signal is true;
	signal G30879: std_logic; attribute dont_touch of G30879: signal is true;
	signal G30880: std_logic; attribute dont_touch of G30880: signal is true;
	signal G30881: std_logic; attribute dont_touch of G30881: signal is true;
	signal G30882: std_logic; attribute dont_touch of G30882: signal is true;
	signal G30883: std_logic; attribute dont_touch of G30883: signal is true;
	signal G30884: std_logic; attribute dont_touch of G30884: signal is true;
	signal G30885: std_logic; attribute dont_touch of G30885: signal is true;
	signal G30886: std_logic; attribute dont_touch of G30886: signal is true;
	signal G30887: std_logic; attribute dont_touch of G30887: signal is true;
	signal G30888: std_logic; attribute dont_touch of G30888: signal is true;
	signal G30889: std_logic; attribute dont_touch of G30889: signal is true;
	signal G30890: std_logic; attribute dont_touch of G30890: signal is true;
	signal G30891: std_logic; attribute dont_touch of G30891: signal is true;
	signal G30892: std_logic; attribute dont_touch of G30892: signal is true;
	signal G30893: std_logic; attribute dont_touch of G30893: signal is true;
	signal G30894: std_logic; attribute dont_touch of G30894: signal is true;
	signal G30895: std_logic; attribute dont_touch of G30895: signal is true;
	signal G30896: std_logic; attribute dont_touch of G30896: signal is true;
	signal G30897: std_logic; attribute dont_touch of G30897: signal is true;
	signal G30898: std_logic; attribute dont_touch of G30898: signal is true;
	signal G30899: std_logic; attribute dont_touch of G30899: signal is true;
	signal G30900: std_logic; attribute dont_touch of G30900: signal is true;
	signal G30901: std_logic; attribute dont_touch of G30901: signal is true;
	signal G30902: std_logic; attribute dont_touch of G30902: signal is true;
	signal G30903: std_logic; attribute dont_touch of G30903: signal is true;
	signal G30904: std_logic; attribute dont_touch of G30904: signal is true;
	signal G30905: std_logic; attribute dont_touch of G30905: signal is true;
	signal G30906: std_logic; attribute dont_touch of G30906: signal is true;
	signal G30907: std_logic; attribute dont_touch of G30907: signal is true;
	signal G30908: std_logic; attribute dont_touch of G30908: signal is true;
	signal G30909: std_logic; attribute dont_touch of G30909: signal is true;
	signal G30910: std_logic; attribute dont_touch of G30910: signal is true;
	signal G30911: std_logic; attribute dont_touch of G30911: signal is true;
	signal G30912: std_logic; attribute dont_touch of G30912: signal is true;
	signal G30913: std_logic; attribute dont_touch of G30913: signal is true;
	signal G30914: std_logic; attribute dont_touch of G30914: signal is true;
	signal G30915: std_logic; attribute dont_touch of G30915: signal is true;
	signal G30916: std_logic; attribute dont_touch of G30916: signal is true;
	signal G30917: std_logic; attribute dont_touch of G30917: signal is true;
	signal G30918: std_logic; attribute dont_touch of G30918: signal is true;
	signal G30919: std_logic; attribute dont_touch of G30919: signal is true;
	signal G30920: std_logic; attribute dont_touch of G30920: signal is true;
	signal G30921: std_logic; attribute dont_touch of G30921: signal is true;
	signal G30922: std_logic; attribute dont_touch of G30922: signal is true;
	signal G30923: std_logic; attribute dont_touch of G30923: signal is true;
	signal G30924: std_logic; attribute dont_touch of G30924: signal is true;
	signal G30925: std_logic; attribute dont_touch of G30925: signal is true;
	signal G30926: std_logic; attribute dont_touch of G30926: signal is true;
	signal G30927: std_logic; attribute dont_touch of G30927: signal is true;
	signal G30928: std_logic; attribute dont_touch of G30928: signal is true;
	signal G30929: std_logic; attribute dont_touch of G30929: signal is true;
	signal G30930: std_logic; attribute dont_touch of G30930: signal is true;
	signal G30931: std_logic; attribute dont_touch of G30931: signal is true;
	signal G30932: std_logic; attribute dont_touch of G30932: signal is true;
	signal G30933: std_logic; attribute dont_touch of G30933: signal is true;
	signal G30934: std_logic; attribute dont_touch of G30934: signal is true;
	signal G30935: std_logic; attribute dont_touch of G30935: signal is true;
	signal G30936: std_logic; attribute dont_touch of G30936: signal is true;
	signal G30937: std_logic; attribute dont_touch of G30937: signal is true;
	signal G30938: std_logic; attribute dont_touch of G30938: signal is true;
	signal G30939: std_logic; attribute dont_touch of G30939: signal is true;
	signal G30940: std_logic; attribute dont_touch of G30940: signal is true;
	signal G30941: std_logic; attribute dont_touch of G30941: signal is true;
	signal G30942: std_logic; attribute dont_touch of G30942: signal is true;
	signal G30943: std_logic; attribute dont_touch of G30943: signal is true;
	signal G30944: std_logic; attribute dont_touch of G30944: signal is true;
	signal G30945: std_logic; attribute dont_touch of G30945: signal is true;
	signal G30946: std_logic; attribute dont_touch of G30946: signal is true;
	signal G30947: std_logic; attribute dont_touch of G30947: signal is true;
	signal G30948: std_logic; attribute dont_touch of G30948: signal is true;
	signal G30949: std_logic; attribute dont_touch of G30949: signal is true;
	signal G30950: std_logic; attribute dont_touch of G30950: signal is true;
	signal G30951: std_logic; attribute dont_touch of G30951: signal is true;
	signal G30952: std_logic; attribute dont_touch of G30952: signal is true;
	signal G30953: std_logic; attribute dont_touch of G30953: signal is true;
	signal G30954: std_logic; attribute dont_touch of G30954: signal is true;
	signal G30955: std_logic; attribute dont_touch of G30955: signal is true;
	signal G30956: std_logic; attribute dont_touch of G30956: signal is true;
	signal G30957: std_logic; attribute dont_touch of G30957: signal is true;
	signal G30958: std_logic; attribute dont_touch of G30958: signal is true;
	signal G30959: std_logic; attribute dont_touch of G30959: signal is true;
	signal G30960: std_logic; attribute dont_touch of G30960: signal is true;
	signal G30961: std_logic; attribute dont_touch of G30961: signal is true;
	signal G30962: std_logic; attribute dont_touch of G30962: signal is true;
	signal G30963: std_logic; attribute dont_touch of G30963: signal is true;
	signal G30964: std_logic; attribute dont_touch of G30964: signal is true;
	signal G30965: std_logic; attribute dont_touch of G30965: signal is true;
	signal G30966: std_logic; attribute dont_touch of G30966: signal is true;
	signal G30967: std_logic; attribute dont_touch of G30967: signal is true;
	signal G30968: std_logic; attribute dont_touch of G30968: signal is true;
	signal G30969: std_logic; attribute dont_touch of G30969: signal is true;
	signal G30970: std_logic; attribute dont_touch of G30970: signal is true;
	signal G30971: std_logic; attribute dont_touch of G30971: signal is true;
	signal G30972: std_logic; attribute dont_touch of G30972: signal is true;
	signal G30973: std_logic; attribute dont_touch of G30973: signal is true;
	signal G30974: std_logic; attribute dont_touch of G30974: signal is true;
	signal G30975: std_logic; attribute dont_touch of G30975: signal is true;
	signal G30976: std_logic; attribute dont_touch of G30976: signal is true;
	signal G30977: std_logic; attribute dont_touch of G30977: signal is true;
	signal G30978: std_logic; attribute dont_touch of G30978: signal is true;
	signal G30979: std_logic; attribute dont_touch of G30979: signal is true;
	signal G30980: std_logic; attribute dont_touch of G30980: signal is true;
	signal G30981: std_logic; attribute dont_touch of G30981: signal is true;
	signal G30982: std_logic; attribute dont_touch of G30982: signal is true;
	signal G30983: std_logic; attribute dont_touch of G30983: signal is true;
	signal G30984: std_logic; attribute dont_touch of G30984: signal is true;
	signal G30985: std_logic; attribute dont_touch of G30985: signal is true;
	signal G30986: std_logic; attribute dont_touch of G30986: signal is true;
	signal G30987: std_logic; attribute dont_touch of G30987: signal is true;
	signal G30988: std_logic; attribute dont_touch of G30988: signal is true;
	signal G30989: std_logic; attribute dont_touch of G30989: signal is true;
	signal I13089: std_logic; attribute dont_touch of I13089: signal is true;
	signal I13092: std_logic; attribute dont_touch of I13092: signal is true;
	signal I13095: std_logic; attribute dont_touch of I13095: signal is true;
	signal I13098: std_logic; attribute dont_touch of I13098: signal is true;
	signal I13101: std_logic; attribute dont_touch of I13101: signal is true;
	signal I13104: std_logic; attribute dont_touch of I13104: signal is true;
	signal I13107: std_logic; attribute dont_touch of I13107: signal is true;
	signal I13110: std_logic; attribute dont_touch of I13110: signal is true;
	signal I13113: std_logic; attribute dont_touch of I13113: signal is true;
	signal I13116: std_logic; attribute dont_touch of I13116: signal is true;
	signal I13119: std_logic; attribute dont_touch of I13119: signal is true;
	signal I13122: std_logic; attribute dont_touch of I13122: signal is true;
	signal I13125: std_logic; attribute dont_touch of I13125: signal is true;
	signal I13128: std_logic; attribute dont_touch of I13128: signal is true;
	signal I13131: std_logic; attribute dont_touch of I13131: signal is true;
	signal I13134: std_logic; attribute dont_touch of I13134: signal is true;
	signal I13137: std_logic; attribute dont_touch of I13137: signal is true;
	signal I13140: std_logic; attribute dont_touch of I13140: signal is true;
	signal I13143: std_logic; attribute dont_touch of I13143: signal is true;
	signal I13146: std_logic; attribute dont_touch of I13146: signal is true;
	signal I13149: std_logic; attribute dont_touch of I13149: signal is true;
	signal I13152: std_logic; attribute dont_touch of I13152: signal is true;
	signal I13155: std_logic; attribute dont_touch of I13155: signal is true;
	signal I13158: std_logic; attribute dont_touch of I13158: signal is true;
	signal I13161: std_logic; attribute dont_touch of I13161: signal is true;
	signal I13165: std_logic; attribute dont_touch of I13165: signal is true;
	signal I13169: std_logic; attribute dont_touch of I13169: signal is true;
	signal I13173: std_logic; attribute dont_touch of I13173: signal is true;
	signal I13176: std_logic; attribute dont_touch of I13176: signal is true;
	signal I13179: std_logic; attribute dont_touch of I13179: signal is true;
	signal I13182: std_logic; attribute dont_touch of I13182: signal is true;
	signal I13186: std_logic; attribute dont_touch of I13186: signal is true;
	signal I13190: std_logic; attribute dont_touch of I13190: signal is true;
	signal I13194: std_logic; attribute dont_touch of I13194: signal is true;
	signal I13197: std_logic; attribute dont_touch of I13197: signal is true;
	signal I13200: std_logic; attribute dont_touch of I13200: signal is true;
	signal I13203: std_logic; attribute dont_touch of I13203: signal is true;
	signal I13207: std_logic; attribute dont_touch of I13207: signal is true;
	signal I13211: std_logic; attribute dont_touch of I13211: signal is true;
	signal I13215: std_logic; attribute dont_touch of I13215: signal is true;
	signal I13218: std_logic; attribute dont_touch of I13218: signal is true;
	signal I13221: std_logic; attribute dont_touch of I13221: signal is true;
	signal I13224: std_logic; attribute dont_touch of I13224: signal is true;
	signal I13228: std_logic; attribute dont_touch of I13228: signal is true;
	signal I13232: std_logic; attribute dont_touch of I13232: signal is true;
	signal I13236: std_logic; attribute dont_touch of I13236: signal is true;
	signal I13239: std_logic; attribute dont_touch of I13239: signal is true;
	signal I13242: std_logic; attribute dont_touch of I13242: signal is true;
	signal I13246: std_logic; attribute dont_touch of I13246: signal is true;
	signal I13275: std_logic; attribute dont_touch of I13275: signal is true;
	signal I13316: std_logic; attribute dont_touch of I13316: signal is true;
	signal I13320: std_logic; attribute dont_touch of I13320: signal is true;
	signal I13366: std_logic; attribute dont_touch of I13366: signal is true;
	signal I13417: std_logic; attribute dont_touch of I13417: signal is true;
	signal I13421: std_logic; attribute dont_touch of I13421: signal is true;
	signal I13430: std_logic; attribute dont_touch of I13430: signal is true;
	signal I13433: std_logic; attribute dont_touch of I13433: signal is true;
	signal I13478: std_logic; attribute dont_touch of I13478: signal is true;
	signal I13501: std_logic; attribute dont_touch of I13501: signal is true;
	signal I13504: std_logic; attribute dont_touch of I13504: signal is true;
	signal I13538: std_logic; attribute dont_touch of I13538: signal is true;
	signal I13575: std_logic; attribute dont_touch of I13575: signal is true;
	signal I13578: std_logic; attribute dont_touch of I13578: signal is true;
	signal I13601: std_logic; attribute dont_touch of I13601: signal is true;
	signal I13604: std_logic; attribute dont_touch of I13604: signal is true;
	signal I13652: std_logic; attribute dont_touch of I13652: signal is true;
	signal I13655: std_logic; attribute dont_touch of I13655: signal is true;
	signal I13677: std_logic; attribute dont_touch of I13677: signal is true;
	signal I13680: std_logic; attribute dont_touch of I13680: signal is true;
	signal I13742: std_logic; attribute dont_touch of I13742: signal is true;
	signal I13745: std_logic; attribute dont_touch of I13745: signal is true;
	signal I13775: std_logic; attribute dont_touch of I13775: signal is true;
	signal I13801: std_logic; attribute dont_touch of I13801: signal is true;
	signal I13804: std_logic; attribute dont_touch of I13804: signal is true;
	signal I13820: std_logic; attribute dont_touch of I13820: signal is true;
	signal I13849: std_logic; attribute dont_touch of I13849: signal is true;
	signal I13868: std_logic; attribute dont_touch of I13868: signal is true;
	signal I13892: std_logic; attribute dont_touch of I13892: signal is true;
	signal I13896: std_logic; attribute dont_touch of I13896: signal is true;
	signal I13901: std_logic; attribute dont_touch of I13901: signal is true;
	signal I13904: std_logic; attribute dont_touch of I13904: signal is true;
	signal I13907: std_logic; attribute dont_touch of I13907: signal is true;
	signal I13910: std_logic; attribute dont_touch of I13910: signal is true;
	signal I13913: std_logic; attribute dont_touch of I13913: signal is true;
	signal I13916: std_logic; attribute dont_touch of I13916: signal is true;
	signal I13919: std_logic; attribute dont_touch of I13919: signal is true;
	signal I13922: std_logic; attribute dont_touch of I13922: signal is true;
	signal I13925: std_logic; attribute dont_touch of I13925: signal is true;
	signal I13928: std_logic; attribute dont_touch of I13928: signal is true;
	signal I13931: std_logic; attribute dont_touch of I13931: signal is true;
	signal I13934: std_logic; attribute dont_touch of I13934: signal is true;
	signal I13937: std_logic; attribute dont_touch of I13937: signal is true;
	signal I13940: std_logic; attribute dont_touch of I13940: signal is true;
	signal I13943: std_logic; attribute dont_touch of I13943: signal is true;
	signal I13947: std_logic; attribute dont_touch of I13947: signal is true;
	signal I13950: std_logic; attribute dont_touch of I13950: signal is true;
	signal I13953: std_logic; attribute dont_touch of I13953: signal is true;
	signal I13956: std_logic; attribute dont_touch of I13956: signal is true;
	signal I13959: std_logic; attribute dont_touch of I13959: signal is true;
	signal I13962: std_logic; attribute dont_touch of I13962: signal is true;
	signal I13965: std_logic; attribute dont_touch of I13965: signal is true;
	signal I13968: std_logic; attribute dont_touch of I13968: signal is true;
	signal I13971: std_logic; attribute dont_touch of I13971: signal is true;
	signal I13974: std_logic; attribute dont_touch of I13974: signal is true;
	signal I13977: std_logic; attribute dont_touch of I13977: signal is true;
	signal I13980: std_logic; attribute dont_touch of I13980: signal is true;
	signal I13984: std_logic; attribute dont_touch of I13984: signal is true;
	signal I13987: std_logic; attribute dont_touch of I13987: signal is true;
	signal I13990: std_logic; attribute dont_touch of I13990: signal is true;
	signal I13993: std_logic; attribute dont_touch of I13993: signal is true;
	signal I13999: std_logic; attribute dont_touch of I13999: signal is true;
	signal I14002: std_logic; attribute dont_touch of I14002: signal is true;
	signal I14006: std_logic; attribute dont_touch of I14006: signal is true;
	signal I14009: std_logic; attribute dont_touch of I14009: signal is true;
	signal I14014: std_logic; attribute dont_touch of I14014: signal is true;
	signal I14017: std_logic; attribute dont_touch of I14017: signal is true;
	signal I14020: std_logic; attribute dont_touch of I14020: signal is true;
	signal I14027: std_logic; attribute dont_touch of I14027: signal is true;
	signal I14030: std_logic; attribute dont_touch of I14030: signal is true;
	signal I14034: std_logic; attribute dont_touch of I14034: signal is true;
	signal I14037: std_logic; attribute dont_touch of I14037: signal is true;
	signal I14040: std_logic; attribute dont_touch of I14040: signal is true;
	signal I14049: std_logic; attribute dont_touch of I14049: signal is true;
	signal I14052: std_logic; attribute dont_touch of I14052: signal is true;
	signal I14056: std_logic; attribute dont_touch of I14056: signal is true;
	signal I14066: std_logic; attribute dont_touch of I14066: signal is true;
	signal I14069: std_logic; attribute dont_touch of I14069: signal is true;
	signal I14073: std_logic; attribute dont_touch of I14073: signal is true;
	signal I14083: std_logic; attribute dont_touch of I14083: signal is true;
	signal I14091: std_logic; attribute dont_touch of I14091: signal is true;
	signal I14094: std_logic; attribute dont_touch of I14094: signal is true;
	signal I14104: std_logic; attribute dont_touch of I14104: signal is true;
	signal I14113: std_logic; attribute dont_touch of I14113: signal is true;
	signal I14134: std_logic; attribute dont_touch of I14134: signal is true;
	signal I14143: std_logic; attribute dont_touch of I14143: signal is true;
	signal I14149: std_logic; attribute dont_touch of I14149: signal is true;
	signal I14163: std_logic; attribute dont_touch of I14163: signal is true;
	signal I14182: std_logic; attribute dont_touch of I14182: signal is true;
	signal I14191: std_logic; attribute dont_touch of I14191: signal is true;
	signal I14195: std_logic; attribute dont_touch of I14195: signal is true;
	signal I14219: std_logic; attribute dont_touch of I14219: signal is true;
	signal I14238: std_logic; attribute dont_touch of I14238: signal is true;
	signal I14243: std_logic; attribute dont_touch of I14243: signal is true;
	signal I14246: std_logic; attribute dont_touch of I14246: signal is true;
	signal I14249: std_logic; attribute dont_touch of I14249: signal is true;
	signal I14280: std_logic; attribute dont_touch of I14280: signal is true;
	signal I14295: std_logic; attribute dont_touch of I14295: signal is true;
	signal I14298: std_logic; attribute dont_touch of I14298: signal is true;
	signal I14306: std_logic; attribute dont_touch of I14306: signal is true;
	signal I14338: std_logic; attribute dont_touch of I14338: signal is true;
	signal I14343: std_logic; attribute dont_touch of I14343: signal is true;
	signal I14357: std_logic; attribute dont_touch of I14357: signal is true;
	signal I14378: std_logic; attribute dont_touch of I14378: signal is true;
	signal I14381: std_logic; attribute dont_touch of I14381: signal is true;
	signal I14384: std_logic; attribute dont_touch of I14384: signal is true;
	signal I14402: std_logic; attribute dont_touch of I14402: signal is true;
	signal I14413: std_logic; attribute dont_touch of I14413: signal is true;
	signal I14416: std_logic; attribute dont_touch of I14416: signal is true;
	signal I14424: std_logic; attribute dont_touch of I14424: signal is true;
	signal I14442: std_logic; attribute dont_touch of I14442: signal is true;
	signal I14446: std_logic; attribute dont_touch of I14446: signal is true;
	signal I14449: std_logic; attribute dont_touch of I14449: signal is true;
	signal I14459: std_logic; attribute dont_touch of I14459: signal is true;
	signal I14472: std_logic; attribute dont_touch of I14472: signal is true;
	signal I14475: std_logic; attribute dont_touch of I14475: signal is true;
	signal I14478: std_logic; attribute dont_touch of I14478: signal is true;
	signal I14489: std_logic; attribute dont_touch of I14489: signal is true;
	signal I14496: std_logic; attribute dont_touch of I14496: signal is true;
	signal I14499: std_logic; attribute dont_touch of I14499: signal is true;
	signal I14502: std_logic; attribute dont_touch of I14502: signal is true;
	signal I14513: std_logic; attribute dont_touch of I14513: signal is true;
	signal I14516: std_logic; attribute dont_touch of I14516: signal is true;
	signal I14519: std_logic; attribute dont_touch of I14519: signal is true;
	signal I14525: std_logic; attribute dont_touch of I14525: signal is true;
	signal I14529: std_logic; attribute dont_touch of I14529: signal is true;
	signal I14532: std_logic; attribute dont_touch of I14532: signal is true;
	signal I14535: std_logic; attribute dont_touch of I14535: signal is true;
	signal I14538: std_logic; attribute dont_touch of I14538: signal is true;
	signal I14541: std_logic; attribute dont_touch of I14541: signal is true;
	signal I14544: std_logic; attribute dont_touch of I14544: signal is true;
	signal I14547: std_logic; attribute dont_touch of I14547: signal is true;
	signal I14550: std_logic; attribute dont_touch of I14550: signal is true;
	signal I14553: std_logic; attribute dont_touch of I14553: signal is true;
	signal I14556: std_logic; attribute dont_touch of I14556: signal is true;
	signal I14559: std_logic; attribute dont_touch of I14559: signal is true;
	signal I14562: std_logic; attribute dont_touch of I14562: signal is true;
	signal I14565: std_logic; attribute dont_touch of I14565: signal is true;
	signal I14568: std_logic; attribute dont_touch of I14568: signal is true;
	signal I14571: std_logic; attribute dont_touch of I14571: signal is true;
	signal I14574: std_logic; attribute dont_touch of I14574: signal is true;
	signal I14577: std_logic; attribute dont_touch of I14577: signal is true;
	signal I14580: std_logic; attribute dont_touch of I14580: signal is true;
	signal I14584: std_logic; attribute dont_touch of I14584: signal is true;
	signal I14587: std_logic; attribute dont_touch of I14587: signal is true;
	signal I14590: std_logic; attribute dont_touch of I14590: signal is true;
	signal I14593: std_logic; attribute dont_touch of I14593: signal is true;
	signal I14596: std_logic; attribute dont_touch of I14596: signal is true;
	signal I14599: std_logic; attribute dont_touch of I14599: signal is true;
	signal I14602: std_logic; attribute dont_touch of I14602: signal is true;
	signal I14605: std_logic; attribute dont_touch of I14605: signal is true;
	signal I14609: std_logic; attribute dont_touch of I14609: signal is true;
	signal I14612: std_logic; attribute dont_touch of I14612: signal is true;
	signal I14615: std_logic; attribute dont_touch of I14615: signal is true;
	signal I14618: std_logic; attribute dont_touch of I14618: signal is true;
	signal I14621: std_logic; attribute dont_touch of I14621: signal is true;
	signal I14624: std_logic; attribute dont_touch of I14624: signal is true;
	signal I14628: std_logic; attribute dont_touch of I14628: signal is true;
	signal I14631: std_logic; attribute dont_touch of I14631: signal is true;
	signal I14634: std_logic; attribute dont_touch of I14634: signal is true;
	signal I14637: std_logic; attribute dont_touch of I14637: signal is true;
	signal I14641: std_logic; attribute dont_touch of I14641: signal is true;
	signal I14644: std_logic; attribute dont_touch of I14644: signal is true;
	signal I14647: std_logic; attribute dont_touch of I14647: signal is true;
	signal I14650: std_logic; attribute dont_touch of I14650: signal is true;
	signal I14654: std_logic; attribute dont_touch of I14654: signal is true;
	signal I14660: std_logic; attribute dont_touch of I14660: signal is true;
	signal I14665: std_logic; attribute dont_touch of I14665: signal is true;
	signal I14668: std_logic; attribute dont_touch of I14668: signal is true;
	signal I14675: std_logic; attribute dont_touch of I14675: signal is true;
	signal I14688: std_logic; attribute dont_touch of I14688: signal is true;
	signal I14704: std_logic; attribute dont_touch of I14704: signal is true;
	signal I14709: std_logic; attribute dont_touch of I14709: signal is true;
	signal I14712: std_logic; attribute dont_touch of I14712: signal is true;
	signal I14715: std_logic; attribute dont_touch of I14715: signal is true;
	signal I14731: std_logic; attribute dont_touch of I14731: signal is true;
	signal I14734: std_logic; attribute dont_touch of I14734: signal is true;
	signal I14739: std_logic; attribute dont_touch of I14739: signal is true;
	signal I14742: std_logic; attribute dont_touch of I14742: signal is true;
	signal I14755: std_logic; attribute dont_touch of I14755: signal is true;
	signal I14760: std_logic; attribute dont_touch of I14760: signal is true;
	signal I14763: std_logic; attribute dont_touch of I14763: signal is true;
	signal I14766: std_logic; attribute dont_touch of I14766: signal is true;
	signal I14769: std_logic; attribute dont_touch of I14769: signal is true;
	signal I14775: std_logic; attribute dont_touch of I14775: signal is true;
	signal I14778: std_logic; attribute dont_touch of I14778: signal is true;
	signal I14783: std_logic; attribute dont_touch of I14783: signal is true;
	signal I14786: std_logic; attribute dont_touch of I14786: signal is true;
	signal I14799: std_logic; attribute dont_touch of I14799: signal is true;
	signal I14802: std_logic; attribute dont_touch of I14802: signal is true;
	signal I14808: std_logic; attribute dont_touch of I14808: signal is true;
	signal I14811: std_logic; attribute dont_touch of I14811: signal is true;
	signal I14816: std_logic; attribute dont_touch of I14816: signal is true;
	signal I14819: std_logic; attribute dont_touch of I14819: signal is true;
	signal I14822: std_logic; attribute dont_touch of I14822: signal is true;
	signal I14825: std_logic; attribute dont_touch of I14825: signal is true;
	signal I14831: std_logic; attribute dont_touch of I14831: signal is true;
	signal I14834: std_logic; attribute dont_touch of I14834: signal is true;
	signal I14839: std_logic; attribute dont_touch of I14839: signal is true;
	signal I14842: std_logic; attribute dont_touch of I14842: signal is true;
	signal I14848: std_logic; attribute dont_touch of I14848: signal is true;
	signal I14857: std_logic; attribute dont_touch of I14857: signal is true;
	signal I14860: std_logic; attribute dont_touch of I14860: signal is true;
	signal I14865: std_logic; attribute dont_touch of I14865: signal is true;
	signal I14868: std_logic; attribute dont_touch of I14868: signal is true;
	signal I14874: std_logic; attribute dont_touch of I14874: signal is true;
	signal I14877: std_logic; attribute dont_touch of I14877: signal is true;
	signal I14882: std_logic; attribute dont_touch of I14882: signal is true;
	signal I14885: std_logic; attribute dont_touch of I14885: signal is true;
	signal I14888: std_logic; attribute dont_touch of I14888: signal is true;
	signal I14891: std_logic; attribute dont_touch of I14891: signal is true;
	signal I14897: std_logic; attribute dont_touch of I14897: signal is true;
	signal I14900: std_logic; attribute dont_touch of I14900: signal is true;
	signal I14917: std_logic; attribute dont_touch of I14917: signal is true;
	signal I14920: std_logic; attribute dont_touch of I14920: signal is true;
	signal I14925: std_logic; attribute dont_touch of I14925: signal is true;
	signal I14928: std_logic; attribute dont_touch of I14928: signal is true;
	signal I14934: std_logic; attribute dont_touch of I14934: signal is true;
	signal I14937: std_logic; attribute dont_touch of I14937: signal is true;
	signal I14942: std_logic; attribute dont_touch of I14942: signal is true;
	signal I14945: std_logic; attribute dont_touch of I14945: signal is true;
	signal I14948: std_logic; attribute dont_touch of I14948: signal is true;
	signal I14951: std_logic; attribute dont_touch of I14951: signal is true;
	signal I14957: std_logic; attribute dont_touch of I14957: signal is true;
	signal I14973: std_logic; attribute dont_touch of I14973: signal is true;
	signal I14976: std_logic; attribute dont_touch of I14976: signal is true;
	signal I14981: std_logic; attribute dont_touch of I14981: signal is true;
	signal I14984: std_logic; attribute dont_touch of I14984: signal is true;
	signal I14990: std_logic; attribute dont_touch of I14990: signal is true;
	signal I14993: std_logic; attribute dont_touch of I14993: signal is true;
	signal I15012: std_logic; attribute dont_touch of I15012: signal is true;
	signal I15015: std_logic; attribute dont_touch of I15015: signal is true;
	signal I15019: std_logic; attribute dont_touch of I15019: signal is true;
	signal I15167: std_logic; attribute dont_touch of I15167: signal is true;
	signal I15168: std_logic; attribute dont_touch of I15168: signal is true;
	signal I15169: std_logic; attribute dont_touch of I15169: signal is true;
	signal I15183: std_logic; attribute dont_touch of I15183: signal is true;
	signal I15184: std_logic; attribute dont_touch of I15184: signal is true;
	signal I15185: std_logic; attribute dont_touch of I15185: signal is true;
	signal I15190: std_logic; attribute dont_touch of I15190: signal is true;
	signal I15191: std_logic; attribute dont_touch of I15191: signal is true;
	signal I15192: std_logic; attribute dont_touch of I15192: signal is true;
	signal I15204: std_logic; attribute dont_touch of I15204: signal is true;
	signal I15205: std_logic; attribute dont_touch of I15205: signal is true;
	signal I15206: std_logic; attribute dont_touch of I15206: signal is true;
	signal I15211: std_logic; attribute dont_touch of I15211: signal is true;
	signal I15212: std_logic; attribute dont_touch of I15212: signal is true;
	signal I15213: std_logic; attribute dont_touch of I15213: signal is true;
	signal I15222: std_logic; attribute dont_touch of I15222: signal is true;
	signal I15226: std_logic; attribute dont_touch of I15226: signal is true;
	signal I15230: std_logic; attribute dont_touch of I15230: signal is true;
	signal I15237: std_logic; attribute dont_touch of I15237: signal is true;
	signal I15238: std_logic; attribute dont_touch of I15238: signal is true;
	signal I15239: std_logic; attribute dont_touch of I15239: signal is true;
	signal I15244: std_logic; attribute dont_touch of I15244: signal is true;
	signal I15245: std_logic; attribute dont_touch of I15245: signal is true;
	signal I15246: std_logic; attribute dont_touch of I15246: signal is true;
	signal I15256: std_logic; attribute dont_touch of I15256: signal is true;
	signal I15262: std_logic; attribute dont_touch of I15262: signal is true;
	signal I15267: std_logic; attribute dont_touch of I15267: signal is true;
	signal I15271: std_logic; attribute dont_touch of I15271: signal is true;
	signal I15276: std_logic; attribute dont_touch of I15276: signal is true;
	signal I15277: std_logic; attribute dont_touch of I15277: signal is true;
	signal I15278: std_logic; attribute dont_touch of I15278: signal is true;
	signal I15288: std_logic; attribute dont_touch of I15288: signal is true;
	signal I15299: std_logic; attribute dont_touch of I15299: signal is true;
	signal I15304: std_logic; attribute dont_touch of I15304: signal is true;
	signal I15308: std_logic; attribute dont_touch of I15308: signal is true;
	signal I15313: std_logic; attribute dont_touch of I15313: signal is true;
	signal I15317: std_logic; attribute dont_touch of I15317: signal is true;
	signal I15326: std_logic; attribute dont_touch of I15326: signal is true;
	signal I15329: std_logic; attribute dont_touch of I15329: signal is true;
	signal I15345: std_logic; attribute dont_touch of I15345: signal is true;
	signal I15350: std_logic; attribute dont_touch of I15350: signal is true;
	signal I15354: std_logic; attribute dont_touch of I15354: signal is true;
	signal I15359: std_logic; attribute dont_touch of I15359: signal is true;
	signal I15369: std_logic; attribute dont_touch of I15369: signal is true;
	signal I15372: std_logic; attribute dont_touch of I15372: signal is true;
	signal I15392: std_logic; attribute dont_touch of I15392: signal is true;
	signal I15398: std_logic; attribute dont_touch of I15398: signal is true;
	signal I15429: std_logic; attribute dont_touch of I15429: signal is true;
	signal I15433: std_logic; attribute dont_touch of I15433: signal is true;
	signal I15442: std_logic; attribute dont_touch of I15442: signal is true;
	signal I15445: std_logic; attribute dont_touch of I15445: signal is true;
	signal I15448: std_logic; attribute dont_touch of I15448: signal is true;
	signal I15451: std_logic; attribute dont_touch of I15451: signal is true;
	signal I15454: std_logic; attribute dont_touch of I15454: signal is true;
	signal I15457: std_logic; attribute dont_touch of I15457: signal is true;
	signal I15460: std_logic; attribute dont_touch of I15460: signal is true;
	signal I15463: std_logic; attribute dont_touch of I15463: signal is true;
	signal I15466: std_logic; attribute dont_touch of I15466: signal is true;
	signal I15469: std_logic; attribute dont_touch of I15469: signal is true;
	signal I15472: std_logic; attribute dont_touch of I15472: signal is true;
	signal I15475: std_logic; attribute dont_touch of I15475: signal is true;
	signal I15478: std_logic; attribute dont_touch of I15478: signal is true;
	signal I15481: std_logic; attribute dont_touch of I15481: signal is true;
	signal I15484: std_logic; attribute dont_touch of I15484: signal is true;
	signal I15487: std_logic; attribute dont_touch of I15487: signal is true;
	signal I15490: std_logic; attribute dont_touch of I15490: signal is true;
	signal I15493: std_logic; attribute dont_touch of I15493: signal is true;
	signal I15499: std_logic; attribute dont_touch of I15499: signal is true;
	signal I15505: std_logic; attribute dont_touch of I15505: signal is true;
	signal I15511: std_logic; attribute dont_touch of I15511: signal is true;
	signal I15517: std_logic; attribute dont_touch of I15517: signal is true;
	signal I15523: std_logic; attribute dont_touch of I15523: signal is true;
	signal I15526: std_logic; attribute dont_touch of I15526: signal is true;
	signal I15532: std_logic; attribute dont_touch of I15532: signal is true;
	signal I15535: std_logic; attribute dont_touch of I15535: signal is true;
	signal I15538: std_logic; attribute dont_touch of I15538: signal is true;
	signal I15543: std_logic; attribute dont_touch of I15543: signal is true;
	signal I15546: std_logic; attribute dont_touch of I15546: signal is true;
	signal I15549: std_logic; attribute dont_touch of I15549: signal is true;
	signal I15553: std_logic; attribute dont_touch of I15553: signal is true;
	signal I15556: std_logic; attribute dont_touch of I15556: signal is true;
	signal I15559: std_logic; attribute dont_touch of I15559: signal is true;
	signal I15562: std_logic; attribute dont_touch of I15562: signal is true;
	signal I15565: std_logic; attribute dont_touch of I15565: signal is true;
	signal I15568: std_logic; attribute dont_touch of I15568: signal is true;
	signal I15571: std_logic; attribute dont_touch of I15571: signal is true;
	signal I15574: std_logic; attribute dont_touch of I15574: signal is true;
	signal I15577: std_logic; attribute dont_touch of I15577: signal is true;
	signal I15580: std_logic; attribute dont_touch of I15580: signal is true;
	signal I15584: std_logic; attribute dont_touch of I15584: signal is true;
	signal I15590: std_logic; attribute dont_touch of I15590: signal is true;
	signal I15593: std_logic; attribute dont_touch of I15593: signal is true;
	signal I15599: std_logic; attribute dont_touch of I15599: signal is true;
	signal I15602: std_logic; attribute dont_touch of I15602: signal is true;
	signal I15605: std_logic; attribute dont_touch of I15605: signal is true;
	signal I15610: std_logic; attribute dont_touch of I15610: signal is true;
	signal I15613: std_logic; attribute dont_touch of I15613: signal is true;
	signal I15616: std_logic; attribute dont_touch of I15616: signal is true;
	signal I15620: std_logic; attribute dont_touch of I15620: signal is true;
	signal I15623: std_logic; attribute dont_touch of I15623: signal is true;
	signal I15626: std_logic; attribute dont_touch of I15626: signal is true;
	signal I15629: std_logic; attribute dont_touch of I15629: signal is true;
	signal I15636: std_logic; attribute dont_touch of I15636: signal is true;
	signal I15642: std_logic; attribute dont_touch of I15642: signal is true;
	signal I15645: std_logic; attribute dont_touch of I15645: signal is true;
	signal I15651: std_logic; attribute dont_touch of I15651: signal is true;
	signal I15654: std_logic; attribute dont_touch of I15654: signal is true;
	signal I15657: std_logic; attribute dont_touch of I15657: signal is true;
	signal I15662: std_logic; attribute dont_touch of I15662: signal is true;
	signal I15671: std_logic; attribute dont_touch of I15671: signal is true;
	signal I15677: std_logic; attribute dont_touch of I15677: signal is true;
	signal I15680: std_logic; attribute dont_touch of I15680: signal is true;
	signal I15696: std_logic; attribute dont_touch of I15696: signal is true;
	signal I15771: std_logic; attribute dont_touch of I15771: signal is true;
	signal I15779: std_logic; attribute dont_touch of I15779: signal is true;
	signal I15784: std_logic; attribute dont_touch of I15784: signal is true;
	signal I15787: std_logic; attribute dont_touch of I15787: signal is true;
	signal I15794: std_logic; attribute dont_touch of I15794: signal is true;
	signal I15800: std_logic; attribute dont_touch of I15800: signal is true;
	signal I15803: std_logic; attribute dont_touch of I15803: signal is true;
	signal I15806: std_logic; attribute dont_touch of I15806: signal is true;
	signal I15810: std_logic; attribute dont_touch of I15810: signal is true;
	signal I15815: std_logic; attribute dont_touch of I15815: signal is true;
	signal I15818: std_logic; attribute dont_touch of I15818: signal is true;
	signal I15822: std_logic; attribute dont_touch of I15822: signal is true;
	signal I15827: std_logic; attribute dont_touch of I15827: signal is true;
	signal I15830: std_logic; attribute dont_touch of I15830: signal is true;
	signal I15833: std_logic; attribute dont_touch of I15833: signal is true;
	signal I15836: std_logic; attribute dont_touch of I15836: signal is true;
	signal I15839: std_logic; attribute dont_touch of I15839: signal is true;
	signal I15843: std_logic; attribute dont_touch of I15843: signal is true;
	signal I15847: std_logic; attribute dont_touch of I15847: signal is true;
	signal I15850: std_logic; attribute dont_touch of I15850: signal is true;
	signal I15853: std_logic; attribute dont_touch of I15853: signal is true;
	signal I15856: std_logic; attribute dont_touch of I15856: signal is true;
	signal I15859: std_logic; attribute dont_touch of I15859: signal is true;
	signal I15863: std_logic; attribute dont_touch of I15863: signal is true;
	signal I15866: std_logic; attribute dont_touch of I15866: signal is true;
	signal I15869: std_logic; attribute dont_touch of I15869: signal is true;
	signal I15873: std_logic; attribute dont_touch of I15873: signal is true;
	signal I15876: std_logic; attribute dont_touch of I15876: signal is true;
	signal I15879: std_logic; attribute dont_touch of I15879: signal is true;
	signal I15882: std_logic; attribute dont_touch of I15882: signal is true;
	signal I15887: std_logic; attribute dont_touch of I15887: signal is true;
	signal I15890: std_logic; attribute dont_touch of I15890: signal is true;
	signal I15893: std_logic; attribute dont_touch of I15893: signal is true;
	signal I15896: std_logic; attribute dont_touch of I15896: signal is true;
	signal I15899: std_logic; attribute dont_touch of I15899: signal is true;
	signal I15902: std_logic; attribute dont_touch of I15902: signal is true;
	signal I15909: std_logic; attribute dont_touch of I15909: signal is true;
	signal I15912: std_logic; attribute dont_touch of I15912: signal is true;
	signal I15915: std_logic; attribute dont_touch of I15915: signal is true;
	signal I15918: std_logic; attribute dont_touch of I15918: signal is true;
	signal I15922: std_logic; attribute dont_touch of I15922: signal is true;
	signal I15925: std_logic; attribute dont_touch of I15925: signal is true;
	signal I15932: std_logic; attribute dont_touch of I15932: signal is true;
	signal I15935: std_logic; attribute dont_touch of I15935: signal is true;
	signal I15938: std_logic; attribute dont_touch of I15938: signal is true;
	signal I15942: std_logic; attribute dont_touch of I15942: signal is true;
	signal I15946: std_logic; attribute dont_touch of I15946: signal is true;
	signal I15949: std_logic; attribute dont_touch of I15949: signal is true;
	signal I15955: std_logic; attribute dont_touch of I15955: signal is true;
	signal I15958: std_logic; attribute dont_touch of I15958: signal is true;
	signal I15961: std_logic; attribute dont_touch of I15961: signal is true;
	signal I15964: std_logic; attribute dont_touch of I15964: signal is true;
	signal I15967: std_logic; attribute dont_touch of I15967: signal is true;
	signal I15971: std_logic; attribute dont_touch of I15971: signal is true;
	signal I15975: std_logic; attribute dont_touch of I15975: signal is true;
	signal I15978: std_logic; attribute dont_touch of I15978: signal is true;
	signal I15983: std_logic; attribute dont_touch of I15983: signal is true;
	signal I15986: std_logic; attribute dont_touch of I15986: signal is true;
	signal I15989: std_logic; attribute dont_touch of I15989: signal is true;
	signal I15992: std_logic; attribute dont_touch of I15992: signal is true;
	signal I15995: std_logic; attribute dont_touch of I15995: signal is true;
	signal I15998: std_logic; attribute dont_touch of I15998: signal is true;
	signal I16002: std_logic; attribute dont_touch of I16002: signal is true;
	signal I16006: std_logic; attribute dont_touch of I16006: signal is true;
	signal I16009: std_logic; attribute dont_touch of I16009: signal is true;
	signal I16012: std_logic; attribute dont_touch of I16012: signal is true;
	signal I16015: std_logic; attribute dont_touch of I16015: signal is true;
	signal I16018: std_logic; attribute dont_touch of I16018: signal is true;
	signal I16021: std_logic; attribute dont_touch of I16021: signal is true;
	signal I16024: std_logic; attribute dont_touch of I16024: signal is true;
	signal I16027: std_logic; attribute dont_touch of I16027: signal is true;
	signal I16031: std_logic; attribute dont_touch of I16031: signal is true;
	signal I16034: std_logic; attribute dont_touch of I16034: signal is true;
	signal I16037: std_logic; attribute dont_touch of I16037: signal is true;
	signal I16041: std_logic; attribute dont_touch of I16041: signal is true;
	signal I16044: std_logic; attribute dont_touch of I16044: signal is true;
	signal I16047: std_logic; attribute dont_touch of I16047: signal is true;
	signal I16050: std_logic; attribute dont_touch of I16050: signal is true;
	signal I16053: std_logic; attribute dont_touch of I16053: signal is true;
	signal I16056: std_logic; attribute dont_touch of I16056: signal is true;
	signal I16059: std_logic; attribute dont_touch of I16059: signal is true;
	signal I16062: std_logic; attribute dont_touch of I16062: signal is true;
	signal I16065: std_logic; attribute dont_touch of I16065: signal is true;
	signal I16068: std_logic; attribute dont_touch of I16068: signal is true;
	signal I16071: std_logic; attribute dont_touch of I16071: signal is true;
	signal I16074: std_logic; attribute dont_touch of I16074: signal is true;
	signal I16079: std_logic; attribute dont_touch of I16079: signal is true;
	signal I16082: std_logic; attribute dont_touch of I16082: signal is true;
	signal I16085: std_logic; attribute dont_touch of I16085: signal is true;
	signal I16089: std_logic; attribute dont_touch of I16089: signal is true;
	signal I16092: std_logic; attribute dont_touch of I16092: signal is true;
	signal I16095: std_logic; attribute dont_touch of I16095: signal is true;
	signal I16098: std_logic; attribute dont_touch of I16098: signal is true;
	signal I16101: std_logic; attribute dont_touch of I16101: signal is true;
	signal I16104: std_logic; attribute dont_touch of I16104: signal is true;
	signal I16107: std_logic; attribute dont_touch of I16107: signal is true;
	signal I16110: std_logic; attribute dont_touch of I16110: signal is true;
	signal I16114: std_logic; attribute dont_touch of I16114: signal is true;
	signal I16117: std_logic; attribute dont_touch of I16117: signal is true;
	signal I16120: std_logic; attribute dont_touch of I16120: signal is true;
	signal I16123: std_logic; attribute dont_touch of I16123: signal is true;
	signal I16128: std_logic; attribute dont_touch of I16128: signal is true;
	signal I16131: std_logic; attribute dont_touch of I16131: signal is true;
	signal I16134: std_logic; attribute dont_touch of I16134: signal is true;
	signal I16138: std_logic; attribute dont_touch of I16138: signal is true;
	signal I16141: std_logic; attribute dont_touch of I16141: signal is true;
	signal I16144: std_logic; attribute dont_touch of I16144: signal is true;
	signal I16147: std_logic; attribute dont_touch of I16147: signal is true;
	signal I16150: std_logic; attribute dont_touch of I16150: signal is true;
	signal I16153: std_logic; attribute dont_touch of I16153: signal is true;
	signal I16156: std_logic; attribute dont_touch of I16156: signal is true;
	signal I16159: std_logic; attribute dont_touch of I16159: signal is true;
	signal I16163: std_logic; attribute dont_touch of I16163: signal is true;
	signal I16166: std_logic; attribute dont_touch of I16166: signal is true;
	signal I16169: std_logic; attribute dont_touch of I16169: signal is true;
	signal I16172: std_logic; attribute dont_touch of I16172: signal is true;
	signal I16176: std_logic; attribute dont_touch of I16176: signal is true;
	signal I16179: std_logic; attribute dont_touch of I16179: signal is true;
	signal I16182: std_logic; attribute dont_touch of I16182: signal is true;
	signal I16185: std_logic; attribute dont_touch of I16185: signal is true;
	signal I16190: std_logic; attribute dont_touch of I16190: signal is true;
	signal I16193: std_logic; attribute dont_touch of I16193: signal is true;
	signal I16196: std_logic; attribute dont_touch of I16196: signal is true;
	signal I16200: std_logic; attribute dont_touch of I16200: signal is true;
	signal I16203: std_logic; attribute dont_touch of I16203: signal is true;
	signal I16206: std_logic; attribute dont_touch of I16206: signal is true;
	signal I16209: std_logic; attribute dont_touch of I16209: signal is true;
	signal I16212: std_logic; attribute dont_touch of I16212: signal is true;
	signal I16215: std_logic; attribute dont_touch of I16215: signal is true;
	signal I16218: std_logic; attribute dont_touch of I16218: signal is true;
	signal I16221: std_logic; attribute dont_touch of I16221: signal is true;
	signal I16225: std_logic; attribute dont_touch of I16225: signal is true;
	signal I16228: std_logic; attribute dont_touch of I16228: signal is true;
	signal I16231: std_logic; attribute dont_touch of I16231: signal is true;
	signal I16234: std_logic; attribute dont_touch of I16234: signal is true;
	signal I16238: std_logic; attribute dont_touch of I16238: signal is true;
	signal I16241: std_logic; attribute dont_touch of I16241: signal is true;
	signal I16244: std_logic; attribute dont_touch of I16244: signal is true;
	signal I16247: std_logic; attribute dont_touch of I16247: signal is true;
	signal I16252: std_logic; attribute dont_touch of I16252: signal is true;
	signal I16255: std_logic; attribute dont_touch of I16255: signal is true;
	signal I16258: std_logic; attribute dont_touch of I16258: signal is true;
	signal I16261: std_logic; attribute dont_touch of I16261: signal is true;
	signal I16264: std_logic; attribute dont_touch of I16264: signal is true;
	signal I16267: std_logic; attribute dont_touch of I16267: signal is true;
	signal I16270: std_logic; attribute dont_touch of I16270: signal is true;
	signal I16273: std_logic; attribute dont_touch of I16273: signal is true;
	signal I16276: std_logic; attribute dont_touch of I16276: signal is true;
	signal I16279: std_logic; attribute dont_touch of I16279: signal is true;
	signal I16283: std_logic; attribute dont_touch of I16283: signal is true;
	signal I16286: std_logic; attribute dont_touch of I16286: signal is true;
	signal I16289: std_logic; attribute dont_touch of I16289: signal is true;
	signal I16292: std_logic; attribute dont_touch of I16292: signal is true;
	signal I16296: std_logic; attribute dont_touch of I16296: signal is true;
	signal I16300: std_logic; attribute dont_touch of I16300: signal is true;
	signal I16303: std_logic; attribute dont_touch of I16303: signal is true;
	signal I16306: std_logic; attribute dont_touch of I16306: signal is true;
	signal I16309: std_logic; attribute dont_touch of I16309: signal is true;
	signal I16312: std_logic; attribute dont_touch of I16312: signal is true;
	signal I16315: std_logic; attribute dont_touch of I16315: signal is true;
	signal I16318: std_logic; attribute dont_touch of I16318: signal is true;
	signal I16321: std_logic; attribute dont_touch of I16321: signal is true;
	signal I16325: std_logic; attribute dont_touch of I16325: signal is true;
	signal I16328: std_logic; attribute dont_touch of I16328: signal is true;
	signal I16332: std_logic; attribute dont_touch of I16332: signal is true;
	signal I16335: std_logic; attribute dont_touch of I16335: signal is true;
	signal I16338: std_logic; attribute dont_touch of I16338: signal is true;
	signal I16341: std_logic; attribute dont_touch of I16341: signal is true;
	signal I16344: std_logic; attribute dont_touch of I16344: signal is true;
	signal I16347: std_logic; attribute dont_touch of I16347: signal is true;
	signal I16354: std_logic; attribute dont_touch of I16354: signal is true;
	signal I16357: std_logic; attribute dont_touch of I16357: signal is true;
	signal I16360: std_logic; attribute dont_touch of I16360: signal is true;
	signal I16363: std_logic; attribute dont_touch of I16363: signal is true;
	signal I16372: std_logic; attribute dont_touch of I16372: signal is true;
	signal I16432: std_logic; attribute dont_touch of I16432: signal is true;
	signal I16438: std_logic; attribute dont_touch of I16438: signal is true;
	signal I16444: std_logic; attribute dont_touch of I16444: signal is true;
	signal I16450: std_logic; attribute dont_touch of I16450: signal is true;
	signal I16453: std_logic; attribute dont_touch of I16453: signal is true;
	signal I16457: std_logic; attribute dont_touch of I16457: signal is true;
	signal I16462: std_logic; attribute dont_touch of I16462: signal is true;
	signal I16465: std_logic; attribute dont_touch of I16465: signal is true;
	signal I16469: std_logic; attribute dont_touch of I16469: signal is true;
	signal I16472: std_logic; attribute dont_touch of I16472: signal is true;
	signal I16476: std_logic; attribute dont_touch of I16476: signal is true;
	signal I16479: std_logic; attribute dont_touch of I16479: signal is true;
	signal I16482: std_logic; attribute dont_touch of I16482: signal is true;
	signal I16486: std_logic; attribute dont_touch of I16486: signal is true;
	signal I16489: std_logic; attribute dont_touch of I16489: signal is true;
	signal I16493: std_logic; attribute dont_touch of I16493: signal is true;
	signal I16499: std_logic; attribute dont_touch of I16499: signal is true;
	signal I16504: std_logic; attribute dont_touch of I16504: signal is true;
	signal I16507: std_logic; attribute dont_touch of I16507: signal is true;
	signal I16511: std_logic; attribute dont_touch of I16511: signal is true;
	signal I16514: std_logic; attribute dont_touch of I16514: signal is true;
	signal I16517: std_logic; attribute dont_touch of I16517: signal is true;
	signal I16521: std_logic; attribute dont_touch of I16521: signal is true;
	signal I16524: std_logic; attribute dont_touch of I16524: signal is true;
	signal I16532: std_logic; attribute dont_touch of I16532: signal is true;
	signal I16538: std_logic; attribute dont_touch of I16538: signal is true;
	signal I16541: std_logic; attribute dont_touch of I16541: signal is true;
	signal I16544: std_logic; attribute dont_touch of I16544: signal is true;
	signal I16549: std_logic; attribute dont_touch of I16549: signal is true;
	signal I16552: std_logic; attribute dont_touch of I16552: signal is true;
	signal I16556: std_logic; attribute dont_touch of I16556: signal is true;
	signal I16559: std_logic; attribute dont_touch of I16559: signal is true;
	signal I16562: std_logic; attribute dont_touch of I16562: signal is true;
	signal I16566: std_logic; attribute dont_touch of I16566: signal is true;
	signal I16569: std_logic; attribute dont_touch of I16569: signal is true;
	signal I16578: std_logic; attribute dont_touch of I16578: signal is true;
	signal I16581: std_logic; attribute dont_touch of I16581: signal is true;
	signal I16587: std_logic; attribute dont_touch of I16587: signal is true;
	signal I16590: std_logic; attribute dont_touch of I16590: signal is true;
	signal I16593: std_logic; attribute dont_touch of I16593: signal is true;
	signal I16598: std_logic; attribute dont_touch of I16598: signal is true;
	signal I16601: std_logic; attribute dont_touch of I16601: signal is true;
	signal I16605: std_logic; attribute dont_touch of I16605: signal is true;
	signal I16608: std_logic; attribute dont_touch of I16608: signal is true;
	signal I16611: std_logic; attribute dont_touch of I16611: signal is true;
	signal I16624: std_logic; attribute dont_touch of I16624: signal is true;
	signal I16627: std_logic; attribute dont_touch of I16627: signal is true;
	signal I16630: std_logic; attribute dont_touch of I16630: signal is true;
	signal I16633: std_logic; attribute dont_touch of I16633: signal is true;
	signal I16641: std_logic; attribute dont_touch of I16641: signal is true;
	signal I16644: std_logic; attribute dont_touch of I16644: signal is true;
	signal I16650: std_logic; attribute dont_touch of I16650: signal is true;
	signal I16653: std_logic; attribute dont_touch of I16653: signal is true;
	signal I16656: std_logic; attribute dont_touch of I16656: signal is true;
	signal I16661: std_logic; attribute dont_touch of I16661: signal is true;
	signal I16664: std_logic; attribute dont_touch of I16664: signal is true;
	signal I16677: std_logic; attribute dont_touch of I16677: signal is true;
	signal I16681: std_logic; attribute dont_touch of I16681: signal is true;
	signal I16684: std_logic; attribute dont_touch of I16684: signal is true;
	signal I16694: std_logic; attribute dont_touch of I16694: signal is true;
	signal I16697: std_logic; attribute dont_touch of I16697: signal is true;
	signal I16700: std_logic; attribute dont_touch of I16700: signal is true;
	signal I16703: std_logic; attribute dont_touch of I16703: signal is true;
	signal I16711: std_logic; attribute dont_touch of I16711: signal is true;
	signal I16714: std_logic; attribute dont_touch of I16714: signal is true;
	signal I16720: std_logic; attribute dont_touch of I16720: signal is true;
	signal I16723: std_logic; attribute dont_touch of I16723: signal is true;
	signal I16726: std_logic; attribute dont_touch of I16726: signal is true;
	signal I16735: std_logic; attribute dont_touch of I16735: signal is true;
	signal I16736: std_logic; attribute dont_touch of I16736: signal is true;
	signal I16741: std_logic; attribute dont_touch of I16741: signal is true;
	signal I16744: std_logic; attribute dont_touch of I16744: signal is true;
	signal I16747: std_logic; attribute dont_touch of I16747: signal is true;
	signal I16759: std_logic; attribute dont_touch of I16759: signal is true;
	signal I16763: std_logic; attribute dont_touch of I16763: signal is true;
	signal I16766: std_logic; attribute dont_touch of I16766: signal is true;
	signal I16776: std_logic; attribute dont_touch of I16776: signal is true;
	signal I16779: std_logic; attribute dont_touch of I16779: signal is true;
	signal I16782: std_logic; attribute dont_touch of I16782: signal is true;
	signal I16785: std_logic; attribute dont_touch of I16785: signal is true;
	signal I16793: std_logic; attribute dont_touch of I16793: signal is true;
	signal I16796: std_logic; attribute dont_touch of I16796: signal is true;
	signal I16811: std_logic; attribute dont_touch of I16811: signal is true;
	signal I16814: std_logic; attribute dont_touch of I16814: signal is true;
	signal I16826: std_logic; attribute dont_touch of I16826: signal is true;
	signal I16827: std_logic; attribute dont_touch of I16827: signal is true;
	signal I16832: std_logic; attribute dont_touch of I16832: signal is true;
	signal I16835: std_logic; attribute dont_touch of I16835: signal is true;
	signal I16838: std_logic; attribute dont_touch of I16838: signal is true;
	signal I16850: std_logic; attribute dont_touch of I16850: signal is true;
	signal I16854: std_logic; attribute dont_touch of I16854: signal is true;
	signal I16857: std_logic; attribute dont_touch of I16857: signal is true;
	signal I16867: std_logic; attribute dont_touch of I16867: signal is true;
	signal I16870: std_logic; attribute dont_touch of I16870: signal is true;
	signal I16873: std_logic; attribute dont_touch of I16873: signal is true;
	signal I16876: std_logic; attribute dont_touch of I16876: signal is true;
	signal I16879: std_logic; attribute dont_touch of I16879: signal is true;
	signal I16880: std_logic; attribute dont_touch of I16880: signal is true;
	signal I16881: std_logic; attribute dont_touch of I16881: signal is true;
	signal I16897: std_logic; attribute dont_touch of I16897: signal is true;
	signal I16900: std_logic; attribute dont_touch of I16900: signal is true;
	signal I16915: std_logic; attribute dont_touch of I16915: signal is true;
	signal I16918: std_logic; attribute dont_touch of I16918: signal is true;
	signal I16930: std_logic; attribute dont_touch of I16930: signal is true;
	signal I16931: std_logic; attribute dont_touch of I16931: signal is true;
	signal I16936: std_logic; attribute dont_touch of I16936: signal is true;
	signal I16939: std_logic; attribute dont_touch of I16939: signal is true;
	signal I16942: std_logic; attribute dont_touch of I16942: signal is true;
	signal I16954: std_logic; attribute dont_touch of I16954: signal is true;
	signal I16958: std_logic; attribute dont_touch of I16958: signal is true;
	signal I16961: std_logic; attribute dont_touch of I16961: signal is true;
	signal I16965: std_logic; attribute dont_touch of I16965: signal is true;
	signal I16966: std_logic; attribute dont_touch of I16966: signal is true;
	signal I16967: std_logic; attribute dont_touch of I16967: signal is true;
	signal I16972: std_logic; attribute dont_touch of I16972: signal is true;
	signal I16984: std_logic; attribute dont_touch of I16984: signal is true;
	signal I16987: std_logic; attribute dont_touch of I16987: signal is true;
	signal I16990: std_logic; attribute dont_touch of I16990: signal is true;
	signal I16993: std_logic; attribute dont_touch of I16993: signal is true;
	signal I17009: std_logic; attribute dont_touch of I17009: signal is true;
	signal I17012: std_logic; attribute dont_touch of I17012: signal is true;
	signal I17027: std_logic; attribute dont_touch of I17027: signal is true;
	signal I17030: std_logic; attribute dont_touch of I17030: signal is true;
	signal I17042: std_logic; attribute dont_touch of I17042: signal is true;
	signal I17043: std_logic; attribute dont_touch of I17043: signal is true;
	signal I17048: std_logic; attribute dont_touch of I17048: signal is true;
	signal I17051: std_logic; attribute dont_touch of I17051: signal is true;
	signal I17054: std_logic; attribute dont_touch of I17054: signal is true;
	signal I17059: std_logic; attribute dont_touch of I17059: signal is true;
	signal I17060: std_logic; attribute dont_touch of I17060: signal is true;
	signal I17061: std_logic; attribute dont_touch of I17061: signal is true;
	signal I17066: std_logic; attribute dont_touch of I17066: signal is true;
	signal I17070: std_logic; attribute dont_touch of I17070: signal is true;
	signal I17081: std_logic; attribute dont_touch of I17081: signal is true;
	signal I17097: std_logic; attribute dont_touch of I17097: signal is true;
	signal I17100: std_logic; attribute dont_touch of I17100: signal is true;
	signal I17103: std_logic; attribute dont_touch of I17103: signal is true;
	signal I17106: std_logic; attribute dont_touch of I17106: signal is true;
	signal I17122: std_logic; attribute dont_touch of I17122: signal is true;
	signal I17125: std_logic; attribute dont_touch of I17125: signal is true;
	signal I17140: std_logic; attribute dont_touch of I17140: signal is true;
	signal I17143: std_logic; attribute dont_touch of I17143: signal is true;
	signal I17149: std_logic; attribute dont_touch of I17149: signal is true;
	signal I17150: std_logic; attribute dont_touch of I17150: signal is true;
	signal I17151: std_logic; attribute dont_touch of I17151: signal is true;
	signal I17156: std_logic; attribute dont_touch of I17156: signal is true;
	signal I17159: std_logic; attribute dont_touch of I17159: signal is true;
	signal I17184: std_logic; attribute dont_touch of I17184: signal is true;
	signal I17200: std_logic; attribute dont_touch of I17200: signal is true;
	signal I17203: std_logic; attribute dont_touch of I17203: signal is true;
	signal I17206: std_logic; attribute dont_touch of I17206: signal is true;
	signal I17209: std_logic; attribute dont_touch of I17209: signal is true;
	signal I17225: std_logic; attribute dont_touch of I17225: signal is true;
	signal I17228: std_logic; attribute dont_touch of I17228: signal is true;
	signal I17235: std_logic; attribute dont_touch of I17235: signal is true;
	signal I17238: std_logic; attribute dont_touch of I17238: signal is true;
	signal I17278: std_logic; attribute dont_touch of I17278: signal is true;
	signal I17294: std_logic; attribute dont_touch of I17294: signal is true;
	signal I17297: std_logic; attribute dont_touch of I17297: signal is true;
	signal I17300: std_logic; attribute dont_touch of I17300: signal is true;
	signal I17303: std_logic; attribute dont_touch of I17303: signal is true;
	signal I17311: std_logic; attribute dont_touch of I17311: signal is true;
	signal I17363: std_logic; attribute dont_touch of I17363: signal is true;
	signal I17370: std_logic; attribute dont_touch of I17370: signal is true;
	signal I17373: std_logic; attribute dont_touch of I17373: signal is true;
	signal I17429: std_logic; attribute dont_touch of I17429: signal is true;
	signal I17433: std_logic; attribute dont_touch of I17433: signal is true;
	signal I17483: std_logic; attribute dont_touch of I17483: signal is true;
	signal I17486: std_logic; attribute dont_touch of I17486: signal is true;
	signal I17527: std_logic; attribute dont_touch of I17527: signal is true;
	signal I17557: std_logic; attribute dont_touch of I17557: signal is true;
	signal I17599: std_logic; attribute dont_touch of I17599: signal is true;
	signal I17627: std_logic; attribute dont_touch of I17627: signal is true;
	signal I17632: std_logic; attribute dont_touch of I17632: signal is true;
	signal I17637: std_logic; attribute dont_touch of I17637: signal is true;
	signal I17641: std_logic; attribute dont_touch of I17641: signal is true;
	signal I17645: std_logic; attribute dont_touch of I17645: signal is true;
	signal I17649: std_logic; attribute dont_touch of I17649: signal is true;
	signal I17653: std_logic; attribute dont_touch of I17653: signal is true;
	signal I17658: std_logic; attribute dont_touch of I17658: signal is true;
	signal I17662: std_logic; attribute dont_touch of I17662: signal is true;
	signal I17666: std_logic; attribute dont_touch of I17666: signal is true;
	signal I17670: std_logic; attribute dont_touch of I17670: signal is true;
	signal I17673: std_logic; attribute dont_touch of I17673: signal is true;
	signal I17677: std_logic; attribute dont_touch of I17677: signal is true;
	signal I17681: std_logic; attribute dont_touch of I17681: signal is true;
	signal I17685: std_logic; attribute dont_touch of I17685: signal is true;
	signal I17689: std_logic; attribute dont_touch of I17689: signal is true;
	signal I17692: std_logic; attribute dont_touch of I17692: signal is true;
	signal I17698: std_logic; attribute dont_touch of I17698: signal is true;
	signal I17701: std_logic; attribute dont_touch of I17701: signal is true;
	signal I17705: std_logic; attribute dont_touch of I17705: signal is true;
	signal I17709: std_logic; attribute dont_touch of I17709: signal is true;
	signal I17712: std_logic; attribute dont_touch of I17712: signal is true;
	signal I17715: std_logic; attribute dont_touch of I17715: signal is true;
	signal I17721: std_logic; attribute dont_touch of I17721: signal is true;
	signal I17724: std_logic; attribute dont_touch of I17724: signal is true;
	signal I17727: std_logic; attribute dont_touch of I17727: signal is true;
	signal I17730: std_logic; attribute dont_touch of I17730: signal is true;
	signal I17734: std_logic; attribute dont_touch of I17734: signal is true;
	signal I17737: std_logic; attribute dont_touch of I17737: signal is true;
	signal I17740: std_logic; attribute dont_touch of I17740: signal is true;
	signal I17743: std_logic; attribute dont_touch of I17743: signal is true;
	signal I17746: std_logic; attribute dont_touch of I17746: signal is true;
	signal I17750: std_logic; attribute dont_touch of I17750: signal is true;
	signal I17753: std_logic; attribute dont_touch of I17753: signal is true;
	signal I17756: std_logic; attribute dont_touch of I17756: signal is true;
	signal I17759: std_logic; attribute dont_touch of I17759: signal is true;
	signal I17762: std_logic; attribute dont_touch of I17762: signal is true;
	signal I17765: std_logic; attribute dont_touch of I17765: signal is true;
	signal I17768: std_logic; attribute dont_touch of I17768: signal is true;
	signal I17771: std_logic; attribute dont_touch of I17771: signal is true;
	signal I17774: std_logic; attribute dont_touch of I17774: signal is true;
	signal I17780: std_logic; attribute dont_touch of I17780: signal is true;
	signal I17783: std_logic; attribute dont_touch of I17783: signal is true;
	signal I17786: std_logic; attribute dont_touch of I17786: signal is true;
	signal I17789: std_logic; attribute dont_touch of I17789: signal is true;
	signal I17792: std_logic; attribute dont_touch of I17792: signal is true;
	signal I17795: std_logic; attribute dont_touch of I17795: signal is true;
	signal I17798: std_logic; attribute dont_touch of I17798: signal is true;
	signal I17801: std_logic; attribute dont_touch of I17801: signal is true;
	signal I17804: std_logic; attribute dont_touch of I17804: signal is true;
	signal I17807: std_logic; attribute dont_touch of I17807: signal is true;
	signal I17813: std_logic; attribute dont_touch of I17813: signal is true;
	signal I17816: std_logic; attribute dont_touch of I17816: signal is true;
	signal I17819: std_logic; attribute dont_touch of I17819: signal is true;
	signal I17822: std_logic; attribute dont_touch of I17822: signal is true;
	signal I17825: std_logic; attribute dont_touch of I17825: signal is true;
	signal I17828: std_logic; attribute dont_touch of I17828: signal is true;
	signal I17831: std_logic; attribute dont_touch of I17831: signal is true;
	signal I17834: std_logic; attribute dont_touch of I17834: signal is true;
	signal I17837: std_logic; attribute dont_touch of I17837: signal is true;
	signal I17840: std_logic; attribute dont_touch of I17840: signal is true;
	signal I17843: std_logic; attribute dont_touch of I17843: signal is true;
	signal I17846: std_logic; attribute dont_touch of I17846: signal is true;
	signal I17849: std_logic; attribute dont_touch of I17849: signal is true;
	signal I17854: std_logic; attribute dont_touch of I17854: signal is true;
	signal I17857: std_logic; attribute dont_touch of I17857: signal is true;
	signal I17860: std_logic; attribute dont_touch of I17860: signal is true;
	signal I17863: std_logic; attribute dont_touch of I17863: signal is true;
	signal I17866: std_logic; attribute dont_touch of I17866: signal is true;
	signal I17869: std_logic; attribute dont_touch of I17869: signal is true;
	signal I17872: std_logic; attribute dont_touch of I17872: signal is true;
	signal I17875: std_logic; attribute dont_touch of I17875: signal is true;
	signal I17878: std_logic; attribute dont_touch of I17878: signal is true;
	signal I17881: std_logic; attribute dont_touch of I17881: signal is true;
	signal I17884: std_logic; attribute dont_touch of I17884: signal is true;
	signal I17889: std_logic; attribute dont_touch of I17889: signal is true;
	signal I17892: std_logic; attribute dont_touch of I17892: signal is true;
	signal I17895: std_logic; attribute dont_touch of I17895: signal is true;
	signal I17898: std_logic; attribute dont_touch of I17898: signal is true;
	signal I17901: std_logic; attribute dont_touch of I17901: signal is true;
	signal I17904: std_logic; attribute dont_touch of I17904: signal is true;
	signal I17907: std_logic; attribute dont_touch of I17907: signal is true;
	signal I17910: std_logic; attribute dont_touch of I17910: signal is true;
	signal I17913: std_logic; attribute dont_touch of I17913: signal is true;
	signal I17916: std_logic; attribute dont_touch of I17916: signal is true;
	signal I17919: std_logic; attribute dont_touch of I17919: signal is true;
	signal I17922: std_logic; attribute dont_touch of I17922: signal is true;
	signal I17925: std_logic; attribute dont_touch of I17925: signal is true;
	signal I17928: std_logic; attribute dont_touch of I17928: signal is true;
	signal I17933: std_logic; attribute dont_touch of I17933: signal is true;
	signal I17936: std_logic; attribute dont_touch of I17936: signal is true;
	signal I17939: std_logic; attribute dont_touch of I17939: signal is true;
	signal I17942: std_logic; attribute dont_touch of I17942: signal is true;
	signal I17945: std_logic; attribute dont_touch of I17945: signal is true;
	signal I17948: std_logic; attribute dont_touch of I17948: signal is true;
	signal I17951: std_logic; attribute dont_touch of I17951: signal is true;
	signal I17954: std_logic; attribute dont_touch of I17954: signal is true;
	signal I17957: std_logic; attribute dont_touch of I17957: signal is true;
	signal I17960: std_logic; attribute dont_touch of I17960: signal is true;
	signal I17963: std_logic; attribute dont_touch of I17963: signal is true;
	signal I17966: std_logic; attribute dont_touch of I17966: signal is true;
	signal I17969: std_logic; attribute dont_touch of I17969: signal is true;
	signal I17972: std_logic; attribute dont_touch of I17972: signal is true;
	signal I17975: std_logic; attribute dont_touch of I17975: signal is true;
	signal I17978: std_logic; attribute dont_touch of I17978: signal is true;
	signal I17981: std_logic; attribute dont_touch of I17981: signal is true;
	signal I17984: std_logic; attribute dont_touch of I17984: signal is true;
	signal I17989: std_logic; attribute dont_touch of I17989: signal is true;
	signal I17992: std_logic; attribute dont_touch of I17992: signal is true;
	signal I17995: std_logic; attribute dont_touch of I17995: signal is true;
	signal I17998: std_logic; attribute dont_touch of I17998: signal is true;
	signal I18001: std_logic; attribute dont_touch of I18001: signal is true;
	signal I18004: std_logic; attribute dont_touch of I18004: signal is true;
	signal I18007: std_logic; attribute dont_touch of I18007: signal is true;
	signal I18010: std_logic; attribute dont_touch of I18010: signal is true;
	signal I18013: std_logic; attribute dont_touch of I18013: signal is true;
	signal I18016: std_logic; attribute dont_touch of I18016: signal is true;
	signal I18019: std_logic; attribute dont_touch of I18019: signal is true;
	signal I18022: std_logic; attribute dont_touch of I18022: signal is true;
	signal I18025: std_logic; attribute dont_touch of I18025: signal is true;
	signal I18028: std_logic; attribute dont_touch of I18028: signal is true;
	signal I18031: std_logic; attribute dont_touch of I18031: signal is true;
	signal I18034: std_logic; attribute dont_touch of I18034: signal is true;
	signal I18037: std_logic; attribute dont_touch of I18037: signal is true;
	signal I18040: std_logic; attribute dont_touch of I18040: signal is true;
	signal I18043: std_logic; attribute dont_touch of I18043: signal is true;
	signal I18046: std_logic; attribute dont_touch of I18046: signal is true;
	signal I18049: std_logic; attribute dont_touch of I18049: signal is true;
	signal I18052: std_logic; attribute dont_touch of I18052: signal is true;
	signal I18055: std_logic; attribute dont_touch of I18055: signal is true;
	signal I18058: std_logic; attribute dont_touch of I18058: signal is true;
	signal I18061: std_logic; attribute dont_touch of I18061: signal is true;
	signal I18064: std_logic; attribute dont_touch of I18064: signal is true;
	signal I18067: std_logic; attribute dont_touch of I18067: signal is true;
	signal I18070: std_logic; attribute dont_touch of I18070: signal is true;
	signal I18073: std_logic; attribute dont_touch of I18073: signal is true;
	signal I18076: std_logic; attribute dont_touch of I18076: signal is true;
	signal I18079: std_logic; attribute dont_touch of I18079: signal is true;
	signal I18082: std_logic; attribute dont_touch of I18082: signal is true;
	signal I18085: std_logic; attribute dont_touch of I18085: signal is true;
	signal I18088: std_logic; attribute dont_touch of I18088: signal is true;
	signal I18091: std_logic; attribute dont_touch of I18091: signal is true;
	signal I18094: std_logic; attribute dont_touch of I18094: signal is true;
	signal I18097: std_logic; attribute dont_touch of I18097: signal is true;
	signal I18100: std_logic; attribute dont_touch of I18100: signal is true;
	signal I18103: std_logic; attribute dont_touch of I18103: signal is true;
	signal I18106: std_logic; attribute dont_touch of I18106: signal is true;
	signal I18107: std_logic; attribute dont_touch of I18107: signal is true;
	signal I18108: std_logic; attribute dont_touch of I18108: signal is true;
	signal I18113: std_logic; attribute dont_touch of I18113: signal is true;
	signal I18114: std_logic; attribute dont_touch of I18114: signal is true;
	signal I18115: std_logic; attribute dont_touch of I18115: signal is true;
	signal I18121: std_logic; attribute dont_touch of I18121: signal is true;
	signal I18124: std_logic; attribute dont_touch of I18124: signal is true;
	signal I18127: std_logic; attribute dont_touch of I18127: signal is true;
	signal I18130: std_logic; attribute dont_touch of I18130: signal is true;
	signal I18133: std_logic; attribute dont_touch of I18133: signal is true;
	signal I18136: std_logic; attribute dont_touch of I18136: signal is true;
	signal I18139: std_logic; attribute dont_touch of I18139: signal is true;
	signal I18142: std_logic; attribute dont_touch of I18142: signal is true;
	signal I18145: std_logic; attribute dont_touch of I18145: signal is true;
	signal I18148: std_logic; attribute dont_touch of I18148: signal is true;
	signal I18151: std_logic; attribute dont_touch of I18151: signal is true;
	signal I18154: std_logic; attribute dont_touch of I18154: signal is true;
	signal I18157: std_logic; attribute dont_touch of I18157: signal is true;
	signal I18160: std_logic; attribute dont_touch of I18160: signal is true;
	signal I18163: std_logic; attribute dont_touch of I18163: signal is true;
	signal I18166: std_logic; attribute dont_touch of I18166: signal is true;
	signal I18169: std_logic; attribute dont_touch of I18169: signal is true;
	signal I18172: std_logic; attribute dont_touch of I18172: signal is true;
	signal I18175: std_logic; attribute dont_touch of I18175: signal is true;
	signal I18178: std_logic; attribute dont_touch of I18178: signal is true;
	signal I18181: std_logic; attribute dont_touch of I18181: signal is true;
	signal I18184: std_logic; attribute dont_touch of I18184: signal is true;
	signal I18187: std_logic; attribute dont_touch of I18187: signal is true;
	signal I18190: std_logic; attribute dont_touch of I18190: signal is true;
	signal I18191: std_logic; attribute dont_touch of I18191: signal is true;
	signal I18192: std_logic; attribute dont_touch of I18192: signal is true;
	signal I18197: std_logic; attribute dont_touch of I18197: signal is true;
	signal I18198: std_logic; attribute dont_touch of I18198: signal is true;
	signal I18199: std_logic; attribute dont_touch of I18199: signal is true;
	signal I18204: std_logic; attribute dont_touch of I18204: signal is true;
	signal I18205: std_logic; attribute dont_touch of I18205: signal is true;
	signal I18206: std_logic; attribute dont_touch of I18206: signal is true;
	signal I18211: std_logic; attribute dont_touch of I18211: signal is true;
	signal I18214: std_logic; attribute dont_touch of I18214: signal is true;
	signal I18217: std_logic; attribute dont_touch of I18217: signal is true;
	signal I18220: std_logic; attribute dont_touch of I18220: signal is true;
	signal I18223: std_logic; attribute dont_touch of I18223: signal is true;
	signal I18226: std_logic; attribute dont_touch of I18226: signal is true;
	signal I18229: std_logic; attribute dont_touch of I18229: signal is true;
	signal I18232: std_logic; attribute dont_touch of I18232: signal is true;
	signal I18235: std_logic; attribute dont_touch of I18235: signal is true;
	signal I18238: std_logic; attribute dont_touch of I18238: signal is true;
	signal I18241: std_logic; attribute dont_touch of I18241: signal is true;
	signal I18244: std_logic; attribute dont_touch of I18244: signal is true;
	signal I18247: std_logic; attribute dont_touch of I18247: signal is true;
	signal I18250: std_logic; attribute dont_touch of I18250: signal is true;
	signal I18253: std_logic; attribute dont_touch of I18253: signal is true;
	signal I18256: std_logic; attribute dont_touch of I18256: signal is true;
	signal I18259: std_logic; attribute dont_touch of I18259: signal is true;
	signal I18262: std_logic; attribute dont_touch of I18262: signal is true;
	signal I18265: std_logic; attribute dont_touch of I18265: signal is true;
	signal I18268: std_logic; attribute dont_touch of I18268: signal is true;
	signal I18271: std_logic; attribute dont_touch of I18271: signal is true;
	signal I18274: std_logic; attribute dont_touch of I18274: signal is true;
	signal I18277: std_logic; attribute dont_touch of I18277: signal is true;
	signal I18280: std_logic; attribute dont_touch of I18280: signal is true;
	signal I18281: std_logic; attribute dont_touch of I18281: signal is true;
	signal I18282: std_logic; attribute dont_touch of I18282: signal is true;
	signal I18287: std_logic; attribute dont_touch of I18287: signal is true;
	signal I18288: std_logic; attribute dont_touch of I18288: signal is true;
	signal I18289: std_logic; attribute dont_touch of I18289: signal is true;
	signal I18295: std_logic; attribute dont_touch of I18295: signal is true;
	signal I18298: std_logic; attribute dont_touch of I18298: signal is true;
	signal I18302: std_logic; attribute dont_touch of I18302: signal is true;
	signal I18305: std_logic; attribute dont_touch of I18305: signal is true;
	signal I18308: std_logic; attribute dont_touch of I18308: signal is true;
	signal I18311: std_logic; attribute dont_touch of I18311: signal is true;
	signal I18314: std_logic; attribute dont_touch of I18314: signal is true;
	signal I18317: std_logic; attribute dont_touch of I18317: signal is true;
	signal I18320: std_logic; attribute dont_touch of I18320: signal is true;
	signal I18323: std_logic; attribute dont_touch of I18323: signal is true;
	signal I18326: std_logic; attribute dont_touch of I18326: signal is true;
	signal I18329: std_logic; attribute dont_touch of I18329: signal is true;
	signal I18332: std_logic; attribute dont_touch of I18332: signal is true;
	signal I18335: std_logic; attribute dont_touch of I18335: signal is true;
	signal I18338: std_logic; attribute dont_touch of I18338: signal is true;
	signal I18341: std_logic; attribute dont_touch of I18341: signal is true;
	signal I18344: std_logic; attribute dont_touch of I18344: signal is true;
	signal I18347: std_logic; attribute dont_touch of I18347: signal is true;
	signal I18350: std_logic; attribute dont_touch of I18350: signal is true;
	signal I18353: std_logic; attribute dont_touch of I18353: signal is true;
	signal I18356: std_logic; attribute dont_touch of I18356: signal is true;
	signal I18359: std_logic; attribute dont_touch of I18359: signal is true;
	signal I18362: std_logic; attribute dont_touch of I18362: signal is true;
	signal I18365: std_logic; attribute dont_touch of I18365: signal is true;
	signal I18368: std_logic; attribute dont_touch of I18368: signal is true;
	signal I18369: std_logic; attribute dont_touch of I18369: signal is true;
	signal I18370: std_logic; attribute dont_touch of I18370: signal is true;
	signal I18375: std_logic; attribute dont_touch of I18375: signal is true;
	signal I18378: std_logic; attribute dont_touch of I18378: signal is true;
	signal I18381: std_logic; attribute dont_touch of I18381: signal is true;
	signal I18386: std_logic; attribute dont_touch of I18386: signal is true;
	signal I18389: std_logic; attribute dont_touch of I18389: signal is true;
	signal I18392: std_logic; attribute dont_touch of I18392: signal is true;
	signal I18396: std_logic; attribute dont_touch of I18396: signal is true;
	signal I18399: std_logic; attribute dont_touch of I18399: signal is true;
	signal I18402: std_logic; attribute dont_touch of I18402: signal is true;
	signal I18405: std_logic; attribute dont_touch of I18405: signal is true;
	signal I18408: std_logic; attribute dont_touch of I18408: signal is true;
	signal I18411: std_logic; attribute dont_touch of I18411: signal is true;
	signal I18414: std_logic; attribute dont_touch of I18414: signal is true;
	signal I18417: std_logic; attribute dont_touch of I18417: signal is true;
	signal I18420: std_logic; attribute dont_touch of I18420: signal is true;
	signal I18423: std_logic; attribute dont_touch of I18423: signal is true;
	signal I18426: std_logic; attribute dont_touch of I18426: signal is true;
	signal I18429: std_logic; attribute dont_touch of I18429: signal is true;
	signal I18432: std_logic; attribute dont_touch of I18432: signal is true;
	signal I18435: std_logic; attribute dont_touch of I18435: signal is true;
	signal I18438: std_logic; attribute dont_touch of I18438: signal is true;
	signal I18441: std_logic; attribute dont_touch of I18441: signal is true;
	signal I18444: std_logic; attribute dont_touch of I18444: signal is true;
	signal I18449: std_logic; attribute dont_touch of I18449: signal is true;
	signal I18452: std_logic; attribute dont_touch of I18452: signal is true;
	signal I18455: std_logic; attribute dont_touch of I18455: signal is true;
	signal I18458: std_logic; attribute dont_touch of I18458: signal is true;
	signal I18461: std_logic; attribute dont_touch of I18461: signal is true;
	signal I18464: std_logic; attribute dont_touch of I18464: signal is true;
	signal I18467: std_logic; attribute dont_touch of I18467: signal is true;
	signal I18470: std_logic; attribute dont_touch of I18470: signal is true;
	signal I18473: std_logic; attribute dont_touch of I18473: signal is true;
	signal I18476: std_logic; attribute dont_touch of I18476: signal is true;
	signal I18479: std_logic; attribute dont_touch of I18479: signal is true;
	signal I18482: std_logic; attribute dont_touch of I18482: signal is true;
	signal I18485: std_logic; attribute dont_touch of I18485: signal is true;
	signal I18488: std_logic; attribute dont_touch of I18488: signal is true;
	signal I18491: std_logic; attribute dont_touch of I18491: signal is true;
	signal I18494: std_logic; attribute dont_touch of I18494: signal is true;
	signal I18497: std_logic; attribute dont_touch of I18497: signal is true;
	signal I18500: std_logic; attribute dont_touch of I18500: signal is true;
	signal I18503: std_logic; attribute dont_touch of I18503: signal is true;
	signal I18506: std_logic; attribute dont_touch of I18506: signal is true;
	signal I18509: std_logic; attribute dont_touch of I18509: signal is true;
	signal I18512: std_logic; attribute dont_touch of I18512: signal is true;
	signal I18515: std_logic; attribute dont_touch of I18515: signal is true;
	signal I18518: std_logic; attribute dont_touch of I18518: signal is true;
	signal I18521: std_logic; attribute dont_touch of I18521: signal is true;
	signal I18524: std_logic; attribute dont_touch of I18524: signal is true;
	signal I18527: std_logic; attribute dont_touch of I18527: signal is true;
	signal I18530: std_logic; attribute dont_touch of I18530: signal is true;
	signal I18533: std_logic; attribute dont_touch of I18533: signal is true;
	signal I18536: std_logic; attribute dont_touch of I18536: signal is true;
	signal I18539: std_logic; attribute dont_touch of I18539: signal is true;
	signal I18542: std_logic; attribute dont_touch of I18542: signal is true;
	signal I18545: std_logic; attribute dont_touch of I18545: signal is true;
	signal I18548: std_logic; attribute dont_touch of I18548: signal is true;
	signal I18551: std_logic; attribute dont_touch of I18551: signal is true;
	signal I18554: std_logic; attribute dont_touch of I18554: signal is true;
	signal I18557: std_logic; attribute dont_touch of I18557: signal is true;
	signal I18560: std_logic; attribute dont_touch of I18560: signal is true;
	signal I18563: std_logic; attribute dont_touch of I18563: signal is true;
	signal I18566: std_logic; attribute dont_touch of I18566: signal is true;
	signal I18569: std_logic; attribute dont_touch of I18569: signal is true;
	signal I18572: std_logic; attribute dont_touch of I18572: signal is true;
	signal I18575: std_logic; attribute dont_touch of I18575: signal is true;
	signal I18578: std_logic; attribute dont_touch of I18578: signal is true;
	signal I18581: std_logic; attribute dont_touch of I18581: signal is true;
	signal I18584: std_logic; attribute dont_touch of I18584: signal is true;
	signal I18587: std_logic; attribute dont_touch of I18587: signal is true;
	signal I18590: std_logic; attribute dont_touch of I18590: signal is true;
	signal I18593: std_logic; attribute dont_touch of I18593: signal is true;
	signal I18596: std_logic; attribute dont_touch of I18596: signal is true;
	signal I18599: std_logic; attribute dont_touch of I18599: signal is true;
	signal I18602: std_logic; attribute dont_touch of I18602: signal is true;
	signal I18605: std_logic; attribute dont_touch of I18605: signal is true;
	signal I18608: std_logic; attribute dont_touch of I18608: signal is true;
	signal I18611: std_logic; attribute dont_touch of I18611: signal is true;
	signal I18614: std_logic; attribute dont_touch of I18614: signal is true;
	signal I18617: std_logic; attribute dont_touch of I18617: signal is true;
	signal I18620: std_logic; attribute dont_touch of I18620: signal is true;
	signal I18623: std_logic; attribute dont_touch of I18623: signal is true;
	signal I18626: std_logic; attribute dont_touch of I18626: signal is true;
	signal I18629: std_logic; attribute dont_touch of I18629: signal is true;
	signal I18632: std_logic; attribute dont_touch of I18632: signal is true;
	signal I18635: std_logic; attribute dont_touch of I18635: signal is true;
	signal I18638: std_logic; attribute dont_touch of I18638: signal is true;
	signal I18641: std_logic; attribute dont_touch of I18641: signal is true;
	signal I18644: std_logic; attribute dont_touch of I18644: signal is true;
	signal I18647: std_logic; attribute dont_touch of I18647: signal is true;
	signal I18650: std_logic; attribute dont_touch of I18650: signal is true;
	signal I18653: std_logic; attribute dont_touch of I18653: signal is true;
	signal I18656: std_logic; attribute dont_touch of I18656: signal is true;
	signal I18659: std_logic; attribute dont_touch of I18659: signal is true;
	signal I18662: std_logic; attribute dont_touch of I18662: signal is true;
	signal I18665: std_logic; attribute dont_touch of I18665: signal is true;
	signal I18668: std_logic; attribute dont_touch of I18668: signal is true;
	signal I18671: std_logic; attribute dont_touch of I18671: signal is true;
	signal I18674: std_logic; attribute dont_touch of I18674: signal is true;
	signal I18677: std_logic; attribute dont_touch of I18677: signal is true;
	signal I18680: std_logic; attribute dont_touch of I18680: signal is true;
	signal I18683: std_logic; attribute dont_touch of I18683: signal is true;
	signal I18686: std_logic; attribute dont_touch of I18686: signal is true;
	signal I18689: std_logic; attribute dont_touch of I18689: signal is true;
	signal I18692: std_logic; attribute dont_touch of I18692: signal is true;
	signal I18695: std_logic; attribute dont_touch of I18695: signal is true;
	signal I18698: std_logic; attribute dont_touch of I18698: signal is true;
	signal I18701: std_logic; attribute dont_touch of I18701: signal is true;
	signal I18704: std_logic; attribute dont_touch of I18704: signal is true;
	signal I18707: std_logic; attribute dont_touch of I18707: signal is true;
	signal I18710: std_logic; attribute dont_touch of I18710: signal is true;
	signal I18713: std_logic; attribute dont_touch of I18713: signal is true;
	signal I18716: std_logic; attribute dont_touch of I18716: signal is true;
	signal I18719: std_logic; attribute dont_touch of I18719: signal is true;
	signal I18722: std_logic; attribute dont_touch of I18722: signal is true;
	signal I18725: std_logic; attribute dont_touch of I18725: signal is true;
	signal I18728: std_logic; attribute dont_touch of I18728: signal is true;
	signal I18731: std_logic; attribute dont_touch of I18731: signal is true;
	signal I18734: std_logic; attribute dont_touch of I18734: signal is true;
	signal I18737: std_logic; attribute dont_touch of I18737: signal is true;
	signal I18740: std_logic; attribute dont_touch of I18740: signal is true;
	signal I18743: std_logic; attribute dont_touch of I18743: signal is true;
	signal I18746: std_logic; attribute dont_touch of I18746: signal is true;
	signal I18749: std_logic; attribute dont_touch of I18749: signal is true;
	signal I18752: std_logic; attribute dont_touch of I18752: signal is true;
	signal I18755: std_logic; attribute dont_touch of I18755: signal is true;
	signal I18758: std_logic; attribute dont_touch of I18758: signal is true;
	signal I18761: std_logic; attribute dont_touch of I18761: signal is true;
	signal I18764: std_logic; attribute dont_touch of I18764: signal is true;
	signal I18767: std_logic; attribute dont_touch of I18767: signal is true;
	signal I18770: std_logic; attribute dont_touch of I18770: signal is true;
	signal I18773: std_logic; attribute dont_touch of I18773: signal is true;
	signal I18777: std_logic; attribute dont_touch of I18777: signal is true;
	signal I18780: std_logic; attribute dont_touch of I18780: signal is true;
	signal I18784: std_logic; attribute dont_touch of I18784: signal is true;
	signal I18787: std_logic; attribute dont_touch of I18787: signal is true;
	signal I18791: std_logic; attribute dont_touch of I18791: signal is true;
	signal I18794: std_logic; attribute dont_touch of I18794: signal is true;
	signal I18799: std_logic; attribute dont_touch of I18799: signal is true;
	signal I18800: std_logic; attribute dont_touch of I18800: signal is true;
	signal I18801: std_logic; attribute dont_touch of I18801: signal is true;
	signal I18810: std_logic; attribute dont_touch of I18810: signal is true;
	signal I18813: std_logic; attribute dont_touch of I18813: signal is true;
	signal I18817: std_logic; attribute dont_touch of I18817: signal is true;
	signal I18820: std_logic; attribute dont_touch of I18820: signal is true;
	signal I18824: std_logic; attribute dont_touch of I18824: signal is true;
	signal I18827: std_logic; attribute dont_touch of I18827: signal is true;
	signal I18835: std_logic; attribute dont_touch of I18835: signal is true;
	signal I18838: std_logic; attribute dont_touch of I18838: signal is true;
	signal I18842: std_logic; attribute dont_touch of I18842: signal is true;
	signal I18845: std_logic; attribute dont_touch of I18845: signal is true;
	signal I18854: std_logic; attribute dont_touch of I18854: signal is true;
	signal I18857: std_logic; attribute dont_touch of I18857: signal is true;
	signal I18866: std_logic; attribute dont_touch of I18866: signal is true;
	signal I18929: std_logic; attribute dont_touch of I18929: signal is true;
	signal I18943: std_logic; attribute dont_touch of I18943: signal is true;
	signal I18962: std_logic; attribute dont_touch of I18962: signal is true;
	signal I18969: std_logic; attribute dont_touch of I18969: signal is true;
	signal I18990: std_logic; attribute dont_touch of I18990: signal is true;
	signal I19025: std_logic; attribute dont_touch of I19025: signal is true;
	signal I19030: std_logic; attribute dont_touch of I19030: signal is true;
	signal I19105: std_logic; attribute dont_touch of I19105: signal is true;
	signal I19119: std_logic; attribute dont_touch of I19119: signal is true;
	signal I19160: std_logic; attribute dont_touch of I19160: signal is true;
	signal I19174: std_logic; attribute dont_touch of I19174: signal is true;
	signal I19195: std_logic; attribute dont_touch of I19195: signal is true;
	signal I19208: std_logic; attribute dont_touch of I19208: signal is true;
	signal I19211: std_logic; attribute dont_touch of I19211: signal is true;
	signal I19226: std_logic; attribute dont_touch of I19226: signal is true;
	signal I19240: std_logic; attribute dont_touch of I19240: signal is true;
	signal I19271: std_logic; attribute dont_touch of I19271: signal is true;
	signal I19274: std_logic; attribute dont_touch of I19274: signal is true;
	signal I19289: std_logic; attribute dont_touch of I19289: signal is true;
	signal I19303: std_logic; attribute dont_touch of I19303: signal is true;
	signal I19307: std_logic; attribute dont_touch of I19307: signal is true;
	signal I19315: std_logic; attribute dont_touch of I19315: signal is true;
	signal I19318: std_logic; attribute dont_touch of I19318: signal is true;
	signal I19321: std_logic; attribute dont_touch of I19321: signal is true;
	signal I19342: std_logic; attribute dont_touch of I19342: signal is true;
	signal I19345: std_logic; attribute dont_touch of I19345: signal is true;
	signal I19360: std_logic; attribute dont_touch of I19360: signal is true;
	signal I19374: std_logic; attribute dont_touch of I19374: signal is true;
	signal I19377: std_logic; attribute dont_touch of I19377: signal is true;
	signal I19380: std_logic; attribute dont_touch of I19380: signal is true;
	signal I19401: std_logic; attribute dont_touch of I19401: signal is true;
	signal I19404: std_logic; attribute dont_touch of I19404: signal is true;
	signal I19412: std_logic; attribute dont_touch of I19412: signal is true;
	signal I19415: std_logic; attribute dont_touch of I19415: signal is true;
	signal I19426: std_logic; attribute dont_touch of I19426: signal is true;
	signal I19429: std_logic; attribute dont_touch of I19429: signal is true;
	signal I19432: std_logic; attribute dont_touch of I19432: signal is true;
	signal I19449: std_logic; attribute dont_touch of I19449: signal is true;
	signal I19452: std_logic; attribute dont_touch of I19452: signal is true;
	signal I19455: std_logic; attribute dont_touch of I19455: signal is true;
	signal I19466: std_logic; attribute dont_touch of I19466: signal is true;
	signal I19469: std_logic; attribute dont_touch of I19469: signal is true;
	signal I19472: std_logic; attribute dont_touch of I19472: signal is true;
	signal I19479: std_logic; attribute dont_touch of I19479: signal is true;
	signal I19482: std_logic; attribute dont_touch of I19482: signal is true;
	signal I19485: std_logic; attribute dont_touch of I19485: signal is true;
	signal I19488: std_logic; attribute dont_touch of I19488: signal is true;
	signal I19500: std_logic; attribute dont_touch of I19500: signal is true;
	signal I19503: std_logic; attribute dont_touch of I19503: signal is true;
	signal I19507: std_logic; attribute dont_touch of I19507: signal is true;
	signal I19510: std_logic; attribute dont_touch of I19510: signal is true;
	signal I19513: std_logic; attribute dont_touch of I19513: signal is true;
	signal I19516: std_logic; attribute dont_touch of I19516: signal is true;
	signal I19523: std_logic; attribute dont_touch of I19523: signal is true;
	signal I19526: std_logic; attribute dont_touch of I19526: signal is true;
	signal I19530: std_logic; attribute dont_touch of I19530: signal is true;
	signal I19533: std_logic; attribute dont_touch of I19533: signal is true;
	signal I19539: std_logic; attribute dont_touch of I19539: signal is true;
	signal I19542: std_logic; attribute dont_touch of I19542: signal is true;
	signal I19545: std_logic; attribute dont_touch of I19545: signal is true;
	signal I19549: std_logic; attribute dont_touch of I19549: signal is true;
	signal I19552: std_logic; attribute dont_touch of I19552: signal is true;
	signal I19557: std_logic; attribute dont_touch of I19557: signal is true;
	signal I19560: std_logic; attribute dont_touch of I19560: signal is true;
	signal I19563: std_logic; attribute dont_touch of I19563: signal is true;
	signal I19569: std_logic; attribute dont_touch of I19569: signal is true;
	signal I19573: std_logic; attribute dont_touch of I19573: signal is true;
	signal I19576: std_logic; attribute dont_touch of I19576: signal is true;
	signal I19582: std_logic; attribute dont_touch of I19582: signal is true;
	signal I19587: std_logic; attribute dont_touch of I19587: signal is true;
	signal I19591: std_logic; attribute dont_touch of I19591: signal is true;
	signal I19595: std_logic; attribute dont_touch of I19595: signal is true;
	signal I19598: std_logic; attribute dont_touch of I19598: signal is true;
	signal I19602: std_logic; attribute dont_touch of I19602: signal is true;
	signal I19605: std_logic; attribute dont_touch of I19605: signal is true;
	signal I19608: std_logic; attribute dont_touch of I19608: signal is true;
	signal I19611: std_logic; attribute dont_touch of I19611: signal is true;
	signal I19615: std_logic; attribute dont_touch of I19615: signal is true;
	signal I19618: std_logic; attribute dont_touch of I19618: signal is true;
	signal I19621: std_logic; attribute dont_touch of I19621: signal is true;
	signal I19624: std_logic; attribute dont_touch of I19624: signal is true;
	signal I19628: std_logic; attribute dont_touch of I19628: signal is true;
	signal I19631: std_logic; attribute dont_touch of I19631: signal is true;
	signal I19634: std_logic; attribute dont_touch of I19634: signal is true;
	signal I19637: std_logic; attribute dont_touch of I19637: signal is true;
	signal I19642: std_logic; attribute dont_touch of I19642: signal is true;
	signal I19645: std_logic; attribute dont_touch of I19645: signal is true;
	signal I19648: std_logic; attribute dont_touch of I19648: signal is true;
	signal I19654: std_logic; attribute dont_touch of I19654: signal is true;
	signal I19657: std_logic; attribute dont_touch of I19657: signal is true;
	signal I19667: std_logic; attribute dont_touch of I19667: signal is true;
	signal I19689: std_logic; attribute dont_touch of I19689: signal is true;
	signal I19702: std_logic; attribute dont_touch of I19702: signal is true;
	signal I19711: std_logic; attribute dont_touch of I19711: signal is true;
	signal I19718: std_logic; attribute dont_touch of I19718: signal is true;
	signal I19722: std_logic; attribute dont_touch of I19722: signal is true;
	signal I19727: std_logic; attribute dont_touch of I19727: signal is true;
	signal I19733: std_logic; attribute dont_touch of I19733: signal is true;
	signal I19736: std_logic; attribute dont_touch of I19736: signal is true;
	signal I19739: std_logic; attribute dont_touch of I19739: signal is true;
	signal I19747: std_logic; attribute dont_touch of I19747: signal is true;
	signal I19750: std_logic; attribute dont_touch of I19750: signal is true;
	signal I19753: std_logic; attribute dont_touch of I19753: signal is true;
	signal I19756: std_logic; attribute dont_touch of I19756: signal is true;
	signal I19759: std_logic; attribute dont_touch of I19759: signal is true;
	signal I19767: std_logic; attribute dont_touch of I19767: signal is true;
	signal I19771: std_logic; attribute dont_touch of I19771: signal is true;
	signal I19774: std_logic; attribute dont_touch of I19774: signal is true;
	signal I19777: std_logic; attribute dont_touch of I19777: signal is true;
	signal I19784: std_logic; attribute dont_touch of I19784: signal is true;
	signal I19787: std_logic; attribute dont_touch of I19787: signal is true;
	signal I19791: std_logic; attribute dont_touch of I19791: signal is true;
	signal I19794: std_logic; attribute dont_touch of I19794: signal is true;
	signal I19797: std_logic; attribute dont_touch of I19797: signal is true;
	signal I19800: std_logic; attribute dont_touch of I19800: signal is true;
	signal I19803: std_logic; attribute dont_touch of I19803: signal is true;
	signal I19808: std_logic; attribute dont_touch of I19808: signal is true;
	signal I19813: std_logic; attribute dont_touch of I19813: signal is true;
	signal I19816: std_logic; attribute dont_touch of I19816: signal is true;
	signal I19820: std_logic; attribute dont_touch of I19820: signal is true;
	signal I19823: std_logic; attribute dont_touch of I19823: signal is true;
	signal I19826: std_logic; attribute dont_touch of I19826: signal is true;
	signal I19829: std_logic; attribute dont_touch of I19829: signal is true;
	signal I19833: std_logic; attribute dont_touch of I19833: signal is true;
	signal I19836: std_logic; attribute dont_touch of I19836: signal is true;
	signal I19844: std_logic; attribute dont_touch of I19844: signal is true;
	signal I19847: std_logic; attribute dont_touch of I19847: signal is true;
	signal I19852: std_logic; attribute dont_touch of I19852: signal is true;
	signal I19855: std_logic; attribute dont_touch of I19855: signal is true;
	signal I19859: std_logic; attribute dont_touch of I19859: signal is true;
	signal I19862: std_logic; attribute dont_touch of I19862: signal is true;
	signal I19865: std_logic; attribute dont_touch of I19865: signal is true;
	signal I19869: std_logic; attribute dont_touch of I19869: signal is true;
	signal I19872: std_logic; attribute dont_touch of I19872: signal is true;
	signal I19877: std_logic; attribute dont_touch of I19877: signal is true;
	signal I19883: std_logic; attribute dont_touch of I19883: signal is true;
	signal I19886: std_logic; attribute dont_touch of I19886: signal is true;
	signal I19891: std_logic; attribute dont_touch of I19891: signal is true;
	signal I19894: std_logic; attribute dont_touch of I19894: signal is true;
	signal I19898: std_logic; attribute dont_touch of I19898: signal is true;
	signal I19901: std_logic; attribute dont_touch of I19901: signal is true;
	signal I19905: std_logic; attribute dont_touch of I19905: signal is true;
	signal I19915: std_logic; attribute dont_touch of I19915: signal is true;
	signal I19921: std_logic; attribute dont_touch of I19921: signal is true;
	signal I19924: std_logic; attribute dont_touch of I19924: signal is true;
	signal I19929: std_logic; attribute dont_touch of I19929: signal is true;
	signal I19932: std_logic; attribute dont_touch of I19932: signal is true;
	signal I19937: std_logic; attribute dont_touch of I19937: signal is true;
	signal I19938: std_logic; attribute dont_touch of I19938: signal is true;
	signal I19952: std_logic; attribute dont_touch of I19952: signal is true;
	signal I19958: std_logic; attribute dont_touch of I19958: signal is true;
	signal I19961: std_logic; attribute dont_touch of I19961: signal is true;
	signal I19971: std_logic; attribute dont_touch of I19971: signal is true;
	signal I19972: std_logic; attribute dont_touch of I19972: signal is true;
	signal I19986: std_logic; attribute dont_touch of I19986: signal is true;
	signal I19996: std_logic; attribute dont_touch of I19996: signal is true;
	signal I19997: std_logic; attribute dont_touch of I19997: signal is true;
	signal I20009: std_logic; attribute dont_touch of I20009: signal is true;
	signal I20021: std_logic; attribute dont_touch of I20021: signal is true;
	signal I20022: std_logic; attribute dont_touch of I20022: signal is true;
	signal I20031: std_logic; attribute dont_touch of I20031: signal is true;
	signal I20032: std_logic; attribute dont_touch of I20032: signal is true;
	signal I20033: std_logic; attribute dont_touch of I20033: signal is true;
	signal I20048: std_logic; attribute dont_touch of I20048: signal is true;
	signal I20049: std_logic; attribute dont_touch of I20049: signal is true;
	signal I20050: std_logic; attribute dont_touch of I20050: signal is true;
	signal I20062: std_logic; attribute dont_touch of I20062: signal is true;
	signal I20100: std_logic; attribute dont_touch of I20100: signal is true;
	signal I20117: std_logic; attribute dont_touch of I20117: signal is true;
	signal I20131: std_logic; attribute dont_touch of I20131: signal is true;
	signal I20132: std_logic; attribute dont_touch of I20132: signal is true;
	signal I20264: std_logic; attribute dont_touch of I20264: signal is true;
	signal I20278: std_logic; attribute dont_touch of I20278: signal is true;
	signal I20283: std_logic; attribute dont_touch of I20283: signal is true;
	signal I20295: std_logic; attribute dont_touch of I20295: signal is true;
	signal I20299: std_logic; attribute dont_touch of I20299: signal is true;
	signal I20305: std_logic; attribute dont_touch of I20305: signal is true;
	signal I20310: std_logic; attribute dont_touch of I20310: signal is true;
	signal I20320: std_logic; attribute dont_touch of I20320: signal is true;
	signal I20324: std_logic; attribute dont_touch of I20324: signal is true;
	signal I20328: std_logic; attribute dont_touch of I20328: signal is true;
	signal I20334: std_logic; attribute dont_touch of I20334: signal is true;
	signal I20339: std_logic; attribute dont_touch of I20339: signal is true;
	signal I20347: std_logic; attribute dont_touch of I20347: signal is true;
	signal I20351: std_logic; attribute dont_touch of I20351: signal is true;
	signal I20355: std_logic; attribute dont_touch of I20355: signal is true;
	signal I20359: std_logic; attribute dont_touch of I20359: signal is true;
	signal I20365: std_logic; attribute dont_touch of I20365: signal is true;
	signal I20376: std_logic; attribute dont_touch of I20376: signal is true;
	signal I20379: std_logic; attribute dont_touch of I20379: signal is true;
	signal I20382: std_logic; attribute dont_touch of I20382: signal is true;
	signal I20386: std_logic; attribute dont_touch of I20386: signal is true;
	signal I20390: std_logic; attribute dont_touch of I20390: signal is true;
	signal I20394: std_logic; attribute dont_touch of I20394: signal is true;
	signal I20398: std_logic; attribute dont_touch of I20398: signal is true;
	signal I20407: std_logic; attribute dont_touch of I20407: signal is true;
	signal I20410: std_logic; attribute dont_touch of I20410: signal is true;
	signal I20414: std_logic; attribute dont_touch of I20414: signal is true;
	signal I20417: std_logic; attribute dont_touch of I20417: signal is true;
	signal I20421: std_logic; attribute dont_touch of I20421: signal is true;
	signal I20425: std_logic; attribute dont_touch of I20425: signal is true;
	signal I20429: std_logic; attribute dont_touch of I20429: signal is true;
	signal I20430: std_logic; attribute dont_touch of I20430: signal is true;
	signal I20431: std_logic; attribute dont_touch of I20431: signal is true;
	signal I20441: std_logic; attribute dont_touch of I20441: signal is true;
	signal I20444: std_logic; attribute dont_touch of I20444: signal is true;
	signal I20448: std_logic; attribute dont_touch of I20448: signal is true;
	signal I20451: std_logic; attribute dont_touch of I20451: signal is true;
	signal I20455: std_logic; attribute dont_touch of I20455: signal is true;
	signal I20458: std_logic; attribute dont_touch of I20458: signal is true;
	signal I20462: std_logic; attribute dont_touch of I20462: signal is true;
	signal I20465: std_logic; attribute dont_touch of I20465: signal is true;
	signal I20466: std_logic; attribute dont_touch of I20466: signal is true;
	signal I20467: std_logic; attribute dont_touch of I20467: signal is true;
	signal I20476: std_logic; attribute dont_touch of I20476: signal is true;
	signal I20479: std_logic; attribute dont_touch of I20479: signal is true;
	signal I20483: std_logic; attribute dont_touch of I20483: signal is true;
	signal I20486: std_logic; attribute dont_touch of I20486: signal is true;
	signal I20490: std_logic; attribute dont_touch of I20490: signal is true;
	signal I20493: std_logic; attribute dont_touch of I20493: signal is true;
	signal I20497: std_logic; attribute dont_touch of I20497: signal is true;
	signal I20500: std_logic; attribute dont_touch of I20500: signal is true;
	signal I20504: std_logic; attribute dont_touch of I20504: signal is true;
	signal I20505: std_logic; attribute dont_touch of I20505: signal is true;
	signal I20506: std_logic; attribute dont_touch of I20506: signal is true;
	signal I20514: std_logic; attribute dont_touch of I20514: signal is true;
	signal I20517: std_logic; attribute dont_touch of I20517: signal is true;
	signal I20520: std_logic; attribute dont_touch of I20520: signal is true;
	signal I20523: std_logic; attribute dont_touch of I20523: signal is true;
	signal I20526: std_logic; attribute dont_touch of I20526: signal is true;
	signal I20529: std_logic; attribute dont_touch of I20529: signal is true;
	signal I20532: std_logic; attribute dont_touch of I20532: signal is true;
	signal I20535: std_logic; attribute dont_touch of I20535: signal is true;
	signal I20538: std_logic; attribute dont_touch of I20538: signal is true;
	signal I20541: std_logic; attribute dont_touch of I20541: signal is true;
	signal I20544: std_logic; attribute dont_touch of I20544: signal is true;
	signal I20547: std_logic; attribute dont_touch of I20547: signal is true;
	signal I20550: std_logic; attribute dont_touch of I20550: signal is true;
	signal I20553: std_logic; attribute dont_touch of I20553: signal is true;
	signal I20556: std_logic; attribute dont_touch of I20556: signal is true;
	signal I20559: std_logic; attribute dont_touch of I20559: signal is true;
	signal I20562: std_logic; attribute dont_touch of I20562: signal is true;
	signal I20565: std_logic; attribute dont_touch of I20565: signal is true;
	signal I20568: std_logic; attribute dont_touch of I20568: signal is true;
	signal I20571: std_logic; attribute dont_touch of I20571: signal is true;
	signal I20574: std_logic; attribute dont_touch of I20574: signal is true;
	signal I20577: std_logic; attribute dont_touch of I20577: signal is true;
	signal I20580: std_logic; attribute dont_touch of I20580: signal is true;
	signal I20583: std_logic; attribute dont_touch of I20583: signal is true;
	signal I20586: std_logic; attribute dont_touch of I20586: signal is true;
	signal I20589: std_logic; attribute dont_touch of I20589: signal is true;
	signal I20592: std_logic; attribute dont_touch of I20592: signal is true;
	signal I20595: std_logic; attribute dont_touch of I20595: signal is true;
	signal I20598: std_logic; attribute dont_touch of I20598: signal is true;
	signal I20601: std_logic; attribute dont_touch of I20601: signal is true;
	signal I20604: std_logic; attribute dont_touch of I20604: signal is true;
	signal I20607: std_logic; attribute dont_touch of I20607: signal is true;
	signal I20610: std_logic; attribute dont_touch of I20610: signal is true;
	signal I20613: std_logic; attribute dont_touch of I20613: signal is true;
	signal I20616: std_logic; attribute dont_touch of I20616: signal is true;
	signal I20619: std_logic; attribute dont_touch of I20619: signal is true;
	signal I20622: std_logic; attribute dont_touch of I20622: signal is true;
	signal I20625: std_logic; attribute dont_touch of I20625: signal is true;
	signal I20628: std_logic; attribute dont_touch of I20628: signal is true;
	signal I20631: std_logic; attribute dont_touch of I20631: signal is true;
	signal I20634: std_logic; attribute dont_touch of I20634: signal is true;
	signal I20637: std_logic; attribute dont_touch of I20637: signal is true;
	signal I20640: std_logic; attribute dont_touch of I20640: signal is true;
	signal I20643: std_logic; attribute dont_touch of I20643: signal is true;
	signal I20646: std_logic; attribute dont_touch of I20646: signal is true;
	signal I20649: std_logic; attribute dont_touch of I20649: signal is true;
	signal I20652: std_logic; attribute dont_touch of I20652: signal is true;
	signal I20655: std_logic; attribute dont_touch of I20655: signal is true;
	signal I20658: std_logic; attribute dont_touch of I20658: signal is true;
	signal I20661: std_logic; attribute dont_touch of I20661: signal is true;
	signal I20664: std_logic; attribute dont_touch of I20664: signal is true;
	signal I20667: std_logic; attribute dont_touch of I20667: signal is true;
	signal I20670: std_logic; attribute dont_touch of I20670: signal is true;
	signal I20673: std_logic; attribute dont_touch of I20673: signal is true;
	signal I20676: std_logic; attribute dont_touch of I20676: signal is true;
	signal I20679: std_logic; attribute dont_touch of I20679: signal is true;
	signal I20682: std_logic; attribute dont_touch of I20682: signal is true;
	signal I20685: std_logic; attribute dont_touch of I20685: signal is true;
	signal I20688: std_logic; attribute dont_touch of I20688: signal is true;
	signal I20691: std_logic; attribute dont_touch of I20691: signal is true;
	signal I20694: std_logic; attribute dont_touch of I20694: signal is true;
	signal I20697: std_logic; attribute dont_touch of I20697: signal is true;
	signal I20700: std_logic; attribute dont_touch of I20700: signal is true;
	signal I20703: std_logic; attribute dont_touch of I20703: signal is true;
	signal I20706: std_logic; attribute dont_touch of I20706: signal is true;
	signal I20709: std_logic; attribute dont_touch of I20709: signal is true;
	signal I20743: std_logic; attribute dont_touch of I20743: signal is true;
	signal I20744: std_logic; attribute dont_touch of I20744: signal is true;
	signal I20745: std_logic; attribute dont_touch of I20745: signal is true;
	signal I20791: std_logic; attribute dont_touch of I20791: signal is true;
	signal I20794: std_logic; attribute dont_touch of I20794: signal is true;
	signal I20799: std_logic; attribute dont_touch of I20799: signal is true;
	signal I20802: std_logic; attribute dont_touch of I20802: signal is true;
	signal I20805: std_logic; attribute dont_touch of I20805: signal is true;
	signal I20810: std_logic; attribute dont_touch of I20810: signal is true;
	signal I20813: std_logic; attribute dont_touch of I20813: signal is true;
	signal I20816: std_logic; attribute dont_touch of I20816: signal is true;
	signal I20820: std_logic; attribute dont_touch of I20820: signal is true;
	signal I20823: std_logic; attribute dont_touch of I20823: signal is true;
	signal I20828: std_logic; attribute dont_touch of I20828: signal is true;
	signal I20832: std_logic; attribute dont_touch of I20832: signal is true;
	signal I20836: std_logic; attribute dont_touch of I20836: signal is true;
	signal I20839: std_logic; attribute dont_touch of I20839: signal is true;
	signal I20844: std_logic; attribute dont_touch of I20844: signal is true;
	signal I20848: std_logic; attribute dont_touch of I20848: signal is true;
	signal I20852: std_logic; attribute dont_touch of I20852: signal is true;
	signal I20858: std_logic; attribute dont_touch of I20858: signal is true;
	signal I20863: std_logic; attribute dont_touch of I20863: signal is true;
	signal I20873: std_logic; attribute dont_touch of I20873: signal is true;
	signal I20886: std_logic; attribute dont_touch of I20886: signal is true;
	signal I20909: std_logic; attribute dont_touch of I20909: signal is true;
	signal I20959: std_logic; attribute dont_touch of I20959: signal is true;
	signal I21012: std_logic; attribute dont_touch of I21012: signal is true;
	signal I21037: std_logic; attribute dont_touch of I21037: signal is true;
	signal I21045: std_logic; attribute dont_touch of I21045: signal is true;
	signal I21064: std_logic; attribute dont_touch of I21064: signal is true;
	signal I21075: std_logic; attribute dont_touch of I21075: signal is true;
	signal I21083: std_logic; attribute dont_touch of I21083: signal is true;
	signal I21096: std_logic; attribute dont_touch of I21096: signal is true;
	signal I21108: std_logic; attribute dont_touch of I21108: signal is true;
	signal I21119: std_logic; attribute dont_touch of I21119: signal is true;
	signal I21127: std_logic; attribute dont_touch of I21127: signal is true;
	signal I21137: std_logic; attribute dont_touch of I21137: signal is true;
	signal I21149: std_logic; attribute dont_touch of I21149: signal is true;
	signal I21160: std_logic; attribute dont_touch of I21160: signal is true;
	signal I21165: std_logic; attribute dont_touch of I21165: signal is true;
	signal I21178: std_logic; attribute dont_touch of I21178: signal is true;
	signal I21190: std_logic; attribute dont_touch of I21190: signal is true;
	signal I21208: std_logic; attribute dont_touch of I21208: signal is true;
	signal I21241: std_logic; attribute dont_touch of I21241: signal is true;
	signal I21246: std_logic; attribute dont_touch of I21246: signal is true;
	signal I21249: std_logic; attribute dont_touch of I21249: signal is true;
	signal I21252: std_logic; attribute dont_touch of I21252: signal is true;
	signal I21256: std_logic; attribute dont_touch of I21256: signal is true;
	signal I21259: std_logic; attribute dont_touch of I21259: signal is true;
	signal I21262: std_logic; attribute dont_touch of I21262: signal is true;
	signal I21267: std_logic; attribute dont_touch of I21267: signal is true;
	signal I21271: std_logic; attribute dont_touch of I21271: signal is true;
	signal I21274: std_logic; attribute dont_touch of I21274: signal is true;
	signal I21277: std_logic; attribute dont_touch of I21277: signal is true;
	signal I21282: std_logic; attribute dont_touch of I21282: signal is true;
	signal I21286: std_logic; attribute dont_touch of I21286: signal is true;
	signal I21289: std_logic; attribute dont_touch of I21289: signal is true;
	signal I21292: std_logic; attribute dont_touch of I21292: signal is true;
	signal I21297: std_logic; attribute dont_touch of I21297: signal is true;
	signal I21301: std_logic; attribute dont_touch of I21301: signal is true;
	signal I21304: std_logic; attribute dont_touch of I21304: signal is true;
	signal I21310: std_logic; attribute dont_touch of I21310: signal is true;
	signal I21313: std_logic; attribute dont_touch of I21313: signal is true;
	signal I21318: std_logic; attribute dont_touch of I21318: signal is true;
	signal I21321: std_logic; attribute dont_touch of I21321: signal is true;
	signal I21326: std_logic; attribute dont_touch of I21326: signal is true;
	signal I21329: std_logic; attribute dont_touch of I21329: signal is true;
	signal I21337: std_logic; attribute dont_touch of I21337: signal is true;
	signal I21340: std_logic; attribute dont_touch of I21340: signal is true;
	signal I21351: std_logic; attribute dont_touch of I21351: signal is true;
	signal I21354: std_logic; attribute dont_touch of I21354: signal is true;
	signal I21361: std_logic; attribute dont_touch of I21361: signal is true;
	signal I21364: std_logic; attribute dont_touch of I21364: signal is true;
	signal I21374: std_logic; attribute dont_touch of I21374: signal is true;
	signal I21377: std_logic; attribute dont_touch of I21377: signal is true;
	signal I21381: std_logic; attribute dont_touch of I21381: signal is true;
	signal I21389: std_logic; attribute dont_touch of I21389: signal is true;
	signal I21392: std_logic; attribute dont_touch of I21392: signal is true;
	signal I21395: std_logic; attribute dont_touch of I21395: signal is true;
	signal I21398: std_logic; attribute dont_touch of I21398: signal is true;
	signal I21404: std_logic; attribute dont_touch of I21404: signal is true;
	signal I21407: std_logic; attribute dont_touch of I21407: signal is true;
	signal I21415: std_logic; attribute dont_touch of I21415: signal is true;
	signal I21420: std_logic; attribute dont_touch of I21420: signal is true;
	signal I21426: std_logic; attribute dont_touch of I21426: signal is true;
	signal I21429: std_logic; attribute dont_touch of I21429: signal is true;
	signal I21432: std_logic; attribute dont_touch of I21432: signal is true;
	signal I21435: std_logic; attribute dont_touch of I21435: signal is true;
	signal I21443: std_logic; attribute dont_touch of I21443: signal is true;
	signal I21446: std_logic; attribute dont_touch of I21446: signal is true;
	signal I21449: std_logic; attribute dont_touch of I21449: signal is true;
	signal I21452: std_logic; attribute dont_touch of I21452: signal is true;
	signal I21458: std_logic; attribute dont_touch of I21458: signal is true;
	signal I21461: std_logic; attribute dont_touch of I21461: signal is true;
	signal I21476: std_logic; attribute dont_touch of I21476: signal is true;
	signal I21479: std_logic; attribute dont_touch of I21479: signal is true;
	signal I21482: std_logic; attribute dont_touch of I21482: signal is true;
	signal I21488: std_logic; attribute dont_touch of I21488: signal is true;
	signal I21491: std_logic; attribute dont_touch of I21491: signal is true;
	signal I21494: std_logic; attribute dont_touch of I21494: signal is true;
	signal I21497: std_logic; attribute dont_touch of I21497: signal is true;
	signal I21505: std_logic; attribute dont_touch of I21505: signal is true;
	signal I21508: std_logic; attribute dont_touch of I21508: signal is true;
	signal I21511: std_logic; attribute dont_touch of I21511: signal is true;
	signal I21514: std_logic; attribute dont_touch of I21514: signal is true;
	signal I21520: std_logic; attribute dont_touch of I21520: signal is true;
	signal I21523: std_logic; attribute dont_touch of I21523: signal is true;
	signal I21531: std_logic; attribute dont_touch of I21531: signal is true;
	signal I21534: std_logic; attribute dont_touch of I21534: signal is true;
	signal I21537: std_logic; attribute dont_touch of I21537: signal is true;
	signal I21548: std_logic; attribute dont_touch of I21548: signal is true;
	signal I21551: std_logic; attribute dont_touch of I21551: signal is true;
	signal I21554: std_logic; attribute dont_touch of I21554: signal is true;
	signal I21560: std_logic; attribute dont_touch of I21560: signal is true;
	signal I21563: std_logic; attribute dont_touch of I21563: signal is true;
	signal I21566: std_logic; attribute dont_touch of I21566: signal is true;
	signal I21569: std_logic; attribute dont_touch of I21569: signal is true;
	signal I21577: std_logic; attribute dont_touch of I21577: signal is true;
	signal I21580: std_logic; attribute dont_touch of I21580: signal is true;
	signal I21583: std_logic; attribute dont_touch of I21583: signal is true;
	signal I21586: std_logic; attribute dont_touch of I21586: signal is true;
	signal I21595: std_logic; attribute dont_touch of I21595: signal is true;
	signal I21598: std_logic; attribute dont_touch of I21598: signal is true;
	signal I21601: std_logic; attribute dont_touch of I21601: signal is true;
	signal I21609: std_logic; attribute dont_touch of I21609: signal is true;
	signal I21612: std_logic; attribute dont_touch of I21612: signal is true;
	signal I21615: std_logic; attribute dont_touch of I21615: signal is true;
	signal I21626: std_logic; attribute dont_touch of I21626: signal is true;
	signal I21629: std_logic; attribute dont_touch of I21629: signal is true;
	signal I21632: std_logic; attribute dont_touch of I21632: signal is true;
	signal I21638: std_logic; attribute dont_touch of I21638: signal is true;
	signal I21641: std_logic; attribute dont_touch of I21641: signal is true;
	signal I21644: std_logic; attribute dont_touch of I21644: signal is true;
	signal I21647: std_logic; attribute dont_touch of I21647: signal is true;
	signal I21655: std_logic; attribute dont_touch of I21655: signal is true;
	signal I21658: std_logic; attribute dont_touch of I21658: signal is true;
	signal I21661: std_logic; attribute dont_touch of I21661: signal is true;
	signal I21666: std_logic; attribute dont_touch of I21666: signal is true;
	signal I21674: std_logic; attribute dont_touch of I21674: signal is true;
	signal I21677: std_logic; attribute dont_touch of I21677: signal is true;
	signal I21680: std_logic; attribute dont_touch of I21680: signal is true;
	signal I21688: std_logic; attribute dont_touch of I21688: signal is true;
	signal I21691: std_logic; attribute dont_touch of I21691: signal is true;
	signal I21694: std_logic; attribute dont_touch of I21694: signal is true;
	signal I21705: std_logic; attribute dont_touch of I21705: signal is true;
	signal I21708: std_logic; attribute dont_touch of I21708: signal is true;
	signal I21711: std_logic; attribute dont_touch of I21711: signal is true;
	signal I21720: std_logic; attribute dont_touch of I21720: signal is true;
	signal I21723: std_logic; attribute dont_touch of I21723: signal is true;
	signal I21726: std_logic; attribute dont_touch of I21726: signal is true;
	signal I21730: std_logic; attribute dont_touch of I21730: signal is true;
	signal I21736: std_logic; attribute dont_touch of I21736: signal is true;
	signal I21739: std_logic; attribute dont_touch of I21739: signal is true;
	signal I21742: std_logic; attribute dont_touch of I21742: signal is true;
	signal I21747: std_logic; attribute dont_touch of I21747: signal is true;
	signal I21755: std_logic; attribute dont_touch of I21755: signal is true;
	signal I21758: std_logic; attribute dont_touch of I21758: signal is true;
	signal I21761: std_logic; attribute dont_touch of I21761: signal is true;
	signal I21769: std_logic; attribute dont_touch of I21769: signal is true;
	signal I21772: std_logic; attribute dont_touch of I21772: signal is true;
	signal I21775: std_logic; attribute dont_touch of I21775: signal is true;
	signal I21780: std_logic; attribute dont_touch of I21780: signal is true;
	signal I21787: std_logic; attribute dont_touch of I21787: signal is true;
	signal I21790: std_logic; attribute dont_touch of I21790: signal is true;
	signal I21793: std_logic; attribute dont_touch of I21793: signal is true;
	signal I21796: std_logic; attribute dont_touch of I21796: signal is true;
	signal I21803: std_logic; attribute dont_touch of I21803: signal is true;
	signal I21806: std_logic; attribute dont_touch of I21806: signal is true;
	signal I21809: std_logic; attribute dont_touch of I21809: signal is true;
	signal I21813: std_logic; attribute dont_touch of I21813: signal is true;
	signal I21819: std_logic; attribute dont_touch of I21819: signal is true;
	signal I21822: std_logic; attribute dont_touch of I21822: signal is true;
	signal I21825: std_logic; attribute dont_touch of I21825: signal is true;
	signal I21830: std_logic; attribute dont_touch of I21830: signal is true;
	signal I21838: std_logic; attribute dont_touch of I21838: signal is true;
	signal I21841: std_logic; attribute dont_touch of I21841: signal is true;
	signal I21844: std_logic; attribute dont_touch of I21844: signal is true;
	signal I21852: std_logic; attribute dont_touch of I21852: signal is true;
	signal I21855: std_logic; attribute dont_touch of I21855: signal is true;
	signal I21862: std_logic; attribute dont_touch of I21862: signal is true;
	signal I21865: std_logic; attribute dont_touch of I21865: signal is true;
	signal I21868: std_logic; attribute dont_touch of I21868: signal is true;
	signal I21871: std_logic; attribute dont_touch of I21871: signal is true;
	signal I21878: std_logic; attribute dont_touch of I21878: signal is true;
	signal I21881: std_logic; attribute dont_touch of I21881: signal is true;
	signal I21884: std_logic; attribute dont_touch of I21884: signal is true;
	signal I21888: std_logic; attribute dont_touch of I21888: signal is true;
	signal I21894: std_logic; attribute dont_touch of I21894: signal is true;
	signal I21897: std_logic; attribute dont_touch of I21897: signal is true;
	signal I21900: std_logic; attribute dont_touch of I21900: signal is true;
	signal I21905: std_logic; attribute dont_touch of I21905: signal is true;
	signal I21908: std_logic; attribute dont_touch of I21908: signal is true;
	signal I21918: std_logic; attribute dont_touch of I21918: signal is true;
	signal I21923: std_logic; attribute dont_touch of I21923: signal is true;
	signal I21926: std_logic; attribute dont_touch of I21926: signal is true;
	signal I21933: std_logic; attribute dont_touch of I21933: signal is true;
	signal I21936: std_logic; attribute dont_touch of I21936: signal is true;
	signal I21939: std_logic; attribute dont_touch of I21939: signal is true;
	signal I21942: std_logic; attribute dont_touch of I21942: signal is true;
	signal I21949: std_logic; attribute dont_touch of I21949: signal is true;
	signal I21952: std_logic; attribute dont_touch of I21952: signal is true;
	signal I21955: std_logic; attribute dont_touch of I21955: signal is true;
	signal I21959: std_logic; attribute dont_touch of I21959: signal is true;
	signal I21962: std_logic; attribute dont_touch of I21962: signal is true;
	signal I21974: std_logic; attribute dont_touch of I21974: signal is true;
	signal I21979: std_logic; attribute dont_touch of I21979: signal is true;
	signal I21982: std_logic; attribute dont_touch of I21982: signal is true;
	signal I21989: std_logic; attribute dont_touch of I21989: signal is true;
	signal I21992: std_logic; attribute dont_touch of I21992: signal is true;
	signal I21995: std_logic; attribute dont_touch of I21995: signal is true;
	signal I21998: std_logic; attribute dont_touch of I21998: signal is true;
	signal I22014: std_logic; attribute dont_touch of I22014: signal is true;
	signal I22019: std_logic; attribute dont_touch of I22019: signal is true;
	signal I22022: std_logic; attribute dont_touch of I22022: signal is true;
	signal I22025: std_logic; attribute dont_touch of I22025: signal is true;
	signal I22028: std_logic; attribute dont_touch of I22028: signal is true;
	signal I22044: std_logic; attribute dont_touch of I22044: signal is true;
	signal I22062: std_logic; attribute dont_touch of I22062: signal is true;
	signal I22063: std_logic; attribute dont_touch of I22063: signal is true;
	signal I22064: std_logic; attribute dont_touch of I22064: signal is true;
	signal I22120: std_logic; attribute dont_touch of I22120: signal is true;
	signal I22136: std_logic; attribute dont_touch of I22136: signal is true;
	signal I22163: std_logic; attribute dont_touch of I22163: signal is true;
	signal I22282: std_logic; attribute dont_touch of I22282: signal is true;
	signal I22283: std_logic; attribute dont_touch of I22283: signal is true;
	signal I22284: std_logic; attribute dont_touch of I22284: signal is true;
	signal I22316: std_logic; attribute dont_touch of I22316: signal is true;
	signal I22317: std_logic; attribute dont_touch of I22317: signal is true;
	signal I22318: std_logic; attribute dont_touch of I22318: signal is true;
	signal I22382: std_logic; attribute dont_touch of I22382: signal is true;
	signal I22414: std_logic; attribute dont_touch of I22414: signal is true;
	signal I22444: std_logic; attribute dont_touch of I22444: signal is true;
	signal I22475: std_logic; attribute dont_touch of I22475: signal is true;
	signal I22503: std_logic; attribute dont_touch of I22503: signal is true;
	signal I22506: std_logic; attribute dont_touch of I22506: signal is true;
	signal I22509: std_logic; attribute dont_touch of I22509: signal is true;
	signal I22512: std_logic; attribute dont_touch of I22512: signal is true;
	signal I22515: std_logic; attribute dont_touch of I22515: signal is true;
	signal I22518: std_logic; attribute dont_touch of I22518: signal is true;
	signal I22521: std_logic; attribute dont_touch of I22521: signal is true;
	signal I22524: std_logic; attribute dont_touch of I22524: signal is true;
	signal I22527: std_logic; attribute dont_touch of I22527: signal is true;
	signal I22530: std_logic; attribute dont_touch of I22530: signal is true;
	signal I22533: std_logic; attribute dont_touch of I22533: signal is true;
	signal I22536: std_logic; attribute dont_touch of I22536: signal is true;
	signal I22539: std_logic; attribute dont_touch of I22539: signal is true;
	signal I22542: std_logic; attribute dont_touch of I22542: signal is true;
	signal I22545: std_logic; attribute dont_touch of I22545: signal is true;
	signal I22548: std_logic; attribute dont_touch of I22548: signal is true;
	signal I22551: std_logic; attribute dont_touch of I22551: signal is true;
	signal I22554: std_logic; attribute dont_touch of I22554: signal is true;
	signal I22557: std_logic; attribute dont_touch of I22557: signal is true;
	signal I22560: std_logic; attribute dont_touch of I22560: signal is true;
	signal I22563: std_logic; attribute dont_touch of I22563: signal is true;
	signal I22566: std_logic; attribute dont_touch of I22566: signal is true;
	signal I22569: std_logic; attribute dont_touch of I22569: signal is true;
	signal I22572: std_logic; attribute dont_touch of I22572: signal is true;
	signal I22575: std_logic; attribute dont_touch of I22575: signal is true;
	signal I22578: std_logic; attribute dont_touch of I22578: signal is true;
	signal I22581: std_logic; attribute dont_touch of I22581: signal is true;
	signal I22584: std_logic; attribute dont_touch of I22584: signal is true;
	signal I22587: std_logic; attribute dont_touch of I22587: signal is true;
	signal I22590: std_logic; attribute dont_touch of I22590: signal is true;
	signal I22593: std_logic; attribute dont_touch of I22593: signal is true;
	signal I22599: std_logic; attribute dont_touch of I22599: signal is true;
	signal I22604: std_logic; attribute dont_touch of I22604: signal is true;
	signal I22611: std_logic; attribute dont_touch of I22611: signal is true;
	signal I22618: std_logic; attribute dont_touch of I22618: signal is true;
	signal I22626: std_logic; attribute dont_touch of I22626: signal is true;
	signal I22630: std_logic; attribute dont_touch of I22630: signal is true;
	signal I22631: std_logic; attribute dont_touch of I22631: signal is true;
	signal I22632: std_logic; attribute dont_touch of I22632: signal is true;
	signal I22640: std_logic; attribute dont_touch of I22640: signal is true;
	signal I22651: std_logic; attribute dont_touch of I22651: signal is true;
	signal I22657: std_logic; attribute dont_touch of I22657: signal is true;
	signal I22663: std_logic; attribute dont_touch of I22663: signal is true;
	signal I22667: std_logic; attribute dont_touch of I22667: signal is true;
	signal I22671: std_logic; attribute dont_touch of I22671: signal is true;
	signal I22676: std_logic; attribute dont_touch of I22676: signal is true;
	signal I22679: std_logic; attribute dont_touch of I22679: signal is true;
	signal I22683: std_logic; attribute dont_touch of I22683: signal is true;
	signal I22687: std_logic; attribute dont_touch of I22687: signal is true;
	signal I22690: std_logic; attribute dont_touch of I22690: signal is true;
	signal I22694: std_logic; attribute dont_touch of I22694: signal is true;
	signal I22699: std_logic; attribute dont_touch of I22699: signal is true;
	signal I22702: std_logic; attribute dont_touch of I22702: signal is true;
	signal I22705: std_logic; attribute dont_touch of I22705: signal is true;
	signal I22706: std_logic; attribute dont_touch of I22706: signal is true;
	signal I22707: std_logic; attribute dont_touch of I22707: signal is true;
	signal I22715: std_logic; attribute dont_touch of I22715: signal is true;
	signal I22718: std_logic; attribute dont_touch of I22718: signal is true;
	signal I22726: std_logic; attribute dont_touch of I22726: signal is true;
	signal I22730: std_logic; attribute dont_touch of I22730: signal is true;
	signal I22737: std_logic; attribute dont_touch of I22737: signal is true;
	signal I22741: std_logic; attribute dont_touch of I22741: signal is true;
	signal I22745: std_logic; attribute dont_touch of I22745: signal is true;
	signal I22752: std_logic; attribute dont_touch of I22752: signal is true;
	signal I22755: std_logic; attribute dont_touch of I22755: signal is true;
	signal I22759: std_logic; attribute dont_touch of I22759: signal is true;
	signal I22763: std_logic; attribute dont_touch of I22763: signal is true;
	signal I22768: std_logic; attribute dont_touch of I22768: signal is true;
	signal I22771: std_logic; attribute dont_touch of I22771: signal is true;
	signal I22775: std_logic; attribute dont_touch of I22775: signal is true;
	signal I22783: std_logic; attribute dont_touch of I22783: signal is true;
	signal I22786: std_logic; attribute dont_touch of I22786: signal is true;
	signal I22789: std_logic; attribute dont_touch of I22789: signal is true;
	signal I22797: std_logic; attribute dont_touch of I22797: signal is true;
	signal I22800: std_logic; attribute dont_touch of I22800: signal is true;
	signal I22803: std_logic; attribute dont_touch of I22803: signal is true;
	signal I22810: std_logic; attribute dont_touch of I22810: signal is true;
	signal I22813: std_logic; attribute dont_touch of I22813: signal is true;
	signal I22820: std_logic; attribute dont_touch of I22820: signal is true;
	signal I22823: std_logic; attribute dont_touch of I22823: signal is true;
	signal I22828: std_logic; attribute dont_touch of I22828: signal is true;
	signal I22836: std_logic; attribute dont_touch of I22836: signal is true;
	signal I22842: std_logic; attribute dont_touch of I22842: signal is true;
	signal I22845: std_logic; attribute dont_touch of I22845: signal is true;
	signal I22852: std_logic; attribute dont_touch of I22852: signal is true;
	signal I22855: std_logic; attribute dont_touch of I22855: signal is true;
	signal I22860: std_logic; attribute dont_touch of I22860: signal is true;
	signal I22866: std_logic; attribute dont_touch of I22866: signal is true;
	signal I22869: std_logic; attribute dont_touch of I22869: signal is true;
	signal I22875: std_logic; attribute dont_touch of I22875: signal is true;
	signal I22881: std_logic; attribute dont_touch of I22881: signal is true;
	signal I22884: std_logic; attribute dont_touch of I22884: signal is true;
	signal I22885: std_logic; attribute dont_touch of I22885: signal is true;
	signal I22886: std_logic; attribute dont_touch of I22886: signal is true;
	signal I22893: std_logic; attribute dont_touch of I22893: signal is true;
	signal I22900: std_logic; attribute dont_touch of I22900: signal is true;
	signal I22901: std_logic; attribute dont_touch of I22901: signal is true;
	signal I22902: std_logic; attribute dont_touch of I22902: signal is true;
	signal I22912: std_logic; attribute dont_touch of I22912: signal is true;
	signal I22917: std_logic; attribute dont_touch of I22917: signal is true;
	signal I22918: std_logic; attribute dont_touch of I22918: signal is true;
	signal I22919: std_logic; attribute dont_touch of I22919: signal is true;
	signal I22924: std_logic; attribute dont_touch of I22924: signal is true;
	signal I22925: std_logic; attribute dont_touch of I22925: signal is true;
	signal I22926: std_logic; attribute dont_touch of I22926: signal is true;
	signal I22936: std_logic; attribute dont_touch of I22936: signal is true;
	signal I22937: std_logic; attribute dont_touch of I22937: signal is true;
	signal I22938: std_logic; attribute dont_touch of I22938: signal is true;
	signal I22945: std_logic; attribute dont_touch of I22945: signal is true;
	signal I22946: std_logic; attribute dont_touch of I22946: signal is true;
	signal I22947: std_logic; attribute dont_touch of I22947: signal is true;
	signal I22952: std_logic; attribute dont_touch of I22952: signal is true;
	signal I22953: std_logic; attribute dont_touch of I22953: signal is true;
	signal I22954: std_logic; attribute dont_touch of I22954: signal is true;
	signal I22962: std_logic; attribute dont_touch of I22962: signal is true;
	signal I22963: std_logic; attribute dont_touch of I22963: signal is true;
	signal I22964: std_logic; attribute dont_touch of I22964: signal is true;
	signal I22972: std_logic; attribute dont_touch of I22972: signal is true;
	signal I22973: std_logic; attribute dont_touch of I22973: signal is true;
	signal I22974: std_logic; attribute dont_touch of I22974: signal is true;
	signal I22981: std_logic; attribute dont_touch of I22981: signal is true;
	signal I22982: std_logic; attribute dont_touch of I22982: signal is true;
	signal I22983: std_logic; attribute dont_touch of I22983: signal is true;
	signal I22988: std_logic; attribute dont_touch of I22988: signal is true;
	signal I22989: std_logic; attribute dont_touch of I22989: signal is true;
	signal I22990: std_logic; attribute dont_touch of I22990: signal is true;
	signal I22998: std_logic; attribute dont_touch of I22998: signal is true;
	signal I22999: std_logic; attribute dont_touch of I22999: signal is true;
	signal I23000: std_logic; attribute dont_touch of I23000: signal is true;
	signal I23008: std_logic; attribute dont_touch of I23008: signal is true;
	signal I23009: std_logic; attribute dont_touch of I23009: signal is true;
	signal I23010: std_logic; attribute dont_touch of I23010: signal is true;
	signal I23018: std_logic; attribute dont_touch of I23018: signal is true;
	signal I23019: std_logic; attribute dont_touch of I23019: signal is true;
	signal I23020: std_logic; attribute dont_touch of I23020: signal is true;
	signal I23027: std_logic; attribute dont_touch of I23027: signal is true;
	signal I23028: std_logic; attribute dont_touch of I23028: signal is true;
	signal I23029: std_logic; attribute dont_touch of I23029: signal is true;
	signal I23034: std_logic; attribute dont_touch of I23034: signal is true;
	signal I23035: std_logic; attribute dont_touch of I23035: signal is true;
	signal I23036: std_logic; attribute dont_touch of I23036: signal is true;
	signal I23045: std_logic; attribute dont_touch of I23045: signal is true;
	signal I23046: std_logic; attribute dont_touch of I23046: signal is true;
	signal I23047: std_logic; attribute dont_touch of I23047: signal is true;
	signal I23055: std_logic; attribute dont_touch of I23055: signal is true;
	signal I23056: std_logic; attribute dont_touch of I23056: signal is true;
	signal I23057: std_logic; attribute dont_touch of I23057: signal is true;
	signal I23065: std_logic; attribute dont_touch of I23065: signal is true;
	signal I23066: std_logic; attribute dont_touch of I23066: signal is true;
	signal I23067: std_logic; attribute dont_touch of I23067: signal is true;
	signal I23074: std_logic; attribute dont_touch of I23074: signal is true;
	signal I23075: std_logic; attribute dont_touch of I23075: signal is true;
	signal I23076: std_logic; attribute dont_touch of I23076: signal is true;
	signal I23082: std_logic; attribute dont_touch of I23082: signal is true;
	signal I23083: std_logic; attribute dont_touch of I23083: signal is true;
	signal I23084: std_logic; attribute dont_touch of I23084: signal is true;
	signal I23093: std_logic; attribute dont_touch of I23093: signal is true;
	signal I23094: std_logic; attribute dont_touch of I23094: signal is true;
	signal I23095: std_logic; attribute dont_touch of I23095: signal is true;
	signal I23103: std_logic; attribute dont_touch of I23103: signal is true;
	signal I23104: std_logic; attribute dont_touch of I23104: signal is true;
	signal I23105: std_logic; attribute dont_touch of I23105: signal is true;
	signal I23113: std_logic; attribute dont_touch of I23113: signal is true;
	signal I23114: std_logic; attribute dont_touch of I23114: signal is true;
	signal I23115: std_logic; attribute dont_touch of I23115: signal is true;
	signal I23123: std_logic; attribute dont_touch of I23123: signal is true;
	signal I23124: std_logic; attribute dont_touch of I23124: signal is true;
	signal I23125: std_logic; attribute dont_touch of I23125: signal is true;
	signal I23131: std_logic; attribute dont_touch of I23131: signal is true;
	signal I23132: std_logic; attribute dont_touch of I23132: signal is true;
	signal I23133: std_logic; attribute dont_touch of I23133: signal is true;
	signal I23142: std_logic; attribute dont_touch of I23142: signal is true;
	signal I23143: std_logic; attribute dont_touch of I23143: signal is true;
	signal I23144: std_logic; attribute dont_touch of I23144: signal is true;
	signal I23152: std_logic; attribute dont_touch of I23152: signal is true;
	signal I23153: std_logic; attribute dont_touch of I23153: signal is true;
	signal I23154: std_logic; attribute dont_touch of I23154: signal is true;
	signal I23161: std_logic; attribute dont_touch of I23161: signal is true;
	signal I23162: std_logic; attribute dont_touch of I23162: signal is true;
	signal I23163: std_logic; attribute dont_touch of I23163: signal is true;
	signal I23171: std_logic; attribute dont_touch of I23171: signal is true;
	signal I23172: std_logic; attribute dont_touch of I23172: signal is true;
	signal I23173: std_logic; attribute dont_touch of I23173: signal is true;
	signal I23179: std_logic; attribute dont_touch of I23179: signal is true;
	signal I23180: std_logic; attribute dont_touch of I23180: signal is true;
	signal I23181: std_logic; attribute dont_touch of I23181: signal is true;
	signal I23190: std_logic; attribute dont_touch of I23190: signal is true;
	signal I23191: std_logic; attribute dont_touch of I23191: signal is true;
	signal I23192: std_logic; attribute dont_touch of I23192: signal is true;
	signal I23198: std_logic; attribute dont_touch of I23198: signal is true;
	signal I23199: std_logic; attribute dont_touch of I23199: signal is true;
	signal I23200: std_logic; attribute dont_touch of I23200: signal is true;
	signal I23207: std_logic; attribute dont_touch of I23207: signal is true;
	signal I23208: std_logic; attribute dont_touch of I23208: signal is true;
	signal I23209: std_logic; attribute dont_touch of I23209: signal is true;
	signal I23217: std_logic; attribute dont_touch of I23217: signal is true;
	signal I23218: std_logic; attribute dont_touch of I23218: signal is true;
	signal I23219: std_logic; attribute dont_touch of I23219: signal is true;
	signal I23225: std_logic; attribute dont_touch of I23225: signal is true;
	signal I23226: std_logic; attribute dont_touch of I23226: signal is true;
	signal I23227: std_logic; attribute dont_touch of I23227: signal is true;
	signal I23233: std_logic; attribute dont_touch of I23233: signal is true;
	signal I23234: std_logic; attribute dont_touch of I23234: signal is true;
	signal I23235: std_logic; attribute dont_touch of I23235: signal is true;
	signal I23242: std_logic; attribute dont_touch of I23242: signal is true;
	signal I23243: std_logic; attribute dont_touch of I23243: signal is true;
	signal I23244: std_logic; attribute dont_touch of I23244: signal is true;
	signal I23253: std_logic; attribute dont_touch of I23253: signal is true;
	signal I23256: std_logic; attribute dont_touch of I23256: signal is true;
	signal I23257: std_logic; attribute dont_touch of I23257: signal is true;
	signal I23258: std_logic; attribute dont_touch of I23258: signal is true;
	signal I23264: std_logic; attribute dont_touch of I23264: signal is true;
	signal I23265: std_logic; attribute dont_touch of I23265: signal is true;
	signal I23266: std_logic; attribute dont_touch of I23266: signal is true;
	signal I23274: std_logic; attribute dont_touch of I23274: signal is true;
	signal I23277: std_logic; attribute dont_touch of I23277: signal is true;
	signal I23278: std_logic; attribute dont_touch of I23278: signal is true;
	signal I23279: std_logic; attribute dont_touch of I23279: signal is true;
	signal I23287: std_logic; attribute dont_touch of I23287: signal is true;
	signal I23292: std_logic; attribute dont_touch of I23292: signal is true;
	signal I23309: std_logic; attribute dont_touch of I23309: signal is true;
	signal I23314: std_logic; attribute dont_touch of I23314: signal is true;
	signal I23317: std_logic; attribute dont_touch of I23317: signal is true;
	signal I23323: std_logic; attribute dont_touch of I23323: signal is true;
	signal I23326: std_logic; attribute dont_touch of I23326: signal is true;
	signal I23329: std_logic; attribute dont_touch of I23329: signal is true;
	signal I23335: std_logic; attribute dont_touch of I23335: signal is true;
	signal I23338: std_logic; attribute dont_touch of I23338: signal is true;
	signal I23341: std_logic; attribute dont_touch of I23341: signal is true;
	signal I23345: std_logic; attribute dont_touch of I23345: signal is true;
	signal I23348: std_logic; attribute dont_touch of I23348: signal is true;
	signal I23351: std_logic; attribute dont_touch of I23351: signal is true;
	signal I23358: std_logic; attribute dont_touch of I23358: signal is true;
	signal I23361: std_logic; attribute dont_touch of I23361: signal is true;
	signal I23364: std_logic; attribute dont_touch of I23364: signal is true;
	signal I23368: std_logic; attribute dont_touch of I23368: signal is true;
	signal I23371: std_logic; attribute dont_touch of I23371: signal is true;
	signal I23374: std_logic; attribute dont_touch of I23374: signal is true;
	signal I23377: std_logic; attribute dont_touch of I23377: signal is true;
	signal I23380: std_logic; attribute dont_touch of I23380: signal is true;
	signal I23383: std_logic; attribute dont_touch of I23383: signal is true;
	signal I23386: std_logic; attribute dont_touch of I23386: signal is true;
	signal I23392: std_logic; attribute dont_touch of I23392: signal is true;
	signal I23395: std_logic; attribute dont_touch of I23395: signal is true;
	signal I23398: std_logic; attribute dont_touch of I23398: signal is true;
	signal I23403: std_logic; attribute dont_touch of I23403: signal is true;
	signal I23406: std_logic; attribute dont_touch of I23406: signal is true;
	signal I23409: std_logic; attribute dont_touch of I23409: signal is true;
	signal I23412: std_logic; attribute dont_touch of I23412: signal is true;
	signal I23415: std_logic; attribute dont_touch of I23415: signal is true;
	signal I23418: std_logic; attribute dont_touch of I23418: signal is true;
	signal I23421: std_logic; attribute dont_touch of I23421: signal is true;
	signal I23424: std_logic; attribute dont_touch of I23424: signal is true;
	signal I23430: std_logic; attribute dont_touch of I23430: signal is true;
	signal I23433: std_logic; attribute dont_touch of I23433: signal is true;
	signal I23436: std_logic; attribute dont_touch of I23436: signal is true;
	signal I23442: std_logic; attribute dont_touch of I23442: signal is true;
	signal I23445: std_logic; attribute dont_touch of I23445: signal is true;
	signal I23448: std_logic; attribute dont_touch of I23448: signal is true;
	signal I23451: std_logic; attribute dont_touch of I23451: signal is true;
	signal I23454: std_logic; attribute dont_touch of I23454: signal is true;
	signal I23457: std_logic; attribute dont_touch of I23457: signal is true;
	signal I23460: std_logic; attribute dont_touch of I23460: signal is true;
	signal I23463: std_logic; attribute dont_touch of I23463: signal is true;
	signal I23466: std_logic; attribute dont_touch of I23466: signal is true;
	signal I23472: std_logic; attribute dont_touch of I23472: signal is true;
	signal I23475: std_logic; attribute dont_touch of I23475: signal is true;
	signal I23478: std_logic; attribute dont_touch of I23478: signal is true;
	signal I23487: std_logic; attribute dont_touch of I23487: signal is true;
	signal I23490: std_logic; attribute dont_touch of I23490: signal is true;
	signal I23493: std_logic; attribute dont_touch of I23493: signal is true;
	signal I23498: std_logic; attribute dont_touch of I23498: signal is true;
	signal I23501: std_logic; attribute dont_touch of I23501: signal is true;
	signal I23504: std_logic; attribute dont_touch of I23504: signal is true;
	signal I23507: std_logic; attribute dont_touch of I23507: signal is true;
	signal I23510: std_logic; attribute dont_touch of I23510: signal is true;
	signal I23513: std_logic; attribute dont_touch of I23513: signal is true;
	signal I23518: std_logic; attribute dont_touch of I23518: signal is true;
	signal I23521: std_logic; attribute dont_touch of I23521: signal is true;
	signal I23524: std_logic; attribute dont_touch of I23524: signal is true;
	signal I23527: std_logic; attribute dont_touch of I23527: signal is true;
	signal I23530: std_logic; attribute dont_touch of I23530: signal is true;
	signal I23539: std_logic; attribute dont_touch of I23539: signal is true;
	signal I23542: std_logic; attribute dont_touch of I23542: signal is true;
	signal I23545: std_logic; attribute dont_touch of I23545: signal is true;
	signal I23553: std_logic; attribute dont_touch of I23553: signal is true;
	signal I23556: std_logic; attribute dont_touch of I23556: signal is true;
	signal I23559: std_logic; attribute dont_touch of I23559: signal is true;
	signal I23564: std_logic; attribute dont_touch of I23564: signal is true;
	signal I23567: std_logic; attribute dont_touch of I23567: signal is true;
	signal I23570: std_logic; attribute dont_touch of I23570: signal is true;
	signal I23575: std_logic; attribute dont_touch of I23575: signal is true;
	signal I23578: std_logic; attribute dont_touch of I23578: signal is true;
	signal I23581: std_logic; attribute dont_touch of I23581: signal is true;
	signal I23584: std_logic; attribute dont_touch of I23584: signal is true;
	signal I23588: std_logic; attribute dont_touch of I23588: signal is true;
	signal I23591: std_logic; attribute dont_touch of I23591: signal is true;
	signal I23599: std_logic; attribute dont_touch of I23599: signal is true;
	signal I23602: std_logic; attribute dont_touch of I23602: signal is true;
	signal I23605: std_logic; attribute dont_touch of I23605: signal is true;
	signal I23608: std_logic; attribute dont_touch of I23608: signal is true;
	signal I23611: std_logic; attribute dont_touch of I23611: signal is true;
	signal I23619: std_logic; attribute dont_touch of I23619: signal is true;
	signal I23622: std_logic; attribute dont_touch of I23622: signal is true;
	signal I23625: std_logic; attribute dont_touch of I23625: signal is true;
	signal I23633: std_logic; attribute dont_touch of I23633: signal is true;
	signal I23636: std_logic; attribute dont_touch of I23636: signal is true;
	signal I23639: std_logic; attribute dont_touch of I23639: signal is true;
	signal I23645: std_logic; attribute dont_touch of I23645: signal is true;
	signal I23648: std_logic; attribute dont_touch of I23648: signal is true;
	signal I23651: std_logic; attribute dont_touch of I23651: signal is true;
	signal I23655: std_logic; attribute dont_touch of I23655: signal is true;
	signal I23658: std_logic; attribute dont_touch of I23658: signal is true;
	signal I23661: std_logic; attribute dont_touch of I23661: signal is true;
	signal I23667: std_logic; attribute dont_touch of I23667: signal is true;
	signal I23670: std_logic; attribute dont_touch of I23670: signal is true;
	signal I23673: std_logic; attribute dont_touch of I23673: signal is true;
	signal I23676: std_logic; attribute dont_touch of I23676: signal is true;
	signal I23679: std_logic; attribute dont_touch of I23679: signal is true;
	signal I23682: std_logic; attribute dont_touch of I23682: signal is true;
	signal I23689: std_logic; attribute dont_touch of I23689: signal is true;
	signal I23692: std_logic; attribute dont_touch of I23692: signal is true;
	signal I23695: std_logic; attribute dont_touch of I23695: signal is true;
	signal I23698: std_logic; attribute dont_touch of I23698: signal is true;
	signal I23701: std_logic; attribute dont_touch of I23701: signal is true;
	signal I23709: std_logic; attribute dont_touch of I23709: signal is true;
	signal I23712: std_logic; attribute dont_touch of I23712: signal is true;
	signal I23715: std_logic; attribute dont_touch of I23715: signal is true;
	signal I23725: std_logic; attribute dont_touch of I23725: signal is true;
	signal I23729: std_logic; attribute dont_touch of I23729: signal is true;
	signal I23733: std_logic; attribute dont_touch of I23733: signal is true;
	signal I23739: std_logic; attribute dont_touch of I23739: signal is true;
	signal I23742: std_logic; attribute dont_touch of I23742: signal is true;
	signal I23745: std_logic; attribute dont_touch of I23745: signal is true;
	signal I23748: std_logic; attribute dont_touch of I23748: signal is true;
	signal I23751: std_logic; attribute dont_touch of I23751: signal is true;
	signal I23754: std_logic; attribute dont_touch of I23754: signal is true;
	signal I23760: std_logic; attribute dont_touch of I23760: signal is true;
	signal I23763: std_logic; attribute dont_touch of I23763: signal is true;
	signal I23766: std_logic; attribute dont_touch of I23766: signal is true;
	signal I23769: std_logic; attribute dont_touch of I23769: signal is true;
	signal I23772: std_logic; attribute dont_touch of I23772: signal is true;
	signal I23775: std_logic; attribute dont_touch of I23775: signal is true;
	signal I23782: std_logic; attribute dont_touch of I23782: signal is true;
	signal I23785: std_logic; attribute dont_touch of I23785: signal is true;
	signal I23788: std_logic; attribute dont_touch of I23788: signal is true;
	signal I23791: std_logic; attribute dont_touch of I23791: signal is true;
	signal I23794: std_logic; attribute dont_touch of I23794: signal is true;
	signal I23806: std_logic; attribute dont_touch of I23806: signal is true;
	signal I23807: std_logic; attribute dont_touch of I23807: signal is true;
	signal I23808: std_logic; attribute dont_touch of I23808: signal is true;
	signal I23817: std_logic; attribute dont_touch of I23817: signal is true;
	signal I23821: std_logic; attribute dont_touch of I23821: signal is true;
	signal I23824: std_logic; attribute dont_touch of I23824: signal is true;
	signal I23830: std_logic; attribute dont_touch of I23830: signal is true;
	signal I23833: std_logic; attribute dont_touch of I23833: signal is true;
	signal I23836: std_logic; attribute dont_touch of I23836: signal is true;
	signal I23839: std_logic; attribute dont_touch of I23839: signal is true;
	signal I23842: std_logic; attribute dont_touch of I23842: signal is true;
	signal I23845: std_logic; attribute dont_touch of I23845: signal is true;
	signal I23851: std_logic; attribute dont_touch of I23851: signal is true;
	signal I23854: std_logic; attribute dont_touch of I23854: signal is true;
	signal I23857: std_logic; attribute dont_touch of I23857: signal is true;
	signal I23860: std_logic; attribute dont_touch of I23860: signal is true;
	signal I23863: std_logic; attribute dont_touch of I23863: signal is true;
	signal I23866: std_logic; attribute dont_touch of I23866: signal is true;
	signal I23874: std_logic; attribute dont_touch of I23874: signal is true;
	signal I23878: std_logic; attribute dont_touch of I23878: signal is true;
	signal I23879: std_logic; attribute dont_touch of I23879: signal is true;
	signal I23880: std_logic; attribute dont_touch of I23880: signal is true;
	signal I23888: std_logic; attribute dont_touch of I23888: signal is true;
	signal I23893: std_logic; attribute dont_touch of I23893: signal is true;
	signal I23894: std_logic; attribute dont_touch of I23894: signal is true;
	signal I23895: std_logic; attribute dont_touch of I23895: signal is true;
	signal I23904: std_logic; attribute dont_touch of I23904: signal is true;
	signal I23908: std_logic; attribute dont_touch of I23908: signal is true;
	signal I23911: std_logic; attribute dont_touch of I23911: signal is true;
	signal I23917: std_logic; attribute dont_touch of I23917: signal is true;
	signal I23920: std_logic; attribute dont_touch of I23920: signal is true;
	signal I23923: std_logic; attribute dont_touch of I23923: signal is true;
	signal I23926: std_logic; attribute dont_touch of I23926: signal is true;
	signal I23929: std_logic; attribute dont_touch of I23929: signal is true;
	signal I23932: std_logic; attribute dont_touch of I23932: signal is true;
	signal I23941: std_logic; attribute dont_touch of I23941: signal is true;
	signal I23942: std_logic; attribute dont_touch of I23942: signal is true;
	signal I23943: std_logic; attribute dont_touch of I23943: signal is true;
	signal I23954: std_logic; attribute dont_touch of I23954: signal is true;
	signal I23958: std_logic; attribute dont_touch of I23958: signal is true;
	signal I23959: std_logic; attribute dont_touch of I23959: signal is true;
	signal I23960: std_logic; attribute dont_touch of I23960: signal is true;
	signal I23966: std_logic; attribute dont_touch of I23966: signal is true;
	signal I23967: std_logic; attribute dont_touch of I23967: signal is true;
	signal I23968: std_logic; attribute dont_touch of I23968: signal is true;
	signal I23976: std_logic; attribute dont_touch of I23976: signal is true;
	signal I23981: std_logic; attribute dont_touch of I23981: signal is true;
	signal I23982: std_logic; attribute dont_touch of I23982: signal is true;
	signal I23983: std_logic; attribute dont_touch of I23983: signal is true;
	signal I23992: std_logic; attribute dont_touch of I23992: signal is true;
	signal I23996: std_logic; attribute dont_touch of I23996: signal is true;
	signal I23999: std_logic; attribute dont_touch of I23999: signal is true;
	signal I24005: std_logic; attribute dont_touch of I24005: signal is true;
	signal I24006: std_logic; attribute dont_touch of I24006: signal is true;
	signal I24007: std_logic; attribute dont_touch of I24007: signal is true;
	signal I24015: std_logic; attribute dont_touch of I24015: signal is true;
	signal I24016: std_logic; attribute dont_touch of I24016: signal is true;
	signal I24017: std_logic; attribute dont_touch of I24017: signal is true;
	signal I24028: std_logic; attribute dont_touch of I24028: signal is true;
	signal I24029: std_logic; attribute dont_touch of I24029: signal is true;
	signal I24030: std_logic; attribute dont_touch of I24030: signal is true;
	signal I24036: std_logic; attribute dont_touch of I24036: signal is true;
	signal I24037: std_logic; attribute dont_touch of I24037: signal is true;
	signal I24038: std_logic; attribute dont_touch of I24038: signal is true;
	signal I24049: std_logic; attribute dont_touch of I24049: signal is true;
	signal I24053: std_logic; attribute dont_touch of I24053: signal is true;
	signal I24054: std_logic; attribute dont_touch of I24054: signal is true;
	signal I24055: std_logic; attribute dont_touch of I24055: signal is true;
	signal I24061: std_logic; attribute dont_touch of I24061: signal is true;
	signal I24062: std_logic; attribute dont_touch of I24062: signal is true;
	signal I24063: std_logic; attribute dont_touch of I24063: signal is true;
	signal I24071: std_logic; attribute dont_touch of I24071: signal is true;
	signal I24076: std_logic; attribute dont_touch of I24076: signal is true;
	signal I24077: std_logic; attribute dont_touch of I24077: signal is true;
	signal I24078: std_logic; attribute dont_touch of I24078: signal is true;
	signal I24091: std_logic; attribute dont_touch of I24091: signal is true;
	signal I24092: std_logic; attribute dont_touch of I24092: signal is true;
	signal I24093: std_logic; attribute dont_touch of I24093: signal is true;
	signal I24102: std_logic; attribute dont_touch of I24102: signal is true;
	signal I24103: std_logic; attribute dont_touch of I24103: signal is true;
	signal I24104: std_logic; attribute dont_touch of I24104: signal is true;
	signal I24110: std_logic; attribute dont_touch of I24110: signal is true;
	signal I24111: std_logic; attribute dont_touch of I24111: signal is true;
	signal I24112: std_logic; attribute dont_touch of I24112: signal is true;
	signal I24123: std_logic; attribute dont_touch of I24123: signal is true;
	signal I24124: std_logic; attribute dont_touch of I24124: signal is true;
	signal I24125: std_logic; attribute dont_touch of I24125: signal is true;
	signal I24131: std_logic; attribute dont_touch of I24131: signal is true;
	signal I24132: std_logic; attribute dont_touch of I24132: signal is true;
	signal I24133: std_logic; attribute dont_touch of I24133: signal is true;
	signal I24144: std_logic; attribute dont_touch of I24144: signal is true;
	signal I24148: std_logic; attribute dont_touch of I24148: signal is true;
	signal I24149: std_logic; attribute dont_touch of I24149: signal is true;
	signal I24150: std_logic; attribute dont_touch of I24150: signal is true;
	signal I24156: std_logic; attribute dont_touch of I24156: signal is true;
	signal I24157: std_logic; attribute dont_touch of I24157: signal is true;
	signal I24158: std_logic; attribute dont_touch of I24158: signal is true;
	signal I24166: std_logic; attribute dont_touch of I24166: signal is true;
	signal I24171: std_logic; attribute dont_touch of I24171: signal is true;
	signal I24178: std_logic; attribute dont_touch of I24178: signal is true;
	signal I24179: std_logic; attribute dont_touch of I24179: signal is true;
	signal I24180: std_logic; attribute dont_touch of I24180: signal is true;
	signal I24186: std_logic; attribute dont_touch of I24186: signal is true;
	signal I24187: std_logic; attribute dont_touch of I24187: signal is true;
	signal I24188: std_logic; attribute dont_touch of I24188: signal is true;
	signal I24194: std_logic; attribute dont_touch of I24194: signal is true;
	signal I24195: std_logic; attribute dont_touch of I24195: signal is true;
	signal I24196: std_logic; attribute dont_touch of I24196: signal is true;
	signal I24205: std_logic; attribute dont_touch of I24205: signal is true;
	signal I24206: std_logic; attribute dont_touch of I24206: signal is true;
	signal I24207: std_logic; attribute dont_touch of I24207: signal is true;
	signal I24213: std_logic; attribute dont_touch of I24213: signal is true;
	signal I24214: std_logic; attribute dont_touch of I24214: signal is true;
	signal I24215: std_logic; attribute dont_touch of I24215: signal is true;
	signal I24226: std_logic; attribute dont_touch of I24226: signal is true;
	signal I24227: std_logic; attribute dont_touch of I24227: signal is true;
	signal I24228: std_logic; attribute dont_touch of I24228: signal is true;
	signal I24234: std_logic; attribute dont_touch of I24234: signal is true;
	signal I24235: std_logic; attribute dont_touch of I24235: signal is true;
	signal I24236: std_logic; attribute dont_touch of I24236: signal is true;
	signal I24247: std_logic; attribute dont_touch of I24247: signal is true;
	signal I24251: std_logic; attribute dont_touch of I24251: signal is true;
	signal I24252: std_logic; attribute dont_touch of I24252: signal is true;
	signal I24253: std_logic; attribute dont_touch of I24253: signal is true;
	signal I24258: std_logic; attribute dont_touch of I24258: signal is true;
	signal I24263: std_logic; attribute dont_touch of I24263: signal is true;
	signal I24264: std_logic; attribute dont_touch of I24264: signal is true;
	signal I24265: std_logic; attribute dont_touch of I24265: signal is true;
	signal I24271: std_logic; attribute dont_touch of I24271: signal is true;
	signal I24272: std_logic; attribute dont_touch of I24272: signal is true;
	signal I24273: std_logic; attribute dont_touch of I24273: signal is true;
	signal I24278: std_logic; attribute dont_touch of I24278: signal is true;
	signal I24279: std_logic; attribute dont_touch of I24279: signal is true;
	signal I24280: std_logic; attribute dont_touch of I24280: signal is true;
	signal I24285: std_logic; attribute dont_touch of I24285: signal is true;
	signal I24290: std_logic; attribute dont_touch of I24290: signal is true;
	signal I24291: std_logic; attribute dont_touch of I24291: signal is true;
	signal I24292: std_logic; attribute dont_touch of I24292: signal is true;
	signal I24298: std_logic; attribute dont_touch of I24298: signal is true;
	signal I24299: std_logic; attribute dont_touch of I24299: signal is true;
	signal I24300: std_logic; attribute dont_touch of I24300: signal is true;
	signal I24306: std_logic; attribute dont_touch of I24306: signal is true;
	signal I24307: std_logic; attribute dont_touch of I24307: signal is true;
	signal I24308: std_logic; attribute dont_touch of I24308: signal is true;
	signal I24317: std_logic; attribute dont_touch of I24317: signal is true;
	signal I24318: std_logic; attribute dont_touch of I24318: signal is true;
	signal I24319: std_logic; attribute dont_touch of I24319: signal is true;
	signal I24325: std_logic; attribute dont_touch of I24325: signal is true;
	signal I24326: std_logic; attribute dont_touch of I24326: signal is true;
	signal I24327: std_logic; attribute dont_touch of I24327: signal is true;
	signal I24338: std_logic; attribute dont_touch of I24338: signal is true;
	signal I24339: std_logic; attribute dont_touch of I24339: signal is true;
	signal I24340: std_logic; attribute dont_touch of I24340: signal is true;
	signal I24346: std_logic; attribute dont_touch of I24346: signal is true;
	signal I24351: std_logic; attribute dont_touch of I24351: signal is true;
	signal I24352: std_logic; attribute dont_touch of I24352: signal is true;
	signal I24353: std_logic; attribute dont_touch of I24353: signal is true;
	signal I24361: std_logic; attribute dont_touch of I24361: signal is true;
	signal I24362: std_logic; attribute dont_touch of I24362: signal is true;
	signal I24363: std_logic; attribute dont_touch of I24363: signal is true;
	signal I24368: std_logic; attribute dont_touch of I24368: signal is true;
	signal I24372: std_logic; attribute dont_touch of I24372: signal is true;
	signal I24373: std_logic; attribute dont_touch of I24373: signal is true;
	signal I24374: std_logic; attribute dont_touch of I24374: signal is true;
	signal I24380: std_logic; attribute dont_touch of I24380: signal is true;
	signal I24381: std_logic; attribute dont_touch of I24381: signal is true;
	signal I24382: std_logic; attribute dont_touch of I24382: signal is true;
	signal I24387: std_logic; attribute dont_touch of I24387: signal is true;
	signal I24388: std_logic; attribute dont_touch of I24388: signal is true;
	signal I24389: std_logic; attribute dont_touch of I24389: signal is true;
	signal I24394: std_logic; attribute dont_touch of I24394: signal is true;
	signal I24399: std_logic; attribute dont_touch of I24399: signal is true;
	signal I24400: std_logic; attribute dont_touch of I24400: signal is true;
	signal I24401: std_logic; attribute dont_touch of I24401: signal is true;
	signal I24407: std_logic; attribute dont_touch of I24407: signal is true;
	signal I24408: std_logic; attribute dont_touch of I24408: signal is true;
	signal I24409: std_logic; attribute dont_touch of I24409: signal is true;
	signal I24415: std_logic; attribute dont_touch of I24415: signal is true;
	signal I24416: std_logic; attribute dont_touch of I24416: signal is true;
	signal I24417: std_logic; attribute dont_touch of I24417: signal is true;
	signal I24426: std_logic; attribute dont_touch of I24426: signal is true;
	signal I24427: std_logic; attribute dont_touch of I24427: signal is true;
	signal I24428: std_logic; attribute dont_touch of I24428: signal is true;
	signal I24436: std_logic; attribute dont_touch of I24436: signal is true;
	signal I24437: std_logic; attribute dont_touch of I24437: signal is true;
	signal I24438: std_logic; attribute dont_touch of I24438: signal is true;
	signal I24443: std_logic; attribute dont_touch of I24443: signal is true;
	signal I24444: std_logic; attribute dont_touch of I24444: signal is true;
	signal I24445: std_logic; attribute dont_touch of I24445: signal is true;
	signal I24452: std_logic; attribute dont_touch of I24452: signal is true;
	signal I24453: std_logic; attribute dont_touch of I24453: signal is true;
	signal I24454: std_logic; attribute dont_touch of I24454: signal is true;
	signal I24459: std_logic; attribute dont_touch of I24459: signal is true;
	signal I24464: std_logic; attribute dont_touch of I24464: signal is true;
	signal I24465: std_logic; attribute dont_touch of I24465: signal is true;
	signal I24466: std_logic; attribute dont_touch of I24466: signal is true;
	signal I24474: std_logic; attribute dont_touch of I24474: signal is true;
	signal I24475: std_logic; attribute dont_touch of I24475: signal is true;
	signal I24476: std_logic; attribute dont_touch of I24476: signal is true;
	signal I24481: std_logic; attribute dont_touch of I24481: signal is true;
	signal I24485: std_logic; attribute dont_touch of I24485: signal is true;
	signal I24486: std_logic; attribute dont_touch of I24486: signal is true;
	signal I24487: std_logic; attribute dont_touch of I24487: signal is true;
	signal I24493: std_logic; attribute dont_touch of I24493: signal is true;
	signal I24494: std_logic; attribute dont_touch of I24494: signal is true;
	signal I24495: std_logic; attribute dont_touch of I24495: signal is true;
	signal I24500: std_logic; attribute dont_touch of I24500: signal is true;
	signal I24501: std_logic; attribute dont_touch of I24501: signal is true;
	signal I24502: std_logic; attribute dont_touch of I24502: signal is true;
	signal I24507: std_logic; attribute dont_touch of I24507: signal is true;
	signal I24512: std_logic; attribute dont_touch of I24512: signal is true;
	signal I24513: std_logic; attribute dont_touch of I24513: signal is true;
	signal I24514: std_logic; attribute dont_touch of I24514: signal is true;
	signal I24520: std_logic; attribute dont_touch of I24520: signal is true;
	signal I24521: std_logic; attribute dont_touch of I24521: signal is true;
	signal I24522: std_logic; attribute dont_touch of I24522: signal is true;
	signal I24530: std_logic; attribute dont_touch of I24530: signal is true;
	signal I24531: std_logic; attribute dont_touch of I24531: signal is true;
	signal I24532: std_logic; attribute dont_touch of I24532: signal is true;
	signal I24537: std_logic; attribute dont_touch of I24537: signal is true;
	signal I24538: std_logic; attribute dont_touch of I24538: signal is true;
	signal I24539: std_logic; attribute dont_touch of I24539: signal is true;
	signal I24544: std_logic; attribute dont_touch of I24544: signal is true;
	signal I24545: std_logic; attribute dont_touch of I24545: signal is true;
	signal I24546: std_logic; attribute dont_touch of I24546: signal is true;
	signal I24553: std_logic; attribute dont_touch of I24553: signal is true;
	signal I24554: std_logic; attribute dont_touch of I24554: signal is true;
	signal I24555: std_logic; attribute dont_touch of I24555: signal is true;
	signal I24560: std_logic; attribute dont_touch of I24560: signal is true;
	signal I24565: std_logic; attribute dont_touch of I24565: signal is true;
	signal I24566: std_logic; attribute dont_touch of I24566: signal is true;
	signal I24567: std_logic; attribute dont_touch of I24567: signal is true;
	signal I24575: std_logic; attribute dont_touch of I24575: signal is true;
	signal I24576: std_logic; attribute dont_touch of I24576: signal is true;
	signal I24577: std_logic; attribute dont_touch of I24577: signal is true;
	signal I24582: std_logic; attribute dont_touch of I24582: signal is true;
	signal I24586: std_logic; attribute dont_touch of I24586: signal is true;
	signal I24587: std_logic; attribute dont_touch of I24587: signal is true;
	signal I24588: std_logic; attribute dont_touch of I24588: signal is true;
	signal I24594: std_logic; attribute dont_touch of I24594: signal is true;
	signal I24595: std_logic; attribute dont_touch of I24595: signal is true;
	signal I24596: std_logic; attribute dont_touch of I24596: signal is true;
	signal I24601: std_logic; attribute dont_touch of I24601: signal is true;
	signal I24602: std_logic; attribute dont_touch of I24602: signal is true;
	signal I24603: std_logic; attribute dont_touch of I24603: signal is true;
	signal I24608: std_logic; attribute dont_touch of I24608: signal is true;
	signal I24611: std_logic; attribute dont_touch of I24611: signal is true;
	signal I24612: std_logic; attribute dont_touch of I24612: signal is true;
	signal I24613: std_logic; attribute dont_touch of I24613: signal is true;
	signal I24619: std_logic; attribute dont_touch of I24619: signal is true;
	signal I24624: std_logic; attribute dont_touch of I24624: signal is true;
	signal I24625: std_logic; attribute dont_touch of I24625: signal is true;
	signal I24626: std_logic; attribute dont_touch of I24626: signal is true;
	signal I24632: std_logic; attribute dont_touch of I24632: signal is true;
	signal I24633: std_logic; attribute dont_touch of I24633: signal is true;
	signal I24634: std_logic; attribute dont_touch of I24634: signal is true;
	signal I24639: std_logic; attribute dont_touch of I24639: signal is true;
	signal I24640: std_logic; attribute dont_touch of I24640: signal is true;
	signal I24641: std_logic; attribute dont_touch of I24641: signal is true;
	signal I24646: std_logic; attribute dont_touch of I24646: signal is true;
	signal I24647: std_logic; attribute dont_touch of I24647: signal is true;
	signal I24648: std_logic; attribute dont_touch of I24648: signal is true;
	signal I24655: std_logic; attribute dont_touch of I24655: signal is true;
	signal I24656: std_logic; attribute dont_touch of I24656: signal is true;
	signal I24657: std_logic; attribute dont_touch of I24657: signal is true;
	signal I24662: std_logic; attribute dont_touch of I24662: signal is true;
	signal I24667: std_logic; attribute dont_touch of I24667: signal is true;
	signal I24668: std_logic; attribute dont_touch of I24668: signal is true;
	signal I24669: std_logic; attribute dont_touch of I24669: signal is true;
	signal I24677: std_logic; attribute dont_touch of I24677: signal is true;
	signal I24678: std_logic; attribute dont_touch of I24678: signal is true;
	signal I24679: std_logic; attribute dont_touch of I24679: signal is true;
	signal I24684: std_logic; attribute dont_touch of I24684: signal is true;
	signal I24689: std_logic; attribute dont_touch of I24689: signal is true;
	signal I24694: std_logic; attribute dont_touch of I24694: signal is true;
	signal I24695: std_logic; attribute dont_touch of I24695: signal is true;
	signal I24696: std_logic; attribute dont_touch of I24696: signal is true;
	signal I24702: std_logic; attribute dont_touch of I24702: signal is true;
	signal I24703: std_logic; attribute dont_touch of I24703: signal is true;
	signal I24704: std_logic; attribute dont_touch of I24704: signal is true;
	signal I24709: std_logic; attribute dont_touch of I24709: signal is true;
	signal I24710: std_logic; attribute dont_touch of I24710: signal is true;
	signal I24711: std_logic; attribute dont_touch of I24711: signal is true;
	signal I24716: std_logic; attribute dont_touch of I24716: signal is true;
	signal I24717: std_logic; attribute dont_touch of I24717: signal is true;
	signal I24718: std_logic; attribute dont_touch of I24718: signal is true;
	signal I24725: std_logic; attribute dont_touch of I24725: signal is true;
	signal I24726: std_logic; attribute dont_touch of I24726: signal is true;
	signal I24727: std_logic; attribute dont_touch of I24727: signal is true;
	signal I24732: std_logic; attribute dont_touch of I24732: signal is true;
	signal I24738: std_logic; attribute dont_touch of I24738: signal is true;
	signal I24743: std_logic; attribute dont_touch of I24743: signal is true;
	signal I24744: std_logic; attribute dont_touch of I24744: signal is true;
	signal I24745: std_logic; attribute dont_touch of I24745: signal is true;
	signal I24751: std_logic; attribute dont_touch of I24751: signal is true;
	signal I24752: std_logic; attribute dont_touch of I24752: signal is true;
	signal I24753: std_logic; attribute dont_touch of I24753: signal is true;
	signal I24758: std_logic; attribute dont_touch of I24758: signal is true;
	signal I24763: std_logic; attribute dont_touch of I24763: signal is true;
	signal I24764: std_logic; attribute dont_touch of I24764: signal is true;
	signal I24765: std_logic; attribute dont_touch of I24765: signal is true;
	signal I24894: std_logic; attribute dont_touch of I24894: signal is true;
	signal I24913: std_logic; attribute dont_touch of I24913: signal is true;
	signal I24916: std_logic; attribute dont_touch of I24916: signal is true;
	signal I24923: std_logic; attribute dont_touch of I24923: signal is true;
	signal I24943: std_logic; attribute dont_touch of I24943: signal is true;
	signal I24950: std_logic; attribute dont_touch of I24950: signal is true;
	signal I24966: std_logic; attribute dont_touch of I24966: signal is true;
	signal I24973: std_logic; attribute dont_touch of I24973: signal is true;
	signal I24982: std_logic; attribute dont_touch of I24982: signal is true;
	signal I24992: std_logic; attribute dont_touch of I24992: signal is true;
	signal I25001: std_logic; attribute dont_touch of I25001: signal is true;
	signal I25004: std_logic; attribute dont_touch of I25004: signal is true;
	signal I25015: std_logic; attribute dont_touch of I25015: signal is true;
	signal I25018: std_logic; attribute dont_touch of I25018: signal is true;
	signal I25021: std_logic; attribute dont_touch of I25021: signal is true;
	signal I25030: std_logic; attribute dont_touch of I25030: signal is true;
	signal I25031: std_logic; attribute dont_touch of I25031: signal is true;
	signal I25032: std_logic; attribute dont_touch of I25032: signal is true;
	signal I25037: std_logic; attribute dont_touch of I25037: signal is true;
	signal I25041: std_logic; attribute dont_touch of I25041: signal is true;
	signal I25044: std_logic; attribute dont_touch of I25044: signal is true;
	signal I25047: std_logic; attribute dont_touch of I25047: signal is true;
	signal I25050: std_logic; attribute dont_touch of I25050: signal is true;
	signal I25054: std_logic; attribute dont_touch of I25054: signal is true;
	signal I25057: std_logic; attribute dont_touch of I25057: signal is true;
	signal I25061: std_logic; attribute dont_touch of I25061: signal is true;
	signal I25064: std_logic; attribute dont_touch of I25064: signal is true;
	signal I25067: std_logic; attribute dont_touch of I25067: signal is true;
	signal I25071: std_logic; attribute dont_touch of I25071: signal is true;
	signal I25074: std_logic; attribute dont_touch of I25074: signal is true;
	signal I25078: std_logic; attribute dont_touch of I25078: signal is true;
	signal I25081: std_logic; attribute dont_touch of I25081: signal is true;
	signal I25084: std_logic; attribute dont_touch of I25084: signal is true;
	signal I25089: std_logic; attribute dont_touch of I25089: signal is true;
	signal I25092: std_logic; attribute dont_touch of I25092: signal is true;
	signal I25096: std_logic; attribute dont_touch of I25096: signal is true;
	signal I25099: std_logic; attribute dont_touch of I25099: signal is true;
	signal I25102: std_logic; attribute dont_touch of I25102: signal is true;
	signal I25105: std_logic; attribute dont_touch of I25105: signal is true;
	signal I25108: std_logic; attribute dont_touch of I25108: signal is true;
	signal I25111: std_logic; attribute dont_touch of I25111: signal is true;
	signal I25114: std_logic; attribute dont_touch of I25114: signal is true;
	signal I25117: std_logic; attribute dont_touch of I25117: signal is true;
	signal I25120: std_logic; attribute dont_touch of I25120: signal is true;
	signal I25123: std_logic; attribute dont_touch of I25123: signal is true;
	signal I25126: std_logic; attribute dont_touch of I25126: signal is true;
	signal I25129: std_logic; attribute dont_touch of I25129: signal is true;
	signal I25132: std_logic; attribute dont_touch of I25132: signal is true;
	signal I25135: std_logic; attribute dont_touch of I25135: signal is true;
	signal I25138: std_logic; attribute dont_touch of I25138: signal is true;
	signal I25141: std_logic; attribute dont_touch of I25141: signal is true;
	signal I25144: std_logic; attribute dont_touch of I25144: signal is true;
	signal I25147: std_logic; attribute dont_touch of I25147: signal is true;
	signal I25150: std_logic; attribute dont_touch of I25150: signal is true;
	signal I25153: std_logic; attribute dont_touch of I25153: signal is true;
	signal I25156: std_logic; attribute dont_touch of I25156: signal is true;
	signal I25159: std_logic; attribute dont_touch of I25159: signal is true;
	signal I25162: std_logic; attribute dont_touch of I25162: signal is true;
	signal I25165: std_logic; attribute dont_touch of I25165: signal is true;
	signal I25168: std_logic; attribute dont_touch of I25168: signal is true;
	signal I25171: std_logic; attribute dont_touch of I25171: signal is true;
	signal I25174: std_logic; attribute dont_touch of I25174: signal is true;
	signal I25177: std_logic; attribute dont_touch of I25177: signal is true;
	signal I25180: std_logic; attribute dont_touch of I25180: signal is true;
	signal I25183: std_logic; attribute dont_touch of I25183: signal is true;
	signal I25186: std_logic; attribute dont_touch of I25186: signal is true;
	signal I25189: std_logic; attribute dont_touch of I25189: signal is true;
	signal I25192: std_logic; attribute dont_touch of I25192: signal is true;
	signal I25195: std_logic; attribute dont_touch of I25195: signal is true;
	signal I25198: std_logic; attribute dont_touch of I25198: signal is true;
	signal I25201: std_logic; attribute dont_touch of I25201: signal is true;
	signal I25204: std_logic; attribute dont_touch of I25204: signal is true;
	signal I25207: std_logic; attribute dont_touch of I25207: signal is true;
	signal I25210: std_logic; attribute dont_touch of I25210: signal is true;
	signal I25213: std_logic; attribute dont_touch of I25213: signal is true;
	signal I25216: std_logic; attribute dont_touch of I25216: signal is true;
	signal I25219: std_logic; attribute dont_touch of I25219: signal is true;
	signal I25222: std_logic; attribute dont_touch of I25222: signal is true;
	signal I25225: std_logic; attribute dont_touch of I25225: signal is true;
	signal I25228: std_logic; attribute dont_touch of I25228: signal is true;
	signal I25231: std_logic; attribute dont_touch of I25231: signal is true;
	signal I25234: std_logic; attribute dont_touch of I25234: signal is true;
	signal I25237: std_logic; attribute dont_touch of I25237: signal is true;
	signal I25240: std_logic; attribute dont_touch of I25240: signal is true;
	signal I25243: std_logic; attribute dont_touch of I25243: signal is true;
	signal I25246: std_logic; attribute dont_touch of I25246: signal is true;
	signal I25249: std_logic; attribute dont_touch of I25249: signal is true;
	signal I25253: std_logic; attribute dont_touch of I25253: signal is true;
	signal I25258: std_logic; attribute dont_touch of I25258: signal is true;
	signal I25264: std_logic; attribute dont_touch of I25264: signal is true;
	signal I25272: std_logic; attribute dont_touch of I25272: signal is true;
	signal I25280: std_logic; attribute dont_touch of I25280: signal is true;
	signal I25283: std_logic; attribute dont_touch of I25283: signal is true;
	signal I25291: std_logic; attribute dont_touch of I25291: signal is true;
	signal I25294: std_logic; attribute dont_touch of I25294: signal is true;
	signal I25300: std_logic; attribute dont_touch of I25300: signal is true;
	signal I25303: std_logic; attribute dont_touch of I25303: signal is true;
	signal I25308: std_logic; attribute dont_touch of I25308: signal is true;
	signal I25311: std_logic; attribute dont_touch of I25311: signal is true;
	signal I25315: std_logic; attribute dont_touch of I25315: signal is true;
	signal I25320: std_logic; attribute dont_touch of I25320: signal is true;
	signal I25325: std_logic; attribute dont_touch of I25325: signal is true;
	signal I25334: std_logic; attribute dont_touch of I25334: signal is true;
	signal I25338: std_logic; attribute dont_touch of I25338: signal is true;
	signal I25344: std_logic; attribute dont_touch of I25344: signal is true;
	signal I25351: std_logic; attribute dont_touch of I25351: signal is true;
	signal I25355: std_logic; attribute dont_touch of I25355: signal is true;
	signal I25358: std_logic; attribute dont_touch of I25358: signal is true;
	signal I25365: std_logic; attribute dont_touch of I25365: signal is true;
	signal I25371: std_logic; attribute dont_touch of I25371: signal is true;
	signal I25374: std_logic; attribute dont_touch of I25374: signal is true;
	signal I25377: std_logic; attribute dont_touch of I25377: signal is true;
	signal I25383: std_logic; attribute dont_touch of I25383: signal is true;
	signal I25386: std_logic; attribute dont_touch of I25386: signal is true;
	signal I25389: std_logic; attribute dont_touch of I25389: signal is true;
	signal I25395: std_logic; attribute dont_touch of I25395: signal is true;
	signal I25399: std_logic; attribute dont_touch of I25399: signal is true;
	signal I25402: std_logic; attribute dont_touch of I25402: signal is true;
	signal I25406: std_logic; attribute dont_touch of I25406: signal is true;
	signal I25412: std_logic; attribute dont_touch of I25412: signal is true;
	signal I25415: std_logic; attribute dont_touch of I25415: signal is true;
	signal I25423: std_logic; attribute dont_touch of I25423: signal is true;
	signal I25426: std_logic; attribute dont_touch of I25426: signal is true;
	signal I25429: std_logic; attribute dont_touch of I25429: signal is true;
	signal I25432: std_logic; attribute dont_touch of I25432: signal is true;
	signal I25442: std_logic; attribute dont_touch of I25442: signal is true;
	signal I25445: std_logic; attribute dont_touch of I25445: signal is true;
	signal I25456: std_logic; attribute dont_touch of I25456: signal is true;
	signal I25459: std_logic; attribute dont_touch of I25459: signal is true;
	signal I25463: std_logic; attribute dont_touch of I25463: signal is true;
	signal I25474: std_logic; attribute dont_touch of I25474: signal is true;
	signal I25477: std_logic; attribute dont_touch of I25477: signal is true;
	signal I25486: std_logic; attribute dont_touch of I25486: signal is true;
	signal I25489: std_logic; attribute dont_touch of I25489: signal is true;
	signal I25492: std_logic; attribute dont_touch of I25492: signal is true;
	signal I25495: std_logic; attribute dont_touch of I25495: signal is true;
	signal I25500: std_logic; attribute dont_touch of I25500: signal is true;
	signal I25506: std_logic; attribute dont_touch of I25506: signal is true;
	signal I25510: std_logic; attribute dont_touch of I25510: signal is true;
	signal I25516: std_logic; attribute dont_touch of I25516: signal is true;
	signal I25521: std_logic; attribute dont_touch of I25521: signal is true;
	signal I25525: std_logic; attribute dont_touch of I25525: signal is true;
	signal I25528: std_logic; attribute dont_touch of I25528: signal is true;
	signal I25532: std_logic; attribute dont_touch of I25532: signal is true;
	signal I25533: std_logic; attribute dont_touch of I25533: signal is true;
	signal I25534: std_logic; attribute dont_touch of I25534: signal is true;
	signal I25539: std_logic; attribute dont_touch of I25539: signal is true;
	signal I25540: std_logic; attribute dont_touch of I25540: signal is true;
	signal I25541: std_logic; attribute dont_touch of I25541: signal is true;
	signal I25549: std_logic; attribute dont_touch of I25549: signal is true;
	signal I25554: std_logic; attribute dont_touch of I25554: signal is true;
	signal I25557: std_logic; attribute dont_touch of I25557: signal is true;
	signal I25560: std_logic; attribute dont_touch of I25560: signal is true;
	signal I25561: std_logic; attribute dont_touch of I25561: signal is true;
	signal I25562: std_logic; attribute dont_touch of I25562: signal is true;
	signal I25567: std_logic; attribute dont_touch of I25567: signal is true;
	signal I25571: std_logic; attribute dont_touch of I25571: signal is true;
	signal I25572: std_logic; attribute dont_touch of I25572: signal is true;
	signal I25573: std_logic; attribute dont_touch of I25573: signal is true;
	signal I25578: std_logic; attribute dont_touch of I25578: signal is true;
	signal I25579: std_logic; attribute dont_touch of I25579: signal is true;
	signal I25580: std_logic; attribute dont_touch of I25580: signal is true;
	signal I25588: std_logic; attribute dont_touch of I25588: signal is true;
	signal I25595: std_logic; attribute dont_touch of I25595: signal is true;
	signal I25596: std_logic; attribute dont_touch of I25596: signal is true;
	signal I25597: std_logic; attribute dont_touch of I25597: signal is true;
	signal I25605: std_logic; attribute dont_touch of I25605: signal is true;
	signal I25606: std_logic; attribute dont_touch of I25606: signal is true;
	signal I25607: std_logic; attribute dont_touch of I25607: signal is true;
	signal I25612: std_logic; attribute dont_touch of I25612: signal is true;
	signal I25616: std_logic; attribute dont_touch of I25616: signal is true;
	signal I25617: std_logic; attribute dont_touch of I25617: signal is true;
	signal I25618: std_logic; attribute dont_touch of I25618: signal is true;
	signal I25623: std_logic; attribute dont_touch of I25623: signal is true;
	signal I25624: std_logic; attribute dont_touch of I25624: signal is true;
	signal I25625: std_logic; attribute dont_touch of I25625: signal is true;
	signal I25633: std_logic; attribute dont_touch of I25633: signal is true;
	signal I25634: std_logic; attribute dont_touch of I25634: signal is true;
	signal I25635: std_logic; attribute dont_touch of I25635: signal is true;
	signal I25643: std_logic; attribute dont_touch of I25643: signal is true;
	signal I25644: std_logic; attribute dont_touch of I25644: signal is true;
	signal I25645: std_logic; attribute dont_touch of I25645: signal is true;
	signal I25653: std_logic; attribute dont_touch of I25653: signal is true;
	signal I25654: std_logic; attribute dont_touch of I25654: signal is true;
	signal I25655: std_logic; attribute dont_touch of I25655: signal is true;
	signal I25660: std_logic; attribute dont_touch of I25660: signal is true;
	signal I25664: std_logic; attribute dont_touch of I25664: signal is true;
	signal I25665: std_logic; attribute dont_touch of I25665: signal is true;
	signal I25666: std_logic; attribute dont_touch of I25666: signal is true;
	signal I25671: std_logic; attribute dont_touch of I25671: signal is true;
	signal I25672: std_logic; attribute dont_touch of I25672: signal is true;
	signal I25673: std_logic; attribute dont_touch of I25673: signal is true;
	signal I25681: std_logic; attribute dont_touch of I25681: signal is true;
	signal I25682: std_logic; attribute dont_touch of I25682: signal is true;
	signal I25683: std_logic; attribute dont_touch of I25683: signal is true;
	signal I25690: std_logic; attribute dont_touch of I25690: signal is true;
	signal I25691: std_logic; attribute dont_touch of I25691: signal is true;
	signal I25692: std_logic; attribute dont_touch of I25692: signal is true;
	signal I25700: std_logic; attribute dont_touch of I25700: signal is true;
	signal I25701: std_logic; attribute dont_touch of I25701: signal is true;
	signal I25702: std_logic; attribute dont_touch of I25702: signal is true;
	signal I25710: std_logic; attribute dont_touch of I25710: signal is true;
	signal I25711: std_logic; attribute dont_touch of I25711: signal is true;
	signal I25712: std_logic; attribute dont_touch of I25712: signal is true;
	signal I25717: std_logic; attribute dont_touch of I25717: signal is true;
	signal I25721: std_logic; attribute dont_touch of I25721: signal is true;
	signal I25722: std_logic; attribute dont_touch of I25722: signal is true;
	signal I25723: std_logic; attribute dont_touch of I25723: signal is true;
	signal I25728: std_logic; attribute dont_touch of I25728: signal is true;
	signal I25731: std_logic; attribute dont_touch of I25731: signal is true;
	signal I25732: std_logic; attribute dont_touch of I25732: signal is true;
	signal I25733: std_logic; attribute dont_touch of I25733: signal is true;
	signal I25740: std_logic; attribute dont_touch of I25740: signal is true;
	signal I25741: std_logic; attribute dont_touch of I25741: signal is true;
	signal I25742: std_logic; attribute dont_touch of I25742: signal is true;
	signal I25750: std_logic; attribute dont_touch of I25750: signal is true;
	signal I25751: std_logic; attribute dont_touch of I25751: signal is true;
	signal I25752: std_logic; attribute dont_touch of I25752: signal is true;
	signal I25761: std_logic; attribute dont_touch of I25761: signal is true;
	signal I25762: std_logic; attribute dont_touch of I25762: signal is true;
	signal I25763: std_logic; attribute dont_touch of I25763: signal is true;
	signal I25768: std_logic; attribute dont_touch of I25768: signal is true;
	signal I25771: std_logic; attribute dont_touch of I25771: signal is true;
	signal I25772: std_logic; attribute dont_touch of I25772: signal is true;
	signal I25773: std_logic; attribute dont_touch of I25773: signal is true;
	signal I25778: std_logic; attribute dont_touch of I25778: signal is true;
	signal I25781: std_logic; attribute dont_touch of I25781: signal is true;
	signal I25782: std_logic; attribute dont_touch of I25782: signal is true;
	signal I25783: std_logic; attribute dont_touch of I25783: signal is true;
	signal I25790: std_logic; attribute dont_touch of I25790: signal is true;
	signal I25791: std_logic; attribute dont_touch of I25791: signal is true;
	signal I25792: std_logic; attribute dont_touch of I25792: signal is true;
	signal I25800: std_logic; attribute dont_touch of I25800: signal is true;
	signal I25801: std_logic; attribute dont_touch of I25801: signal is true;
	signal I25802: std_logic; attribute dont_touch of I25802: signal is true;
	signal I25809: std_logic; attribute dont_touch of I25809: signal is true;
	signal I25810: std_logic; attribute dont_touch of I25810: signal is true;
	signal I25811: std_logic; attribute dont_touch of I25811: signal is true;
	signal I25816: std_logic; attribute dont_touch of I25816: signal is true;
	signal I25819: std_logic; attribute dont_touch of I25819: signal is true;
	signal I25820: std_logic; attribute dont_touch of I25820: signal is true;
	signal I25821: std_logic; attribute dont_touch of I25821: signal is true;
	signal I25826: std_logic; attribute dont_touch of I25826: signal is true;
	signal I25829: std_logic; attribute dont_touch of I25829: signal is true;
	signal I25830: std_logic; attribute dont_touch of I25830: signal is true;
	signal I25831: std_logic; attribute dont_touch of I25831: signal is true;
	signal I25838: std_logic; attribute dont_touch of I25838: signal is true;
	signal I25839: std_logic; attribute dont_touch of I25839: signal is true;
	signal I25840: std_logic; attribute dont_touch of I25840: signal is true;
	signal I25846: std_logic; attribute dont_touch of I25846: signal is true;
	signal I25847: std_logic; attribute dont_touch of I25847: signal is true;
	signal I25848: std_logic; attribute dont_touch of I25848: signal is true;
	signal I25855: std_logic; attribute dont_touch of I25855: signal is true;
	signal I25856: std_logic; attribute dont_touch of I25856: signal is true;
	signal I25857: std_logic; attribute dont_touch of I25857: signal is true;
	signal I25862: std_logic; attribute dont_touch of I25862: signal is true;
	signal I25865: std_logic; attribute dont_touch of I25865: signal is true;
	signal I25866: std_logic; attribute dont_touch of I25866: signal is true;
	signal I25867: std_logic; attribute dont_touch of I25867: signal is true;
	signal I25872: std_logic; attribute dont_touch of I25872: signal is true;
	signal I25880: std_logic; attribute dont_touch of I25880: signal is true;
	signal I25881: std_logic; attribute dont_touch of I25881: signal is true;
	signal I25882: std_logic; attribute dont_touch of I25882: signal is true;
	signal I25888: std_logic; attribute dont_touch of I25888: signal is true;
	signal I25889: std_logic; attribute dont_touch of I25889: signal is true;
	signal I25890: std_logic; attribute dont_touch of I25890: signal is true;
	signal I25897: std_logic; attribute dont_touch of I25897: signal is true;
	signal I25898: std_logic; attribute dont_touch of I25898: signal is true;
	signal I25899: std_logic; attribute dont_touch of I25899: signal is true;
	signal I25904: std_logic; attribute dont_touch of I25904: signal is true;
	signal I25913: std_logic; attribute dont_touch of I25913: signal is true;
	signal I25914: std_logic; attribute dont_touch of I25914: signal is true;
	signal I25915: std_logic; attribute dont_touch of I25915: signal is true;
	signal I25921: std_logic; attribute dont_touch of I25921: signal is true;
	signal I25922: std_logic; attribute dont_touch of I25922: signal is true;
	signal I25923: std_logic; attribute dont_touch of I25923: signal is true;
	signal I25938: std_logic; attribute dont_touch of I25938: signal is true;
	signal I25939: std_logic; attribute dont_touch of I25939: signal is true;
	signal I25940: std_logic; attribute dont_touch of I25940: signal is true;
	signal I25966: std_logic; attribute dont_touch of I25966: signal is true;
	signal I25971: std_logic; attribute dont_touch of I25971: signal is true;
	signal I25977: std_logic; attribute dont_touch of I25977: signal is true;
	signal I25985: std_logic; attribute dont_touch of I25985: signal is true;
	signal I25994: std_logic; attribute dont_touch of I25994: signal is true;
	signal I26006: std_logic; attribute dont_touch of I26006: signal is true;
	signal I26025: std_logic; attribute dont_touch of I26025: signal is true;
	signal I26028: std_logic; attribute dont_touch of I26028: signal is true;
	signal I26051: std_logic; attribute dont_touch of I26051: signal is true;
	signal I26078: std_logic; attribute dont_touch of I26078: signal is true;
	signal I26085: std_logic; attribute dont_touch of I26085: signal is true;
	signal I26112: std_logic; attribute dont_touch of I26112: signal is true;
	signal I26115: std_logic; attribute dont_touch of I26115: signal is true;
	signal I26123: std_logic; attribute dont_touch of I26123: signal is true;
	signal I26134: std_logic; attribute dont_touch of I26134: signal is true;
	signal I26154: std_logic; attribute dont_touch of I26154: signal is true;
	signal I26171: std_logic; attribute dont_touch of I26171: signal is true;
	signal I26182: std_logic; attribute dont_touch of I26182: signal is true;
	signal I26195: std_logic; attribute dont_touch of I26195: signal is true;
	signal I26198: std_logic; attribute dont_touch of I26198: signal is true;
	signal I26220: std_logic; attribute dont_touch of I26220: signal is true;
	signal I26231: std_logic; attribute dont_touch of I26231: signal is true;
	signal I26237: std_logic; attribute dont_touch of I26237: signal is true;
	signal I26240: std_logic; attribute dont_touch of I26240: signal is true;
	signal I26266: std_logic; attribute dont_touch of I26266: signal is true;
	signal I26276: std_logic; attribute dont_touch of I26276: signal is true;
	signal I26282: std_logic; attribute dont_touch of I26282: signal is true;
	signal I26285: std_logic; attribute dont_touch of I26285: signal is true;
	signal I26311: std_logic; attribute dont_touch of I26311: signal is true;
	signal I26317: std_logic; attribute dont_touch of I26317: signal is true;
	signal I26320: std_logic; attribute dont_touch of I26320: signal is true;
	signal I26334: std_logic; attribute dont_touch of I26334: signal is true;
	signal I26337: std_logic; attribute dont_touch of I26337: signal is true;
	signal I26340: std_logic; attribute dont_touch of I26340: signal is true;
	signal I26348: std_logic; attribute dont_touch of I26348: signal is true;
	signal I26354: std_logic; attribute dont_touch of I26354: signal is true;
	signal I26357: std_logic; attribute dont_touch of I26357: signal is true;
	signal I26365: std_logic; attribute dont_touch of I26365: signal is true;
	signal I26369: std_logic; attribute dont_touch of I26369: signal is true;
	signal I26377: std_logic; attribute dont_touch of I26377: signal is true;
	signal I26383: std_logic; attribute dont_touch of I26383: signal is true;
	signal I26388: std_logic; attribute dont_touch of I26388: signal is true;
	signal I26396: std_logic; attribute dont_touch of I26396: signal is true;
	signal I26401: std_logic; attribute dont_touch of I26401: signal is true;
	signal I26407: std_logic; attribute dont_touch of I26407: signal is true;
	signal I26413: std_logic; attribute dont_touch of I26413: signal is true;
	signal I26416: std_logic; attribute dont_touch of I26416: signal is true;
	signal I26420: std_logic; attribute dont_touch of I26420: signal is true;
	signal I26426: std_logic; attribute dont_touch of I26426: signal is true;
	signal I26429: std_logic; attribute dont_touch of I26429: signal is true;
	signal I26432: std_logic; attribute dont_touch of I26432: signal is true;
	signal I26437: std_logic; attribute dont_touch of I26437: signal is true;
	signal I26440: std_logic; attribute dont_touch of I26440: signal is true;
	signal I26444: std_logic; attribute dont_touch of I26444: signal is true;
	signal I26455: std_logic; attribute dont_touch of I26455: signal is true;
	signal I26458: std_logic; attribute dont_touch of I26458: signal is true;
	signal I26461: std_logic; attribute dont_touch of I26461: signal is true;
	signal I26464: std_logic; attribute dont_touch of I26464: signal is true;
	signal I26469: std_logic; attribute dont_touch of I26469: signal is true;
	signal I26472: std_logic; attribute dont_touch of I26472: signal is true;
	signal I26476: std_logic; attribute dont_touch of I26476: signal is true;
	signal I26481: std_logic; attribute dont_touch of I26481: signal is true;
	signal I26491: std_logic; attribute dont_touch of I26491: signal is true;
	signal I26494: std_logic; attribute dont_touch of I26494: signal is true;
	signal I26497: std_logic; attribute dont_touch of I26497: signal is true;
	signal I26500: std_logic; attribute dont_touch of I26500: signal is true;
	signal I26505: std_logic; attribute dont_touch of I26505: signal is true;
	signal I26508: std_logic; attribute dont_touch of I26508: signal is true;
	signal I26512: std_logic; attribute dont_touch of I26512: signal is true;
	signal I26525: std_logic; attribute dont_touch of I26525: signal is true;
	signal I26528: std_logic; attribute dont_touch of I26528: signal is true;
	signal I26532: std_logic; attribute dont_touch of I26532: signal is true;
	signal I26535: std_logic; attribute dont_touch of I26535: signal is true;
	signal I26538: std_logic; attribute dont_touch of I26538: signal is true;
	signal I26541: std_logic; attribute dont_touch of I26541: signal is true;
	signal I26545: std_logic; attribute dont_touch of I26545: signal is true;
	signal I26558: std_logic; attribute dont_touch of I26558: signal is true;
	signal I26561: std_logic; attribute dont_touch of I26561: signal is true;
	signal I26564: std_logic; attribute dont_touch of I26564: signal is true;
	signal I26567: std_logic; attribute dont_touch of I26567: signal is true;
	signal I26571: std_logic; attribute dont_touch of I26571: signal is true;
	signal I26574: std_logic; attribute dont_touch of I26574: signal is true;
	signal I26590: std_logic; attribute dont_touch of I26590: signal is true;
	signal I26593: std_logic; attribute dont_touch of I26593: signal is true;
	signal I26596: std_logic; attribute dont_touch of I26596: signal is true;
	signal I26599: std_logic; attribute dont_touch of I26599: signal is true;
	signal I26612: std_logic; attribute dont_touch of I26612: signal is true;
	signal I26615: std_logic; attribute dont_touch of I26615: signal is true;
	signal I26621: std_logic; attribute dont_touch of I26621: signal is true;
	signal I26624: std_logic; attribute dont_touch of I26624: signal is true;
	signal I26627: std_logic; attribute dont_touch of I26627: signal is true;
	signal I26630: std_logic; attribute dont_touch of I26630: signal is true;
	signal I26639: std_logic; attribute dont_touch of I26639: signal is true;
	signal I26642: std_logic; attribute dont_touch of I26642: signal is true;
	signal I26645: std_logic; attribute dont_touch of I26645: signal is true;
	signal I26651: std_logic; attribute dont_touch of I26651: signal is true;
	signal I26654: std_logic; attribute dont_touch of I26654: signal is true;
	signal I26661: std_logic; attribute dont_touch of I26661: signal is true;
	signal I26664: std_logic; attribute dont_touch of I26664: signal is true;
	signal I26667: std_logic; attribute dont_touch of I26667: signal is true;
	signal I26676: std_logic; attribute dont_touch of I26676: signal is true;
	signal I26679: std_logic; attribute dont_touch of I26679: signal is true;
	signal I26682: std_logic; attribute dont_touch of I26682: signal is true;
	signal I26690: std_logic; attribute dont_touch of I26690: signal is true;
	signal I26695: std_logic; attribute dont_touch of I26695: signal is true;
	signal I26708: std_logic; attribute dont_touch of I26708: signal is true;
	signal I26714: std_logic; attribute dont_touch of I26714: signal is true;
	signal I26726: std_logic; attribute dont_touch of I26726: signal is true;
	signal I26745: std_logic; attribute dont_touch of I26745: signal is true;
	signal I26777: std_logic; attribute dont_touch of I26777: signal is true;
	signal I26796: std_logic; attribute dont_touch of I26796: signal is true;
	signal I26816: std_logic; attribute dont_touch of I26816: signal is true;
	signal I26819: std_logic; attribute dont_touch of I26819: signal is true;
	signal I26843: std_logic; attribute dont_touch of I26843: signal is true;
	signal I26846: std_logic; attribute dont_touch of I26846: signal is true;
	signal I26868: std_logic; attribute dont_touch of I26868: signal is true;
	signal I26871: std_logic; attribute dont_touch of I26871: signal is true;
	signal I26874: std_logic; attribute dont_touch of I26874: signal is true;
	signal I26892: std_logic; attribute dont_touch of I26892: signal is true;
	signal I26895: std_logic; attribute dont_touch of I26895: signal is true;
	signal I26898: std_logic; attribute dont_touch of I26898: signal is true;
	signal I26910: std_logic; attribute dont_touch of I26910: signal is true;
	signal I26913: std_logic; attribute dont_touch of I26913: signal is true;
	signal I26916: std_logic; attribute dont_touch of I26916: signal is true;
	signal I26923: std_logic; attribute dont_touch of I26923: signal is true;
	signal I26926: std_logic; attribute dont_touch of I26926: signal is true;
	signal I26931: std_logic; attribute dont_touch of I26931: signal is true;
	signal I26934: std_logic; attribute dont_touch of I26934: signal is true;
	signal I26940: std_logic; attribute dont_touch of I26940: signal is true;
	signal I26947: std_logic; attribute dont_touch of I26947: signal is true;
	signal I26960: std_logic; attribute dont_touch of I26960: signal is true;
	signal I26966: std_logic; attribute dont_touch of I26966: signal is true;
	signal I26972: std_logic; attribute dont_touch of I26972: signal is true;
	signal I26980: std_logic; attribute dont_touch of I26980: signal is true;
	signal I26985: std_logic; attribute dont_touch of I26985: signal is true;
	signal I26990: std_logic; attribute dont_touch of I26990: signal is true;
	signal I26993: std_logic; attribute dont_touch of I26993: signal is true;
	signal I26996: std_logic; attribute dont_touch of I26996: signal is true;
	signal I26999: std_logic; attribute dont_touch of I26999: signal is true;
	signal I27002: std_logic; attribute dont_touch of I27002: signal is true;
	signal I27005: std_logic; attribute dont_touch of I27005: signal is true;
	signal I27008: std_logic; attribute dont_touch of I27008: signal is true;
	signal I27011: std_logic; attribute dont_touch of I27011: signal is true;
	signal I27014: std_logic; attribute dont_touch of I27014: signal is true;
	signal I27017: std_logic; attribute dont_touch of I27017: signal is true;
	signal I27020: std_logic; attribute dont_touch of I27020: signal is true;
	signal I27023: std_logic; attribute dont_touch of I27023: signal is true;
	signal I27026: std_logic; attribute dont_touch of I27026: signal is true;
	signal I27029: std_logic; attribute dont_touch of I27029: signal is true;
	signal I27032: std_logic; attribute dont_touch of I27032: signal is true;
	signal I27035: std_logic; attribute dont_touch of I27035: signal is true;
	signal I27038: std_logic; attribute dont_touch of I27038: signal is true;
	signal I27041: std_logic; attribute dont_touch of I27041: signal is true;
	signal I27044: std_logic; attribute dont_touch of I27044: signal is true;
	signal I27047: std_logic; attribute dont_touch of I27047: signal is true;
	signal I27050: std_logic; attribute dont_touch of I27050: signal is true;
	signal I27053: std_logic; attribute dont_touch of I27053: signal is true;
	signal I27056: std_logic; attribute dont_touch of I27056: signal is true;
	signal I27059: std_logic; attribute dont_touch of I27059: signal is true;
	signal I27062: std_logic; attribute dont_touch of I27062: signal is true;
	signal I27065: std_logic; attribute dont_touch of I27065: signal is true;
	signal I27068: std_logic; attribute dont_touch of I27068: signal is true;
	signal I27071: std_logic; attribute dont_touch of I27071: signal is true;
	signal I27074: std_logic; attribute dont_touch of I27074: signal is true;
	signal I27077: std_logic; attribute dont_touch of I27077: signal is true;
	signal I27080: std_logic; attribute dont_touch of I27080: signal is true;
	signal I27083: std_logic; attribute dont_touch of I27083: signal is true;
	signal I27086: std_logic; attribute dont_touch of I27086: signal is true;
	signal I27089: std_logic; attribute dont_touch of I27089: signal is true;
	signal I27092: std_logic; attribute dont_touch of I27092: signal is true;
	signal I27095: std_logic; attribute dont_touch of I27095: signal is true;
	signal I27098: std_logic; attribute dont_touch of I27098: signal is true;
	signal I27101: std_logic; attribute dont_touch of I27101: signal is true;
	signal I27104: std_logic; attribute dont_touch of I27104: signal is true;
	signal I27107: std_logic; attribute dont_touch of I27107: signal is true;
	signal I27110: std_logic; attribute dont_touch of I27110: signal is true;
	signal I27113: std_logic; attribute dont_touch of I27113: signal is true;
	signal I27116: std_logic; attribute dont_touch of I27116: signal is true;
	signal I27119: std_logic; attribute dont_touch of I27119: signal is true;
	signal I27122: std_logic; attribute dont_touch of I27122: signal is true;
	signal I27125: std_logic; attribute dont_touch of I27125: signal is true;
	signal I27128: std_logic; attribute dont_touch of I27128: signal is true;
	signal I27131: std_logic; attribute dont_touch of I27131: signal is true;
	signal I27134: std_logic; attribute dont_touch of I27134: signal is true;
	signal I27137: std_logic; attribute dont_touch of I27137: signal is true;
	signal I27140: std_logic; attribute dont_touch of I27140: signal is true;
	signal I27143: std_logic; attribute dont_touch of I27143: signal is true;
	signal I27146: std_logic; attribute dont_touch of I27146: signal is true;
	signal I27149: std_logic; attribute dont_touch of I27149: signal is true;
	signal I27152: std_logic; attribute dont_touch of I27152: signal is true;
	signal I27155: std_logic; attribute dont_touch of I27155: signal is true;
	signal I27158: std_logic; attribute dont_touch of I27158: signal is true;
	signal I27161: std_logic; attribute dont_touch of I27161: signal is true;
	signal I27164: std_logic; attribute dont_touch of I27164: signal is true;
	signal I27167: std_logic; attribute dont_touch of I27167: signal is true;
	signal I27170: std_logic; attribute dont_touch of I27170: signal is true;
	signal I27173: std_logic; attribute dont_touch of I27173: signal is true;
	signal I27176: std_logic; attribute dont_touch of I27176: signal is true;
	signal I27179: std_logic; attribute dont_touch of I27179: signal is true;
	signal I27182: std_logic; attribute dont_touch of I27182: signal is true;
	signal I27185: std_logic; attribute dont_touch of I27185: signal is true;
	signal I27188: std_logic; attribute dont_touch of I27188: signal is true;
	signal I27191: std_logic; attribute dont_touch of I27191: signal is true;
	signal I27194: std_logic; attribute dont_touch of I27194: signal is true;
	signal I27197: std_logic; attribute dont_touch of I27197: signal is true;
	signal I27200: std_logic; attribute dont_touch of I27200: signal is true;
	signal I27203: std_logic; attribute dont_touch of I27203: signal is true;
	signal I27206: std_logic; attribute dont_touch of I27206: signal is true;
	signal I27209: std_logic; attribute dont_touch of I27209: signal is true;
	signal I27212: std_logic; attribute dont_touch of I27212: signal is true;
	signal I27215: std_logic; attribute dont_touch of I27215: signal is true;
	signal I27218: std_logic; attribute dont_touch of I27218: signal is true;
	signal I27221: std_logic; attribute dont_touch of I27221: signal is true;
	signal I27225: std_logic; attribute dont_touch of I27225: signal is true;
	signal I27228: std_logic; attribute dont_touch of I27228: signal is true;
	signal I27232: std_logic; attribute dont_touch of I27232: signal is true;
	signal I27235: std_logic; attribute dont_touch of I27235: signal is true;
	signal I27240: std_logic; attribute dont_touch of I27240: signal is true;
	signal I27243: std_logic; attribute dont_touch of I27243: signal is true;
	signal I27246: std_logic; attribute dont_touch of I27246: signal is true;
	signal I27250: std_logic; attribute dont_touch of I27250: signal is true;
	signal I27253: std_logic; attribute dont_touch of I27253: signal is true;
	signal I27257: std_logic; attribute dont_touch of I27257: signal is true;
	signal I27260: std_logic; attribute dont_touch of I27260: signal is true;
	signal I27264: std_logic; attribute dont_touch of I27264: signal is true;
	signal I27267: std_logic; attribute dont_touch of I27267: signal is true;
	signal I27270: std_logic; attribute dont_touch of I27270: signal is true;
	signal I27275: std_logic; attribute dont_touch of I27275: signal is true;
	signal I27278: std_logic; attribute dont_touch of I27278: signal is true;
	signal I27281: std_logic; attribute dont_touch of I27281: signal is true;
	signal I27285: std_logic; attribute dont_touch of I27285: signal is true;
	signal I27288: std_logic; attribute dont_touch of I27288: signal is true;
	signal I27293: std_logic; attribute dont_touch of I27293: signal is true;
	signal I27297: std_logic; attribute dont_touch of I27297: signal is true;
	signal I27300: std_logic; attribute dont_touch of I27300: signal is true;
	signal I27303: std_logic; attribute dont_touch of I27303: signal is true;
	signal I27308: std_logic; attribute dont_touch of I27308: signal is true;
	signal I27311: std_logic; attribute dont_touch of I27311: signal is true;
	signal I27314: std_logic; attribute dont_touch of I27314: signal is true;
	signal I27318: std_logic; attribute dont_touch of I27318: signal is true;
	signal I27321: std_logic; attribute dont_touch of I27321: signal is true;
	signal I27324: std_logic; attribute dont_touch of I27324: signal is true;
	signal I27328: std_logic; attribute dont_touch of I27328: signal is true;
	signal I27332: std_logic; attribute dont_touch of I27332: signal is true;
	signal I27335: std_logic; attribute dont_touch of I27335: signal is true;
	signal I27338: std_logic; attribute dont_touch of I27338: signal is true;
	signal I27343: std_logic; attribute dont_touch of I27343: signal is true;
	signal I27346: std_logic; attribute dont_touch of I27346: signal is true;
	signal I27349: std_logic; attribute dont_touch of I27349: signal is true;
	signal I27352: std_logic; attribute dont_touch of I27352: signal is true;
	signal I27355: std_logic; attribute dont_touch of I27355: signal is true;
	signal I27358: std_logic; attribute dont_touch of I27358: signal is true;
	signal I27361: std_logic; attribute dont_touch of I27361: signal is true;
	signal I27365: std_logic; attribute dont_touch of I27365: signal is true;
	signal I27369: std_logic; attribute dont_touch of I27369: signal is true;
	signal I27372: std_logic; attribute dont_touch of I27372: signal is true;
	signal I27375: std_logic; attribute dont_touch of I27375: signal is true;
	signal I27379: std_logic; attribute dont_touch of I27379: signal is true;
	signal I27382: std_logic; attribute dont_touch of I27382: signal is true;
	signal I27385: std_logic; attribute dont_touch of I27385: signal is true;
	signal I27388: std_logic; attribute dont_touch of I27388: signal is true;
	signal I27391: std_logic; attribute dont_touch of I27391: signal is true;
	signal I27395: std_logic; attribute dont_touch of I27395: signal is true;
	signal I27399: std_logic; attribute dont_touch of I27399: signal is true;
	signal I27402: std_logic; attribute dont_touch of I27402: signal is true;
	signal I27405: std_logic; attribute dont_touch of I27405: signal is true;
	signal I27408: std_logic; attribute dont_touch of I27408: signal is true;
	signal I27411: std_logic; attribute dont_touch of I27411: signal is true;
	signal I27416: std_logic; attribute dont_touch of I27416: signal is true;
	signal I27419: std_logic; attribute dont_touch of I27419: signal is true;
	signal I27422: std_logic; attribute dont_touch of I27422: signal is true;
	signal I27426: std_logic; attribute dont_touch of I27426: signal is true;
	signal I27488: std_logic; attribute dont_touch of I27488: signal is true;
	signal I27491: std_logic; attribute dont_touch of I27491: signal is true;
	signal I27516: std_logic; attribute dont_touch of I27516: signal is true;
	signal I27531: std_logic; attribute dont_touch of I27531: signal is true;
	signal I27534: std_logic; attribute dont_touch of I27534: signal is true;
	signal I27537: std_logic; attribute dont_touch of I27537: signal is true;
	signal I27549: std_logic; attribute dont_touch of I27549: signal is true;
	signal I27565: std_logic; attribute dont_touch of I27565: signal is true;
	signal I27577: std_logic; attribute dont_touch of I27577: signal is true;
	signal I27585: std_logic; attribute dont_touch of I27585: signal is true;
	signal I27593: std_logic; attribute dont_touch of I27593: signal is true;
	signal I27614: std_logic; attribute dont_touch of I27614: signal is true;
	signal I27621: std_logic; attribute dont_touch of I27621: signal is true;
	signal I27646: std_logic; attribute dont_touch of I27646: signal is true;
	signal I27658: std_logic; attribute dont_touch of I27658: signal is true;
	signal I27667: std_logic; attribute dont_touch of I27667: signal is true;
	signal I27672: std_logic; attribute dont_touch of I27672: signal is true;
	signal I27684: std_logic; attribute dont_touch of I27684: signal is true;
	signal I27689: std_logic; attribute dont_touch of I27689: signal is true;
	signal I27695: std_logic; attribute dont_touch of I27695: signal is true;
	signal I27705: std_logic; attribute dont_touch of I27705: signal is true;
	signal I27711: std_logic; attribute dont_touch of I27711: signal is true;
	signal I27717: std_logic; attribute dont_touch of I27717: signal is true;
	signal I27727: std_logic; attribute dont_touch of I27727: signal is true;
	signal I27733: std_logic; attribute dont_touch of I27733: signal is true;
	signal I27739: std_logic; attribute dont_touch of I27739: signal is true;
	signal I27749: std_logic; attribute dont_touch of I27749: signal is true;
	signal I27755: std_logic; attribute dont_touch of I27755: signal is true;
	signal I27761: std_logic; attribute dont_touch of I27761: signal is true;
	signal I27766: std_logic; attribute dont_touch of I27766: signal is true;
	signal I27772: std_logic; attribute dont_touch of I27772: signal is true;
	signal I27779: std_logic; attribute dont_touch of I27779: signal is true;
	signal I27785: std_logic; attribute dont_touch of I27785: signal is true;
	signal I27822: std_logic; attribute dont_touch of I27822: signal is true;
	signal I27827: std_logic; attribute dont_touch of I27827: signal is true;
	signal I27832: std_logic; attribute dont_touch of I27832: signal is true;
	signal I27838: std_logic; attribute dont_touch of I27838: signal is true;
	signal I27868: std_logic; attribute dont_touch of I27868: signal is true;
	signal I27897: std_logic; attribute dont_touch of I27897: signal is true;
	signal I27900: std_logic; attribute dont_touch of I27900: signal is true;
	signal I27917: std_logic; attribute dont_touch of I27917: signal is true;
	signal I27920: std_logic; attribute dont_touch of I27920: signal is true;
	signal I27927: std_logic; attribute dont_touch of I27927: signal is true;
	signal I27942: std_logic; attribute dont_touch of I27942: signal is true;
	signal I27949: std_logic; attribute dont_touch of I27949: signal is true;
	signal I27958: std_logic; attribute dont_touch of I27958: signal is true;
	signal I27969: std_logic; attribute dont_touch of I27969: signal is true;
	signal I27972: std_logic; attribute dont_touch of I27972: signal is true;
	signal I27976: std_logic; attribute dont_touch of I27976: signal is true;
	signal I27984: std_logic; attribute dont_touch of I27984: signal is true;
	signal I27992: std_logic; attribute dont_touch of I27992: signal is true;
	signal I28000: std_logic; attribute dont_touch of I28000: signal is true;
	signal I28003: std_logic; attribute dont_touch of I28003: signal is true;
	signal I28009: std_logic; attribute dont_touch of I28009: signal is true;
	signal I28013: std_logic; attribute dont_touch of I28013: signal is true;
	signal I28019: std_logic; attribute dont_touch of I28019: signal is true;
	signal I28027: std_logic; attribute dont_touch of I28027: signal is true;
	signal I28031: std_logic; attribute dont_touch of I28031: signal is true;
	signal I28034: std_logic; attribute dont_touch of I28034: signal is true;
	signal I28038: std_logic; attribute dont_touch of I28038: signal is true;
	signal I28043: std_logic; attribute dont_touch of I28043: signal is true;
	signal I28047: std_logic; attribute dont_touch of I28047: signal is true;
	signal I28051: std_logic; attribute dont_touch of I28051: signal is true;
	signal I28057: std_logic; attribute dont_touch of I28057: signal is true;
	signal I28061: std_logic; attribute dont_touch of I28061: signal is true;
	signal I28065: std_logic; attribute dont_touch of I28065: signal is true;
	signal I28068: std_logic; attribute dont_touch of I28068: signal is true;
	signal I28072: std_logic; attribute dont_touch of I28072: signal is true;
	signal I28076: std_logic; attribute dont_touch of I28076: signal is true;
	signal I28080: std_logic; attribute dont_touch of I28080: signal is true;
	signal I28084: std_logic; attribute dont_touch of I28084: signal is true;
	signal I28087: std_logic; attribute dont_touch of I28087: signal is true;
	signal I28090: std_logic; attribute dont_touch of I28090: signal is true;
	signal I28093: std_logic; attribute dont_touch of I28093: signal is true;
	signal I28096: std_logic; attribute dont_touch of I28096: signal is true;
	signal I28100: std_logic; attribute dont_touch of I28100: signal is true;
	signal I28103: std_logic; attribute dont_touch of I28103: signal is true;
	signal I28107: std_logic; attribute dont_touch of I28107: signal is true;
	signal I28111: std_logic; attribute dont_touch of I28111: signal is true;
	signal I28115: std_logic; attribute dont_touch of I28115: signal is true;
	signal I28119: std_logic; attribute dont_touch of I28119: signal is true;
	signal I28123: std_logic; attribute dont_touch of I28123: signal is true;
	signal I28126: std_logic; attribute dont_touch of I28126: signal is true;
	signal I28130: std_logic; attribute dont_touch of I28130: signal is true;
	signal I28133: std_logic; attribute dont_touch of I28133: signal is true;
	signal I28137: std_logic; attribute dont_touch of I28137: signal is true;
	signal I28143: std_logic; attribute dont_touch of I28143: signal is true;
	signal I28148: std_logic; attribute dont_touch of I28148: signal is true;
	signal I28152: std_logic; attribute dont_touch of I28152: signal is true;
	signal I28155: std_logic; attribute dont_touch of I28155: signal is true;
	signal I28159: std_logic; attribute dont_touch of I28159: signal is true;
	signal I28162: std_logic; attribute dont_touch of I28162: signal is true;
	signal I28169: std_logic; attribute dont_touch of I28169: signal is true;
	signal I28174: std_logic; attribute dont_touch of I28174: signal is true;
	signal I28178: std_logic; attribute dont_touch of I28178: signal is true;
	signal I28181: std_logic; attribute dont_touch of I28181: signal is true;
	signal I28184: std_logic; attribute dont_touch of I28184: signal is true;
	signal I28189: std_logic; attribute dont_touch of I28189: signal is true;
	signal I28190: std_logic; attribute dont_touch of I28190: signal is true;
	signal I28191: std_logic; attribute dont_touch of I28191: signal is true;
	signal I28201: std_logic; attribute dont_touch of I28201: signal is true;
	signal I28206: std_logic; attribute dont_touch of I28206: signal is true;
	signal I28210: std_logic; attribute dont_touch of I28210: signal is true;
	signal I28217: std_logic; attribute dont_touch of I28217: signal is true;
	signal I28218: std_logic; attribute dont_touch of I28218: signal is true;
	signal I28219: std_logic; attribute dont_touch of I28219: signal is true;
	signal I28229: std_logic; attribute dont_touch of I28229: signal is true;
	signal I28235: std_logic; attribute dont_touch of I28235: signal is true;
	signal I28247: std_logic; attribute dont_touch of I28247: signal is true;
	signal I28248: std_logic; attribute dont_touch of I28248: signal is true;
	signal I28249: std_logic; attribute dont_touch of I28249: signal is true;
	signal I28271: std_logic; attribute dont_touch of I28271: signal is true;
	signal I28272: std_logic; attribute dont_touch of I28272: signal is true;
	signal I28273: std_logic; attribute dont_touch of I28273: signal is true;
	signal I28305: std_logic; attribute dont_touch of I28305: signal is true;
	signal I28314: std_logic; attribute dont_touch of I28314: signal is true;
	signal I28318: std_logic; attribute dont_touch of I28318: signal is true;
	signal I28323: std_logic; attribute dont_touch of I28323: signal is true;
	signal I28330: std_logic; attribute dont_touch of I28330: signal is true;
	signal I28335: std_logic; attribute dont_touch of I28335: signal is true;
	signal I28341: std_logic; attribute dont_touch of I28341: signal is true;
	signal I28346: std_logic; attribute dont_touch of I28346: signal is true;
	signal I28351: std_logic; attribute dont_touch of I28351: signal is true;
	signal I28357: std_logic; attribute dont_touch of I28357: signal is true;
	signal I28360: std_logic; attribute dont_touch of I28360: signal is true;
	signal I28365: std_logic; attribute dont_touch of I28365: signal is true;
	signal I28369: std_logic; attribute dont_touch of I28369: signal is true;
	signal I28374: std_logic; attribute dont_touch of I28374: signal is true;
	signal I28380: std_logic; attribute dont_touch of I28380: signal is true;
	signal I28432: std_logic; attribute dont_touch of I28432: signal is true;
	signal I28435: std_logic; attribute dont_touch of I28435: signal is true;
	signal I28443: std_logic; attribute dont_touch of I28443: signal is true;
	signal I28447: std_logic; attribute dont_touch of I28447: signal is true;
	signal I28450: std_logic; attribute dont_touch of I28450: signal is true;
	signal I28455: std_logic; attribute dont_touch of I28455: signal is true;
	signal I28458: std_logic; attribute dont_touch of I28458: signal is true;
	signal I28461: std_logic; attribute dont_touch of I28461: signal is true;
	signal I28464: std_logic; attribute dont_touch of I28464: signal is true;
	signal I28467: std_logic; attribute dont_touch of I28467: signal is true;
	signal I28470: std_logic; attribute dont_touch of I28470: signal is true;
	signal I28473: std_logic; attribute dont_touch of I28473: signal is true;
	signal I28476: std_logic; attribute dont_touch of I28476: signal is true;
	signal I28479: std_logic; attribute dont_touch of I28479: signal is true;
	signal I28482: std_logic; attribute dont_touch of I28482: signal is true;
	signal I28485: std_logic; attribute dont_touch of I28485: signal is true;
	signal I28488: std_logic; attribute dont_touch of I28488: signal is true;
	signal I28491: std_logic; attribute dont_touch of I28491: signal is true;
	signal I28494: std_logic; attribute dont_touch of I28494: signal is true;
	signal I28497: std_logic; attribute dont_touch of I28497: signal is true;
	signal I28500: std_logic; attribute dont_touch of I28500: signal is true;
	signal I28503: std_logic; attribute dont_touch of I28503: signal is true;
	signal I28506: std_logic; attribute dont_touch of I28506: signal is true;
	signal I28509: std_logic; attribute dont_touch of I28509: signal is true;
	signal I28512: std_logic; attribute dont_touch of I28512: signal is true;
	signal I28515: std_logic; attribute dont_touch of I28515: signal is true;
	signal I28518: std_logic; attribute dont_touch of I28518: signal is true;
	signal I28521: std_logic; attribute dont_touch of I28521: signal is true;
	signal I28524: std_logic; attribute dont_touch of I28524: signal is true;
	signal I28527: std_logic; attribute dont_touch of I28527: signal is true;
	signal I28541: std_logic; attribute dont_touch of I28541: signal is true;
	signal I28550: std_logic; attribute dont_touch of I28550: signal is true;
	signal I28557: std_logic; attribute dont_touch of I28557: signal is true;
	signal I28564: std_logic; attribute dont_touch of I28564: signal is true;
	signal I28582: std_logic; attribute dont_touch of I28582: signal is true;
	signal I28594: std_logic; attribute dont_touch of I28594: signal is true;
	signal I28609: std_logic; attribute dont_touch of I28609: signal is true;
	signal I28628: std_logic; attribute dont_touch of I28628: signal is true;
	signal I28649: std_logic; attribute dont_touch of I28649: signal is true;
	signal I28671: std_logic; attribute dont_touch of I28671: signal is true;
	signal I28693: std_logic; attribute dont_touch of I28693: signal is true;
	signal I28712: std_logic; attribute dont_touch of I28712: signal is true;
	signal I28726: std_logic; attribute dont_touch of I28726: signal is true;
	signal I28727: std_logic; attribute dont_touch of I28727: signal is true;
	signal I28728: std_logic; attribute dont_touch of I28728: signal is true;
	signal I28741: std_logic; attribute dont_touch of I28741: signal is true;
	signal I28742: std_logic; attribute dont_touch of I28742: signal is true;
	signal I28743: std_logic; attribute dont_touch of I28743: signal is true;
	signal I28753: std_logic; attribute dont_touch of I28753: signal is true;
	signal I28754: std_logic; attribute dont_touch of I28754: signal is true;
	signal I28755: std_logic; attribute dont_touch of I28755: signal is true;
	signal I28765: std_logic; attribute dont_touch of I28765: signal is true;
	signal I28766: std_logic; attribute dont_touch of I28766: signal is true;
	signal I28767: std_logic; attribute dont_touch of I28767: signal is true;
	signal I28781: std_logic; attribute dont_touch of I28781: signal is true;
	signal I28789: std_logic; attribute dont_touch of I28789: signal is true;
	signal I28792: std_logic; attribute dont_touch of I28792: signal is true;
	signal I28800: std_logic; attribute dont_touch of I28800: signal is true;
	signal I28813: std_logic; attribute dont_touch of I28813: signal is true;
	signal I28825: std_logic; attribute dont_touch of I28825: signal is true;
	signal I28833: std_logic; attribute dont_touch of I28833: signal is true;
	signal I28876: std_logic; attribute dont_touch of I28876: signal is true;
	signal I28896: std_logic; attribute dont_touch of I28896: signal is true;
	signal I28913: std_logic; attribute dont_touch of I28913: signal is true;
	signal I28928: std_logic; attribute dont_touch of I28928: signal is true;
	signal I28949: std_logic; attribute dont_touch of I28949: signal is true;
	signal I28953: std_logic; attribute dont_touch of I28953: signal is true;
	signal I28956: std_logic; attribute dont_touch of I28956: signal is true;
	signal I28959: std_logic; attribute dont_touch of I28959: signal is true;
	signal I28962: std_logic; attribute dont_touch of I28962: signal is true;
	signal I28966: std_logic; attribute dont_touch of I28966: signal is true;
	signal I28969: std_logic; attribute dont_touch of I28969: signal is true;
	signal I28972: std_logic; attribute dont_touch of I28972: signal is true;
	signal I28975: std_logic; attribute dont_touch of I28975: signal is true;
	signal I28978: std_logic; attribute dont_touch of I28978: signal is true;
	signal I28981: std_logic; attribute dont_touch of I28981: signal is true;
	signal I28984: std_logic; attribute dont_touch of I28984: signal is true;
	signal I28988: std_logic; attribute dont_touch of I28988: signal is true;
	signal I28991: std_logic; attribute dont_touch of I28991: signal is true;
	signal I28994: std_logic; attribute dont_touch of I28994: signal is true;
	signal I28997: std_logic; attribute dont_touch of I28997: signal is true;
	signal I29001: std_logic; attribute dont_touch of I29001: signal is true;
	signal I29004: std_logic; attribute dont_touch of I29004: signal is true;
	signal I29007: std_logic; attribute dont_touch of I29007: signal is true;
	signal I29010: std_logic; attribute dont_touch of I29010: signal is true;
	signal I29013: std_logic; attribute dont_touch of I29013: signal is true;
	signal I29016: std_logic; attribute dont_touch of I29016: signal is true;
	signal I29019: std_logic; attribute dont_touch of I29019: signal is true;
	signal I29023: std_logic; attribute dont_touch of I29023: signal is true;
	signal I29026: std_logic; attribute dont_touch of I29026: signal is true;
	signal I29030: std_logic; attribute dont_touch of I29030: signal is true;
	signal I29033: std_logic; attribute dont_touch of I29033: signal is true;
	signal I29036: std_logic; attribute dont_touch of I29036: signal is true;
	signal I29040: std_logic; attribute dont_touch of I29040: signal is true;
	signal I29043: std_logic; attribute dont_touch of I29043: signal is true;
	signal I29046: std_logic; attribute dont_touch of I29046: signal is true;
	signal I29049: std_logic; attribute dont_touch of I29049: signal is true;
	signal I29052: std_logic; attribute dont_touch of I29052: signal is true;
	signal I29055: std_logic; attribute dont_touch of I29055: signal is true;
	signal I29058: std_logic; attribute dont_touch of I29058: signal is true;
	signal I29064: std_logic; attribute dont_touch of I29064: signal is true;
	signal I29067: std_logic; attribute dont_touch of I29067: signal is true;
	signal I29070: std_logic; attribute dont_touch of I29070: signal is true;
	signal I29073: std_logic; attribute dont_touch of I29073: signal is true;
	signal I29077: std_logic; attribute dont_touch of I29077: signal is true;
	signal I29080: std_logic; attribute dont_touch of I29080: signal is true;
	signal I29083: std_logic; attribute dont_touch of I29083: signal is true;
	signal I29087: std_logic; attribute dont_touch of I29087: signal is true;
	signal I29090: std_logic; attribute dont_touch of I29090: signal is true;
	signal I29093: std_logic; attribute dont_touch of I29093: signal is true;
	signal I29098: std_logic; attribute dont_touch of I29098: signal is true;
	signal I29101: std_logic; attribute dont_touch of I29101: signal is true;
	signal I29104: std_logic; attribute dont_touch of I29104: signal is true;
	signal I29107: std_logic; attribute dont_touch of I29107: signal is true;
	signal I29110: std_logic; attribute dont_touch of I29110: signal is true;
	signal I29116: std_logic; attribute dont_touch of I29116: signal is true;
	signal I29119: std_logic; attribute dont_touch of I29119: signal is true;
	signal I29122: std_logic; attribute dont_touch of I29122: signal is true;
	signal I29125: std_logic; attribute dont_touch of I29125: signal is true;
	signal I29129: std_logic; attribute dont_touch of I29129: signal is true;
	signal I29132: std_logic; attribute dont_touch of I29132: signal is true;
	signal I29135: std_logic; attribute dont_touch of I29135: signal is true;
	signal I29142: std_logic; attribute dont_touch of I29142: signal is true;
	signal I29145: std_logic; attribute dont_touch of I29145: signal is true;
	signal I29148: std_logic; attribute dont_touch of I29148: signal is true;
	signal I29151: std_logic; attribute dont_touch of I29151: signal is true;
	signal I29154: std_logic; attribute dont_touch of I29154: signal is true;
	signal I29159: std_logic; attribute dont_touch of I29159: signal is true;
	signal I29162: std_logic; attribute dont_touch of I29162: signal is true;
	signal I29165: std_logic; attribute dont_touch of I29165: signal is true;
	signal I29168: std_logic; attribute dont_touch of I29168: signal is true;
	signal I29174: std_logic; attribute dont_touch of I29174: signal is true;
	signal I29177: std_logic; attribute dont_touch of I29177: signal is true;
	signal I29180: std_logic; attribute dont_touch of I29180: signal is true;
	signal I29183: std_logic; attribute dont_touch of I29183: signal is true;
	signal I29191: std_logic; attribute dont_touch of I29191: signal is true;
	signal I29194: std_logic; attribute dont_touch of I29194: signal is true;
	signal I29197: std_logic; attribute dont_touch of I29197: signal is true;
	signal I29203: std_logic; attribute dont_touch of I29203: signal is true;
	signal I29206: std_logic; attribute dont_touch of I29206: signal is true;
	signal I29209: std_logic; attribute dont_touch of I29209: signal is true;
	signal I29212: std_logic; attribute dont_touch of I29212: signal is true;
	signal I29215: std_logic; attribute dont_touch of I29215: signal is true;
	signal I29220: std_logic; attribute dont_touch of I29220: signal is true;
	signal I29223: std_logic; attribute dont_touch of I29223: signal is true;
	signal I29226: std_logic; attribute dont_touch of I29226: signal is true;
	signal I29229: std_logic; attribute dont_touch of I29229: signal is true;
	signal I29235: std_logic; attribute dont_touch of I29235: signal is true;
	signal I29238: std_logic; attribute dont_touch of I29238: signal is true;
	signal I29243: std_logic; attribute dont_touch of I29243: signal is true;
	signal I29246: std_logic; attribute dont_touch of I29246: signal is true;
	signal I29249: std_logic; attribute dont_touch of I29249: signal is true;
	signal I29252: std_logic; attribute dont_touch of I29252: signal is true;
	signal I29259: std_logic; attribute dont_touch of I29259: signal is true;
	signal I29262: std_logic; attribute dont_touch of I29262: signal is true;
	signal I29265: std_logic; attribute dont_touch of I29265: signal is true;
	signal I29271: std_logic; attribute dont_touch of I29271: signal is true;
	signal I29274: std_logic; attribute dont_touch of I29274: signal is true;
	signal I29277: std_logic; attribute dont_touch of I29277: signal is true;
	signal I29280: std_logic; attribute dont_touch of I29280: signal is true;
	signal I29283: std_logic; attribute dont_touch of I29283: signal is true;
	signal I29288: std_logic; attribute dont_touch of I29288: signal is true;
	signal I29291: std_logic; attribute dont_touch of I29291: signal is true;
	signal I29294: std_logic; attribute dont_touch of I29294: signal is true;
	signal I29301: std_logic; attribute dont_touch of I29301: signal is true;
	signal I29304: std_logic; attribute dont_touch of I29304: signal is true;
	signal I29307: std_logic; attribute dont_touch of I29307: signal is true;
	signal I29310: std_logic; attribute dont_touch of I29310: signal is true;
	signal I29313: std_logic; attribute dont_touch of I29313: signal is true;
	signal I29317: std_logic; attribute dont_touch of I29317: signal is true;
	signal I29320: std_logic; attribute dont_touch of I29320: signal is true;
	signal I29323: std_logic; attribute dont_touch of I29323: signal is true;
	signal I29326: std_logic; attribute dont_touch of I29326: signal is true;
	signal I29333: std_logic; attribute dont_touch of I29333: signal is true;
	signal I29336: std_logic; attribute dont_touch of I29336: signal is true;
	signal I29339: std_logic; attribute dont_touch of I29339: signal is true;
	signal I29345: std_logic; attribute dont_touch of I29345: signal is true;
	signal I29348: std_logic; attribute dont_touch of I29348: signal is true;
	signal I29351: std_logic; attribute dont_touch of I29351: signal is true;
	signal I29354: std_logic; attribute dont_touch of I29354: signal is true;
	signal I29357: std_logic; attribute dont_touch of I29357: signal is true;
	signal I29360: std_logic; attribute dont_touch of I29360: signal is true;
	signal I29366: std_logic; attribute dont_touch of I29366: signal is true;
	signal I29369: std_logic; attribute dont_touch of I29369: signal is true;
	signal I29372: std_logic; attribute dont_touch of I29372: signal is true;
	signal I29375: std_logic; attribute dont_touch of I29375: signal is true;
	signal I29378: std_logic; attribute dont_touch of I29378: signal is true;
	signal I29383: std_logic; attribute dont_touch of I29383: signal is true;
	signal I29386: std_logic; attribute dont_touch of I29386: signal is true;
	signal I29389: std_logic; attribute dont_touch of I29389: signal is true;
	signal I29392: std_logic; attribute dont_touch of I29392: signal is true;
	signal I29395: std_logic; attribute dont_touch of I29395: signal is true;
	signal I29399: std_logic; attribute dont_touch of I29399: signal is true;
	signal I29402: std_logic; attribute dont_touch of I29402: signal is true;
	signal I29405: std_logic; attribute dont_touch of I29405: signal is true;
	signal I29408: std_logic; attribute dont_touch of I29408: signal is true;
	signal I29415: std_logic; attribute dont_touch of I29415: signal is true;
	signal I29418: std_logic; attribute dont_touch of I29418: signal is true;
	signal I29421: std_logic; attribute dont_touch of I29421: signal is true;
	signal I29426: std_logic; attribute dont_touch of I29426: signal is true;
	signal I29429: std_logic; attribute dont_touch of I29429: signal is true;
	signal I29432: std_logic; attribute dont_touch of I29432: signal is true;
	signal I29435: std_logic; attribute dont_touch of I29435: signal is true;
	signal I29439: std_logic; attribute dont_touch of I29439: signal is true;
	signal I29442: std_logic; attribute dont_touch of I29442: signal is true;
	signal I29445: std_logic; attribute dont_touch of I29445: signal is true;
	signal I29448: std_logic; attribute dont_touch of I29448: signal is true;
	signal I29451: std_logic; attribute dont_touch of I29451: signal is true;
	signal I29456: std_logic; attribute dont_touch of I29456: signal is true;
	signal I29459: std_logic; attribute dont_touch of I29459: signal is true;
	signal I29462: std_logic; attribute dont_touch of I29462: signal is true;
	signal I29465: std_logic; attribute dont_touch of I29465: signal is true;
	signal I29468: std_logic; attribute dont_touch of I29468: signal is true;
	signal I29472: std_logic; attribute dont_touch of I29472: signal is true;
	signal I29475: std_logic; attribute dont_touch of I29475: signal is true;
	signal I29478: std_logic; attribute dont_touch of I29478: signal is true;
	signal I29481: std_logic; attribute dont_touch of I29481: signal is true;
	signal I29484: std_logic; attribute dont_touch of I29484: signal is true;
	signal I29490: std_logic; attribute dont_touch of I29490: signal is true;
	signal I29493: std_logic; attribute dont_touch of I29493: signal is true;
	signal I29496: std_logic; attribute dont_touch of I29496: signal is true;
	signal I29500: std_logic; attribute dont_touch of I29500: signal is true;
	signal I29503: std_logic; attribute dont_touch of I29503: signal is true;
	signal I29506: std_logic; attribute dont_touch of I29506: signal is true;
	signal I29509: std_logic; attribute dont_touch of I29509: signal is true;
	signal I29513: std_logic; attribute dont_touch of I29513: signal is true;
	signal I29516: std_logic; attribute dont_touch of I29516: signal is true;
	signal I29519: std_logic; attribute dont_touch of I29519: signal is true;
	signal I29522: std_logic; attribute dont_touch of I29522: signal is true;
	signal I29525: std_logic; attribute dont_touch of I29525: signal is true;
	signal I29530: std_logic; attribute dont_touch of I29530: signal is true;
	signal I29533: std_logic; attribute dont_touch of I29533: signal is true;
	signal I29536: std_logic; attribute dont_touch of I29536: signal is true;
	signal I29539: std_logic; attribute dont_touch of I29539: signal is true;
	signal I29542: std_logic; attribute dont_touch of I29542: signal is true;
	signal I29547: std_logic; attribute dont_touch of I29547: signal is true;
	signal I29550: std_logic; attribute dont_touch of I29550: signal is true;
	signal I29556: std_logic; attribute dont_touch of I29556: signal is true;
	signal I29559: std_logic; attribute dont_touch of I29559: signal is true;
	signal I29562: std_logic; attribute dont_touch of I29562: signal is true;
	signal I29566: std_logic; attribute dont_touch of I29566: signal is true;
	signal I29569: std_logic; attribute dont_touch of I29569: signal is true;
	signal I29572: std_logic; attribute dont_touch of I29572: signal is true;
	signal I29575: std_logic; attribute dont_touch of I29575: signal is true;
	signal I29579: std_logic; attribute dont_touch of I29579: signal is true;
	signal I29582: std_logic; attribute dont_touch of I29582: signal is true;
	signal I29585: std_logic; attribute dont_touch of I29585: signal is true;
	signal I29588: std_logic; attribute dont_touch of I29588: signal is true;
	signal I29591: std_logic; attribute dont_touch of I29591: signal is true;
	signal I29600: std_logic; attribute dont_touch of I29600: signal is true;
	signal I29603: std_logic; attribute dont_touch of I29603: signal is true;
	signal I29606: std_logic; attribute dont_touch of I29606: signal is true;
	signal I29610: std_logic; attribute dont_touch of I29610: signal is true;
	signal I29613: std_logic; attribute dont_touch of I29613: signal is true;
	signal I29619: std_logic; attribute dont_touch of I29619: signal is true;
	signal I29622: std_logic; attribute dont_touch of I29622: signal is true;
	signal I29625: std_logic; attribute dont_touch of I29625: signal is true;
	signal I29629: std_logic; attribute dont_touch of I29629: signal is true;
	signal I29632: std_logic; attribute dont_touch of I29632: signal is true;
	signal I29635: std_logic; attribute dont_touch of I29635: signal is true;
	signal I29638: std_logic; attribute dont_touch of I29638: signal is true;
	signal I29641: std_logic; attribute dont_touch of I29641: signal is true;
	signal I29653: std_logic; attribute dont_touch of I29653: signal is true;
	signal I29656: std_logic; attribute dont_touch of I29656: signal is true;
	signal I29660: std_logic; attribute dont_touch of I29660: signal is true;
	signal I29663: std_logic; attribute dont_touch of I29663: signal is true;
	signal I29669: std_logic; attribute dont_touch of I29669: signal is true;
	signal I29672: std_logic; attribute dont_touch of I29672: signal is true;
	signal I29675: std_logic; attribute dont_touch of I29675: signal is true;
	signal I29687: std_logic; attribute dont_touch of I29687: signal is true;
	signal I29690: std_logic; attribute dont_touch of I29690: signal is true;
	signal I29694: std_logic; attribute dont_touch of I29694: signal is true;
	signal I29697: std_logic; attribute dont_touch of I29697: signal is true;
	signal I29700: std_logic; attribute dont_touch of I29700: signal is true;
	signal I29712: std_logic; attribute dont_touch of I29712: signal is true;
	signal I29715: std_logic; attribute dont_touch of I29715: signal is true;
	signal I29724: std_logic; attribute dont_touch of I29724: signal is true;
	signal I29727: std_logic; attribute dont_touch of I29727: signal is true;
	signal I29736: std_logic; attribute dont_touch of I29736: signal is true;
	signal I29741: std_logic; attribute dont_touch of I29741: signal is true;
	signal I29797: std_logic; attribute dont_touch of I29797: signal is true;
	signal I29802: std_logic; attribute dont_touch of I29802: signal is true;
	signal I29812: std_logic; attribute dont_touch of I29812: signal is true;
	signal I29817: std_logic; attribute dont_touch of I29817: signal is true;
	signal I29827: std_logic; attribute dont_touch of I29827: signal is true;
	signal I29841: std_logic; attribute dont_touch of I29841: signal is true;
	signal I29852: std_logic; attribute dont_touch of I29852: signal is true;
	signal I29863: std_logic; attribute dont_touch of I29863: signal is true;
	signal I29872: std_logic; attribute dont_touch of I29872: signal is true;
	signal I29881: std_logic; attribute dont_touch of I29881: signal is true;
	signal I29897: std_logic; attribute dont_touch of I29897: signal is true;
	signal I29900: std_logic; attribute dont_touch of I29900: signal is true;
	signal I29903: std_logic; attribute dont_touch of I29903: signal is true;
	signal I29906: std_logic; attribute dont_touch of I29906: signal is true;
	signal I29909: std_logic; attribute dont_touch of I29909: signal is true;
	signal I29912: std_logic; attribute dont_touch of I29912: signal is true;
	signal I29915: std_logic; attribute dont_touch of I29915: signal is true;
	signal I29918: std_logic; attribute dont_touch of I29918: signal is true;
	signal I29921: std_logic; attribute dont_touch of I29921: signal is true;
	signal I29924: std_logic; attribute dont_touch of I29924: signal is true;
	signal I29927: std_logic; attribute dont_touch of I29927: signal is true;
	signal I29930: std_logic; attribute dont_touch of I29930: signal is true;
	signal I29933: std_logic; attribute dont_touch of I29933: signal is true;
	signal I29936: std_logic; attribute dont_touch of I29936: signal is true;
	signal I29939: std_logic; attribute dont_touch of I29939: signal is true;
	signal I29942: std_logic; attribute dont_touch of I29942: signal is true;
	signal I29945: std_logic; attribute dont_touch of I29945: signal is true;
	signal I29948: std_logic; attribute dont_touch of I29948: signal is true;
	signal I29951: std_logic; attribute dont_touch of I29951: signal is true;
	signal I29954: std_logic; attribute dont_touch of I29954: signal is true;
	signal I29957: std_logic; attribute dont_touch of I29957: signal is true;
	signal I29960: std_logic; attribute dont_touch of I29960: signal is true;
	signal I29963: std_logic; attribute dont_touch of I29963: signal is true;
	signal I29966: std_logic; attribute dont_touch of I29966: signal is true;
	signal I29969: std_logic; attribute dont_touch of I29969: signal is true;
	signal I29972: std_logic; attribute dont_touch of I29972: signal is true;
	signal I29975: std_logic; attribute dont_touch of I29975: signal is true;
	signal I29978: std_logic; attribute dont_touch of I29978: signal is true;
	signal I29981: std_logic; attribute dont_touch of I29981: signal is true;
	signal I29984: std_logic; attribute dont_touch of I29984: signal is true;
	signal I29987: std_logic; attribute dont_touch of I29987: signal is true;
	signal I29990: std_logic; attribute dont_touch of I29990: signal is true;
	signal I29993: std_logic; attribute dont_touch of I29993: signal is true;
	signal I29996: std_logic; attribute dont_touch of I29996: signal is true;
	signal I29999: std_logic; attribute dont_touch of I29999: signal is true;
	signal I30002: std_logic; attribute dont_touch of I30002: signal is true;
	signal I30005: std_logic; attribute dont_touch of I30005: signal is true;
	signal I30008: std_logic; attribute dont_touch of I30008: signal is true;
	signal I30011: std_logic; attribute dont_touch of I30011: signal is true;
	signal I30014: std_logic; attribute dont_touch of I30014: signal is true;
	signal I30017: std_logic; attribute dont_touch of I30017: signal is true;
	signal I30020: std_logic; attribute dont_touch of I30020: signal is true;
	signal I30023: std_logic; attribute dont_touch of I30023: signal is true;
	signal I30026: std_logic; attribute dont_touch of I30026: signal is true;
	signal I30029: std_logic; attribute dont_touch of I30029: signal is true;
	signal I30032: std_logic; attribute dont_touch of I30032: signal is true;
	signal I30035: std_logic; attribute dont_touch of I30035: signal is true;
	signal I30038: std_logic; attribute dont_touch of I30038: signal is true;
	signal I30041: std_logic; attribute dont_touch of I30041: signal is true;
	signal I30044: std_logic; attribute dont_touch of I30044: signal is true;
	signal I30047: std_logic; attribute dont_touch of I30047: signal is true;
	signal I30050: std_logic; attribute dont_touch of I30050: signal is true;
	signal I30053: std_logic; attribute dont_touch of I30053: signal is true;
	signal I30056: std_logic; attribute dont_touch of I30056: signal is true;
	signal I30059: std_logic; attribute dont_touch of I30059: signal is true;
	signal I30062: std_logic; attribute dont_touch of I30062: signal is true;
	signal I30065: std_logic; attribute dont_touch of I30065: signal is true;
	signal I30068: std_logic; attribute dont_touch of I30068: signal is true;
	signal I30071: std_logic; attribute dont_touch of I30071: signal is true;
	signal I30074: std_logic; attribute dont_touch of I30074: signal is true;
	signal I30077: std_logic; attribute dont_touch of I30077: signal is true;
	signal I30080: std_logic; attribute dont_touch of I30080: signal is true;
	signal I30083: std_logic; attribute dont_touch of I30083: signal is true;
	signal I30086: std_logic; attribute dont_touch of I30086: signal is true;
	signal I30089: std_logic; attribute dont_touch of I30089: signal is true;
	signal I30092: std_logic; attribute dont_touch of I30092: signal is true;
	signal I30095: std_logic; attribute dont_touch of I30095: signal is true;
	signal I30098: std_logic; attribute dont_touch of I30098: signal is true;
	signal I30101: std_logic; attribute dont_touch of I30101: signal is true;
	signal I30104: std_logic; attribute dont_touch of I30104: signal is true;
	signal I30107: std_logic; attribute dont_touch of I30107: signal is true;
	signal I30110: std_logic; attribute dont_touch of I30110: signal is true;
	signal I30113: std_logic; attribute dont_touch of I30113: signal is true;
	signal I30116: std_logic; attribute dont_touch of I30116: signal is true;
	signal I30119: std_logic; attribute dont_touch of I30119: signal is true;
	signal I30122: std_logic; attribute dont_touch of I30122: signal is true;
	signal I30125: std_logic; attribute dont_touch of I30125: signal is true;
	signal I30128: std_logic; attribute dont_touch of I30128: signal is true;
	signal I30131: std_logic; attribute dont_touch of I30131: signal is true;
	signal I30134: std_logic; attribute dont_touch of I30134: signal is true;
	signal I30137: std_logic; attribute dont_touch of I30137: signal is true;
	signal I30140: std_logic; attribute dont_touch of I30140: signal is true;
	signal I30143: std_logic; attribute dont_touch of I30143: signal is true;
	signal I30146: std_logic; attribute dont_touch of I30146: signal is true;
	signal I30149: std_logic; attribute dont_touch of I30149: signal is true;
	signal I30152: std_logic; attribute dont_touch of I30152: signal is true;
	signal I30155: std_logic; attribute dont_touch of I30155: signal is true;
	signal I30158: std_logic; attribute dont_touch of I30158: signal is true;
	signal I30161: std_logic; attribute dont_touch of I30161: signal is true;
	signal I30164: std_logic; attribute dont_touch of I30164: signal is true;
	signal I30167: std_logic; attribute dont_touch of I30167: signal is true;
	signal I30170: std_logic; attribute dont_touch of I30170: signal is true;
	signal I30173: std_logic; attribute dont_touch of I30173: signal is true;
	signal I30176: std_logic; attribute dont_touch of I30176: signal is true;
	signal I30179: std_logic; attribute dont_touch of I30179: signal is true;
	signal I30182: std_logic; attribute dont_touch of I30182: signal is true;
	signal I30185: std_logic; attribute dont_touch of I30185: signal is true;
	signal I30188: std_logic; attribute dont_touch of I30188: signal is true;
	signal I30191: std_logic; attribute dont_touch of I30191: signal is true;
	signal I30194: std_logic; attribute dont_touch of I30194: signal is true;
	signal I30197: std_logic; attribute dont_touch of I30197: signal is true;
	signal I30200: std_logic; attribute dont_touch of I30200: signal is true;
	signal I30203: std_logic; attribute dont_touch of I30203: signal is true;
	signal I30206: std_logic; attribute dont_touch of I30206: signal is true;
	signal I30209: std_logic; attribute dont_touch of I30209: signal is true;
	signal I30212: std_logic; attribute dont_touch of I30212: signal is true;
	signal I30215: std_logic; attribute dont_touch of I30215: signal is true;
	signal I30218: std_logic; attribute dont_touch of I30218: signal is true;
	signal I30221: std_logic; attribute dont_touch of I30221: signal is true;
	signal I30224: std_logic; attribute dont_touch of I30224: signal is true;
	signal I30227: std_logic; attribute dont_touch of I30227: signal is true;
	signal I30230: std_logic; attribute dont_touch of I30230: signal is true;
	signal I30233: std_logic; attribute dont_touch of I30233: signal is true;
	signal I30236: std_logic; attribute dont_touch of I30236: signal is true;
	signal I30239: std_logic; attribute dont_touch of I30239: signal is true;
	signal I30242: std_logic; attribute dont_touch of I30242: signal is true;
	signal I30245: std_logic; attribute dont_touch of I30245: signal is true;
	signal I30248: std_logic; attribute dont_touch of I30248: signal is true;
	signal I30251: std_logic; attribute dont_touch of I30251: signal is true;
	signal I30254: std_logic; attribute dont_touch of I30254: signal is true;
	signal I30257: std_logic; attribute dont_touch of I30257: signal is true;
	signal I30260: std_logic; attribute dont_touch of I30260: signal is true;
	signal I30263: std_logic; attribute dont_touch of I30263: signal is true;
	signal I30266: std_logic; attribute dont_touch of I30266: signal is true;
	signal I30269: std_logic; attribute dont_touch of I30269: signal is true;
	signal I30272: std_logic; attribute dont_touch of I30272: signal is true;
	signal I30275: std_logic; attribute dont_touch of I30275: signal is true;
	signal I30278: std_logic; attribute dont_touch of I30278: signal is true;
	signal I30281: std_logic; attribute dont_touch of I30281: signal is true;
	signal I30284: std_logic; attribute dont_touch of I30284: signal is true;
	signal I30287: std_logic; attribute dont_touch of I30287: signal is true;
	signal I30290: std_logic; attribute dont_touch of I30290: signal is true;
	signal I30293: std_logic; attribute dont_touch of I30293: signal is true;
	signal I30296: std_logic; attribute dont_touch of I30296: signal is true;
	signal I30299: std_logic; attribute dont_touch of I30299: signal is true;
	signal I30302: std_logic; attribute dont_touch of I30302: signal is true;
	signal I30305: std_logic; attribute dont_touch of I30305: signal is true;
	signal I30308: std_logic; attribute dont_touch of I30308: signal is true;
	signal I30311: std_logic; attribute dont_touch of I30311: signal is true;
	signal I30314: std_logic; attribute dont_touch of I30314: signal is true;
	signal I30317: std_logic; attribute dont_touch of I30317: signal is true;
	signal I30320: std_logic; attribute dont_touch of I30320: signal is true;
	signal I30323: std_logic; attribute dont_touch of I30323: signal is true;
	signal I30326: std_logic; attribute dont_touch of I30326: signal is true;
	signal I30329: std_logic; attribute dont_touch of I30329: signal is true;
	signal I30332: std_logic; attribute dont_touch of I30332: signal is true;
	signal I30335: std_logic; attribute dont_touch of I30335: signal is true;
	signal I30338: std_logic; attribute dont_touch of I30338: signal is true;
	signal I30341: std_logic; attribute dont_touch of I30341: signal is true;
	signal I30344: std_logic; attribute dont_touch of I30344: signal is true;
	signal I30347: std_logic; attribute dont_touch of I30347: signal is true;
	signal I30350: std_logic; attribute dont_touch of I30350: signal is true;
	signal I30353: std_logic; attribute dont_touch of I30353: signal is true;
	signal I30356: std_logic; attribute dont_touch of I30356: signal is true;
	signal I30359: std_logic; attribute dont_touch of I30359: signal is true;
	signal I30362: std_logic; attribute dont_touch of I30362: signal is true;
	signal I30365: std_logic; attribute dont_touch of I30365: signal is true;
	signal I30368: std_logic; attribute dont_touch of I30368: signal is true;
	signal I30371: std_logic; attribute dont_touch of I30371: signal is true;
	signal I30374: std_logic; attribute dont_touch of I30374: signal is true;
	signal I30377: std_logic; attribute dont_touch of I30377: signal is true;
	signal I30380: std_logic; attribute dont_touch of I30380: signal is true;
	signal I30383: std_logic; attribute dont_touch of I30383: signal is true;
	signal I30386: std_logic; attribute dont_touch of I30386: signal is true;
	signal I30389: std_logic; attribute dont_touch of I30389: signal is true;
	signal I30392: std_logic; attribute dont_touch of I30392: signal is true;
	signal I30395: std_logic; attribute dont_touch of I30395: signal is true;
	signal I30398: std_logic; attribute dont_touch of I30398: signal is true;
	signal I30401: std_logic; attribute dont_touch of I30401: signal is true;
	signal I30404: std_logic; attribute dont_touch of I30404: signal is true;
	signal I30407: std_logic; attribute dont_touch of I30407: signal is true;
	signal I30467: std_logic; attribute dont_touch of I30467: signal is true;
	signal I30470: std_logic; attribute dont_touch of I30470: signal is true;
	signal I30476: std_logic; attribute dont_touch of I30476: signal is true;
	signal I30480: std_logic; attribute dont_touch of I30480: signal is true;
	signal I30483: std_logic; attribute dont_touch of I30483: signal is true;
	signal I30486: std_logic; attribute dont_touch of I30486: signal is true;
	signal I30489: std_logic; attribute dont_touch of I30489: signal is true;
	signal I30493: std_logic; attribute dont_touch of I30493: signal is true;
	signal I30496: std_logic; attribute dont_touch of I30496: signal is true;
	signal I30501: std_logic; attribute dont_touch of I30501: signal is true;
	signal I30504: std_logic; attribute dont_touch of I30504: signal is true;
	signal I30508: std_logic; attribute dont_touch of I30508: signal is true;
	signal I30511: std_logic; attribute dont_touch of I30511: signal is true;
	signal I30516: std_logic; attribute dont_touch of I30516: signal is true;
	signal I30519: std_logic; attribute dont_touch of I30519: signal is true;
	signal I30525: std_logic; attribute dont_touch of I30525: signal is true;
	signal I30531: std_logic; attribute dont_touch of I30531: signal is true;
	signal I30536: std_logic; attribute dont_touch of I30536: signal is true;
	signal I30544: std_logic; attribute dont_touch of I30544: signal is true;
	signal I30547: std_logic; attribute dont_touch of I30547: signal is true;
	signal I30552: std_logic; attribute dont_touch of I30552: signal is true;
	signal I30560: std_logic; attribute dont_touch of I30560: signal is true;
	signal I30563: std_logic; attribute dont_touch of I30563: signal is true;
	signal I30568: std_logic; attribute dont_touch of I30568: signal is true;
	signal I30575: std_logic; attribute dont_touch of I30575: signal is true;
	signal I30578: std_logic; attribute dont_touch of I30578: signal is true;
	signal I30586: std_logic; attribute dont_touch of I30586: signal is true;
	signal I30589: std_logic; attribute dont_touch of I30589: signal is true;
	signal I30594: std_logic; attribute dont_touch of I30594: signal is true;
	signal I30598: std_logic; attribute dont_touch of I30598: signal is true;
	signal I30601: std_logic; attribute dont_touch of I30601: signal is true;
	signal I30607: std_logic; attribute dont_touch of I30607: signal is true;
	signal I30611: std_logic; attribute dont_touch of I30611: signal is true;
	signal I30614: std_logic; attribute dont_touch of I30614: signal is true;
	signal I30617: std_logic; attribute dont_touch of I30617: signal is true;
	signal I30623: std_logic; attribute dont_touch of I30623: signal is true;
	signal I30626: std_logic; attribute dont_touch of I30626: signal is true;
	signal I30632: std_logic; attribute dont_touch of I30632: signal is true;
	signal I30636: std_logic; attribute dont_touch of I30636: signal is true;
	signal I30639: std_logic; attribute dont_touch of I30639: signal is true;
	signal I30642: std_logic; attribute dont_touch of I30642: signal is true;
	signal I30648: std_logic; attribute dont_touch of I30648: signal is true;
	signal I30651: std_logic; attribute dont_touch of I30651: signal is true;
	signal I30654: std_logic; attribute dont_touch of I30654: signal is true;
	signal I30660: std_logic; attribute dont_touch of I30660: signal is true;
	signal I30663: std_logic; attribute dont_touch of I30663: signal is true;
	signal I30669: std_logic; attribute dont_touch of I30669: signal is true;
	signal I30673: std_logic; attribute dont_touch of I30673: signal is true;
	signal I30676: std_logic; attribute dont_touch of I30676: signal is true;
	signal I30679: std_logic; attribute dont_touch of I30679: signal is true;
	signal I30686: std_logic; attribute dont_touch of I30686: signal is true;
	signal I30689: std_logic; attribute dont_touch of I30689: signal is true;
	signal I30692: std_logic; attribute dont_touch of I30692: signal is true;
	signal I30695: std_logic; attribute dont_touch of I30695: signal is true;
	signal I30701: std_logic; attribute dont_touch of I30701: signal is true;
	signal I30704: std_logic; attribute dont_touch of I30704: signal is true;
	signal I30707: std_logic; attribute dont_touch of I30707: signal is true;
	signal I30713: std_logic; attribute dont_touch of I30713: signal is true;
	signal I30716: std_logic; attribute dont_touch of I30716: signal is true;
	signal I30722: std_logic; attribute dont_touch of I30722: signal is true;
	signal I30725: std_logic; attribute dont_touch of I30725: signal is true;
	signal I30728: std_logic; attribute dont_touch of I30728: signal is true;
	signal I30735: std_logic; attribute dont_touch of I30735: signal is true;
	signal I30738: std_logic; attribute dont_touch of I30738: signal is true;
	signal I30741: std_logic; attribute dont_touch of I30741: signal is true;
	signal I30748: std_logic; attribute dont_touch of I30748: signal is true;
	signal I30751: std_logic; attribute dont_touch of I30751: signal is true;
	signal I30754: std_logic; attribute dont_touch of I30754: signal is true;
	signal I30757: std_logic; attribute dont_touch of I30757: signal is true;
	signal I30763: std_logic; attribute dont_touch of I30763: signal is true;
	signal I30766: std_logic; attribute dont_touch of I30766: signal is true;
	signal I30769: std_logic; attribute dont_touch of I30769: signal is true;
	signal I30776: std_logic; attribute dont_touch of I30776: signal is true;
	signal I30779: std_logic; attribute dont_touch of I30779: signal is true;
	signal I30782: std_logic; attribute dont_touch of I30782: signal is true;
	signal I30786: std_logic; attribute dont_touch of I30786: signal is true;
	signal I30790: std_logic; attribute dont_touch of I30790: signal is true;
	signal I30791: std_logic; attribute dont_touch of I30791: signal is true;
	signal I30792: std_logic; attribute dont_touch of I30792: signal is true;
	signal I30797: std_logic; attribute dont_touch of I30797: signal is true;
	signal I30800: std_logic; attribute dont_touch of I30800: signal is true;
	signal I30803: std_logic; attribute dont_touch of I30803: signal is true;
	signal I30810: std_logic; attribute dont_touch of I30810: signal is true;
	signal I30813: std_logic; attribute dont_touch of I30813: signal is true;
	signal I30816: std_logic; attribute dont_touch of I30816: signal is true;
	signal I30823: std_logic; attribute dont_touch of I30823: signal is true;
	signal I30826: std_logic; attribute dont_touch of I30826: signal is true;
	signal I30829: std_logic; attribute dont_touch of I30829: signal is true;
	signal I30832: std_logic; attribute dont_touch of I30832: signal is true;
	signal I30838: std_logic; attribute dont_touch of I30838: signal is true;
	signal I30841: std_logic; attribute dont_touch of I30841: signal is true;
	signal I30844: std_logic; attribute dont_touch of I30844: signal is true;
	signal I30847: std_logic; attribute dont_touch of I30847: signal is true;
	signal I30854: std_logic; attribute dont_touch of I30854: signal is true;
	signal I30857: std_logic; attribute dont_touch of I30857: signal is true;
	signal I30860: std_logic; attribute dont_touch of I30860: signal is true;
	signal I30864: std_logic; attribute dont_touch of I30864: signal is true;
	signal I30868: std_logic; attribute dont_touch of I30868: signal is true;
	signal I30869: std_logic; attribute dont_touch of I30869: signal is true;
	signal I30870: std_logic; attribute dont_touch of I30870: signal is true;
	signal I30875: std_logic; attribute dont_touch of I30875: signal is true;
	signal I30878: std_logic; attribute dont_touch of I30878: signal is true;
	signal I30881: std_logic; attribute dont_touch of I30881: signal is true;
	signal I30888: std_logic; attribute dont_touch of I30888: signal is true;
	signal I30891: std_logic; attribute dont_touch of I30891: signal is true;
	signal I30894: std_logic; attribute dont_touch of I30894: signal is true;
	signal I30901: std_logic; attribute dont_touch of I30901: signal is true;
	signal I30905: std_logic; attribute dont_touch of I30905: signal is true;
	signal I30908: std_logic; attribute dont_touch of I30908: signal is true;
	signal I30911: std_logic; attribute dont_touch of I30911: signal is true;
	signal I30914: std_logic; attribute dont_touch of I30914: signal is true;
	signal I30917: std_logic; attribute dont_touch of I30917: signal is true;
	signal I30922: std_logic; attribute dont_touch of I30922: signal is true;
	signal I30925: std_logic; attribute dont_touch of I30925: signal is true;
	signal I30928: std_logic; attribute dont_touch of I30928: signal is true;
	signal I30931: std_logic; attribute dont_touch of I30931: signal is true;
	signal I30938: std_logic; attribute dont_touch of I30938: signal is true;
	signal I30941: std_logic; attribute dont_touch of I30941: signal is true;
	signal I30944: std_logic; attribute dont_touch of I30944: signal is true;
	signal I30948: std_logic; attribute dont_touch of I30948: signal is true;
	signal I30952: std_logic; attribute dont_touch of I30952: signal is true;
	signal I30953: std_logic; attribute dont_touch of I30953: signal is true;
	signal I30954: std_logic; attribute dont_touch of I30954: signal is true;
	signal I30959: std_logic; attribute dont_touch of I30959: signal is true;
	signal I30962: std_logic; attribute dont_touch of I30962: signal is true;
	signal I30965: std_logic; attribute dont_touch of I30965: signal is true;
	signal I30973: std_logic; attribute dont_touch of I30973: signal is true;
	signal I30976: std_logic; attribute dont_touch of I30976: signal is true;
	signal I30979: std_logic; attribute dont_touch of I30979: signal is true;
	signal I30985: std_logic; attribute dont_touch of I30985: signal is true;
	signal I30988: std_logic; attribute dont_touch of I30988: signal is true;
	signal I30991: std_logic; attribute dont_touch of I30991: signal is true;
	signal I30994: std_logic; attribute dont_touch of I30994: signal is true;
	signal I30997: std_logic; attribute dont_touch of I30997: signal is true;
	signal I31000: std_logic; attribute dont_touch of I31000: signal is true;
	signal I31005: std_logic; attribute dont_touch of I31005: signal is true;
	signal I31008: std_logic; attribute dont_touch of I31008: signal is true;
	signal I31011: std_logic; attribute dont_touch of I31011: signal is true;
	signal I31014: std_logic; attribute dont_touch of I31014: signal is true;
	signal I31021: std_logic; attribute dont_touch of I31021: signal is true;
	signal I31024: std_logic; attribute dont_touch of I31024: signal is true;
	signal I31027: std_logic; attribute dont_touch of I31027: signal is true;
	signal I31031: std_logic; attribute dont_touch of I31031: signal is true;
	signal I31035: std_logic; attribute dont_touch of I31035: signal is true;
	signal I31036: std_logic; attribute dont_touch of I31036: signal is true;
	signal I31037: std_logic; attribute dont_touch of I31037: signal is true;
	signal I31043: std_logic; attribute dont_touch of I31043: signal is true;
	signal I31050: std_logic; attribute dont_touch of I31050: signal is true;
	signal I31053: std_logic; attribute dont_touch of I31053: signal is true;
	signal I31056: std_logic; attribute dont_touch of I31056: signal is true;
	signal I31062: std_logic; attribute dont_touch of I31062: signal is true;
	signal I31065: std_logic; attribute dont_touch of I31065: signal is true;
	signal I31068: std_logic; attribute dont_touch of I31068: signal is true;
	signal I31071: std_logic; attribute dont_touch of I31071: signal is true;
	signal I31074: std_logic; attribute dont_touch of I31074: signal is true;
	signal I31077: std_logic; attribute dont_touch of I31077: signal is true;
	signal I31082: std_logic; attribute dont_touch of I31082: signal is true;
	signal I31085: std_logic; attribute dont_touch of I31085: signal is true;
	signal I31088: std_logic; attribute dont_touch of I31088: signal is true;
	signal I31091: std_logic; attribute dont_touch of I31091: signal is true;
	signal I31102: std_logic; attribute dont_touch of I31102: signal is true;
	signal I31109: std_logic; attribute dont_touch of I31109: signal is true;
	signal I31112: std_logic; attribute dont_touch of I31112: signal is true;
	signal I31115: std_logic; attribute dont_touch of I31115: signal is true;
	signal I31121: std_logic; attribute dont_touch of I31121: signal is true;
	signal I31124: std_logic; attribute dont_touch of I31124: signal is true;
	signal I31127: std_logic; attribute dont_touch of I31127: signal is true;
	signal I31130: std_logic; attribute dont_touch of I31130: signal is true;
	signal I31133: std_logic; attribute dont_touch of I31133: signal is true;
	signal I31136: std_logic; attribute dont_touch of I31136: signal is true;
	signal I31141: std_logic; attribute dont_touch of I31141: signal is true;
	signal I31144: std_logic; attribute dont_touch of I31144: signal is true;
	signal I31152: std_logic; attribute dont_touch of I31152: signal is true;
	signal I31159: std_logic; attribute dont_touch of I31159: signal is true;
	signal I31162: std_logic; attribute dont_touch of I31162: signal is true;
	signal I31165: std_logic; attribute dont_touch of I31165: signal is true;
	signal I31171: std_logic; attribute dont_touch of I31171: signal is true;
	signal I31181: std_logic; attribute dont_touch of I31181: signal is true;
	signal I31188: std_logic; attribute dont_touch of I31188: signal is true;
	signal I31195: std_logic; attribute dont_touch of I31195: signal is true;
	signal I31205: std_logic; attribute dont_touch of I31205: signal is true;
	signal I31213: std_logic; attribute dont_touch of I31213: signal is true;
	signal I31226: std_logic; attribute dont_touch of I31226: signal is true;
	signal I31232: std_logic; attribute dont_touch of I31232: signal is true;
	signal I31235: std_logic; attribute dont_touch of I31235: signal is true;
	signal I31244: std_logic; attribute dont_touch of I31244: signal is true;
	signal I31250: std_logic; attribute dont_touch of I31250: signal is true;
	signal I31253: std_logic; attribute dont_touch of I31253: signal is true;
	signal I31257: std_logic; attribute dont_touch of I31257: signal is true;
	signal I31266: std_logic; attribute dont_touch of I31266: signal is true;
	signal I31270: std_logic; attribute dont_touch of I31270: signal is true;
	signal I31274: std_logic; attribute dont_touch of I31274: signal is true;
	signal I31282: std_logic; attribute dont_touch of I31282: signal is true;
	signal I31286: std_logic; attribute dont_touch of I31286: signal is true;
	signal I31290: std_logic; attribute dont_touch of I31290: signal is true;
	signal I31298: std_logic; attribute dont_touch of I31298: signal is true;
	signal I31302: std_logic; attribute dont_touch of I31302: signal is true;
	signal I31310: std_logic; attribute dont_touch of I31310: signal is true;
	signal I31387: std_logic; attribute dont_touch of I31387: signal is true;
	signal I31417: std_logic; attribute dont_touch of I31417: signal is true;
	signal I31426: std_logic; attribute dont_touch of I31426: signal is true;
	signal I31436: std_logic; attribute dont_touch of I31436: signal is true;
	signal I31445: std_logic; attribute dont_touch of I31445: signal is true;
	signal I31451: std_logic; attribute dont_touch of I31451: signal is true;
	signal I31454: std_logic; attribute dont_touch of I31454: signal is true;
	signal I31457: std_logic; attribute dont_touch of I31457: signal is true;
	signal I31460: std_logic; attribute dont_touch of I31460: signal is true;
	signal I31463: std_logic; attribute dont_touch of I31463: signal is true;
	signal I31466: std_logic; attribute dont_touch of I31466: signal is true;
	signal I31469: std_logic; attribute dont_touch of I31469: signal is true;
	signal I31472: std_logic; attribute dont_touch of I31472: signal is true;
	signal I31475: std_logic; attribute dont_touch of I31475: signal is true;
	signal I31478: std_logic; attribute dont_touch of I31478: signal is true;
	signal I31481: std_logic; attribute dont_touch of I31481: signal is true;
	signal I31484: std_logic; attribute dont_touch of I31484: signal is true;
	signal I31487: std_logic; attribute dont_touch of I31487: signal is true;
	signal I31490: std_logic; attribute dont_touch of I31490: signal is true;
	signal I31493: std_logic; attribute dont_touch of I31493: signal is true;
	signal I31496: std_logic; attribute dont_touch of I31496: signal is true;
	signal I31499: std_logic; attribute dont_touch of I31499: signal is true;
	signal I31502: std_logic; attribute dont_touch of I31502: signal is true;
	signal I31505: std_logic; attribute dont_touch of I31505: signal is true;
	signal I31508: std_logic; attribute dont_touch of I31508: signal is true;
	signal I31511: std_logic; attribute dont_touch of I31511: signal is true;
	signal I31514: std_logic; attribute dont_touch of I31514: signal is true;
	signal I31517: std_logic; attribute dont_touch of I31517: signal is true;
	signal I31520: std_logic; attribute dont_touch of I31520: signal is true;
	signal I31523: std_logic; attribute dont_touch of I31523: signal is true;
	signal I31526: std_logic; attribute dont_touch of I31526: signal is true;
	signal I31529: std_logic; attribute dont_touch of I31529: signal is true;
	signal I31532: std_logic; attribute dont_touch of I31532: signal is true;
	signal I31535: std_logic; attribute dont_touch of I31535: signal is true;
	signal I31538: std_logic; attribute dont_touch of I31538: signal is true;
	signal I31541: std_logic; attribute dont_touch of I31541: signal is true;
	signal I31544: std_logic; attribute dont_touch of I31544: signal is true;
	signal I31547: std_logic; attribute dont_touch of I31547: signal is true;
	signal I31550: std_logic; attribute dont_touch of I31550: signal is true;
	signal I31553: std_logic; attribute dont_touch of I31553: signal is true;
	signal I31556: std_logic; attribute dont_touch of I31556: signal is true;
	signal I31559: std_logic; attribute dont_touch of I31559: signal is true;
	signal I31562: std_logic; attribute dont_touch of I31562: signal is true;
	signal I31565: std_logic; attribute dont_touch of I31565: signal is true;
	signal I31568: std_logic; attribute dont_touch of I31568: signal is true;
	signal I31571: std_logic; attribute dont_touch of I31571: signal is true;
	signal I31574: std_logic; attribute dont_touch of I31574: signal is true;
	signal I31577: std_logic; attribute dont_touch of I31577: signal is true;
	signal I31580: std_logic; attribute dont_touch of I31580: signal is true;
	signal I31583: std_logic; attribute dont_touch of I31583: signal is true;
	signal I31586: std_logic; attribute dont_touch of I31586: signal is true;
	signal I31589: std_logic; attribute dont_touch of I31589: signal is true;
	signal I31592: std_logic; attribute dont_touch of I31592: signal is true;
	signal I31595: std_logic; attribute dont_touch of I31595: signal is true;
	signal I31598: std_logic; attribute dont_touch of I31598: signal is true;
	signal I31601: std_logic; attribute dont_touch of I31601: signal is true;
	signal I31604: std_logic; attribute dont_touch of I31604: signal is true;
	signal I31607: std_logic; attribute dont_touch of I31607: signal is true;
	signal I31610: std_logic; attribute dont_touch of I31610: signal is true;
	signal I31613: std_logic; attribute dont_touch of I31613: signal is true;
	signal I31616: std_logic; attribute dont_touch of I31616: signal is true;
	signal I31619: std_logic; attribute dont_touch of I31619: signal is true;
	signal I31622: std_logic; attribute dont_touch of I31622: signal is true;
	signal I31625: std_logic; attribute dont_touch of I31625: signal is true;
	signal I31628: std_logic; attribute dont_touch of I31628: signal is true;
	signal I31631: std_logic; attribute dont_touch of I31631: signal is true;
	signal I31634: std_logic; attribute dont_touch of I31634: signal is true;
	signal I31637: std_logic; attribute dont_touch of I31637: signal is true;
	signal I31640: std_logic; attribute dont_touch of I31640: signal is true;
	signal I31643: std_logic; attribute dont_touch of I31643: signal is true;
	signal I31646: std_logic; attribute dont_touch of I31646: signal is true;
	signal I31649: std_logic; attribute dont_touch of I31649: signal is true;
	signal I31652: std_logic; attribute dont_touch of I31652: signal is true;
	signal I31655: std_logic; attribute dont_touch of I31655: signal is true;
	signal I31658: std_logic; attribute dont_touch of I31658: signal is true;
	signal I31661: std_logic; attribute dont_touch of I31661: signal is true;
	signal I31664: std_logic; attribute dont_touch of I31664: signal is true;
	signal I31667: std_logic; attribute dont_touch of I31667: signal is true;
	signal I31670: std_logic; attribute dont_touch of I31670: signal is true;
	signal I31673: std_logic; attribute dont_touch of I31673: signal is true;
	signal I31676: std_logic; attribute dont_touch of I31676: signal is true;
	signal I31679: std_logic; attribute dont_touch of I31679: signal is true;
	signal I31682: std_logic; attribute dont_touch of I31682: signal is true;
	signal I31685: std_logic; attribute dont_touch of I31685: signal is true;
	signal I31688: std_logic; attribute dont_touch of I31688: signal is true;
	signal I31691: std_logic; attribute dont_touch of I31691: signal is true;
	signal I31694: std_logic; attribute dont_touch of I31694: signal is true;
	signal I31697: std_logic; attribute dont_touch of I31697: signal is true;
	signal I31700: std_logic; attribute dont_touch of I31700: signal is true;
	signal I31703: std_logic; attribute dont_touch of I31703: signal is true;
	signal I31706: std_logic; attribute dont_touch of I31706: signal is true;
	signal I31709: std_logic; attribute dont_touch of I31709: signal is true;
	signal I31712: std_logic; attribute dont_touch of I31712: signal is true;
	signal I31715: std_logic; attribute dont_touch of I31715: signal is true;
	signal I31718: std_logic; attribute dont_touch of I31718: signal is true;
	signal I31721: std_logic; attribute dont_touch of I31721: signal is true;
	signal I31724: std_logic; attribute dont_touch of I31724: signal is true;
	signal I31727: std_logic; attribute dont_touch of I31727: signal is true;
	signal I31730: std_logic; attribute dont_touch of I31730: signal is true;
	signal I31733: std_logic; attribute dont_touch of I31733: signal is true;
	signal I31736: std_logic; attribute dont_touch of I31736: signal is true;
	signal I31739: std_logic; attribute dont_touch of I31739: signal is true;
	signal I31742: std_logic; attribute dont_touch of I31742: signal is true;
	signal I31745: std_logic; attribute dont_touch of I31745: signal is true;
	signal I31748: std_logic; attribute dont_touch of I31748: signal is true;
	signal I31751: std_logic; attribute dont_touch of I31751: signal is true;
	signal I31754: std_logic; attribute dont_touch of I31754: signal is true;
	signal I31757: std_logic; attribute dont_touch of I31757: signal is true;
	signal I31760: std_logic; attribute dont_touch of I31760: signal is true;
	signal I31763: std_logic; attribute dont_touch of I31763: signal is true;
	signal I31766: std_logic; attribute dont_touch of I31766: signal is true;
	signal I31769: std_logic; attribute dont_touch of I31769: signal is true;
	signal I31772: std_logic; attribute dont_touch of I31772: signal is true;
	signal I31775: std_logic; attribute dont_touch of I31775: signal is true;
	signal I31778: std_logic; attribute dont_touch of I31778: signal is true;
	signal I31781: std_logic; attribute dont_touch of I31781: signal is true;
	signal I31784: std_logic; attribute dont_touch of I31784: signal is true;
	signal I31787: std_logic; attribute dont_touch of I31787: signal is true;
	signal I31790: std_logic; attribute dont_touch of I31790: signal is true;
	signal I31793: std_logic; attribute dont_touch of I31793: signal is true;
	signal I31796: std_logic; attribute dont_touch of I31796: signal is true;
	signal I31799: std_logic; attribute dont_touch of I31799: signal is true;
	signal I31802: std_logic; attribute dont_touch of I31802: signal is true;
	signal I31805: std_logic; attribute dont_touch of I31805: signal is true;
	signal I31808: std_logic; attribute dont_touch of I31808: signal is true;
	signal I31811: std_logic; attribute dont_touch of I31811: signal is true;
	signal I31814: std_logic; attribute dont_touch of I31814: signal is true;
	signal I31817: std_logic; attribute dont_touch of I31817: signal is true;
	signal I31820: std_logic; attribute dont_touch of I31820: signal is true;
	signal I31823: std_logic; attribute dont_touch of I31823: signal is true;
	signal I31826: std_logic; attribute dont_touch of I31826: signal is true;
	signal I31829: std_logic; attribute dont_touch of I31829: signal is true;
	signal I31832: std_logic; attribute dont_touch of I31832: signal is true;
	signal I31835: std_logic; attribute dont_touch of I31835: signal is true;
	signal I31838: std_logic; attribute dont_touch of I31838: signal is true;
	signal I31841: std_logic; attribute dont_touch of I31841: signal is true;
	signal I31844: std_logic; attribute dont_touch of I31844: signal is true;
	signal I31847: std_logic; attribute dont_touch of I31847: signal is true;
	signal I31850: std_logic; attribute dont_touch of I31850: signal is true;
	signal I31853: std_logic; attribute dont_touch of I31853: signal is true;
	signal I31856: std_logic; attribute dont_touch of I31856: signal is true;
	signal I31859: std_logic; attribute dont_touch of I31859: signal is true;
	signal I31862: std_logic; attribute dont_touch of I31862: signal is true;
	signal I31865: std_logic; attribute dont_touch of I31865: signal is true;
	signal I31868: std_logic; attribute dont_touch of I31868: signal is true;
	signal I31871: std_logic; attribute dont_touch of I31871: signal is true;
	signal I31874: std_logic; attribute dont_touch of I31874: signal is true;
	signal I31877: std_logic; attribute dont_touch of I31877: signal is true;
	signal I31880: std_logic; attribute dont_touch of I31880: signal is true;
	signal I31883: std_logic; attribute dont_touch of I31883: signal is true;
	signal I31886: std_logic; attribute dont_touch of I31886: signal is true;
	signal I31889: std_logic; attribute dont_touch of I31889: signal is true;
	signal I31892: std_logic; attribute dont_touch of I31892: signal is true;
	signal I31895: std_logic; attribute dont_touch of I31895: signal is true;
	signal I31898: std_logic; attribute dont_touch of I31898: signal is true;
	signal I31901: std_logic; attribute dont_touch of I31901: signal is true;
	signal I31904: std_logic; attribute dont_touch of I31904: signal is true;
	signal I31907: std_logic; attribute dont_touch of I31907: signal is true;
	signal I31910: std_logic; attribute dont_touch of I31910: signal is true;
	signal I31913: std_logic; attribute dont_touch of I31913: signal is true;
	signal I31916: std_logic; attribute dont_touch of I31916: signal is true;
	signal I31919: std_logic; attribute dont_touch of I31919: signal is true;
	signal I31922: std_logic; attribute dont_touch of I31922: signal is true;
	signal I31925: std_logic; attribute dont_touch of I31925: signal is true;
	signal I31928: std_logic; attribute dont_touch of I31928: signal is true;
	signal I31931: std_logic; attribute dont_touch of I31931: signal is true;
	signal I31934: std_logic; attribute dont_touch of I31934: signal is true;
	signal I31937: std_logic; attribute dont_touch of I31937: signal is true;
	signal I31940: std_logic; attribute dont_touch of I31940: signal is true;
	signal I31943: std_logic; attribute dont_touch of I31943: signal is true;
	signal I31946: std_logic; attribute dont_touch of I31946: signal is true;
	signal I31949: std_logic; attribute dont_touch of I31949: signal is true;
	signal I32042: std_logic; attribute dont_touch of I32042: signal is true;
	signal I32057: std_logic; attribute dont_touch of I32057: signal is true;
	signal I32067: std_logic; attribute dont_touch of I32067: signal is true;
	signal I32074: std_logic; attribute dont_touch of I32074: signal is true;
	signal I32081: std_logic; attribute dont_touch of I32081: signal is true;
	signal I32085: std_logic; attribute dont_touch of I32085: signal is true;
	signal I32092: std_logic; attribute dont_touch of I32092: signal is true;
	signal I32098: std_logic; attribute dont_touch of I32098: signal is true;
	signal I32102: std_logic; attribute dont_touch of I32102: signal is true;
	signal I32109: std_logic; attribute dont_touch of I32109: signal is true;
	signal I32112: std_logic; attribute dont_touch of I32112: signal is true;
	signal I32116: std_logic; attribute dont_touch of I32116: signal is true;
	signal I32120: std_logic; attribute dont_touch of I32120: signal is true;
	signal I32126: std_logic; attribute dont_touch of I32126: signal is true;
	signal I32129: std_logic; attribute dont_touch of I32129: signal is true;
	signal I32133: std_logic; attribute dont_touch of I32133: signal is true;
	signal I32137: std_logic; attribute dont_touch of I32137: signal is true;
	signal I32140: std_logic; attribute dont_touch of I32140: signal is true;
	signal I32143: std_logic; attribute dont_touch of I32143: signal is true;
	signal I32146: std_logic; attribute dont_touch of I32146: signal is true;
	signal I32150: std_logic; attribute dont_touch of I32150: signal is true;
	signal I32153: std_logic; attribute dont_touch of I32153: signal is true;
	signal I32156: std_logic; attribute dont_touch of I32156: signal is true;
	signal I32159: std_logic; attribute dont_touch of I32159: signal is true;
	signal I32164: std_logic; attribute dont_touch of I32164: signal is true;
	signal I32167: std_logic; attribute dont_touch of I32167: signal is true;
	signal I32170: std_logic; attribute dont_touch of I32170: signal is true;
	signal I32175: std_logic; attribute dont_touch of I32175: signal is true;
	signal I32178: std_logic; attribute dont_touch of I32178: signal is true;
	signal I32181: std_logic; attribute dont_touch of I32181: signal is true;
	signal I32184: std_logic; attribute dont_touch of I32184: signal is true;
	signal I32189: std_logic; attribute dont_touch of I32189: signal is true;
	signal I32193: std_logic; attribute dont_touch of I32193: signal is true;
	signal I32198: std_logic; attribute dont_touch of I32198: signal is true;
	signal I32203: std_logic; attribute dont_touch of I32203: signal is true;
	signal I32210: std_logic; attribute dont_touch of I32210: signal is true;
	signal I32248: std_logic; attribute dont_touch of I32248: signal is true;
	signal I32251: std_logic; attribute dont_touch of I32251: signal is true;
	signal I32265: std_logic; attribute dont_touch of I32265: signal is true;
	signal I32266: std_logic; attribute dont_touch of I32266: signal is true;
	signal I32267: std_logic; attribute dont_touch of I32267: signal is true;
	signal I32281: std_logic; attribute dont_touch of I32281: signal is true;
	signal I32284: std_logic; attribute dont_touch of I32284: signal is true;
	signal I32285: std_logic; attribute dont_touch of I32285: signal is true;
	signal I32286: std_logic; attribute dont_touch of I32286: signal is true;
	signal I32295: std_logic; attribute dont_touch of I32295: signal is true;
	signal I32296: std_logic; attribute dont_touch of I32296: signal is true;
	signal I32297: std_logic; attribute dont_touch of I32297: signal is true;
	signal I32308: std_logic; attribute dont_touch of I32308: signal is true;
	signal I32309: std_logic; attribute dont_touch of I32309: signal is true;
	signal I32310: std_logic; attribute dont_touch of I32310: signal is true;
	signal I32320: std_logic; attribute dont_touch of I32320: signal is true;
	signal I32323: std_logic; attribute dont_touch of I32323: signal is true;
	signal I32324: std_logic; attribute dont_touch of I32324: signal is true;
	signal I32325: std_logic; attribute dont_touch of I32325: signal is true;
	signal I32333: std_logic; attribute dont_touch of I32333: signal is true;
	signal I32334: std_logic; attribute dont_touch of I32334: signal is true;
	signal I32335: std_logic; attribute dont_touch of I32335: signal is true;
	signal I32345: std_logic; attribute dont_touch of I32345: signal is true;
	signal I32346: std_logic; attribute dont_touch of I32346: signal is true;
	signal I32347: std_logic; attribute dont_touch of I32347: signal is true;
	signal I32355: std_logic; attribute dont_touch of I32355: signal is true;
	signal I32356: std_logic; attribute dont_touch of I32356: signal is true;
	signal I32357: std_logic; attribute dont_touch of I32357: signal is true;
	signal I32365: std_logic; attribute dont_touch of I32365: signal is true;
	signal I32368: std_logic; attribute dont_touch of I32368: signal is true;
	signal I32369: std_logic; attribute dont_touch of I32369: signal is true;
	signal I32370: std_logic; attribute dont_touch of I32370: signal is true;
	signal I32378: std_logic; attribute dont_touch of I32378: signal is true;
	signal I32379: std_logic; attribute dont_touch of I32379: signal is true;
	signal I32380: std_logic; attribute dont_touch of I32380: signal is true;
	signal I32388: std_logic; attribute dont_touch of I32388: signal is true;
	signal I32391: std_logic; attribute dont_touch of I32391: signal is true;
	signal I32392: std_logic; attribute dont_touch of I32392: signal is true;
	signal I32393: std_logic; attribute dont_touch of I32393: signal is true;
	signal I32400: std_logic; attribute dont_touch of I32400: signal is true;
	signal I32401: std_logic; attribute dont_touch of I32401: signal is true;
	signal I32402: std_logic; attribute dont_touch of I32402: signal is true;
	signal I32409: std_logic; attribute dont_touch of I32409: signal is true;
	signal I32410: std_logic; attribute dont_touch of I32410: signal is true;
	signal I32411: std_logic; attribute dont_touch of I32411: signal is true;
	signal I32419: std_logic; attribute dont_touch of I32419: signal is true;
	signal I32422: std_logic; attribute dont_touch of I32422: signal is true;
	signal I32423: std_logic; attribute dont_touch of I32423: signal is true;
	signal I32424: std_logic; attribute dont_touch of I32424: signal is true;
	signal I32430: std_logic; attribute dont_touch of I32430: signal is true;
	signal I32431: std_logic; attribute dont_touch of I32431: signal is true;
	signal I32432: std_logic; attribute dont_touch of I32432: signal is true;
	signal I32439: std_logic; attribute dont_touch of I32439: signal is true;
	signal I32443: std_logic; attribute dont_touch of I32443: signal is true;
	signal I32444: std_logic; attribute dont_touch of I32444: signal is true;
	signal I32445: std_logic; attribute dont_touch of I32445: signal is true;
	signal I32451: std_logic; attribute dont_touch of I32451: signal is true;
	signal I32452: std_logic; attribute dont_touch of I32452: signal is true;
	signal I32453: std_logic; attribute dont_touch of I32453: signal is true;
	signal I32460: std_logic; attribute dont_touch of I32460: signal is true;
	signal I32461: std_logic; attribute dont_touch of I32461: signal is true;
	signal I32462: std_logic; attribute dont_touch of I32462: signal is true;
	signal I32468: std_logic; attribute dont_touch of I32468: signal is true;
	signal I32469: std_logic; attribute dont_touch of I32469: signal is true;
	signal I32470: std_logic; attribute dont_touch of I32470: signal is true;
	signal I32478: std_logic; attribute dont_touch of I32478: signal is true;
	signal I32479: std_logic; attribute dont_touch of I32479: signal is true;
	signal I32480: std_logic; attribute dont_touch of I32480: signal is true;
	signal I32487: std_logic; attribute dont_touch of I32487: signal is true;
	signal I32490: std_logic; attribute dont_touch of I32490: signal is true;
	signal I32491: std_logic; attribute dont_touch of I32491: signal is true;
	signal I32492: std_logic; attribute dont_touch of I32492: signal is true;
	signal I32498: std_logic; attribute dont_touch of I32498: signal is true;
	signal I32499: std_logic; attribute dont_touch of I32499: signal is true;
	signal I32500: std_logic; attribute dont_touch of I32500: signal is true;
	signal I32506: std_logic; attribute dont_touch of I32506: signal is true;
	signal I32509: std_logic; attribute dont_touch of I32509: signal is true;
	signal I32510: std_logic; attribute dont_touch of I32510: signal is true;
	signal I32511: std_logic; attribute dont_touch of I32511: signal is true;
	signal I32518: std_logic; attribute dont_touch of I32518: signal is true;
	signal I32519: std_logic; attribute dont_touch of I32519: signal is true;
	signal I32520: std_logic; attribute dont_touch of I32520: signal is true;
	signal I32526: std_logic; attribute dont_touch of I32526: signal is true;
	signal I32527: std_logic; attribute dont_touch of I32527: signal is true;
	signal I32528: std_logic; attribute dont_touch of I32528: signal is true;
	signal I32535: std_logic; attribute dont_touch of I32535: signal is true;
	signal I32538: std_logic; attribute dont_touch of I32538: signal is true;
	signal I32539: std_logic; attribute dont_touch of I32539: signal is true;
	signal I32540: std_logic; attribute dont_touch of I32540: signal is true;
	signal I32546: std_logic; attribute dont_touch of I32546: signal is true;
	signal I32547: std_logic; attribute dont_touch of I32547: signal is true;
	signal I32548: std_logic; attribute dont_touch of I32548: signal is true;
	signal I32556: std_logic; attribute dont_touch of I32556: signal is true;
	signal I32559: std_logic; attribute dont_touch of I32559: signal is true;
	signal I32560: std_logic; attribute dont_touch of I32560: signal is true;
	signal I32561: std_logic; attribute dont_touch of I32561: signal is true;
	signal I32567: std_logic; attribute dont_touch of I32567: signal is true;
	signal I32568: std_logic; attribute dont_touch of I32568: signal is true;
	signal I32569: std_logic; attribute dont_touch of I32569: signal is true;
	signal I32575: std_logic; attribute dont_touch of I32575: signal is true;
	signal I32576: std_logic; attribute dont_touch of I32576: signal is true;
	signal I32577: std_logic; attribute dont_touch of I32577: signal is true;
	signal I32583: std_logic; attribute dont_touch of I32583: signal is true;
	signal I32586: std_logic; attribute dont_touch of I32586: signal is true;
	signal I32587: std_logic; attribute dont_touch of I32587: signal is true;
	signal I32588: std_logic; attribute dont_touch of I32588: signal is true;
	signal I32595: std_logic; attribute dont_touch of I32595: signal is true;
	signal I32596: std_logic; attribute dont_touch of I32596: signal is true;
	signal I32597: std_logic; attribute dont_touch of I32597: signal is true;
	signal I32604: std_logic; attribute dont_touch of I32604: signal is true;
	signal I32607: std_logic; attribute dont_touch of I32607: signal is true;
	signal I32608: std_logic; attribute dont_touch of I32608: signal is true;
	signal I32609: std_logic; attribute dont_touch of I32609: signal is true;
	signal I32615: std_logic; attribute dont_touch of I32615: signal is true;
	signal I32616: std_logic; attribute dont_touch of I32616: signal is true;
	signal I32617: std_logic; attribute dont_touch of I32617: signal is true;
	signal I32624: std_logic; attribute dont_touch of I32624: signal is true;
	signal I32625: std_logic; attribute dont_touch of I32625: signal is true;
	signal I32626: std_logic; attribute dont_touch of I32626: signal is true;
	signal I32633: std_logic; attribute dont_touch of I32633: signal is true;
	signal I32634: std_logic; attribute dont_touch of I32634: signal is true;
	signal I32635: std_logic; attribute dont_touch of I32635: signal is true;
	signal I32642: std_logic; attribute dont_touch of I32642: signal is true;
	signal I32645: std_logic; attribute dont_touch of I32645: signal is true;
	signal I32646: std_logic; attribute dont_touch of I32646: signal is true;
	signal I32647: std_logic; attribute dont_touch of I32647: signal is true;
	signal I32659: std_logic; attribute dont_touch of I32659: signal is true;
	signal I32660: std_logic; attribute dont_touch of I32660: signal is true;
	signal I32661: std_logic; attribute dont_touch of I32661: signal is true;
	signal I32668: std_logic; attribute dont_touch of I32668: signal is true;
	signal I32669: std_logic; attribute dont_touch of I32669: signal is true;
	signal I32670: std_logic; attribute dont_touch of I32670: signal is true;
	signal I32677: std_logic; attribute dont_touch of I32677: signal is true;
	signal I32678: std_logic; attribute dont_touch of I32678: signal is true;
	signal I32679: std_logic; attribute dont_touch of I32679: signal is true;
	signal I32686: std_logic; attribute dont_touch of I32686: signal is true;
	signal I32687: std_logic; attribute dont_touch of I32687: signal is true;
	signal I32688: std_logic; attribute dont_touch of I32688: signal is true;
	signal I32695: std_logic; attribute dont_touch of I32695: signal is true;
	signal I32696: std_logic; attribute dont_touch of I32696: signal is true;
	signal I32697: std_logic; attribute dont_touch of I32697: signal is true;
	signal I32704: std_logic; attribute dont_touch of I32704: signal is true;
	signal I32708: std_logic; attribute dont_touch of I32708: signal is true;
	signal I32709: std_logic; attribute dont_touch of I32709: signal is true;
	signal I32710: std_logic; attribute dont_touch of I32710: signal is true;
	signal I32716: std_logic; attribute dont_touch of I32716: signal is true;
	signal I32719: std_logic; attribute dont_touch of I32719: signal is true;
	signal I32724: std_logic; attribute dont_touch of I32724: signal is true;
	signal I32725: std_logic; attribute dont_touch of I32725: signal is true;
	signal I32726: std_logic; attribute dont_touch of I32726: signal is true;
	signal I32829: std_logic; attribute dont_touch of I32829: signal is true;
	signal I32835: std_logic; attribute dont_touch of I32835: signal is true;
	signal I32844: std_logic; attribute dont_touch of I32844: signal is true;
	signal I32847: std_logic; attribute dont_touch of I32847: signal is true;
	signal I32851: std_logic; attribute dont_touch of I32851: signal is true;
	signal I32854: std_logic; attribute dont_touch of I32854: signal is true;
	signal I32857: std_logic; attribute dont_touch of I32857: signal is true;
	signal I32860: std_logic; attribute dont_touch of I32860: signal is true;
	signal I32868: std_logic; attribute dont_touch of I32868: signal is true;
	signal I32871: std_logic; attribute dont_touch of I32871: signal is true;
	signal I32874: std_logic; attribute dont_touch of I32874: signal is true;
	signal I32877: std_logic; attribute dont_touch of I32877: signal is true;
	signal I32880: std_logic; attribute dont_touch of I32880: signal is true;
	signal I32883: std_logic; attribute dont_touch of I32883: signal is true;
	signal I32886: std_logic; attribute dont_touch of I32886: signal is true;
	signal I32889: std_logic; attribute dont_touch of I32889: signal is true;
	signal I32892: std_logic; attribute dont_touch of I32892: signal is true;
	signal I32895: std_logic; attribute dont_touch of I32895: signal is true;
	signal I32898: std_logic; attribute dont_touch of I32898: signal is true;
	signal I32901: std_logic; attribute dont_touch of I32901: signal is true;
	signal I32904: std_logic; attribute dont_touch of I32904: signal is true;
	signal I32907: std_logic; attribute dont_touch of I32907: signal is true;
	signal I32910: std_logic; attribute dont_touch of I32910: signal is true;
	signal I32913: std_logic; attribute dont_touch of I32913: signal is true;
	signal I32916: std_logic; attribute dont_touch of I32916: signal is true;
	signal I32919: std_logic; attribute dont_touch of I32919: signal is true;
	signal I32922: std_logic; attribute dont_touch of I32922: signal is true;
	signal I32925: std_logic; attribute dont_touch of I32925: signal is true;
	signal I32928: std_logic; attribute dont_touch of I32928: signal is true;
	signal I32931: std_logic; attribute dont_touch of I32931: signal is true;
	signal I32934: std_logic; attribute dont_touch of I32934: signal is true;
	signal I32937: std_logic; attribute dont_touch of I32937: signal is true;
	signal I32940: std_logic; attribute dont_touch of I32940: signal is true;
	signal I32943: std_logic; attribute dont_touch of I32943: signal is true;
	signal I32946: std_logic; attribute dont_touch of I32946: signal is true;
	signal I32949: std_logic; attribute dont_touch of I32949: signal is true;
	signal I32952: std_logic; attribute dont_touch of I32952: signal is true;
	signal I32955: std_logic; attribute dont_touch of I32955: signal is true;
	signal I32958: std_logic; attribute dont_touch of I32958: signal is true;
	signal I32961: std_logic; attribute dont_touch of I32961: signal is true;
	signal I32964: std_logic; attribute dont_touch of I32964: signal is true;
	signal I32967: std_logic; attribute dont_touch of I32967: signal is true;
	signal I32970: std_logic; attribute dont_touch of I32970: signal is true;
	signal I32973: std_logic; attribute dont_touch of I32973: signal is true;
	signal I32976: std_logic; attribute dont_touch of I32976: signal is true;
	signal I32979: std_logic; attribute dont_touch of I32979: signal is true;
	signal I32982: std_logic; attribute dont_touch of I32982: signal is true;
	signal I32985: std_logic; attribute dont_touch of I32985: signal is true;
	signal I32988: std_logic; attribute dont_touch of I32988: signal is true;
	signal I32991: std_logic; attribute dont_touch of I32991: signal is true;
	signal I32994: std_logic; attribute dont_touch of I32994: signal is true;
	signal I32997: std_logic; attribute dont_touch of I32997: signal is true;
	signal I33000: std_logic; attribute dont_touch of I33000: signal is true;
	signal I33003: std_logic; attribute dont_touch of I33003: signal is true;
	signal I33006: std_logic; attribute dont_touch of I33006: signal is true;
	signal I33009: std_logic; attribute dont_touch of I33009: signal is true;
	signal I33013: std_logic; attribute dont_touch of I33013: signal is true;
	signal I33016: std_logic; attribute dont_touch of I33016: signal is true;
	signal I33128: std_logic; attribute dont_touch of I33128: signal is true;
	signal I33136: std_logic; attribute dont_touch of I33136: signal is true;
	signal I33145: std_logic; attribute dont_touch of I33145: signal is true;
	signal I33154: std_logic; attribute dont_touch of I33154: signal is true;
	signal I33157: std_logic; attribute dont_touch of I33157: signal is true;
	signal I33168: std_logic; attribute dont_touch of I33168: signal is true;
	signal I33182: std_logic; attribute dont_touch of I33182: signal is true;
	signal I33188: std_logic; attribute dont_touch of I33188: signal is true;
	signal I33198: std_logic; attribute dont_touch of I33198: signal is true;
	signal I33205: std_logic; attribute dont_touch of I33205: signal is true;
	signal I33219: std_logic; attribute dont_touch of I33219: signal is true;
	signal I33232: std_logic; attribute dont_touch of I33232: signal is true;
	signal I33246: std_logic; attribute dont_touch of I33246: signal is true;
	signal I33249: std_logic; attribute dont_touch of I33249: signal is true;
	signal I33257: std_logic; attribute dont_touch of I33257: signal is true;
	signal I33260: std_logic; attribute dont_touch of I33260: signal is true;
	signal I33265: std_logic; attribute dont_touch of I33265: signal is true;
	signal I33268: std_logic; attribute dont_touch of I33268: signal is true;
	signal I33278: std_logic; attribute dont_touch of I33278: signal is true;
	signal I33282: std_logic; attribute dont_touch of I33282: signal is true;
	signal I33286: std_logic; attribute dont_touch of I33286: signal is true;
	signal I33289: std_logic; attribute dont_touch of I33289: signal is true;
	signal I33293: std_logic; attribute dont_touch of I33293: signal is true;
	signal I33297: std_logic; attribute dont_touch of I33297: signal is true;
	signal I33300: std_logic; attribute dont_touch of I33300: signal is true;
	signal I33304: std_logic; attribute dont_touch of I33304: signal is true;
	signal I33307: std_logic; attribute dont_touch of I33307: signal is true;
	signal I33312: std_logic; attribute dont_touch of I33312: signal is true;
	signal I33316: std_logic; attribute dont_touch of I33316: signal is true;
	signal I33321: std_logic; attribute dont_touch of I33321: signal is true;
	signal I33324: std_logic; attribute dont_touch of I33324: signal is true;
	signal I33327: std_logic; attribute dont_touch of I33327: signal is true;
	signal I33330: std_logic; attribute dont_touch of I33330: signal is true;
	signal I33335: std_logic; attribute dont_touch of I33335: signal is true;
	signal I33338: std_logic; attribute dont_touch of I33338: signal is true;
	signal I33343: std_logic; attribute dont_touch of I33343: signal is true;
	signal I33347: std_logic; attribute dont_touch of I33347: signal is true;
	signal I33352: std_logic; attribute dont_touch of I33352: signal is true;
	signal I33355: std_logic; attribute dont_touch of I33355: signal is true;
	signal I33358: std_logic; attribute dont_touch of I33358: signal is true;
	signal I33361: std_logic; attribute dont_touch of I33361: signal is true;
	signal I33364: std_logic; attribute dont_touch of I33364: signal is true;
	signal I33368: std_logic; attribute dont_touch of I33368: signal is true;
	signal I33371: std_logic; attribute dont_touch of I33371: signal is true;
	signal I33374: std_logic; attribute dont_touch of I33374: signal is true;
	signal I33377: std_logic; attribute dont_touch of I33377: signal is true;
	signal I33382: std_logic; attribute dont_touch of I33382: signal is true;
	signal I33385: std_logic; attribute dont_touch of I33385: signal is true;
	signal I33390: std_logic; attribute dont_touch of I33390: signal is true;
	signal I33396: std_logic; attribute dont_touch of I33396: signal is true;
	signal I33399: std_logic; attribute dont_touch of I33399: signal is true;
	signal I33402: std_logic; attribute dont_touch of I33402: signal is true;
	signal I33405: std_logic; attribute dont_touch of I33405: signal is true;
	signal I33408: std_logic; attribute dont_touch of I33408: signal is true;
	signal I33411: std_logic; attribute dont_touch of I33411: signal is true;
	signal I33415: std_logic; attribute dont_touch of I33415: signal is true;
	signal I33418: std_logic; attribute dont_touch of I33418: signal is true;
	signal I33421: std_logic; attribute dont_touch of I33421: signal is true;
	signal I33424: std_logic; attribute dont_touch of I33424: signal is true;
	signal I33427: std_logic; attribute dont_touch of I33427: signal is true;
	signal I33431: std_logic; attribute dont_touch of I33431: signal is true;
	signal I33434: std_logic; attribute dont_touch of I33434: signal is true;
	signal I33437: std_logic; attribute dont_touch of I33437: signal is true;
	signal I33440: std_logic; attribute dont_touch of I33440: signal is true;
	signal I33445: std_logic; attribute dont_touch of I33445: signal is true;
	signal I33448: std_logic; attribute dont_touch of I33448: signal is true;
	signal I33457: std_logic; attribute dont_touch of I33457: signal is true;
	signal I33460: std_logic; attribute dont_touch of I33460: signal is true;
	signal I33463: std_logic; attribute dont_touch of I33463: signal is true;
	signal I33466: std_logic; attribute dont_touch of I33466: signal is true;
	signal I33469: std_logic; attribute dont_touch of I33469: signal is true;
	signal I33472: std_logic; attribute dont_touch of I33472: signal is true;
	signal I33476: std_logic; attribute dont_touch of I33476: signal is true;
	signal I33479: std_logic; attribute dont_touch of I33479: signal is true;
	signal I33482: std_logic; attribute dont_touch of I33482: signal is true;
	signal I33485: std_logic; attribute dont_touch of I33485: signal is true;
	signal I33488: std_logic; attribute dont_touch of I33488: signal is true;
	signal I33491: std_logic; attribute dont_touch of I33491: signal is true;
	signal I33495: std_logic; attribute dont_touch of I33495: signal is true;
	signal I33498: std_logic; attribute dont_touch of I33498: signal is true;
	signal I33501: std_logic; attribute dont_touch of I33501: signal is true;
	signal I33504: std_logic; attribute dont_touch of I33504: signal is true;
	signal I33507: std_logic; attribute dont_touch of I33507: signal is true;
	signal I33511: std_logic; attribute dont_touch of I33511: signal is true;
	signal I33514: std_logic; attribute dont_touch of I33514: signal is true;
	signal I33517: std_logic; attribute dont_touch of I33517: signal is true;
	signal I33520: std_logic; attribute dont_touch of I33520: signal is true;
	signal I33526: std_logic; attribute dont_touch of I33526: signal is true;
	signal I33529: std_logic; attribute dont_touch of I33529: signal is true;
	signal I33532: std_logic; attribute dont_touch of I33532: signal is true;
	signal I33535: std_logic; attribute dont_touch of I33535: signal is true;
	signal I33539: std_logic; attribute dont_touch of I33539: signal is true;
	signal I33542: std_logic; attribute dont_touch of I33542: signal is true;
	signal I33545: std_logic; attribute dont_touch of I33545: signal is true;
	signal I33548: std_logic; attribute dont_touch of I33548: signal is true;
	signal I33551: std_logic; attribute dont_touch of I33551: signal is true;
	signal I33554: std_logic; attribute dont_touch of I33554: signal is true;
	signal I33558: std_logic; attribute dont_touch of I33558: signal is true;
	signal I33561: std_logic; attribute dont_touch of I33561: signal is true;
	signal I33564: std_logic; attribute dont_touch of I33564: signal is true;
	signal I33567: std_logic; attribute dont_touch of I33567: signal is true;
	signal I33570: std_logic; attribute dont_touch of I33570: signal is true;
	signal I33573: std_logic; attribute dont_touch of I33573: signal is true;
	signal I33577: std_logic; attribute dont_touch of I33577: signal is true;
	signal I33580: std_logic; attribute dont_touch of I33580: signal is true;
	signal I33583: std_logic; attribute dont_touch of I33583: signal is true;
	signal I33586: std_logic; attribute dont_touch of I33586: signal is true;
	signal I33589: std_logic; attribute dont_touch of I33589: signal is true;
	signal I33593: std_logic; attribute dont_touch of I33593: signal is true;
	signal I33596: std_logic; attribute dont_touch of I33596: signal is true;
	signal I33600: std_logic; attribute dont_touch of I33600: signal is true;
	signal I33603: std_logic; attribute dont_touch of I33603: signal is true;
	signal I33608: std_logic; attribute dont_touch of I33608: signal is true;
	signal I33611: std_logic; attribute dont_touch of I33611: signal is true;
	signal I33614: std_logic; attribute dont_touch of I33614: signal is true;
	signal I33617: std_logic; attribute dont_touch of I33617: signal is true;
	signal I33621: std_logic; attribute dont_touch of I33621: signal is true;
	signal I33624: std_logic; attribute dont_touch of I33624: signal is true;
	signal I33627: std_logic; attribute dont_touch of I33627: signal is true;
	signal I33630: std_logic; attribute dont_touch of I33630: signal is true;
	signal I33633: std_logic; attribute dont_touch of I33633: signal is true;
	signal I33636: std_logic; attribute dont_touch of I33636: signal is true;
	signal I33640: std_logic; attribute dont_touch of I33640: signal is true;
	signal I33643: std_logic; attribute dont_touch of I33643: signal is true;
	signal I33646: std_logic; attribute dont_touch of I33646: signal is true;
	signal I33649: std_logic; attribute dont_touch of I33649: signal is true;
	signal I33652: std_logic; attribute dont_touch of I33652: signal is true;
	signal I33655: std_logic; attribute dont_touch of I33655: signal is true;
	signal I33659: std_logic; attribute dont_touch of I33659: signal is true;
	signal I33662: std_logic; attribute dont_touch of I33662: signal is true;
	signal I33667: std_logic; attribute dont_touch of I33667: signal is true;
	signal I33670: std_logic; attribute dont_touch of I33670: signal is true;
	signal I33673: std_logic; attribute dont_touch of I33673: signal is true;
	signal I33676: std_logic; attribute dont_touch of I33676: signal is true;
	signal I33680: std_logic; attribute dont_touch of I33680: signal is true;
	signal I33683: std_logic; attribute dont_touch of I33683: signal is true;
	signal I33686: std_logic; attribute dont_touch of I33686: signal is true;
	signal I33689: std_logic; attribute dont_touch of I33689: signal is true;
	signal I33692: std_logic; attribute dont_touch of I33692: signal is true;
	signal I33695: std_logic; attribute dont_touch of I33695: signal is true;
	signal I33700: std_logic; attribute dont_touch of I33700: signal is true;
	signal I33703: std_logic; attribute dont_touch of I33703: signal is true;
	signal I33708: std_logic; attribute dont_touch of I33708: signal is true;
	signal I33711: std_logic; attribute dont_touch of I33711: signal is true;
	signal I33714: std_logic; attribute dont_touch of I33714: signal is true;
	signal I33717: std_logic; attribute dont_touch of I33717: signal is true;
	signal I33723: std_logic; attribute dont_touch of I33723: signal is true;
	signal I33726: std_logic; attribute dont_touch of I33726: signal is true;
	signal I33732: std_logic; attribute dont_touch of I33732: signal is true;
	signal I33737: std_logic; attribute dont_touch of I33737: signal is true;
	signal I33790: std_logic; attribute dont_touch of I33790: signal is true;
	signal I33798: std_logic; attribute dont_touch of I33798: signal is true;
	signal I33801: std_logic; attribute dont_touch of I33801: signal is true;
	signal I33804: std_logic; attribute dont_touch of I33804: signal is true;
	signal I33807: std_logic; attribute dont_touch of I33807: signal is true;
	signal I33810: std_logic; attribute dont_touch of I33810: signal is true;
	signal I33813: std_logic; attribute dont_touch of I33813: signal is true;
	signal I33816: std_logic; attribute dont_touch of I33816: signal is true;
	signal I33819: std_logic; attribute dont_touch of I33819: signal is true;
	signal I33822: std_logic; attribute dont_touch of I33822: signal is true;
	signal I33825: std_logic; attribute dont_touch of I33825: signal is true;
	signal I33828: std_logic; attribute dont_touch of I33828: signal is true;
	signal I33831: std_logic; attribute dont_touch of I33831: signal is true;
	signal I33834: std_logic; attribute dont_touch of I33834: signal is true;
	signal I33837: std_logic; attribute dont_touch of I33837: signal is true;
	signal I33840: std_logic; attribute dont_touch of I33840: signal is true;
	signal I33843: std_logic; attribute dont_touch of I33843: signal is true;
	signal I33846: std_logic; attribute dont_touch of I33846: signal is true;
	signal I33849: std_logic; attribute dont_touch of I33849: signal is true;
	signal I33852: std_logic; attribute dont_touch of I33852: signal is true;
	signal I33855: std_logic; attribute dont_touch of I33855: signal is true;
	signal I33858: std_logic; attribute dont_touch of I33858: signal is true;
	signal I33861: std_logic; attribute dont_touch of I33861: signal is true;
	signal I33864: std_logic; attribute dont_touch of I33864: signal is true;
	signal I33867: std_logic; attribute dont_touch of I33867: signal is true;
	signal I33870: std_logic; attribute dont_touch of I33870: signal is true;
	signal I33873: std_logic; attribute dont_touch of I33873: signal is true;
	signal I33876: std_logic; attribute dont_touch of I33876: signal is true;
	signal I33879: std_logic; attribute dont_touch of I33879: signal is true;
	signal I33882: std_logic; attribute dont_touch of I33882: signal is true;
	signal I33885: std_logic; attribute dont_touch of I33885: signal is true;
	signal I33888: std_logic; attribute dont_touch of I33888: signal is true;
	signal I33891: std_logic; attribute dont_touch of I33891: signal is true;
	signal I33894: std_logic; attribute dont_touch of I33894: signal is true;
	signal I33897: std_logic; attribute dont_touch of I33897: signal is true;
	signal I33900: std_logic; attribute dont_touch of I33900: signal is true;
	signal I33903: std_logic; attribute dont_touch of I33903: signal is true;
	signal I33906: std_logic; attribute dont_touch of I33906: signal is true;
	signal I33909: std_logic; attribute dont_touch of I33909: signal is true;
	signal I33912: std_logic; attribute dont_touch of I33912: signal is true;
	signal I33915: std_logic; attribute dont_touch of I33915: signal is true;
	signal I33918: std_logic; attribute dont_touch of I33918: signal is true;
	signal I33954: std_logic; attribute dont_touch of I33954: signal is true;
	signal I33961: std_logic; attribute dont_touch of I33961: signal is true;
	signal I33968: std_logic; attribute dont_touch of I33968: signal is true;
	signal I33974: std_logic; attribute dont_touch of I33974: signal is true;
	signal I33984: std_logic; attribute dont_touch of I33984: signal is true;
	signal I33990: std_logic; attribute dont_touch of I33990: signal is true;
	signal I33995: std_logic; attribute dont_touch of I33995: signal is true;
	signal I33999: std_logic; attribute dont_touch of I33999: signal is true;
	signal I34002: std_logic; attribute dont_touch of I34002: signal is true;
	signal I34009: std_logic; attribute dont_touch of I34009: signal is true;
	signal I34012: std_logic; attribute dont_touch of I34012: signal is true;
	signal I34017: std_logic; attribute dont_touch of I34017: signal is true;
	signal I34020: std_logic; attribute dont_touch of I34020: signal is true;
	signal I34026: std_logic; attribute dont_touch of I34026: signal is true;
	signal I34029: std_logic; attribute dont_touch of I34029: signal is true;
	signal I34032: std_logic; attribute dont_touch of I34032: signal is true;
	signal I34041: std_logic; attribute dont_touch of I34041: signal is true;
	signal I34044: std_logic; attribute dont_touch of I34044: signal is true;
	signal I34051: std_logic; attribute dont_touch of I34051: signal is true;
	signal I34056: std_logic; attribute dont_touch of I34056: signal is true;
	signal I34059: std_logic; attribute dont_touch of I34059: signal is true;
	signal I34063: std_logic; attribute dont_touch of I34063: signal is true;
	signal I34068: std_logic; attribute dont_touch of I34068: signal is true;
	signal I34071: std_logic; attribute dont_touch of I34071: signal is true;
	signal I34074: std_logic; attribute dont_touch of I34074: signal is true;
	signal I34077: std_logic; attribute dont_touch of I34077: signal is true;
	signal I34080: std_logic; attribute dont_touch of I34080: signal is true;
	signal I34083: std_logic; attribute dont_touch of I34083: signal is true;
	signal I34086: std_logic; attribute dont_touch of I34086: signal is true;
	signal I34091: std_logic; attribute dont_touch of I34091: signal is true;
	signal I34096: std_logic; attribute dont_touch of I34096: signal is true;
	signal I34099: std_logic; attribute dont_touch of I34099: signal is true;
	signal I34102: std_logic; attribute dont_touch of I34102: signal is true;
	signal I34105: std_logic; attribute dont_touch of I34105: signal is true;
	signal I34108: std_logic; attribute dont_touch of I34108: signal is true;
	signal I34111: std_logic; attribute dont_touch of I34111: signal is true;
	signal I34114: std_logic; attribute dont_touch of I34114: signal is true;
	signal I34118: std_logic; attribute dont_touch of I34118: signal is true;
	signal I34121: std_logic; attribute dont_touch of I34121: signal is true;
	signal I34124: std_logic; attribute dont_touch of I34124: signal is true;
	signal I34128: std_logic; attribute dont_touch of I34128: signal is true;
	signal I34132: std_logic; attribute dont_touch of I34132: signal is true;
	signal I34135: std_logic; attribute dont_touch of I34135: signal is true;
	signal I34140: std_logic; attribute dont_touch of I34140: signal is true;
	signal I34143: std_logic; attribute dont_touch of I34143: signal is true;
	signal I34146: std_logic; attribute dont_touch of I34146: signal is true;
	signal I34150: std_logic; attribute dont_touch of I34150: signal is true;
	signal I34153: std_logic; attribute dont_touch of I34153: signal is true;
	signal I34156: std_logic; attribute dont_touch of I34156: signal is true;
	signal I34159: std_logic; attribute dont_touch of I34159: signal is true;
	signal I34162: std_logic; attribute dont_touch of I34162: signal is true;
	signal I34165: std_logic; attribute dont_touch of I34165: signal is true;
	signal I34168: std_logic; attribute dont_touch of I34168: signal is true;
	signal I34172: std_logic; attribute dont_touch of I34172: signal is true;
	signal I34180: std_logic; attribute dont_touch of I34180: signal is true;
	signal I34183: std_logic; attribute dont_touch of I34183: signal is true;
	signal I34189: std_logic; attribute dont_touch of I34189: signal is true;
	signal I34192: std_logic; attribute dont_touch of I34192: signal is true;
	signal I34195: std_logic; attribute dont_touch of I34195: signal is true;
	signal I34198: std_logic; attribute dont_touch of I34198: signal is true;
	signal I34201: std_logic; attribute dont_touch of I34201: signal is true;
	signal I34204: std_logic; attribute dont_touch of I34204: signal is true;
	signal I34207: std_logic; attribute dont_touch of I34207: signal is true;
	signal I34210: std_logic; attribute dont_touch of I34210: signal is true;
	signal I34220: std_logic; attribute dont_touch of I34220: signal is true;
	signal I34230: std_logic; attribute dont_touch of I34230: signal is true;
	signal I34233: std_logic; attribute dont_touch of I34233: signal is true;
	signal I34238: std_logic; attribute dont_touch of I34238: signal is true;
	signal I34241: std_logic; attribute dont_touch of I34241: signal is true;
	signal I34244: std_logic; attribute dont_touch of I34244: signal is true;
	signal I34254: std_logic; attribute dont_touch of I34254: signal is true;
	signal I34266: std_logic; attribute dont_touch of I34266: signal is true;
	signal I34274: std_logic; attribute dont_touch of I34274: signal is true;
	signal I34277: std_logic; attribute dont_touch of I34277: signal is true;
	signal I34296: std_logic; attribute dont_touch of I34296: signal is true;
	signal I34306: std_logic; attribute dont_touch of I34306: signal is true;
	signal I34313: std_logic; attribute dont_touch of I34313: signal is true;
	signal I34316: std_logic; attribute dont_touch of I34316: signal is true;
	signal I34321: std_logic; attribute dont_touch of I34321: signal is true;
	signal I34327: std_logic; attribute dont_touch of I34327: signal is true;
	signal I34343: std_logic; attribute dont_touch of I34343: signal is true;
	signal I34353: std_logic; attribute dont_touch of I34353: signal is true;
	signal I34358: std_logic; attribute dont_touch of I34358: signal is true;
	signal I34363: std_logic; attribute dont_touch of I34363: signal is true;
	signal I34369: std_logic; attribute dont_touch of I34369: signal is true;
	signal I34385: std_logic; attribute dont_touch of I34385: signal is true;
	signal I34388: std_logic; attribute dont_touch of I34388: signal is true;
	signal I34392: std_logic; attribute dont_touch of I34392: signal is true;
	signal I34395: std_logic; attribute dont_touch of I34395: signal is true;
	signal I34400: std_logic; attribute dont_touch of I34400: signal is true;
	signal I34405: std_logic; attribute dont_touch of I34405: signal is true;
	signal I34411: std_logic; attribute dont_touch of I34411: signal is true;
	signal I34421: std_logic; attribute dont_touch of I34421: signal is true;
	signal I34425: std_logic; attribute dont_touch of I34425: signal is true;
	signal I34428: std_logic; attribute dont_touch of I34428: signal is true;
	signal I34433: std_logic; attribute dont_touch of I34433: signal is true;
	signal I34438: std_logic; attribute dont_touch of I34438: signal is true;
	signal I34444: std_logic; attribute dont_touch of I34444: signal is true;
	signal I34449: std_logic; attribute dont_touch of I34449: signal is true;
	signal I34453: std_logic; attribute dont_touch of I34453: signal is true;
	signal I34456: std_logic; attribute dont_touch of I34456: signal is true;
	signal I34461: std_logic; attribute dont_touch of I34461: signal is true;
	signal I34464: std_logic; attribute dont_touch of I34464: signal is true;
	signal I34469: std_logic; attribute dont_touch of I34469: signal is true;
	signal I34473: std_logic; attribute dont_touch of I34473: signal is true;
	signal I34476: std_logic; attribute dont_touch of I34476: signal is true;
	signal I34479: std_logic; attribute dont_touch of I34479: signal is true;
	signal I34505: std_logic; attribute dont_touch of I34505: signal is true;
	signal I34535: std_logic; attribute dont_touch of I34535: signal is true;
	signal I34579: std_logic; attribute dont_touch of I34579: signal is true;
	signal I34641: std_logic; attribute dont_touch of I34641: signal is true;
	signal I34644: std_logic; attribute dont_touch of I34644: signal is true;
	signal I34647: std_logic; attribute dont_touch of I34647: signal is true;
	signal I34650: std_logic; attribute dont_touch of I34650: signal is true;
	signal I34653: std_logic; attribute dont_touch of I34653: signal is true;
	signal I34656: std_logic; attribute dont_touch of I34656: signal is true;
	signal I34659: std_logic; attribute dont_touch of I34659: signal is true;
	signal I34662: std_logic; attribute dont_touch of I34662: signal is true;
	signal I34665: std_logic; attribute dont_touch of I34665: signal is true;
	signal I34668: std_logic; attribute dont_touch of I34668: signal is true;
	signal I34671: std_logic; attribute dont_touch of I34671: signal is true;
	signal I34674: std_logic; attribute dont_touch of I34674: signal is true;
	signal I34677: std_logic; attribute dont_touch of I34677: signal is true;
	signal I34680: std_logic; attribute dont_touch of I34680: signal is true;
	signal I34683: std_logic; attribute dont_touch of I34683: signal is true;
	signal I34686: std_logic; attribute dont_touch of I34686: signal is true;
	signal I34689: std_logic; attribute dont_touch of I34689: signal is true;
	signal I34692: std_logic; attribute dont_touch of I34692: signal is true;
	signal I34695: std_logic; attribute dont_touch of I34695: signal is true;
	signal I34698: std_logic; attribute dont_touch of I34698: signal is true;
	signal I34701: std_logic; attribute dont_touch of I34701: signal is true;
	signal I34704: std_logic; attribute dont_touch of I34704: signal is true;
	signal I34707: std_logic; attribute dont_touch of I34707: signal is true;
	signal I34710: std_logic; attribute dont_touch of I34710: signal is true;
	signal I34713: std_logic; attribute dont_touch of I34713: signal is true;
	signal I34716: std_logic; attribute dont_touch of I34716: signal is true;
	signal I34719: std_logic; attribute dont_touch of I34719: signal is true;
	signal I34722: std_logic; attribute dont_touch of I34722: signal is true;
	signal I34725: std_logic; attribute dont_touch of I34725: signal is true;
	signal I34728: std_logic; attribute dont_touch of I34728: signal is true;
	signal I34731: std_logic; attribute dont_touch of I34731: signal is true;
	signal I34734: std_logic; attribute dont_touch of I34734: signal is true;
	signal I34737: std_logic; attribute dont_touch of I34737: signal is true;
	signal I34740: std_logic; attribute dont_touch of I34740: signal is true;
	signal I34743: std_logic; attribute dont_touch of I34743: signal is true;
	signal I34746: std_logic; attribute dont_touch of I34746: signal is true;
	signal I34749: std_logic; attribute dont_touch of I34749: signal is true;
	signal I34752: std_logic; attribute dont_touch of I34752: signal is true;
	signal I34755: std_logic; attribute dont_touch of I34755: signal is true;
	signal I34758: std_logic; attribute dont_touch of I34758: signal is true;
	signal I34761: std_logic; attribute dont_touch of I34761: signal is true;
	signal I34764: std_logic; attribute dont_touch of I34764: signal is true;
	signal I34767: std_logic; attribute dont_touch of I34767: signal is true;
	signal I34770: std_logic; attribute dont_touch of I34770: signal is true;
	signal I34773: std_logic; attribute dont_touch of I34773: signal is true;
	signal I34776: std_logic; attribute dont_touch of I34776: signal is true;
	signal I34779: std_logic; attribute dont_touch of I34779: signal is true;
	signal I34782: std_logic; attribute dont_touch of I34782: signal is true;
	signal I34785: std_logic; attribute dont_touch of I34785: signal is true;
	signal I34788: std_logic; attribute dont_touch of I34788: signal is true;
	signal I34791: std_logic; attribute dont_touch of I34791: signal is true;
	signal I34794: std_logic; attribute dont_touch of I34794: signal is true;
	signal I34797: std_logic; attribute dont_touch of I34797: signal is true;
	signal I34800: std_logic; attribute dont_touch of I34800: signal is true;
	signal I34803: std_logic; attribute dont_touch of I34803: signal is true;
	signal I34806: std_logic; attribute dont_touch of I34806: signal is true;
	signal I34809: std_logic; attribute dont_touch of I34809: signal is true;
	signal I34812: std_logic; attribute dont_touch of I34812: signal is true;
	signal I34815: std_logic; attribute dont_touch of I34815: signal is true;
	signal I34818: std_logic; attribute dont_touch of I34818: signal is true;
	signal I34821: std_logic; attribute dont_touch of I34821: signal is true;
	signal I34824: std_logic; attribute dont_touch of I34824: signal is true;
	signal I34827: std_logic; attribute dont_touch of I34827: signal is true;
	signal I34830: std_logic; attribute dont_touch of I34830: signal is true;
	signal I34833: std_logic; attribute dont_touch of I34833: signal is true;
	signal I34836: std_logic; attribute dont_touch of I34836: signal is true;
	signal I34839: std_logic; attribute dont_touch of I34839: signal is true;
	signal I34842: std_logic; attribute dont_touch of I34842: signal is true;
	signal I34845: std_logic; attribute dont_touch of I34845: signal is true;
	signal I34848: std_logic; attribute dont_touch of I34848: signal is true;
	signal I34851: std_logic; attribute dont_touch of I34851: signal is true;
	signal I34854: std_logic; attribute dont_touch of I34854: signal is true;
	signal I34857: std_logic; attribute dont_touch of I34857: signal is true;
	signal I34860: std_logic; attribute dont_touch of I34860: signal is true;
	signal I34863: std_logic; attribute dont_touch of I34863: signal is true;
	signal I34866: std_logic; attribute dont_touch of I34866: signal is true;
	signal I34872: std_logic; attribute dont_touch of I34872: signal is true;
	signal I34879: std_logic; attribute dont_touch of I34879: signal is true;
	signal I34901: std_logic; attribute dont_touch of I34901: signal is true;
	signal I34909: std_logic; attribute dont_touch of I34909: signal is true;
	signal I34916: std_logic; attribute dont_touch of I34916: signal is true;
	signal I34921: std_logic; attribute dont_touch of I34921: signal is true;
	signal I34946: std_logic; attribute dont_touch of I34946: signal is true;
	signal I34957: std_logic; attribute dont_touch of I34957: signal is true;
	signal I34961: std_logic; attribute dont_touch of I34961: signal is true;
	signal I34964: std_logic; attribute dont_touch of I34964: signal is true;
	signal I34967: std_logic; attribute dont_touch of I34967: signal is true;
	signal I34971: std_logic; attribute dont_touch of I34971: signal is true;
	signal I34974: std_logic; attribute dont_touch of I34974: signal is true;
	signal I34977: std_logic; attribute dont_touch of I34977: signal is true;
	signal I34980: std_logic; attribute dont_touch of I34980: signal is true;
	signal I34983: std_logic; attribute dont_touch of I34983: signal is true;
	signal I34986: std_logic; attribute dont_touch of I34986: signal is true;
	signal I34990: std_logic; attribute dont_touch of I34990: signal is true;
	signal I34993: std_logic; attribute dont_touch of I34993: signal is true;
	signal I34997: std_logic; attribute dont_touch of I34997: signal is true;
	signal I35000: std_logic; attribute dont_touch of I35000: signal is true;
	signal I35003: std_logic; attribute dont_touch of I35003: signal is true;
	signal I35007: std_logic; attribute dont_touch of I35007: signal is true;
	signal I35011: std_logic; attribute dont_touch of I35011: signal is true;
	signal I35014: std_logic; attribute dont_touch of I35014: signal is true;
	signal I35017: std_logic; attribute dont_touch of I35017: signal is true;
	signal I35020: std_logic; attribute dont_touch of I35020: signal is true;
	signal I35021: std_logic; attribute dont_touch of I35021: signal is true;
	signal I35022: std_logic; attribute dont_touch of I35022: signal is true;
	signal I35028: std_logic; attribute dont_touch of I35028: signal is true;
	signal I35031: std_logic; attribute dont_touch of I35031: signal is true;
	signal I35034: std_logic; attribute dont_touch of I35034: signal is true;
	signal I35035: std_logic; attribute dont_touch of I35035: signal is true;
	signal I35036: std_logic; attribute dont_touch of I35036: signal is true;
	signal I35042: std_logic; attribute dont_touch of I35042: signal is true;
	signal I35043: std_logic; attribute dont_touch of I35043: signal is true;
	signal I35044: std_logic; attribute dont_touch of I35044: signal is true;
	signal I35049: std_logic; attribute dont_touch of I35049: signal is true;
	signal I35053: std_logic; attribute dont_touch of I35053: signal is true;
	signal I35057: std_logic; attribute dont_touch of I35057: signal is true;
	signal I35058: std_logic; attribute dont_touch of I35058: signal is true;
	signal I35059: std_logic; attribute dont_touch of I35059: signal is true;
	signal I35064: std_logic; attribute dont_touch of I35064: signal is true;
	signal I35067: std_logic; attribute dont_touch of I35067: signal is true;
	signal I35072: std_logic; attribute dont_touch of I35072: signal is true;
	signal I35076: std_logic; attribute dont_touch of I35076: signal is true;
	signal I35079: std_logic; attribute dont_touch of I35079: signal is true;
	signal I35083: std_logic; attribute dont_touch of I35083: signal is true;
	signal I35087: std_logic; attribute dont_touch of I35087: signal is true;
	signal I35092: std_logic; attribute dont_touch of I35092: signal is true;
	signal I35095: std_logic; attribute dont_touch of I35095: signal is true;
	signal I35099: std_logic; attribute dont_touch of I35099: signal is true;
	signal I35106: std_logic; attribute dont_touch of I35106: signal is true;
	signal I35109: std_logic; attribute dont_touch of I35109: signal is true;
	signal I35116: std_logic; attribute dont_touch of I35116: signal is true;
	signal I35123: std_logic; attribute dont_touch of I35123: signal is true;
	signal I35124: std_logic; attribute dont_touch of I35124: signal is true;
	signal I35125: std_logic; attribute dont_touch of I35125: signal is true;
	signal I35136: std_logic; attribute dont_touch of I35136: signal is true;
	signal I35141: std_logic; attribute dont_touch of I35141: signal is true;
	signal I35146: std_logic; attribute dont_touch of I35146: signal is true;
	signal I35153: std_logic; attribute dont_touch of I35153: signal is true;
	signal I35172: std_logic; attribute dont_touch of I35172: signal is true;
	signal I35254: std_logic; attribute dont_touch of I35254: signal is true;
	signal I35283: std_logic; attribute dont_touch of I35283: signal is true;
	signal I35297: std_logic; attribute dont_touch of I35297: signal is true;
	signal I35301: std_logic; attribute dont_touch of I35301: signal is true;
	signal I35313: std_logic; attribute dont_touch of I35313: signal is true;
	signal I35319: std_logic; attribute dont_touch of I35319: signal is true;
	signal I35334: std_logic; attribute dont_touch of I35334: signal is true;
	signal I35341: std_logic; attribute dont_touch of I35341: signal is true;
	signal I35347: std_logic; attribute dont_touch of I35347: signal is true;
	signal I35351: std_logic; attribute dont_touch of I35351: signal is true;
	signal I35355: std_logic; attribute dont_touch of I35355: signal is true;
	signal I35360: std_logic; attribute dont_touch of I35360: signal is true;
	signal I35364: std_logic; attribute dont_touch of I35364: signal is true;
	signal I35369: std_logic; attribute dont_touch of I35369: signal is true;
	signal I35373: std_logic; attribute dont_touch of I35373: signal is true;
	signal I35376: std_logic; attribute dont_touch of I35376: signal is true;
	signal I35383: std_logic; attribute dont_touch of I35383: signal is true;
	signal I35389: std_logic; attribute dont_touch of I35389: signal is true;
	signal I35394: std_logic; attribute dont_touch of I35394: signal is true;
	signal I35399: std_logic; attribute dont_touch of I35399: signal is true;
	signal I35404: std_logic; attribute dont_touch of I35404: signal is true;
	signal I35407: std_logic; attribute dont_touch of I35407: signal is true;
	signal I35410: std_logic; attribute dont_touch of I35410: signal is true;
	signal I35413: std_logic; attribute dont_touch of I35413: signal is true;
	signal I35416: std_logic; attribute dont_touch of I35416: signal is true;
	signal I35419: std_logic; attribute dont_touch of I35419: signal is true;
	signal I35422: std_logic; attribute dont_touch of I35422: signal is true;
	signal I35425: std_logic; attribute dont_touch of I35425: signal is true;
	signal I35428: std_logic; attribute dont_touch of I35428: signal is true;
	signal I35431: std_logic; attribute dont_touch of I35431: signal is true;
	signal I35434: std_logic; attribute dont_touch of I35434: signal is true;
	signal I35437: std_logic; attribute dont_touch of I35437: signal is true;
	signal I35440: std_logic; attribute dont_touch of I35440: signal is true;
	signal I35443: std_logic; attribute dont_touch of I35443: signal is true;
	signal I35446: std_logic; attribute dont_touch of I35446: signal is true;
	signal I35449: std_logic; attribute dont_touch of I35449: signal is true;
	signal I35452: std_logic; attribute dont_touch of I35452: signal is true;
	signal I35455: std_logic; attribute dont_touch of I35455: signal is true;
	signal I35458: std_logic; attribute dont_touch of I35458: signal is true;
	signal I35461: std_logic; attribute dont_touch of I35461: signal is true;
	signal I35464: std_logic; attribute dont_touch of I35464: signal is true;
	signal I35467: std_logic; attribute dont_touch of I35467: signal is true;
	signal I35470: std_logic; attribute dont_touch of I35470: signal is true;
	signal I35473: std_logic; attribute dont_touch of I35473: signal is true;
	signal I35476: std_logic; attribute dont_touch of I35476: signal is true;
	signal I35479: std_logic; attribute dont_touch of I35479: signal is true;
	signal I35482: std_logic; attribute dont_touch of I35482: signal is true;
	signal I35485: std_logic; attribute dont_touch of I35485: signal is true;
	signal I35488: std_logic; attribute dont_touch of I35488: signal is true;
	signal I35491: std_logic; attribute dont_touch of I35491: signal is true;
	signal I35494: std_logic; attribute dont_touch of I35494: signal is true;
	signal I35497: std_logic; attribute dont_touch of I35497: signal is true;
	signal I35500: std_logic; attribute dont_touch of I35500: signal is true;
	signal I35503: std_logic; attribute dont_touch of I35503: signal is true;
	signal I35506: std_logic; attribute dont_touch of I35506: signal is true;
	signal I35509: std_logic; attribute dont_touch of I35509: signal is true;
	signal I35512: std_logic; attribute dont_touch of I35512: signal is true;
	signal I35515: std_logic; attribute dont_touch of I35515: signal is true;
	signal I35518: std_logic; attribute dont_touch of I35518: signal is true;
	signal I35521: std_logic; attribute dont_touch of I35521: signal is true;
	signal I35524: std_logic; attribute dont_touch of I35524: signal is true;
	signal I35527: std_logic; attribute dont_touch of I35527: signal is true;
	signal I35530: std_logic; attribute dont_touch of I35530: signal is true;
	signal I35533: std_logic; attribute dont_touch of I35533: signal is true;
	signal I35536: std_logic; attribute dont_touch of I35536: signal is true;
	signal I35539: std_logic; attribute dont_touch of I35539: signal is true;
	signal I35542: std_logic; attribute dont_touch of I35542: signal is true;
	signal I35545: std_logic; attribute dont_touch of I35545: signal is true;
	signal I35548: std_logic; attribute dont_touch of I35548: signal is true;
	signal I35551: std_logic; attribute dont_touch of I35551: signal is true;
	signal I35554: std_logic; attribute dont_touch of I35554: signal is true;
	signal I35667: std_logic; attribute dont_touch of I35667: signal is true;
	signal I35673: std_logic; attribute dont_touch of I35673: signal is true;
	signal I35678: std_logic; attribute dont_touch of I35678: signal is true;
	signal I35681: std_logic; attribute dont_touch of I35681: signal is true;
	signal I35686: std_logic; attribute dont_touch of I35686: signal is true;
	signal I35689: std_logic; attribute dont_touch of I35689: signal is true;
	signal I35695: std_logic; attribute dont_touch of I35695: signal is true;
	signal I35698: std_logic; attribute dont_touch of I35698: signal is true;
	signal I35701: std_logic; attribute dont_touch of I35701: signal is true;
	signal I35702: std_logic; attribute dont_touch of I35702: signal is true;
	signal I35703: std_logic; attribute dont_touch of I35703: signal is true;
	signal I35708: std_logic; attribute dont_touch of I35708: signal is true;
	signal I35711: std_logic; attribute dont_touch of I35711: signal is true;
	signal I35714: std_logic; attribute dont_touch of I35714: signal is true;
	signal I35715: std_logic; attribute dont_touch of I35715: signal is true;
	signal I35716: std_logic; attribute dont_touch of I35716: signal is true;
	signal I35723: std_logic; attribute dont_touch of I35723: signal is true;
	signal I35727: std_logic; attribute dont_touch of I35727: signal is true;
	signal I35731: std_logic; attribute dont_touch of I35731: signal is true;
	signal I35737: std_logic; attribute dont_touch of I35737: signal is true;
	signal I35741: std_logic; attribute dont_touch of I35741: signal is true;
	signal I35744: std_logic; attribute dont_touch of I35744: signal is true;
	signal I35750: std_logic; attribute dont_touch of I35750: signal is true;
	signal I35756: std_logic; attribute dont_touch of I35756: signal is true;
	signal I35759: std_logic; attribute dont_touch of I35759: signal is true;
	signal I35762: std_logic; attribute dont_touch of I35762: signal is true;
	signal I35768: std_logic; attribute dont_touch of I35768: signal is true;
	signal I35772: std_logic; attribute dont_touch of I35772: signal is true;
	signal I35777: std_logic; attribute dont_touch of I35777: signal is true;
	signal I35780: std_logic; attribute dont_touch of I35780: signal is true;
	signal I35783: std_logic; attribute dont_touch of I35783: signal is true;
	signal I35791: std_logic; attribute dont_touch of I35791: signal is true;
	signal I35796: std_logic; attribute dont_touch of I35796: signal is true;
	signal I35799: std_logic; attribute dont_touch of I35799: signal is true;
	signal I35803: std_logic; attribute dont_touch of I35803: signal is true;
	signal I35809: std_logic; attribute dont_touch of I35809: signal is true;
	signal I35814: std_logic; attribute dont_touch of I35814: signal is true;
	signal I35817: std_logic; attribute dont_touch of I35817: signal is true;
	signal I35821: std_logic; attribute dont_touch of I35821: signal is true;
	signal I35824: std_logic; attribute dont_touch of I35824: signal is true;
	signal I35829: std_logic; attribute dont_touch of I35829: signal is true;
	signal I35834: std_logic; attribute dont_touch of I35834: signal is true;
	signal I35837: std_logic; attribute dont_touch of I35837: signal is true;
	signal I35841: std_logic; attribute dont_touch of I35841: signal is true;
	signal I35844: std_logic; attribute dont_touch of I35844: signal is true;
	signal I35849: std_logic; attribute dont_touch of I35849: signal is true;
	signal I35852: std_logic; attribute dont_touch of I35852: signal is true;
	signal I35856: std_logic; attribute dont_touch of I35856: signal is true;
	signal I35859: std_logic; attribute dont_touch of I35859: signal is true;
	signal I35863: std_logic; attribute dont_touch of I35863: signal is true;
	signal I35868: std_logic; attribute dont_touch of I35868: signal is true;
	signal I35872: std_logic; attribute dont_touch of I35872: signal is true;
	signal I35876: std_logic; attribute dont_touch of I35876: signal is true;
	signal I35879: std_logic; attribute dont_touch of I35879: signal is true;
	signal I35883: std_logic; attribute dont_touch of I35883: signal is true;
	signal I35886: std_logic; attribute dont_touch of I35886: signal is true;
	signal I35890: std_logic; attribute dont_touch of I35890: signal is true;
	signal I35893: std_logic; attribute dont_touch of I35893: signal is true;
	signal I35897: std_logic; attribute dont_touch of I35897: signal is true;
	signal I35900: std_logic; attribute dont_touch of I35900: signal is true;
	signal I35904: std_logic; attribute dont_touch of I35904: signal is true;
	signal I35905: std_logic; attribute dont_touch of I35905: signal is true;
	signal I35906: std_logic; attribute dont_touch of I35906: signal is true;
	signal I35915: std_logic; attribute dont_touch of I35915: signal is true;
	signal I35919: std_logic; attribute dont_touch of I35919: signal is true;
	signal I35923: std_logic; attribute dont_touch of I35923: signal is true;
	signal I35926: std_logic; attribute dont_touch of I35926: signal is true;
	signal I35930: std_logic; attribute dont_touch of I35930: signal is true;
	signal I35933: std_logic; attribute dont_touch of I35933: signal is true;
	signal I35937: std_logic; attribute dont_touch of I35937: signal is true;
	signal I35940: std_logic; attribute dont_touch of I35940: signal is true;
	signal I35944: std_logic; attribute dont_touch of I35944: signal is true;
	signal I35945: std_logic; attribute dont_touch of I35945: signal is true;
	signal I35946: std_logic; attribute dont_touch of I35946: signal is true;
	signal I35953: std_logic; attribute dont_touch of I35953: signal is true;
	signal I35957: std_logic; attribute dont_touch of I35957: signal is true;
	signal I35961: std_logic; attribute dont_touch of I35961: signal is true;
	signal I35964: std_logic; attribute dont_touch of I35964: signal is true;
	signal I35968: std_logic; attribute dont_touch of I35968: signal is true;
	signal I35974: std_logic; attribute dont_touch of I35974: signal is true;
	signal I35975: std_logic; attribute dont_touch of I35975: signal is true;
	signal I35976: std_logic; attribute dont_touch of I35976: signal is true;
	signal I35983: std_logic; attribute dont_touch of I35983: signal is true;
	signal I35992: std_logic; attribute dont_touch of I35992: signal is true;
	signal I35993: std_logic; attribute dont_touch of I35993: signal is true;
	signal I35994: std_logic; attribute dont_touch of I35994: signal is true;
	signal I36008: std_logic; attribute dont_touch of I36008: signal is true;
	signal I36032: std_logic; attribute dont_touch of I36032: signal is true;
	signal I36042: std_logic; attribute dont_touch of I36042: signal is true;
	signal I36046: std_logic; attribute dont_touch of I36046: signal is true;
	signal I36052: std_logic; attribute dont_touch of I36052: signal is true;
	signal I36060: std_logic; attribute dont_touch of I36060: signal is true;
	signal I36063: std_logic; attribute dont_touch of I36063: signal is true;
	signal I36066: std_logic; attribute dont_touch of I36066: signal is true;
	signal I36069: std_logic; attribute dont_touch of I36069: signal is true;
	signal I36072: std_logic; attribute dont_touch of I36072: signal is true;
	signal I36075: std_logic; attribute dont_touch of I36075: signal is true;
	signal I36078: std_logic; attribute dont_touch of I36078: signal is true;
	signal I36081: std_logic; attribute dont_touch of I36081: signal is true;
	signal I36084: std_logic; attribute dont_touch of I36084: signal is true;
	signal I36087: std_logic; attribute dont_touch of I36087: signal is true;
	signal I36090: std_logic; attribute dont_touch of I36090: signal is true;
	signal I36093: std_logic; attribute dont_touch of I36093: signal is true;
	signal I36096: std_logic; attribute dont_touch of I36096: signal is true;
	signal I36099: std_logic; attribute dont_touch of I36099: signal is true;
	signal I36102: std_logic; attribute dont_touch of I36102: signal is true;
	signal I36105: std_logic; attribute dont_touch of I36105: signal is true;
	signal I36108: std_logic; attribute dont_touch of I36108: signal is true;
	signal I36111: std_logic; attribute dont_touch of I36111: signal is true;
	signal I36114: std_logic; attribute dont_touch of I36114: signal is true;
	signal I36117: std_logic; attribute dont_touch of I36117: signal is true;
	signal I36120: std_logic; attribute dont_touch of I36120: signal is true;
	signal I36123: std_logic; attribute dont_touch of I36123: signal is true;
	signal I36126: std_logic; attribute dont_touch of I36126: signal is true;
	signal I36129: std_logic; attribute dont_touch of I36129: signal is true;
	signal I36132: std_logic; attribute dont_touch of I36132: signal is true;
	signal I36135: std_logic; attribute dont_touch of I36135: signal is true;
	signal I36138: std_logic; attribute dont_touch of I36138: signal is true;
	signal I36141: std_logic; attribute dont_touch of I36141: signal is true;
	signal I36144: std_logic; attribute dont_touch of I36144: signal is true;
	signal I36147: std_logic; attribute dont_touch of I36147: signal is true;
	signal I36150: std_logic; attribute dont_touch of I36150: signal is true;
	signal I36153: std_logic; attribute dont_touch of I36153: signal is true;
	signal I36156: std_logic; attribute dont_touch of I36156: signal is true;
	signal I36159: std_logic; attribute dont_touch of I36159: signal is true;
	signal I36162: std_logic; attribute dont_touch of I36162: signal is true;
	signal I36213: std_logic; attribute dont_touch of I36213: signal is true;
	signal I36217: std_logic; attribute dont_touch of I36217: signal is true;
	signal I36221: std_logic; attribute dont_touch of I36221: signal is true;
	signal I36224: std_logic; attribute dont_touch of I36224: signal is true;
	signal I36227: std_logic; attribute dont_touch of I36227: signal is true;
	signal I36230: std_logic; attribute dont_touch of I36230: signal is true;
	signal I36234: std_logic; attribute dont_touch of I36234: signal is true;
	signal I36237: std_logic; attribute dont_touch of I36237: signal is true;
	signal I36240: std_logic; attribute dont_touch of I36240: signal is true;
	signal I36243: std_logic; attribute dont_touch of I36243: signal is true;
	signal I36246: std_logic; attribute dont_touch of I36246: signal is true;
	signal I36250: std_logic; attribute dont_touch of I36250: signal is true;
	signal I36253: std_logic; attribute dont_touch of I36253: signal is true;
	signal I36256: std_logic; attribute dont_touch of I36256: signal is true;
	signal I36257: std_logic; attribute dont_touch of I36257: signal is true;
	signal I36258: std_logic; attribute dont_touch of I36258: signal is true;
	signal I36264: std_logic; attribute dont_touch of I36264: signal is true;
	signal I36267: std_logic; attribute dont_touch of I36267: signal is true;
	signal I36270: std_logic; attribute dont_touch of I36270: signal is true;
	signal I36271: std_logic; attribute dont_touch of I36271: signal is true;
	signal I36272: std_logic; attribute dont_touch of I36272: signal is true;
	signal I36280: std_logic; attribute dont_touch of I36280: signal is true;
	signal I36283: std_logic; attribute dont_touch of I36283: signal is true;
	signal I36289: std_logic; attribute dont_touch of I36289: signal is true;
	signal I36290: std_logic; attribute dont_touch of I36290: signal is true;
	signal I36291: std_logic; attribute dont_touch of I36291: signal is true;
	signal I36296: std_logic; attribute dont_touch of I36296: signal is true;
	signal I36300: std_logic; attribute dont_touch of I36300: signal is true;
	signal I36301: std_logic; attribute dont_touch of I36301: signal is true;
	signal I36302: std_logic; attribute dont_touch of I36302: signal is true;
	signal I36307: std_logic; attribute dont_touch of I36307: signal is true;
	signal I36311: std_logic; attribute dont_touch of I36311: signal is true;
	signal I36314: std_logic; attribute dont_touch of I36314: signal is true;
	signal I36315: std_logic; attribute dont_touch of I36315: signal is true;
	signal I36316: std_logic; attribute dont_touch of I36316: signal is true;
	signal I36321: std_logic; attribute dont_touch of I36321: signal is true;
	signal I36327: std_logic; attribute dont_touch of I36327: signal is true;
	signal I36330: std_logic; attribute dont_touch of I36330: signal is true;
	signal I36337: std_logic; attribute dont_touch of I36337: signal is true;
	signal I36341: std_logic; attribute dont_touch of I36341: signal is true;
	signal I36347: std_logic; attribute dont_touch of I36347: signal is true;
	signal I36354: std_logic; attribute dont_touch of I36354: signal is true;
	signal I36358: std_logic; attribute dont_touch of I36358: signal is true;
	signal I36362: std_logic; attribute dont_touch of I36362: signal is true;
	signal I36367: std_logic; attribute dont_touch of I36367: signal is true;
	signal I36371: std_logic; attribute dont_touch of I36371: signal is true;
	signal I36379: std_logic; attribute dont_touch of I36379: signal is true;
	signal I36382: std_logic; attribute dont_touch of I36382: signal is true;
	signal I36390: std_logic; attribute dont_touch of I36390: signal is true;
	signal I36393: std_logic; attribute dont_touch of I36393: signal is true;
	signal I36397: std_logic; attribute dont_touch of I36397: signal is true;
	signal I36404: std_logic; attribute dont_touch of I36404: signal is true;
	signal I36407: std_logic; attribute dont_touch of I36407: signal is true;
	signal I36411: std_logic; attribute dont_touch of I36411: signal is true;
	signal I36417: std_logic; attribute dont_touch of I36417: signal is true;
	signal I36420: std_logic; attribute dont_touch of I36420: signal is true;
	signal I36423: std_logic; attribute dont_touch of I36423: signal is true;
	signal I36426: std_logic; attribute dont_touch of I36426: signal is true;
	signal I36432: std_logic; attribute dont_touch of I36432: signal is true;
	signal I36438: std_logic; attribute dont_touch of I36438: signal is true;
	signal I36441: std_logic; attribute dont_touch of I36441: signal is true;
	signal I36444: std_logic; attribute dont_touch of I36444: signal is true;
	signal I36447: std_logic; attribute dont_touch of I36447: signal is true;
	signal I36450: std_logic; attribute dont_touch of I36450: signal is true;
	signal I36454: std_logic; attribute dont_touch of I36454: signal is true;
	signal I36459: std_logic; attribute dont_touch of I36459: signal is true;
	signal I36462: std_logic; attribute dont_touch of I36462: signal is true;
	signal I36465: std_logic; attribute dont_touch of I36465: signal is true;
	signal I36468: std_logic; attribute dont_touch of I36468: signal is true;
	signal I36473: std_logic; attribute dont_touch of I36473: signal is true;
	signal I36476: std_logic; attribute dont_touch of I36476: signal is true;
	signal I36479: std_logic; attribute dont_touch of I36479: signal is true;
	signal I36483: std_logic; attribute dont_touch of I36483: signal is true;
	signal I36486: std_logic; attribute dont_touch of I36486: signal is true;
	signal I36490: std_logic; attribute dont_touch of I36490: signal is true;
	signal I36493: std_logic; attribute dont_touch of I36493: signal is true;
	signal I36496: std_logic; attribute dont_touch of I36496: signal is true;
	signal I36499: std_logic; attribute dont_touch of I36499: signal is true;
	signal I36502: std_logic; attribute dont_touch of I36502: signal is true;
	signal I36507: std_logic; attribute dont_touch of I36507: signal is true;
	signal I36510: std_logic; attribute dont_touch of I36510: signal is true;
	signal I36513: std_logic; attribute dont_touch of I36513: signal is true;
	signal I36516: std_logic; attribute dont_touch of I36516: signal is true;
	signal I36521: std_logic; attribute dont_touch of I36521: signal is true;
	signal I36524: std_logic; attribute dont_touch of I36524: signal is true;
	signal I36527: std_logic; attribute dont_touch of I36527: signal is true;
	signal I36530: std_logic; attribute dont_touch of I36530: signal is true;
	signal I36533: std_logic; attribute dont_touch of I36533: signal is true;
	signal I36536: std_logic; attribute dont_touch of I36536: signal is true;
	signal I36539: std_logic; attribute dont_touch of I36539: signal is true;
	signal I36542: std_logic; attribute dont_touch of I36542: signal is true;
	signal I36545: std_logic; attribute dont_touch of I36545: signal is true;
	signal I36551: std_logic; attribute dont_touch of I36551: signal is true;
	signal I36554: std_logic; attribute dont_touch of I36554: signal is true;
	signal I36557: std_logic; attribute dont_touch of I36557: signal is true;
	signal I36560: std_logic; attribute dont_touch of I36560: signal is true;
	signal I36563: std_logic; attribute dont_touch of I36563: signal is true;
	signal I36568: std_logic; attribute dont_touch of I36568: signal is true;
	signal I36571: std_logic; attribute dont_touch of I36571: signal is true;
	signal I36574: std_logic; attribute dont_touch of I36574: signal is true;
	signal I36577: std_logic; attribute dont_touch of I36577: signal is true;
	signal I36582: std_logic; attribute dont_touch of I36582: signal is true;
	signal I36585: std_logic; attribute dont_touch of I36585: signal is true;
	signal I36588: std_logic; attribute dont_touch of I36588: signal is true;
	signal I36591: std_logic; attribute dont_touch of I36591: signal is true;
	signal I36592: std_logic; attribute dont_touch of I36592: signal is true;
	signal I36593: std_logic; attribute dont_touch of I36593: signal is true;
	signal I36598: std_logic; attribute dont_touch of I36598: signal is true;
	signal I36601: std_logic; attribute dont_touch of I36601: signal is true;
	signal I36604: std_logic; attribute dont_touch of I36604: signal is true;
	signal I36609: std_logic; attribute dont_touch of I36609: signal is true;
	signal I36612: std_logic; attribute dont_touch of I36612: signal is true;
	signal I36615: std_logic; attribute dont_touch of I36615: signal is true;
	signal I36618: std_logic; attribute dont_touch of I36618: signal is true;
	signal I36621: std_logic; attribute dont_touch of I36621: signal is true;
	signal I36627: std_logic; attribute dont_touch of I36627: signal is true;
	signal I36630: std_logic; attribute dont_touch of I36630: signal is true;
	signal I36633: std_logic; attribute dont_touch of I36633: signal is true;
	signal I36636: std_logic; attribute dont_touch of I36636: signal is true;
	signal I36639: std_logic; attribute dont_touch of I36639: signal is true;
	signal I36644: std_logic; attribute dont_touch of I36644: signal is true;
	signal I36647: std_logic; attribute dont_touch of I36647: signal is true;
	signal I36650: std_logic; attribute dont_touch of I36650: signal is true;
	signal I36653: std_logic; attribute dont_touch of I36653: signal is true;
	signal I36656: std_logic; attribute dont_touch of I36656: signal is true;
	signal I36659: std_logic; attribute dont_touch of I36659: signal is true;
	signal I36663: std_logic; attribute dont_touch of I36663: signal is true;
	signal I36666: std_logic; attribute dont_touch of I36666: signal is true;
	signal I36667: std_logic; attribute dont_touch of I36667: signal is true;
	signal I36668: std_logic; attribute dont_touch of I36668: signal is true;
	signal I36673: std_logic; attribute dont_touch of I36673: signal is true;
	signal I36676: std_logic; attribute dont_touch of I36676: signal is true;
	signal I36679: std_logic; attribute dont_touch of I36679: signal is true;
	signal I36684: std_logic; attribute dont_touch of I36684: signal is true;
	signal I36687: std_logic; attribute dont_touch of I36687: signal is true;
	signal I36690: std_logic; attribute dont_touch of I36690: signal is true;
	signal I36693: std_logic; attribute dont_touch of I36693: signal is true;
	signal I36696: std_logic; attribute dont_touch of I36696: signal is true;
	signal I36702: std_logic; attribute dont_touch of I36702: signal is true;
	signal I36705: std_logic; attribute dont_touch of I36705: signal is true;
	signal I36708: std_logic; attribute dont_touch of I36708: signal is true;
	signal I36711: std_logic; attribute dont_touch of I36711: signal is true;
	signal I36714: std_logic; attribute dont_touch of I36714: signal is true;
	signal I36718: std_logic; attribute dont_touch of I36718: signal is true;
	signal I36721: std_logic; attribute dont_touch of I36721: signal is true;
	signal I36724: std_logic; attribute dont_touch of I36724: signal is true;
	signal I36728: std_logic; attribute dont_touch of I36728: signal is true;
	signal I36731: std_logic; attribute dont_touch of I36731: signal is true;
	signal I36732: std_logic; attribute dont_touch of I36732: signal is true;
	signal I36733: std_logic; attribute dont_touch of I36733: signal is true;
	signal I36738: std_logic; attribute dont_touch of I36738: signal is true;
	signal I36741: std_logic; attribute dont_touch of I36741: signal is true;
	signal I36744: std_logic; attribute dont_touch of I36744: signal is true;
	signal I36749: std_logic; attribute dont_touch of I36749: signal is true;
	signal I36752: std_logic; attribute dont_touch of I36752: signal is true;
	signal I36755: std_logic; attribute dont_touch of I36755: signal is true;
	signal I36758: std_logic; attribute dont_touch of I36758: signal is true;
	signal I36761: std_logic; attribute dont_touch of I36761: signal is true;
	signal I36766: std_logic; attribute dont_touch of I36766: signal is true;
	signal I36769: std_logic; attribute dont_touch of I36769: signal is true;
	signal I36772: std_logic; attribute dont_touch of I36772: signal is true;
	signal I36776: std_logic; attribute dont_touch of I36776: signal is true;
	signal I36779: std_logic; attribute dont_touch of I36779: signal is true;
	signal I36780: std_logic; attribute dont_touch of I36780: signal is true;
	signal I36781: std_logic; attribute dont_touch of I36781: signal is true;
	signal I36786: std_logic; attribute dont_touch of I36786: signal is true;
	signal I36789: std_logic; attribute dont_touch of I36789: signal is true;
	signal I36792: std_logic; attribute dont_touch of I36792: signal is true;
	signal I36797: std_logic; attribute dont_touch of I36797: signal is true;
	signal I36800: std_logic; attribute dont_touch of I36800: signal is true;
	signal I36803: std_logic; attribute dont_touch of I36803: signal is true;
	signal I36808: std_logic; attribute dont_touch of I36808: signal is true;
	signal I36848: std_logic; attribute dont_touch of I36848: signal is true;
	signal I36860: std_logic; attribute dont_touch of I36860: signal is true;
	signal I36864: std_logic; attribute dont_touch of I36864: signal is true;
	signal I36867: std_logic; attribute dont_touch of I36867: signal is true;
	signal I36870: std_logic; attribute dont_touch of I36870: signal is true;
	signal I36873: std_logic; attribute dont_touch of I36873: signal is true;
	signal I36876: std_logic; attribute dont_touch of I36876: signal is true;
	signal I36879: std_logic; attribute dont_touch of I36879: signal is true;
	signal I36882: std_logic; attribute dont_touch of I36882: signal is true;
	signal I36885: std_logic; attribute dont_touch of I36885: signal is true;
	signal I36888: std_logic; attribute dont_touch of I36888: signal is true;
	signal I36891: std_logic; attribute dont_touch of I36891: signal is true;
	signal I36894: std_logic; attribute dont_touch of I36894: signal is true;
	signal I36897: std_logic; attribute dont_touch of I36897: signal is true;
	signal I36900: std_logic; attribute dont_touch of I36900: signal is true;
	signal I36903: std_logic; attribute dont_touch of I36903: signal is true;
	signal I36906: std_logic; attribute dont_touch of I36906: signal is true;
	signal I36909: std_logic; attribute dont_touch of I36909: signal is true;
	signal I36912: std_logic; attribute dont_touch of I36912: signal is true;
	signal I36915: std_logic; attribute dont_touch of I36915: signal is true;
	signal I36918: std_logic; attribute dont_touch of I36918: signal is true;
	signal I36921: std_logic; attribute dont_touch of I36921: signal is true;
	signal I36924: std_logic; attribute dont_touch of I36924: signal is true;
	signal I36927: std_logic; attribute dont_touch of I36927: signal is true;
	signal I36930: std_logic; attribute dont_touch of I36930: signal is true;
	signal I36933: std_logic; attribute dont_touch of I36933: signal is true;
	signal I36936: std_logic; attribute dont_touch of I36936: signal is true;
	signal I36939: std_logic; attribute dont_touch of I36939: signal is true;
	signal I36942: std_logic; attribute dont_touch of I36942: signal is true;
	signal I36945: std_logic; attribute dont_touch of I36945: signal is true;
	signal I36948: std_logic; attribute dont_touch of I36948: signal is true;
	signal I36951: std_logic; attribute dont_touch of I36951: signal is true;
	signal I36954: std_logic; attribute dont_touch of I36954: signal is true;
	signal I36957: std_logic; attribute dont_touch of I36957: signal is true;
	signal I36960: std_logic; attribute dont_touch of I36960: signal is true;
	signal I36963: std_logic; attribute dont_touch of I36963: signal is true;
	signal I36966: std_logic; attribute dont_touch of I36966: signal is true;
	signal I36969: std_logic; attribute dont_touch of I36969: signal is true;
	signal I36972: std_logic; attribute dont_touch of I36972: signal is true;
	signal I36975: std_logic; attribute dont_touch of I36975: signal is true;
	signal I36978: std_logic; attribute dont_touch of I36978: signal is true;
	signal I36981: std_logic; attribute dont_touch of I36981: signal is true;
	signal I36984: std_logic; attribute dont_touch of I36984: signal is true;
	signal I36987: std_logic; attribute dont_touch of I36987: signal is true;
	signal I36990: std_logic; attribute dont_touch of I36990: signal is true;
	signal I36993: std_logic; attribute dont_touch of I36993: signal is true;
	signal I36996: std_logic; attribute dont_touch of I36996: signal is true;
	signal I36999: std_logic; attribute dont_touch of I36999: signal is true;
	signal I37002: std_logic; attribute dont_touch of I37002: signal is true;
	signal I37005: std_logic; attribute dont_touch of I37005: signal is true;
	signal I37008: std_logic; attribute dont_touch of I37008: signal is true;
	signal I37011: std_logic; attribute dont_touch of I37011: signal is true;
	signal I37014: std_logic; attribute dont_touch of I37014: signal is true;
	signal I37017: std_logic; attribute dont_touch of I37017: signal is true;
	signal I37020: std_logic; attribute dont_touch of I37020: signal is true;
	signal I37023: std_logic; attribute dont_touch of I37023: signal is true;
	signal I37026: std_logic; attribute dont_touch of I37026: signal is true;
	signal I37029: std_logic; attribute dont_touch of I37029: signal is true;
	signal I37032: std_logic; attribute dont_touch of I37032: signal is true;
	signal I37035: std_logic; attribute dont_touch of I37035: signal is true;
	signal I37038: std_logic; attribute dont_touch of I37038: signal is true;
	signal I37041: std_logic; attribute dont_touch of I37041: signal is true;
	signal I37044: std_logic; attribute dont_touch of I37044: signal is true;
	signal I37047: std_logic; attribute dont_touch of I37047: signal is true;
	signal I37050: std_logic; attribute dont_touch of I37050: signal is true;
	signal I37053: std_logic; attribute dont_touch of I37053: signal is true;
	signal I37056: std_logic; attribute dont_touch of I37056: signal is true;
	signal I37059: std_logic; attribute dont_touch of I37059: signal is true;
	signal I37062: std_logic; attribute dont_touch of I37062: signal is true;
	signal I37065: std_logic; attribute dont_touch of I37065: signal is true;
	signal I37068: std_logic; attribute dont_touch of I37068: signal is true;
	signal I37071: std_logic; attribute dont_touch of I37071: signal is true;
	signal I37074: std_logic; attribute dont_touch of I37074: signal is true;
	signal I37077: std_logic; attribute dont_touch of I37077: signal is true;
	signal I37080: std_logic; attribute dont_touch of I37080: signal is true;
	signal I37083: std_logic; attribute dont_touch of I37083: signal is true;
	signal I37086: std_logic; attribute dont_touch of I37086: signal is true;
	signal I37089: std_logic; attribute dont_touch of I37089: signal is true;
	signal I37092: std_logic; attribute dont_touch of I37092: signal is true;
	signal I37095: std_logic; attribute dont_touch of I37095: signal is true;
	signal I37098: std_logic; attribute dont_touch of I37098: signal is true;
	signal I37101: std_logic; attribute dont_touch of I37101: signal is true;
	signal I37104: std_logic; attribute dont_touch of I37104: signal is true;
	signal I37107: std_logic; attribute dont_touch of I37107: signal is true;
	signal I37110: std_logic; attribute dont_touch of I37110: signal is true;
	signal I37113: std_logic; attribute dont_touch of I37113: signal is true;
	signal I37116: std_logic; attribute dont_touch of I37116: signal is true;
	signal I37119: std_logic; attribute dont_touch of I37119: signal is true;
	signal I37122: std_logic; attribute dont_touch of I37122: signal is true;
	signal I37125: std_logic; attribute dont_touch of I37125: signal is true;
	signal I37128: std_logic; attribute dont_touch of I37128: signal is true;
	signal I37131: std_logic; attribute dont_touch of I37131: signal is true;
	signal I37134: std_logic; attribute dont_touch of I37134: signal is true;
	signal I37137: std_logic; attribute dont_touch of I37137: signal is true;
	signal I37140: std_logic; attribute dont_touch of I37140: signal is true;
	signal I37143: std_logic; attribute dont_touch of I37143: signal is true;
	signal I37146: std_logic; attribute dont_touch of I37146: signal is true;
	signal I37149: std_logic; attribute dont_touch of I37149: signal is true;
	signal I37152: std_logic; attribute dont_touch of I37152: signal is true;
	signal I37155: std_logic; attribute dont_touch of I37155: signal is true;
	signal I37158: std_logic; attribute dont_touch of I37158: signal is true;
	signal I37161: std_logic; attribute dont_touch of I37161: signal is true;
	signal I37164: std_logic; attribute dont_touch of I37164: signal is true;
	signal I37167: std_logic; attribute dont_touch of I37167: signal is true;
	signal I37170: std_logic; attribute dont_touch of I37170: signal is true;
	signal I37173: std_logic; attribute dont_touch of I37173: signal is true;
	signal I37176: std_logic; attribute dont_touch of I37176: signal is true;
	signal I37179: std_logic; attribute dont_touch of I37179: signal is true;
	signal I37182: std_logic; attribute dont_touch of I37182: signal is true;
	signal I37185: std_logic; attribute dont_touch of I37185: signal is true;
	signal I37188: std_logic; attribute dont_touch of I37188: signal is true;
	signal I37191: std_logic; attribute dont_touch of I37191: signal is true;
	signal I37194: std_logic; attribute dont_touch of I37194: signal is true;
	signal I37197: std_logic; attribute dont_touch of I37197: signal is true;
	signal I37200: std_logic; attribute dont_touch of I37200: signal is true;
	signal I37203: std_logic; attribute dont_touch of I37203: signal is true;
	signal I37228: std_logic; attribute dont_touch of I37228: signal is true;
	signal I37232: std_logic; attribute dont_touch of I37232: signal is true;
	signal I37238: std_logic; attribute dont_touch of I37238: signal is true;
	signal I37252: std_logic; attribute dont_touch of I37252: signal is true;
	signal I37260: std_logic; attribute dont_touch of I37260: signal is true;
	signal I37266: std_logic; attribute dont_touch of I37266: signal is true;
	signal I37269: std_logic; attribute dont_touch of I37269: signal is true;
	signal I37273: std_logic; attribute dont_touch of I37273: signal is true;
	signal I37277: std_logic; attribute dont_touch of I37277: signal is true;
	signal I37280: std_logic; attribute dont_touch of I37280: signal is true;
	signal I37284: std_logic; attribute dont_touch of I37284: signal is true;
	signal I37291: std_logic; attribute dont_touch of I37291: signal is true;
	signal I37295: std_logic; attribute dont_touch of I37295: signal is true;
	signal I37296: std_logic; attribute dont_touch of I37296: signal is true;
	signal I37297: std_logic; attribute dont_touch of I37297: signal is true;
	signal I37303: std_logic; attribute dont_touch of I37303: signal is true;
	signal I37304: std_logic; attribute dont_touch of I37304: signal is true;
	signal I37305: std_logic; attribute dont_touch of I37305: signal is true;
	signal I37311: std_logic; attribute dont_touch of I37311: signal is true;
	signal I37312: std_logic; attribute dont_touch of I37312: signal is true;
	signal I37313: std_logic; attribute dont_touch of I37313: signal is true;
	signal I37319: std_logic; attribute dont_touch of I37319: signal is true;
	signal I37322: std_logic; attribute dont_touch of I37322: signal is true;
	signal I37323: std_logic; attribute dont_touch of I37323: signal is true;
	signal I37324: std_logic; attribute dont_touch of I37324: signal is true;
	signal I37330: std_logic; attribute dont_touch of I37330: signal is true;
	signal I37334: std_logic; attribute dont_touch of I37334: signal is true;
	signal I37356: std_logic; attribute dont_touch of I37356: signal is true;
	signal I37357: std_logic; attribute dont_touch of I37357: signal is true;
	signal I37358: std_logic; attribute dont_touch of I37358: signal is true;
	signal I37379: std_logic; attribute dont_touch of I37379: signal is true;
	signal I37386: std_logic; attribute dont_touch of I37386: signal is true;
	signal I37394: std_logic; attribute dont_touch of I37394: signal is true;
	signal I37400: std_logic; attribute dont_touch of I37400: signal is true;
	signal I37410: std_logic; attribute dont_touch of I37410: signal is true;
	signal I37415: std_logic; attribute dont_touch of I37415: signal is true;
	signal I37426: std_logic; attribute dont_touch of I37426: signal is true;
	signal I37459: std_logic; attribute dont_touch of I37459: signal is true;
	signal I37467: std_logic; attribute dont_touch of I37467: signal is true;
	signal I37471: std_logic; attribute dont_touch of I37471: signal is true;
	signal I37474: std_logic; attribute dont_touch of I37474: signal is true;
	signal I37481: std_logic; attribute dont_touch of I37481: signal is true;
	signal I37484: std_logic; attribute dont_touch of I37484: signal is true;
	signal I37488: std_logic; attribute dont_touch of I37488: signal is true;
	signal I37494: std_logic; attribute dont_touch of I37494: signal is true;
	signal I37497: std_logic; attribute dont_touch of I37497: signal is true;
	signal I37502: std_logic; attribute dont_touch of I37502: signal is true;
	signal I37508: std_logic; attribute dont_touch of I37508: signal is true;
	signal I37514: std_logic; attribute dont_touch of I37514: signal is true;
	signal I37566: std_logic; attribute dont_touch of I37566: signal is true;
	signal I37569: std_logic; attribute dont_touch of I37569: signal is true;
	signal I37572: std_logic; attribute dont_touch of I37572: signal is true;
	signal I37575: std_logic; attribute dont_touch of I37575: signal is true;
	signal I37578: std_logic; attribute dont_touch of I37578: signal is true;
	signal I37581: std_logic; attribute dont_touch of I37581: signal is true;
	signal I37584: std_logic; attribute dont_touch of I37584: signal is true;
	signal I37587: std_logic; attribute dont_touch of I37587: signal is true;
	signal I37590: std_logic; attribute dont_touch of I37590: signal is true;
	signal I37593: std_logic; attribute dont_touch of I37593: signal is true;
	signal I37596: std_logic; attribute dont_touch of I37596: signal is true;
	signal I37599: std_logic; attribute dont_touch of I37599: signal is true;
	signal I37602: std_logic; attribute dont_touch of I37602: signal is true;
	signal I37605: std_logic; attribute dont_touch of I37605: signal is true;
	signal I37608: std_logic; attribute dont_touch of I37608: signal is true;
	signal I37611: std_logic; attribute dont_touch of I37611: signal is true;
	signal I37614: std_logic; attribute dont_touch of I37614: signal is true;
	signal I37617: std_logic; attribute dont_touch of I37617: signal is true;
	signal I37620: std_logic; attribute dont_touch of I37620: signal is true;
	signal I37623: std_logic; attribute dont_touch of I37623: signal is true;
	signal I37626: std_logic; attribute dont_touch of I37626: signal is true;
	signal I37629: std_logic; attribute dont_touch of I37629: signal is true;
	signal I37632: std_logic; attribute dont_touch of I37632: signal is true;
	signal I37635: std_logic; attribute dont_touch of I37635: signal is true;
	signal I37638: std_logic; attribute dont_touch of I37638: signal is true;
	signal I37641: std_logic; attribute dont_touch of I37641: signal is true;
	signal I37644: std_logic; attribute dont_touch of I37644: signal is true;
	signal I37647: std_logic; attribute dont_touch of I37647: signal is true;
	signal I37650: std_logic; attribute dont_touch of I37650: signal is true;
	signal I37653: std_logic; attribute dont_touch of I37653: signal is true;
	signal I37656: std_logic; attribute dont_touch of I37656: signal is true;
	signal I37659: std_logic; attribute dont_touch of I37659: signal is true;
	signal I37662: std_logic; attribute dont_touch of I37662: signal is true;
	signal I37665: std_logic; attribute dont_touch of I37665: signal is true;
	signal I37702: std_logic; attribute dont_touch of I37702: signal is true;
	signal I37712: std_logic; attribute dont_touch of I37712: signal is true;
	signal I37716: std_logic; attribute dont_touch of I37716: signal is true;
	signal I37725: std_logic; attribute dont_touch of I37725: signal is true;
	signal I37729: std_logic; attribute dont_touch of I37729: signal is true;
	signal I37736: std_logic; attribute dont_touch of I37736: signal is true;
	signal I37740: std_logic; attribute dont_touch of I37740: signal is true;
	signal I37746: std_logic; attribute dont_touch of I37746: signal is true;
	signal I37752: std_logic; attribute dont_touch of I37752: signal is true;
	signal I37757: std_logic; attribute dont_touch of I37757: signal is true;
	signal I37760: std_logic; attribute dont_touch of I37760: signal is true;
	signal I37765: std_logic; attribute dont_touch of I37765: signal is true;
	signal I37768: std_logic; attribute dont_touch of I37768: signal is true;
	signal I37771: std_logic; attribute dont_touch of I37771: signal is true;
	signal I37775: std_logic; attribute dont_touch of I37775: signal is true;
	signal I37778: std_logic; attribute dont_touch of I37778: signal is true;
	signal I37781: std_logic; attribute dont_touch of I37781: signal is true;
	signal I37784: std_logic; attribute dont_touch of I37784: signal is true;
	signal I37787: std_logic; attribute dont_touch of I37787: signal is true;
	signal I37790: std_logic; attribute dont_touch of I37790: signal is true;
	signal I37793: std_logic; attribute dont_touch of I37793: signal is true;
	signal I37796: std_logic; attribute dont_touch of I37796: signal is true;
	signal I37800: std_logic; attribute dont_touch of I37800: signal is true;
	signal I37804: std_logic; attribute dont_touch of I37804: signal is true;
	signal I37808: std_logic; attribute dont_touch of I37808: signal is true;
	signal I37813: std_logic; attribute dont_touch of I37813: signal is true;
	signal I37814: std_logic; attribute dont_touch of I37814: signal is true;
	signal I37815: std_logic; attribute dont_touch of I37815: signal is true;
	signal I37822: std_logic; attribute dont_touch of I37822: signal is true;
	signal I37823: std_logic; attribute dont_touch of I37823: signal is true;
	signal I37824: std_logic; attribute dont_touch of I37824: signal is true;
	signal I37842: std_logic; attribute dont_touch of I37842: signal is true;
	signal I37846: std_logic; attribute dont_touch of I37846: signal is true;
	signal I37851: std_logic; attribute dont_touch of I37851: signal is true;
	signal I37854: std_logic; attribute dont_touch of I37854: signal is true;
	signal I37858: std_logic; attribute dont_touch of I37858: signal is true;
	signal I37863: std_logic; attribute dont_touch of I37863: signal is true;
	signal I37868: std_logic; attribute dont_touch of I37868: signal is true;
	signal I37871: std_logic; attribute dont_touch of I37871: signal is true;
	signal I37875: std_logic; attribute dont_touch of I37875: signal is true;
	signal I37880: std_logic; attribute dont_touch of I37880: signal is true;
	signal I37885: std_logic; attribute dont_touch of I37885: signal is true;
	signal I37891: std_logic; attribute dont_touch of I37891: signal is true;
	signal I37894: std_logic; attribute dont_touch of I37894: signal is true;
	signal I37897: std_logic; attribute dont_touch of I37897: signal is true;
	signal I37901: std_logic; attribute dont_touch of I37901: signal is true;
	signal I37906: std_logic; attribute dont_touch of I37906: signal is true;
	signal I37912: std_logic; attribute dont_touch of I37912: signal is true;
	signal I37917: std_logic; attribute dont_touch of I37917: signal is true;
	signal I37920: std_logic; attribute dont_touch of I37920: signal is true;
	signal I37924: std_logic; attribute dont_touch of I37924: signal is true;
	signal I37928: std_logic; attribute dont_touch of I37928: signal is true;
	signal I37934: std_logic; attribute dont_touch of I37934: signal is true;
	signal I37939: std_logic; attribute dont_touch of I37939: signal is true;
	signal I37942: std_logic; attribute dont_touch of I37942: signal is true;
	signal I37946: std_logic; attribute dont_touch of I37946: signal is true;
	signal I37950: std_logic; attribute dont_touch of I37950: signal is true;
	signal I37956: std_logic; attribute dont_touch of I37956: signal is true;
	signal I37961: std_logic; attribute dont_touch of I37961: signal is true;
	signal I37965: std_logic; attribute dont_touch of I37965: signal is true;
	signal I37968: std_logic; attribute dont_touch of I37968: signal is true;
	signal I37973: std_logic; attribute dont_touch of I37973: signal is true;
	signal I37978: std_logic; attribute dont_touch of I37978: signal is true;
	signal I37982: std_logic; attribute dont_touch of I37982: signal is true;
	signal I37986: std_logic; attribute dont_touch of I37986: signal is true;
	signal I37991: std_logic; attribute dont_touch of I37991: signal is true;
	signal I37994: std_logic; attribute dont_touch of I37994: signal is true;
	signal I37999: std_logic; attribute dont_touch of I37999: signal is true;
	signal I38003: std_logic; attribute dont_touch of I38003: signal is true;
	signal I38007: std_logic; attribute dont_touch of I38007: signal is true;
	signal I38011: std_logic; attribute dont_touch of I38011: signal is true;
	signal I38014: std_logic; attribute dont_touch of I38014: signal is true;
	signal I38018: std_logic; attribute dont_touch of I38018: signal is true;
	signal I38024: std_logic; attribute dont_touch of I38024: signal is true;
	signal I38028: std_logic; attribute dont_touch of I38028: signal is true;
	signal I38032: std_logic; attribute dont_touch of I38032: signal is true;
	signal I38035: std_logic; attribute dont_touch of I38035: signal is true;
	signal I38038: std_logic; attribute dont_touch of I38038: signal is true;
	signal I38042: std_logic; attribute dont_touch of I38042: signal is true;
	signal I38046: std_logic; attribute dont_touch of I38046: signal is true;
	signal I38049: std_logic; attribute dont_touch of I38049: signal is true;
	signal I38053: std_logic; attribute dont_touch of I38053: signal is true;
	signal I38056: std_logic; attribute dont_touch of I38056: signal is true;
	signal I38059: std_logic; attribute dont_touch of I38059: signal is true;
	signal I38064: std_logic; attribute dont_touch of I38064: signal is true;
	signal I38068: std_logic; attribute dont_touch of I38068: signal is true;
	signal I38071: std_logic; attribute dont_touch of I38071: signal is true;
	signal I38074: std_logic; attribute dont_touch of I38074: signal is true;
	signal I38077: std_logic; attribute dont_touch of I38077: signal is true;
	signal I38080: std_logic; attribute dont_touch of I38080: signal is true;
	signal I38085: std_logic; attribute dont_touch of I38085: signal is true;
	signal I38088: std_logic; attribute dont_touch of I38088: signal is true;
	signal I38091: std_logic; attribute dont_touch of I38091: signal is true;
	signal I38094: std_logic; attribute dont_touch of I38094: signal is true;
	signal I38097: std_logic; attribute dont_touch of I38097: signal is true;
	signal I38101: std_logic; attribute dont_touch of I38101: signal is true;
	signal I38104: std_logic; attribute dont_touch of I38104: signal is true;
	signal I38107: std_logic; attribute dont_touch of I38107: signal is true;
	signal I38111: std_logic; attribute dont_touch of I38111: signal is true;
	signal I38119: std_logic; attribute dont_touch of I38119: signal is true;
	signal I38122: std_logic; attribute dont_touch of I38122: signal is true;
	signal I38125: std_logic; attribute dont_touch of I38125: signal is true;
	signal I38128: std_logic; attribute dont_touch of I38128: signal is true;
	signal I38136: std_logic; attribute dont_touch of I38136: signal is true;
	signal I38139: std_logic; attribute dont_touch of I38139: signal is true;
	signal I38142: std_logic; attribute dont_touch of I38142: signal is true;
	signal I38145: std_logic; attribute dont_touch of I38145: signal is true;
	signal I38148: std_logic; attribute dont_touch of I38148: signal is true;
	signal I38151: std_logic; attribute dont_touch of I38151: signal is true;
	signal I38154: std_logic; attribute dont_touch of I38154: signal is true;
	signal I38157: std_logic; attribute dont_touch of I38157: signal is true;
	signal I38160: std_logic; attribute dont_touch of I38160: signal is true;
	signal I38163: std_logic; attribute dont_touch of I38163: signal is true;
	signal I38166: std_logic; attribute dont_touch of I38166: signal is true;
	signal I38169: std_logic; attribute dont_touch of I38169: signal is true;
	signal I38172: std_logic; attribute dont_touch of I38172: signal is true;
	signal I38175: std_logic; attribute dont_touch of I38175: signal is true;
	signal I38178: std_logic; attribute dont_touch of I38178: signal is true;
	signal I38181: std_logic; attribute dont_touch of I38181: signal is true;
	signal I38184: std_logic; attribute dont_touch of I38184: signal is true;
	signal I38187: std_logic; attribute dont_touch of I38187: signal is true;
	signal I38190: std_logic; attribute dont_touch of I38190: signal is true;
	signal I38193: std_logic; attribute dont_touch of I38193: signal is true;
	signal I38196: std_logic; attribute dont_touch of I38196: signal is true;
	signal I38199: std_logic; attribute dont_touch of I38199: signal is true;
	signal I38202: std_logic; attribute dont_touch of I38202: signal is true;
	signal I38205: std_logic; attribute dont_touch of I38205: signal is true;
	signal I38208: std_logic; attribute dont_touch of I38208: signal is true;
	signal I38211: std_logic; attribute dont_touch of I38211: signal is true;
	signal I38214: std_logic; attribute dont_touch of I38214: signal is true;
	signal I38217: std_logic; attribute dont_touch of I38217: signal is true;
	signal I38220: std_logic; attribute dont_touch of I38220: signal is true;
	signal I38223: std_logic; attribute dont_touch of I38223: signal is true;
	signal I38226: std_logic; attribute dont_touch of I38226: signal is true;
	signal I38229: std_logic; attribute dont_touch of I38229: signal is true;
	signal I38232: std_logic; attribute dont_touch of I38232: signal is true;
	signal I38235: std_logic; attribute dont_touch of I38235: signal is true;
	signal I38238: std_logic; attribute dont_touch of I38238: signal is true;
	signal I38241: std_logic; attribute dont_touch of I38241: signal is true;
	signal I38245: std_logic; attribute dont_touch of I38245: signal is true;
	signal I38250: std_logic; attribute dont_touch of I38250: signal is true;
	signal I38258: std_logic; attribute dont_touch of I38258: signal is true;
	signal I38272: std_logic; attribute dont_touch of I38272: signal is true;
	signal I38275: std_logic; attribute dont_touch of I38275: signal is true;
	signal I38278: std_logic; attribute dont_touch of I38278: signal is true;
	signal I38282: std_logic; attribute dont_touch of I38282: signal is true;
	signal I38321: std_logic; attribute dont_touch of I38321: signal is true;
	signal I38330: std_logic; attribute dont_touch of I38330: signal is true;
	signal I38339: std_logic; attribute dont_touch of I38339: signal is true;
	signal I38342: std_logic; attribute dont_touch of I38342: signal is true;
	signal I38345: std_logic; attribute dont_touch of I38345: signal is true;
	signal I38348: std_logic; attribute dont_touch of I38348: signal is true;
	signal I38352: std_logic; attribute dont_touch of I38352: signal is true;
	signal I38355: std_logic; attribute dont_touch of I38355: signal is true;
	signal I38360: std_logic; attribute dont_touch of I38360: signal is true;
	signal I38363: std_logic; attribute dont_touch of I38363: signal is true;
	signal I38369: std_logic; attribute dont_touch of I38369: signal is true;
	signal I38378: std_logic; attribute dont_touch of I38378: signal is true;
	signal I38379: std_logic; attribute dont_touch of I38379: signal is true;
	signal I38380: std_logic; attribute dont_touch of I38380: signal is true;
	signal I38386: std_logic; attribute dont_touch of I38386: signal is true;
	signal I38391: std_logic; attribute dont_touch of I38391: signal is true;
	signal I38396: std_logic; attribute dont_touch of I38396: signal is true;
	signal I38401: std_logic; attribute dont_touch of I38401: signal is true;
	signal I38405: std_logic; attribute dont_touch of I38405: signal is true;
	signal I38408: std_logic; attribute dont_touch of I38408: signal is true;
	signal I38412: std_logic; attribute dont_touch of I38412: signal is true;
	signal I38421: std_logic; attribute dont_touch of I38421: signal is true;
	signal I38428: std_logic; attribute dont_touch of I38428: signal is true;
	signal I38434: std_logic; attribute dont_touch of I38434: signal is true;
	signal I38437: std_logic; attribute dont_touch of I38437: signal is true;
	signal I38440: std_logic; attribute dont_touch of I38440: signal is true;
	signal I38447: std_logic; attribute dont_touch of I38447: signal is true;
	signal I38450: std_logic; attribute dont_touch of I38450: signal is true;
	signal I38453: std_logic; attribute dont_touch of I38453: signal is true;
	signal I38456: std_logic; attribute dont_touch of I38456: signal is true;
	signal I38459: std_logic; attribute dont_touch of I38459: signal is true;
	signal I38462: std_logic; attribute dont_touch of I38462: signal is true;
	signal I38466: std_logic; attribute dont_touch of I38466: signal is true;
	signal I38471: std_logic; attribute dont_touch of I38471: signal is true;
	signal I38474: std_logic; attribute dont_touch of I38474: signal is true;
	signal I38477: std_logic; attribute dont_touch of I38477: signal is true;
	signal I38480: std_logic; attribute dont_touch of I38480: signal is true;
	signal I38483: std_logic; attribute dont_touch of I38483: signal is true;
	signal I38486: std_logic; attribute dont_touch of I38486: signal is true;
	signal I38491: std_logic; attribute dont_touch of I38491: signal is true;
	signal I38496: std_logic; attribute dont_touch of I38496: signal is true;
	signal I38499: std_logic; attribute dont_touch of I38499: signal is true;
	signal I38502: std_logic; attribute dont_touch of I38502: signal is true;
	signal I38505: std_logic; attribute dont_touch of I38505: signal is true;
	signal I38510: std_logic; attribute dont_touch of I38510: signal is true;
	signal I38515: std_logic; attribute dont_touch of I38515: signal is true;
	signal I38518: std_logic; attribute dont_touch of I38518: signal is true;
	signal I38524: std_logic; attribute dont_touch of I38524: signal is true;
	signal I38536: std_logic; attribute dont_touch of I38536: signal is true;
	signal I38539: std_logic; attribute dont_touch of I38539: signal is true;
	signal I38548: std_logic; attribute dont_touch of I38548: signal is true;
	signal I38591: std_logic; attribute dont_touch of I38591: signal is true;
	signal I38594: std_logic; attribute dont_touch of I38594: signal is true;
	signal I38599: std_logic; attribute dont_touch of I38599: signal is true;
	signal I38602: std_logic; attribute dont_touch of I38602: signal is true;
	signal I38606: std_logic; attribute dont_touch of I38606: signal is true;
	signal I38609: std_logic; attribute dont_touch of I38609: signal is true;
	signal I38613: std_logic; attribute dont_touch of I38613: signal is true;
	signal I38617: std_logic; attribute dont_touch of I38617: signal is true;
	signal I38620: std_logic; attribute dont_touch of I38620: signal is true;
	signal I38623: std_logic; attribute dont_touch of I38623: signal is true;
	signal I38626: std_logic; attribute dont_touch of I38626: signal is true;
	signal I38629: std_logic; attribute dont_touch of I38629: signal is true;
	signal I38632: std_logic; attribute dont_touch of I38632: signal is true;
	signal I38635: std_logic; attribute dont_touch of I38635: signal is true;
	signal I38638: std_logic; attribute dont_touch of I38638: signal is true;
	signal I38641: std_logic; attribute dont_touch of I38641: signal is true;
	signal I38644: std_logic; attribute dont_touch of I38644: signal is true;
	signal I38647: std_logic; attribute dont_touch of I38647: signal is true;
	signal I38650: std_logic; attribute dont_touch of I38650: signal is true;
	signal I38653: std_logic; attribute dont_touch of I38653: signal is true;
	signal I38656: std_logic; attribute dont_touch of I38656: signal is true;
	signal I38659: std_logic; attribute dont_touch of I38659: signal is true;
	signal I38662: std_logic; attribute dont_touch of I38662: signal is true;
	signal I38665: std_logic; attribute dont_touch of I38665: signal is true;
	signal I38668: std_logic; attribute dont_touch of I38668: signal is true;
	signal I38671: std_logic; attribute dont_touch of I38671: signal is true;
	signal I38674: std_logic; attribute dont_touch of I38674: signal is true;
	signal I38677: std_logic; attribute dont_touch of I38677: signal is true;
	signal I38680: std_logic; attribute dont_touch of I38680: signal is true;
	signal I38683: std_logic; attribute dont_touch of I38683: signal is true;
	signal I38686: std_logic; attribute dont_touch of I38686: signal is true;
	signal I38689: std_logic; attribute dont_touch of I38689: signal is true;
	signal I38692: std_logic; attribute dont_touch of I38692: signal is true;
	signal I38695: std_logic; attribute dont_touch of I38695: signal is true;
	signal I38698: std_logic; attribute dont_touch of I38698: signal is true;
	signal I38701: std_logic; attribute dont_touch of I38701: signal is true;
	signal I38704: std_logic; attribute dont_touch of I38704: signal is true;
	signal I38707: std_logic; attribute dont_touch of I38707: signal is true;
	signal I38710: std_logic; attribute dont_touch of I38710: signal is true;
	signal I38713: std_logic; attribute dont_touch of I38713: signal is true;
	signal I38716: std_logic; attribute dont_touch of I38716: signal is true;
	signal I38719: std_logic; attribute dont_touch of I38719: signal is true;
	signal I38722: std_logic; attribute dont_touch of I38722: signal is true;
	signal I38725: std_logic; attribute dont_touch of I38725: signal is true;
	signal I38728: std_logic; attribute dont_touch of I38728: signal is true;
	signal I38731: std_logic; attribute dont_touch of I38731: signal is true;
	signal I38734: std_logic; attribute dont_touch of I38734: signal is true;
	signal I38737: std_logic; attribute dont_touch of I38737: signal is true;
	signal I38740: std_logic; attribute dont_touch of I38740: signal is true;
	signal I38743: std_logic; attribute dont_touch of I38743: signal is true;
	signal I38746: std_logic; attribute dont_touch of I38746: signal is true;
	signal I38749: std_logic; attribute dont_touch of I38749: signal is true;
	signal I38752: std_logic; attribute dont_touch of I38752: signal is true;
	signal I38755: std_logic; attribute dont_touch of I38755: signal is true;
	signal I38758: std_logic; attribute dont_touch of I38758: signal is true;
	signal I38761: std_logic; attribute dont_touch of I38761: signal is true;
	signal I38764: std_logic; attribute dont_touch of I38764: signal is true;
	signal I38767: std_logic; attribute dont_touch of I38767: signal is true;
	signal I38770: std_logic; attribute dont_touch of I38770: signal is true;
	signal I38801: std_logic; attribute dont_touch of I38801: signal is true;
	signal I38804: std_logic; attribute dont_touch of I38804: signal is true;
	signal I38807: std_logic; attribute dont_touch of I38807: signal is true;
	signal I38810: std_logic; attribute dont_touch of I38810: signal is true;
	signal I38811: std_logic; attribute dont_touch of I38811: signal is true;
	signal I38812: std_logic; attribute dont_touch of I38812: signal is true;
	signal I38817: std_logic; attribute dont_touch of I38817: signal is true;
	signal I38820: std_logic; attribute dont_touch of I38820: signal is true;
	signal I38821: std_logic; attribute dont_touch of I38821: signal is true;
	signal I38822: std_logic; attribute dont_touch of I38822: signal is true;
	signal I38827: std_logic; attribute dont_touch of I38827: signal is true;
	signal I38831: std_logic; attribute dont_touch of I38831: signal is true;
	signal I38832: std_logic; attribute dont_touch of I38832: signal is true;
	signal I38833: std_logic; attribute dont_touch of I38833: signal is true;
	signal I38838: std_logic; attribute dont_touch of I38838: signal is true;
	signal I38841: std_logic; attribute dont_touch of I38841: signal is true;
	signal I38842: std_logic; attribute dont_touch of I38842: signal is true;
	signal I38843: std_logic; attribute dont_touch of I38843: signal is true;
	signal I38848: std_logic; attribute dont_touch of I38848: signal is true;
	signal I38851: std_logic; attribute dont_touch of I38851: signal is true;
	signal I38854: std_logic; attribute dont_touch of I38854: signal is true;
	signal I38857: std_logic; attribute dont_touch of I38857: signal is true;
	signal I38860: std_logic; attribute dont_touch of I38860: signal is true;
	signal I38863: std_logic; attribute dont_touch of I38863: signal is true;
	signal I38866: std_logic; attribute dont_touch of I38866: signal is true;
	signal I38869: std_logic; attribute dont_touch of I38869: signal is true;
	signal I38872: std_logic; attribute dont_touch of I38872: signal is true;
	signal I38875: std_logic; attribute dont_touch of I38875: signal is true;
	signal I38878: std_logic; attribute dont_touch of I38878: signal is true;
	signal I38881: std_logic; attribute dont_touch of I38881: signal is true;
	signal I38885: std_logic; attribute dont_touch of I38885: signal is true;
	signal I38898: std_logic; attribute dont_touch of I38898: signal is true;
	signal I38905: std_logic; attribute dont_touch of I38905: signal is true;
	signal I38909: std_logic; attribute dont_touch of I38909: signal is true;
	signal I38916: std_logic; attribute dont_touch of I38916: signal is true;
	signal I38920: std_logic; attribute dont_touch of I38920: signal is true;
	signal I38924: std_logic; attribute dont_touch of I38924: signal is true;
	signal I38931: std_logic; attribute dont_touch of I38931: signal is true;
	signal I38936: std_logic; attribute dont_touch of I38936: signal is true;
	signal I38940: std_logic; attribute dont_touch of I38940: signal is true;
	signal I38947: std_logic; attribute dont_touch of I38947: signal is true;
	signal I38951: std_logic; attribute dont_touch of I38951: signal is true;
	signal I38958: std_logic; attribute dont_touch of I38958: signal is true;
	signal I38975: std_logic; attribute dont_touch of I38975: signal is true;
	signal I38999: std_logic; attribute dont_touch of I38999: signal is true;
	signal I39002: std_logic; attribute dont_touch of I39002: signal is true;
	signal I39005: std_logic; attribute dont_touch of I39005: signal is true;
	signal I39008: std_logic; attribute dont_touch of I39008: signal is true;
	signal I39011: std_logic; attribute dont_touch of I39011: signal is true;
	signal I39014: std_logic; attribute dont_touch of I39014: signal is true;
	signal I39017: std_logic; attribute dont_touch of I39017: signal is true;
	signal I39020: std_logic; attribute dont_touch of I39020: signal is true;
	signal I39023: std_logic; attribute dont_touch of I39023: signal is true;
	signal I39026: std_logic; attribute dont_touch of I39026: signal is true;
	signal I39029: std_logic; attribute dont_touch of I39029: signal is true;
	signal I39032: std_logic; attribute dont_touch of I39032: signal is true;
	signal I39035: std_logic; attribute dont_touch of I39035: signal is true;
	signal I39038: std_logic; attribute dont_touch of I39038: signal is true;
	signal I39041: std_logic; attribute dont_touch of I39041: signal is true;
	signal I39044: std_logic; attribute dont_touch of I39044: signal is true;
	signal I39047: std_logic; attribute dont_touch of I39047: signal is true;
	signal I39050: std_logic; attribute dont_touch of I39050: signal is true;
	signal I39053: std_logic; attribute dont_touch of I39053: signal is true;
	signal I39056: std_logic; attribute dont_touch of I39056: signal is true;
	signal I39059: std_logic; attribute dont_touch of I39059: signal is true;
	signal I39062: std_logic; attribute dont_touch of I39062: signal is true;
	signal I39065: std_logic; attribute dont_touch of I39065: signal is true;
	signal I39068: std_logic; attribute dont_touch of I39068: signal is true;
	signal I39071: std_logic; attribute dont_touch of I39071: signal is true;
	signal I39074: std_logic; attribute dont_touch of I39074: signal is true;
	signal I39077: std_logic; attribute dont_touch of I39077: signal is true;
	signal I39080: std_logic; attribute dont_touch of I39080: signal is true;
	signal I39083: std_logic; attribute dont_touch of I39083: signal is true;
	signal I39086: std_logic; attribute dont_touch of I39086: signal is true;
	signal I39089: std_logic; attribute dont_touch of I39089: signal is true;
	signal I39121: std_logic; attribute dont_touch of I39121: signal is true;
	signal I39124: std_logic; attribute dont_touch of I39124: signal is true;
	signal I39127: std_logic; attribute dont_touch of I39127: signal is true;
	signal I39130: std_logic; attribute dont_touch of I39130: signal is true;
	signal I39133: std_logic; attribute dont_touch of I39133: signal is true;
	signal I39136: std_logic; attribute dont_touch of I39136: signal is true;
	signal I39139: std_logic; attribute dont_touch of I39139: signal is true;
	signal I39142: std_logic; attribute dont_touch of I39142: signal is true;
	signal I39145: std_logic; attribute dont_touch of I39145: signal is true;
	signal I39148: std_logic; attribute dont_touch of I39148: signal is true;
	signal I39151: std_logic; attribute dont_touch of I39151: signal is true;
	signal I39154: std_logic; attribute dont_touch of I39154: signal is true;
	signal I39157: std_logic; attribute dont_touch of I39157: signal is true;
	signal I39160: std_logic; attribute dont_touch of I39160: signal is true;
	signal I39164: std_logic; attribute dont_touch of I39164: signal is true;
	signal I39168: std_logic; attribute dont_touch of I39168: signal is true;
	signal I39234: std_logic; attribute dont_touch of I39234: signal is true;
	signal I39237: std_logic; attribute dont_touch of I39237: signal is true;
	signal I39240: std_logic; attribute dont_touch of I39240: signal is true;
	signal I39243: std_logic; attribute dont_touch of I39243: signal is true;
	signal I39246: std_logic; attribute dont_touch of I39246: signal is true;
	signal I39249: std_logic; attribute dont_touch of I39249: signal is true;
	signal I39252: std_logic; attribute dont_touch of I39252: signal is true;
	signal I39255: std_logic; attribute dont_touch of I39255: signal is true;
	signal I39258: std_logic; attribute dont_touch of I39258: signal is true;
	signal I39261: std_logic; attribute dont_touch of I39261: signal is true;
	signal I39264: std_logic; attribute dont_touch of I39264: signal is true;
	signal I39267: std_logic; attribute dont_touch of I39267: signal is true;
	signal I39270: std_logic; attribute dont_touch of I39270: signal is true;
	signal I39273: std_logic; attribute dont_touch of I39273: signal is true;
	signal I39276: std_logic; attribute dont_touch of I39276: signal is true;
	signal I39279: std_logic; attribute dont_touch of I39279: signal is true;
	signal I39323: std_logic; attribute dont_touch of I39323: signal is true;
	signal I39324: std_logic; attribute dont_touch of I39324: signal is true;
	signal I39325: std_logic; attribute dont_touch of I39325: signal is true;
	signal I39331: std_logic; attribute dont_touch of I39331: signal is true;
	signal I39332: std_logic; attribute dont_touch of I39332: signal is true;
	signal I39333: std_logic; attribute dont_touch of I39333: signal is true;
	signal I39339: std_logic; attribute dont_touch of I39339: signal is true;
	signal I39340: std_logic; attribute dont_touch of I39340: signal is true;
	signal I39341: std_logic; attribute dont_touch of I39341: signal is true;
	signal I39347: std_logic; attribute dont_touch of I39347: signal is true;
	signal I39348: std_logic; attribute dont_touch of I39348: signal is true;
	signal I39349: std_logic; attribute dont_touch of I39349: signal is true;
	signal I39359: std_logic; attribute dont_touch of I39359: signal is true;
	signal I39360: std_logic; attribute dont_touch of I39360: signal is true;
	signal I39361: std_logic; attribute dont_touch of I39361: signal is true;
	signal I39367: std_logic; attribute dont_touch of I39367: signal is true;
	signal I39368: std_logic; attribute dont_touch of I39368: signal is true;
	signal I39369: std_logic; attribute dont_touch of I39369: signal is true;
	signal I39375: std_logic; attribute dont_touch of I39375: signal is true;
	signal I39376: std_logic; attribute dont_touch of I39376: signal is true;
	signal I39377: std_logic; attribute dont_touch of I39377: signal is true;
	signal I39384: std_logic; attribute dont_touch of I39384: signal is true;
	signal I39385: std_logic; attribute dont_touch of I39385: signal is true;
	signal I39386: std_logic; attribute dont_touch of I39386: signal is true;
	signal I39391: std_logic; attribute dont_touch of I39391: signal is true;
	signal I39392: std_logic; attribute dont_touch of I39392: signal is true;
	signal I39393: std_logic; attribute dont_touch of I39393: signal is true;
	signal I39398: std_logic; attribute dont_touch of I39398: signal is true;
	signal I39401: std_logic; attribute dont_touch of I39401: signal is true;
	signal I39404: std_logic; attribute dont_touch of I39404: signal is true;
	signal I39407: std_logic; attribute dont_touch of I39407: signal is true;
	signal I39411: std_logic; attribute dont_touch of I39411: signal is true;
	signal I39414: std_logic; attribute dont_touch of I39414: signal is true;
	signal I39418: std_logic; attribute dont_touch of I39418: signal is true;
	signal I39423: std_logic; attribute dont_touch of I39423: signal is true;
	signal I39454: std_logic; attribute dont_touch of I39454: signal is true;
	signal I39457: std_logic; attribute dont_touch of I39457: signal is true;
	signal I39460: std_logic; attribute dont_touch of I39460: signal is true;
	signal I39463: std_logic; attribute dont_touch of I39463: signal is true;
	signal I39466: std_logic; attribute dont_touch of I39466: signal is true;
	signal I39469: std_logic; attribute dont_touch of I39469: signal is true;
	signal I39472: std_logic; attribute dont_touch of I39472: signal is true;
	signal I39475: std_logic; attribute dont_touch of I39475: signal is true;
	signal I39532: std_logic; attribute dont_touch of I39532: signal is true;
	signal I39533: std_logic; attribute dont_touch of I39533: signal is true;
	signal I39534: std_logic; attribute dont_touch of I39534: signal is true;
	signal I39539: std_logic; attribute dont_touch of I39539: signal is true;
	signal I39540: std_logic; attribute dont_touch of I39540: signal is true;
	signal I39541: std_logic; attribute dont_touch of I39541: signal is true;
	signal I39550: std_logic; attribute dont_touch of I39550: signal is true;
	signal I39573: std_logic; attribute dont_touch of I39573: signal is true;
	signal I39577: std_logic; attribute dont_touch of I39577: signal is true;
	signal I39585: std_logic; attribute dont_touch of I39585: signal is true;
	signal I39622: std_logic; attribute dont_touch of I39622: signal is true;
	signal I39625: std_logic; attribute dont_touch of I39625: signal is true;
	signal I39628: std_logic; attribute dont_touch of I39628: signal is true;
	signal I39631: std_logic; attribute dont_touch of I39631: signal is true;
	signal I39635: std_logic; attribute dont_touch of I39635: signal is true;
	signal I39638: std_logic; attribute dont_touch of I39638: signal is true;
	signal I39641: std_logic; attribute dont_touch of I39641: signal is true;
	signal I39647: std_logic; attribute dont_touch of I39647: signal is true;
	signal I39674: std_logic; attribute dont_touch of I39674: signal is true;
	signal I39689: std_logic; attribute dont_touch of I39689: signal is true;
	signal I39690: std_logic; attribute dont_touch of I39690: signal is true;
	signal I39691: std_logic; attribute dont_touch of I39691: signal is true;
	signal I39761: std_logic; attribute dont_touch of I39761: signal is true;
	signal I39764: std_logic; attribute dont_touch of I39764: signal is true;
	signal I39767: std_logic; attribute dont_touch of I39767: signal is true;
	signal I39770: std_logic; attribute dont_touch of I39770: signal is true;
	signal I39773: std_logic; attribute dont_touch of I39773: signal is true;
	signal I39776: std_logic; attribute dont_touch of I39776: signal is true;
	signal I39779: std_logic; attribute dont_touch of I39779: signal is true;
	signal I39782: std_logic; attribute dont_touch of I39782: signal is true;
	signal I39785: std_logic; attribute dont_touch of I39785: signal is true;
	signal I39788: std_logic; attribute dont_touch of I39788: signal is true;
	signal I39791: std_logic; attribute dont_touch of I39791: signal is true;
	signal I39794: std_logic; attribute dont_touch of I39794: signal is true;
	signal I39797: std_logic; attribute dont_touch of I39797: signal is true;
	signal I39800: std_logic; attribute dont_touch of I39800: signal is true;
	signal I39803: std_logic; attribute dont_touch of I39803: signal is true;
	signal I39806: std_logic; attribute dont_touch of I39806: signal is true;
	signal I39809: std_logic; attribute dont_touch of I39809: signal is true;
	signal I39812: std_logic; attribute dont_touch of I39812: signal is true;
	signal I39815: std_logic; attribute dont_touch of I39815: signal is true;
	signal I39818: std_logic; attribute dont_touch of I39818: signal is true;
	signal I39821: std_logic; attribute dont_touch of I39821: signal is true;
	signal I39825: std_logic; attribute dont_touch of I39825: signal is true;
	signal I39828: std_logic; attribute dont_touch of I39828: signal is true;
	signal I39832: std_logic; attribute dont_touch of I39832: signal is true;
	signal I39835: std_logic; attribute dont_touch of I39835: signal is true;
	signal I39840: std_logic; attribute dont_touch of I39840: signal is true;
	signal I39843: std_logic; attribute dont_touch of I39843: signal is true;
	signal I39848: std_logic; attribute dont_touch of I39848: signal is true;
	signal I39853: std_logic; attribute dont_touch of I39853: signal is true;
	signal I39856: std_logic; attribute dont_touch of I39856: signal is true;
	signal I39859: std_logic; attribute dont_touch of I39859: signal is true;
	signal I39863: std_logic; attribute dont_touch of I39863: signal is true;
	signal I39866: std_logic; attribute dont_touch of I39866: signal is true;
	signal I39870: std_logic; attribute dont_touch of I39870: signal is true;
	signal I39873: std_logic; attribute dont_touch of I39873: signal is true;
	signal I39878: std_logic; attribute dont_touch of I39878: signal is true;
	signal I39881: std_logic; attribute dont_touch of I39881: signal is true;
	signal I39886: std_logic; attribute dont_touch of I39886: signal is true;
	signal I39889: std_logic; attribute dont_touch of I39889: signal is true;
	signal I39892: std_logic; attribute dont_touch of I39892: signal is true;
	signal I39895: std_logic; attribute dont_touch of I39895: signal is true;
	signal I39899: std_logic; attribute dont_touch of I39899: signal is true;
	signal I39902: std_logic; attribute dont_touch of I39902: signal is true;
	signal I39906: std_logic; attribute dont_touch of I39906: signal is true;
	signal I39909: std_logic; attribute dont_touch of I39909: signal is true;
	signal I39913: std_logic; attribute dont_touch of I39913: signal is true;
	signal I39916: std_logic; attribute dont_touch of I39916: signal is true;
	signal I39919: std_logic; attribute dont_touch of I39919: signal is true;
	signal I39922: std_logic; attribute dont_touch of I39922: signal is true;
	signal I39926: std_logic; attribute dont_touch of I39926: signal is true;
	signal I39930: std_logic; attribute dont_touch of I39930: signal is true;
	signal I39933: std_logic; attribute dont_touch of I39933: signal is true;
	signal I39936: std_logic; attribute dont_touch of I39936: signal is true;
	signal I39939: std_logic; attribute dont_touch of I39939: signal is true;
	signal I39942: std_logic; attribute dont_touch of I39942: signal is true;
	signal I39945: std_logic; attribute dont_touch of I39945: signal is true;
	signal I39948: std_logic; attribute dont_touch of I39948: signal is true;
	signal I39951: std_logic; attribute dont_touch of I39951: signal is true;
	signal I39976: std_logic; attribute dont_touch of I39976: signal is true;
	signal I39982: std_logic; attribute dont_touch of I39982: signal is true;
	signal I39985: std_logic; attribute dont_touch of I39985: signal is true;
	signal I39991: std_logic; attribute dont_touch of I39991: signal is true;
	signal I39997: std_logic; attribute dont_touch of I39997: signal is true;
	signal I40002: std_logic; attribute dont_touch of I40002: signal is true;
	signal I40008: std_logic; attribute dont_touch of I40008: signal is true;
	signal I40016: std_logic; attribute dont_touch of I40016: signal is true;
	signal I40021: std_logic; attribute dont_touch of I40021: signal is true;
	signal I40027: std_logic; attribute dont_touch of I40027: signal is true;
	signal I40032: std_logic; attribute dont_touch of I40032: signal is true;
	signal I40039: std_logic; attribute dont_touch of I40039: signal is true;
	signal I40044: std_logic; attribute dont_touch of I40044: signal is true;
	signal I40051: std_logic; attribute dont_touch of I40051: signal is true;
	signal I40054: std_logic; attribute dont_touch of I40054: signal is true;
	signal I40059: std_logic; attribute dont_touch of I40059: signal is true;
	signal I40066: std_logic; attribute dont_touch of I40066: signal is true;
	signal I40071: std_logic; attribute dont_touch of I40071: signal is true;
	signal I40075: std_logic; attribute dont_touch of I40075: signal is true;
	signal I40078: std_logic; attribute dont_touch of I40078: signal is true;
	signal I40083: std_logic; attribute dont_touch of I40083: signal is true;
	signal I40086: std_logic; attribute dont_touch of I40086: signal is true;
	signal I40091: std_logic; attribute dont_touch of I40091: signal is true;
	signal I40098: std_logic; attribute dont_touch of I40098: signal is true;
	signal I40101: std_logic; attribute dont_touch of I40101: signal is true;
	signal I40104: std_logic; attribute dont_touch of I40104: signal is true;
	signal I40107: std_logic; attribute dont_touch of I40107: signal is true;
	signal I40110: std_logic; attribute dont_touch of I40110: signal is true;
	signal I40113: std_logic; attribute dont_touch of I40113: signal is true;
	signal I40116: std_logic; attribute dont_touch of I40116: signal is true;
	signal I40119: std_logic; attribute dont_touch of I40119: signal is true;
	signal I40122: std_logic; attribute dont_touch of I40122: signal is true;
	signal I40125: std_logic; attribute dont_touch of I40125: signal is true;
	signal I40128: std_logic; attribute dont_touch of I40128: signal is true;
	signal I40131: std_logic; attribute dont_touch of I40131: signal is true;
	signal I40134: std_logic; attribute dont_touch of I40134: signal is true;
	signal I40137: std_logic; attribute dont_touch of I40137: signal is true;
	signal I40140: std_logic; attribute dont_touch of I40140: signal is true;
	signal I40143: std_logic; attribute dont_touch of I40143: signal is true;
	signal I40146: std_logic; attribute dont_touch of I40146: signal is true;
	signal I40149: std_logic; attribute dont_touch of I40149: signal is true;
	signal I40152: std_logic; attribute dont_touch of I40152: signal is true;
	signal I40155: std_logic; attribute dont_touch of I40155: signal is true;
	signal I40158: std_logic; attribute dont_touch of I40158: signal is true;
	signal I40161: std_logic; attribute dont_touch of I40161: signal is true;
	signal I40164: std_logic; attribute dont_touch of I40164: signal is true;
	signal I40167: std_logic; attribute dont_touch of I40167: signal is true;
	signal I40170: std_logic; attribute dont_touch of I40170: signal is true;
	signal I40173: std_logic; attribute dont_touch of I40173: signal is true;
	signal I40176: std_logic; attribute dont_touch of I40176: signal is true;
	signal I40179: std_logic; attribute dont_touch of I40179: signal is true;
	signal I40182: std_logic; attribute dont_touch of I40182: signal is true;
	signal I40185: std_logic; attribute dont_touch of I40185: signal is true;
	signal I40188: std_logic; attribute dont_touch of I40188: signal is true;
	signal I40191: std_logic; attribute dont_touch of I40191: signal is true;
	signal I40194: std_logic; attribute dont_touch of I40194: signal is true;
	signal I40197: std_logic; attribute dont_touch of I40197: signal is true;
	signal I40200: std_logic; attribute dont_touch of I40200: signal is true;
	signal I40203: std_logic; attribute dont_touch of I40203: signal is true;
	signal I40206: std_logic; attribute dont_touch of I40206: signal is true;
	signal I40209: std_logic; attribute dont_touch of I40209: signal is true;
	signal I40212: std_logic; attribute dont_touch of I40212: signal is true;
	signal I40215: std_logic; attribute dont_touch of I40215: signal is true;
	signal I40218: std_logic; attribute dont_touch of I40218: signal is true;
	signal I40221: std_logic; attribute dont_touch of I40221: signal is true;
	signal I40224: std_logic; attribute dont_touch of I40224: signal is true;
	signal I40227: std_logic; attribute dont_touch of I40227: signal is true;
	signal I40230: std_logic; attribute dont_touch of I40230: signal is true;
	signal I40233: std_logic; attribute dont_touch of I40233: signal is true;
	signal I40236: std_logic; attribute dont_touch of I40236: signal is true;
	signal I40239: std_logic; attribute dont_touch of I40239: signal is true;
	signal I40242: std_logic; attribute dont_touch of I40242: signal is true;
	signal I40245: std_logic; attribute dont_touch of I40245: signal is true;
	signal I40248: std_logic; attribute dont_touch of I40248: signal is true;
	signal I40251: std_logic; attribute dont_touch of I40251: signal is true;
	signal I40254: std_logic; attribute dont_touch of I40254: signal is true;
	signal I40257: std_logic; attribute dont_touch of I40257: signal is true;
	signal I40260: std_logic; attribute dont_touch of I40260: signal is true;
	signal I40263: std_logic; attribute dont_touch of I40263: signal is true;
	signal I40266: std_logic; attribute dont_touch of I40266: signal is true;
	signal I40269: std_logic; attribute dont_touch of I40269: signal is true;
	signal I40272: std_logic; attribute dont_touch of I40272: signal is true;
	signal I40275: std_logic; attribute dont_touch of I40275: signal is true;
	signal I40288: std_logic; attribute dont_touch of I40288: signal is true;
	signal I40291: std_logic; attribute dont_touch of I40291: signal is true;
	signal I40294: std_logic; attribute dont_touch of I40294: signal is true;
	signal I40297: std_logic; attribute dont_touch of I40297: signal is true;
	signal I40300: std_logic; attribute dont_touch of I40300: signal is true;
	signal I40303: std_logic; attribute dont_touch of I40303: signal is true;
	signal I40307: std_logic; attribute dont_touch of I40307: signal is true;
	signal I40310: std_logic; attribute dont_touch of I40310: signal is true;
	signal I40313: std_logic; attribute dont_touch of I40313: signal is true;
	signal I40317: std_logic; attribute dont_touch of I40317: signal is true;
	signal I40320: std_logic; attribute dont_touch of I40320: signal is true;
	signal I40326: std_logic; attribute dont_touch of I40326: signal is true;
	signal I40420: std_logic; attribute dont_touch of I40420: signal is true;
	signal I40423: std_logic; attribute dont_touch of I40423: signal is true;
	signal I40426: std_logic; attribute dont_touch of I40426: signal is true;
	signal I40429: std_logic; attribute dont_touch of I40429: signal is true;
	signal I40432: std_logic; attribute dont_touch of I40432: signal is true;
	signal I40435: std_logic; attribute dont_touch of I40435: signal is true;
	signal I40438: std_logic; attribute dont_touch of I40438: signal is true;
	signal I40441: std_logic; attribute dont_touch of I40441: signal is true;
	signal I40444: std_logic; attribute dont_touch of I40444: signal is true;
	signal I40447: std_logic; attribute dont_touch of I40447: signal is true;
	signal I40450: std_logic; attribute dont_touch of I40450: signal is true;
	signal I40453: std_logic; attribute dont_touch of I40453: signal is true;
	signal I40456: std_logic; attribute dont_touch of I40456: signal is true;
	signal I40459: std_logic; attribute dont_touch of I40459: signal is true;
	signal I40462: std_logic; attribute dont_touch of I40462: signal is true;
	signal I40465: std_logic; attribute dont_touch of I40465: signal is true;
	signal I40468: std_logic; attribute dont_touch of I40468: signal is true;
	signal I40471: std_logic; attribute dont_touch of I40471: signal is true;
	signal I40475: std_logic; attribute dont_touch of I40475: signal is true;
	signal I40478: std_logic; attribute dont_touch of I40478: signal is true;
	signal I40481: std_logic; attribute dont_touch of I40481: signal is true;
	signal I40484: std_logic; attribute dont_touch of I40484: signal is true;
	signal I40487: std_logic; attribute dont_touch of I40487: signal is true;
	signal I40490: std_logic; attribute dont_touch of I40490: signal is true;
	signal I40495: std_logic; attribute dont_touch of I40495: signal is true;
	signal I40498: std_logic; attribute dont_touch of I40498: signal is true;
	signal I40501: std_logic; attribute dont_touch of I40501: signal is true;
	signal I40504: std_logic; attribute dont_touch of I40504: signal is true;
	signal I40507: std_logic; attribute dont_touch of I40507: signal is true;
	signal I40510: std_logic; attribute dont_touch of I40510: signal is true;
	signal I40515: std_logic; attribute dont_touch of I40515: signal is true;
	signal I40518: std_logic; attribute dont_touch of I40518: signal is true;
	signal I40521: std_logic; attribute dont_touch of I40521: signal is true;
	signal I40524: std_logic; attribute dont_touch of I40524: signal is true;
	signal I40527: std_logic; attribute dont_touch of I40527: signal is true;
	signal I40531: std_logic; attribute dont_touch of I40531: signal is true;
	signal I40534: std_logic; attribute dont_touch of I40534: signal is true;
	signal I40537: std_logic; attribute dont_touch of I40537: signal is true;
	signal I40542: std_logic; attribute dont_touch of I40542: signal is true;
	signal I40555: std_logic; attribute dont_touch of I40555: signal is true;
	signal I40558: std_logic; attribute dont_touch of I40558: signal is true;
	signal I40559: std_logic; attribute dont_touch of I40559: signal is true;
	signal I40560: std_logic; attribute dont_touch of I40560: signal is true;
	signal I40565: std_logic; attribute dont_touch of I40565: signal is true;
	signal I40568: std_logic; attribute dont_touch of I40568: signal is true;
	signal I40571: std_logic; attribute dont_touch of I40571: signal is true;
	signal I40572: std_logic; attribute dont_touch of I40572: signal is true;
	signal I40573: std_logic; attribute dont_touch of I40573: signal is true;
	signal I40578: std_logic; attribute dont_touch of I40578: signal is true;
	signal I40581: std_logic; attribute dont_touch of I40581: signal is true;
	signal I40584: std_logic; attribute dont_touch of I40584: signal is true;
	signal I40587: std_logic; attribute dont_touch of I40587: signal is true;
	signal I40588: std_logic; attribute dont_touch of I40588: signal is true;
	signal I40589: std_logic; attribute dont_touch of I40589: signal is true;
	signal I40594: std_logic; attribute dont_touch of I40594: signal is true;
	signal I40597: std_logic; attribute dont_touch of I40597: signal is true;
	signal I40600: std_logic; attribute dont_touch of I40600: signal is true;
	signal I40603: std_logic; attribute dont_touch of I40603: signal is true;
	signal I40604: std_logic; attribute dont_touch of I40604: signal is true;
	signal I40605: std_logic; attribute dont_touch of I40605: signal is true;
	signal I40611: std_logic; attribute dont_touch of I40611: signal is true;
	signal I40614: std_logic; attribute dont_touch of I40614: signal is true;
	signal I40618: std_logic; attribute dont_touch of I40618: signal is true;
	signal I40627: std_logic; attribute dont_touch of I40627: signal is true;
	signal I40628: std_logic; attribute dont_touch of I40628: signal is true;
	signal I40629: std_logic; attribute dont_touch of I40629: signal is true;
	signal I40634: std_logic; attribute dont_touch of I40634: signal is true;
	signal I40637: std_logic; attribute dont_touch of I40637: signal is true;
	signal I40640: std_logic; attribute dont_touch of I40640: signal is true;
	signal I40643: std_logic; attribute dont_touch of I40643: signal is true;
	signal I40647: std_logic; attribute dont_touch of I40647: signal is true;
	signal I40651: std_logic; attribute dont_touch of I40651: signal is true;
	signal I40654: std_logic; attribute dont_touch of I40654: signal is true;
	signal I40658: std_logic; attribute dont_touch of I40658: signal is true;
	signal I40661: std_logic; attribute dont_touch of I40661: signal is true;
	signal I40664: std_logic; attribute dont_touch of I40664: signal is true;
	signal I40667: std_logic; attribute dont_touch of I40667: signal is true;
	signal I40670: std_logic; attribute dont_touch of I40670: signal is true;
	signal I40673: std_logic; attribute dont_touch of I40673: signal is true;
	signal I40676: std_logic; attribute dont_touch of I40676: signal is true;
	signal I40679: std_logic; attribute dont_touch of I40679: signal is true;
	signal I40682: std_logic; attribute dont_touch of I40682: signal is true;
	signal I40685: std_logic; attribute dont_touch of I40685: signal is true;
	signal I40688: std_logic; attribute dont_touch of I40688: signal is true;
	signal I40691: std_logic; attribute dont_touch of I40691: signal is true;
	signal I40694: std_logic; attribute dont_touch of I40694: signal is true;
	signal I40697: std_logic; attribute dont_touch of I40697: signal is true;
	signal I40700: std_logic; attribute dont_touch of I40700: signal is true;
	signal I40703: std_logic; attribute dont_touch of I40703: signal is true;
	signal I40706: std_logic; attribute dont_touch of I40706: signal is true;
	signal I40709: std_logic; attribute dont_touch of I40709: signal is true;
	signal I40712: std_logic; attribute dont_touch of I40712: signal is true;
	signal I40715: std_logic; attribute dont_touch of I40715: signal is true;
	signal I40718: std_logic; attribute dont_touch of I40718: signal is true;
	signal I40721: std_logic; attribute dont_touch of I40721: signal is true;
	signal I40724: std_logic; attribute dont_touch of I40724: signal is true;
	signal I40727: std_logic; attribute dont_touch of I40727: signal is true;
	signal I40730: std_logic; attribute dont_touch of I40730: signal is true;
	signal I40733: std_logic; attribute dont_touch of I40733: signal is true;
	signal I40736: std_logic; attribute dont_touch of I40736: signal is true;
	signal I40739: std_logic; attribute dont_touch of I40739: signal is true;
	signal I40742: std_logic; attribute dont_touch of I40742: signal is true;
	signal I40745: std_logic; attribute dont_touch of I40745: signal is true;
	signal I40748: std_logic; attribute dont_touch of I40748: signal is true;
	signal I40751: std_logic; attribute dont_touch of I40751: signal is true;
	signal I40754: std_logic; attribute dont_touch of I40754: signal is true;
	signal I40757: std_logic; attribute dont_touch of I40757: signal is true;
	signal I40760: std_logic; attribute dont_touch of I40760: signal is true;
	signal I40763: std_logic; attribute dont_touch of I40763: signal is true;
	signal I40766: std_logic; attribute dont_touch of I40766: signal is true;
	signal I40769: std_logic; attribute dont_touch of I40769: signal is true;
	signal I40772: std_logic; attribute dont_touch of I40772: signal is true;
	signal I40775: std_logic; attribute dont_touch of I40775: signal is true;
	signal I40778: std_logic; attribute dont_touch of I40778: signal is true;
	signal I40781: std_logic; attribute dont_touch of I40781: signal is true;
	signal I40784: std_logic; attribute dont_touch of I40784: signal is true;
	signal I40787: std_logic; attribute dont_touch of I40787: signal is true;
	signal I40790: std_logic; attribute dont_touch of I40790: signal is true;
	signal I40793: std_logic; attribute dont_touch of I40793: signal is true;
	signal I40796: std_logic; attribute dont_touch of I40796: signal is true;
	signal I40799: std_logic; attribute dont_touch of I40799: signal is true;
	signal I40802: std_logic; attribute dont_touch of I40802: signal is true;
	signal I40805: std_logic; attribute dont_touch of I40805: signal is true;
	signal I40808: std_logic; attribute dont_touch of I40808: signal is true;
	signal I40811: std_logic; attribute dont_touch of I40811: signal is true;
	signal I40814: std_logic; attribute dont_touch of I40814: signal is true;
	signal I40817: std_logic; attribute dont_touch of I40817: signal is true;
	signal I40820: std_logic; attribute dont_touch of I40820: signal is true;
	signal I40823: std_logic; attribute dont_touch of I40823: signal is true;
	signal I40826: std_logic; attribute dont_touch of I40826: signal is true;
	signal I40829: std_logic; attribute dont_touch of I40829: signal is true;
	signal I40832: std_logic; attribute dont_touch of I40832: signal is true;
	signal I40835: std_logic; attribute dont_touch of I40835: signal is true;
	signal I40838: std_logic; attribute dont_touch of I40838: signal is true;
	signal I40841: std_logic; attribute dont_touch of I40841: signal is true;
	signal I40844: std_logic; attribute dont_touch of I40844: signal is true;
	signal I40847: std_logic; attribute dont_touch of I40847: signal is true;
	signal I40850: std_logic; attribute dont_touch of I40850: signal is true;
	signal I40853: std_logic; attribute dont_touch of I40853: signal is true;
	signal I40856: std_logic; attribute dont_touch of I40856: signal is true;
	signal I40859: std_logic; attribute dont_touch of I40859: signal is true;
	signal I40862: std_logic; attribute dont_touch of I40862: signal is true;
	signal I40865: std_logic; attribute dont_touch of I40865: signal is true;
	signal I40868: std_logic; attribute dont_touch of I40868: signal is true;
	signal I40871: std_logic; attribute dont_touch of I40871: signal is true;
	signal I40874: std_logic; attribute dont_touch of I40874: signal is true;
	signal I40877: std_logic; attribute dont_touch of I40877: signal is true;
	signal I40880: std_logic; attribute dont_touch of I40880: signal is true;
	signal I40883: std_logic; attribute dont_touch of I40883: signal is true;
	signal I40886: std_logic; attribute dont_touch of I40886: signal is true;
	signal I40889: std_logic; attribute dont_touch of I40889: signal is true;
	signal I40892: std_logic; attribute dont_touch of I40892: signal is true;
	signal I40895: std_logic; attribute dont_touch of I40895: signal is true;
	signal I40898: std_logic; attribute dont_touch of I40898: signal is true;
	signal I40901: std_logic; attribute dont_touch of I40901: signal is true;
	signal I40904: std_logic; attribute dont_touch of I40904: signal is true;
	signal I40907: std_logic; attribute dont_touch of I40907: signal is true;
	signal I40910: std_logic; attribute dont_touch of I40910: signal is true;
	signal I40913: std_logic; attribute dont_touch of I40913: signal is true;
	signal I40916: std_logic; attribute dont_touch of I40916: signal is true;
	signal I40919: std_logic; attribute dont_touch of I40919: signal is true;
	signal I40922: std_logic; attribute dont_touch of I40922: signal is true;
	signal I40925: std_logic; attribute dont_touch of I40925: signal is true;
	signal I40928: std_logic; attribute dont_touch of I40928: signal is true;
	signal I40931: std_logic; attribute dont_touch of I40931: signal is true;
	signal I40934: std_logic; attribute dont_touch of I40934: signal is true;
	signal I40937: std_logic; attribute dont_touch of I40937: signal is true;
	signal I40940: std_logic; attribute dont_touch of I40940: signal is true;
	signal I40943: std_logic; attribute dont_touch of I40943: signal is true;
	signal I40946: std_logic; attribute dont_touch of I40946: signal is true;
	signal I40949: std_logic; attribute dont_touch of I40949: signal is true;
	signal I40952: std_logic; attribute dont_touch of I40952: signal is true;
	signal I40955: std_logic; attribute dont_touch of I40955: signal is true;
	signal I40958: std_logic; attribute dont_touch of I40958: signal is true;
	signal I40961: std_logic; attribute dont_touch of I40961: signal is true;
	signal I40964: std_logic; attribute dont_touch of I40964: signal is true;
	signal I40967: std_logic; attribute dont_touch of I40967: signal is true;
	signal I40970: std_logic; attribute dont_touch of I40970: signal is true;
	signal I40973: std_logic; attribute dont_touch of I40973: signal is true;
	signal I40976: std_logic; attribute dont_touch of I40976: signal is true;
	signal I40979: std_logic; attribute dont_touch of I40979: signal is true;
	signal I40982: std_logic; attribute dont_touch of I40982: signal is true;
	signal I40985: std_logic; attribute dont_touch of I40985: signal is true;
	signal I40988: std_logic; attribute dont_touch of I40988: signal is true;
	signal I40991: std_logic; attribute dont_touch of I40991: signal is true;
	signal I40994: std_logic; attribute dont_touch of I40994: signal is true;
	signal I40997: std_logic; attribute dont_touch of I40997: signal is true;
	signal I41010: std_logic; attribute dont_touch of I41010: signal is true;
	signal I41011: std_logic; attribute dont_touch of I41011: signal is true;
	signal I41012: std_logic; attribute dont_touch of I41012: signal is true;
	signal I41017: std_logic; attribute dont_touch of I41017: signal is true;
	signal I41018: std_logic; attribute dont_touch of I41018: signal is true;
	signal I41019: std_logic; attribute dont_touch of I41019: signal is true;
	signal I41024: std_logic; attribute dont_touch of I41024: signal is true;
	signal I41035: std_logic; attribute dont_touch of I41035: signal is true;
	signal I41038: std_logic; attribute dont_touch of I41038: signal is true;
	signal I41041: std_logic; attribute dont_touch of I41041: signal is true;
	signal I41044: std_logic; attribute dont_touch of I41044: signal is true;
	signal I41047: std_logic; attribute dont_touch of I41047: signal is true;
	signal I41050: std_logic; attribute dont_touch of I41050: signal is true;
	signal I41053: std_logic; attribute dont_touch of I41053: signal is true;
	signal I41064: std_logic; attribute dont_touch of I41064: signal is true;
	signal I41065: std_logic; attribute dont_touch of I41065: signal is true;
	signal I41066: std_logic; attribute dont_touch of I41066: signal is true;
	signal I41090: std_logic; attribute dont_touch of I41090: signal is true;
	signal I41093: std_logic; attribute dont_touch of I41093: signal is true;
	signal I41096: std_logic; attribute dont_touch of I41096: signal is true;
	signal I41099: std_logic; attribute dont_touch of I41099: signal is true;
	signal I41102: std_logic; attribute dont_touch of I41102: signal is true;
	signal I41105: std_logic; attribute dont_touch of I41105: signal is true;
	signal I41108: std_logic; attribute dont_touch of I41108: signal is true;
	signal I41111: std_logic; attribute dont_touch of I41111: signal is true;
	signal I41114: std_logic; attribute dont_touch of I41114: signal is true;
	signal I41117: std_logic; attribute dont_touch of I41117: signal is true;
	signal I41120: std_logic; attribute dont_touch of I41120: signal is true;
	signal I41123: std_logic; attribute dont_touch of I41123: signal is true;
	signal I41126: std_logic; attribute dont_touch of I41126: signal is true;
	signal I41129: std_logic; attribute dont_touch of I41129: signal is true;
	signal I41132: std_logic; attribute dont_touch of I41132: signal is true;
	signal I41135: std_logic; attribute dont_touch of I41135: signal is true;
	signal I41138: std_logic; attribute dont_touch of I41138: signal is true;
	signal I41141: std_logic; attribute dont_touch of I41141: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			G1<=G20594;
			G2<=G20592;
			G5<=G20590;
			G8<=G20591;
			G11<=G20608;
			G14<=G20589;
			G17<=G20607;
			G20<=G20606;
			G23<=G20605;
			G26<=G20604;
			G27<=G20599;
			G30<=G20600;
			G33<=G20601;
			G36<=G20602;
			G39<=G20598;
			G42<=G20597;
			G45<=G20596;
			G48<=G20595;
			G52<=G29794;
			G56<=G29627;
			G61<=G29413;
			G65<=G29131;
			G70<=G28673;
			G74<=G28206;
			G79<=G27683;
			G83<=G27189;
			G88<=G26678;
			G92<=G25983;
			G97<=G2854;
			G101<=G2851;
			G105<=G2848;
			G109<=G2845;
			G113<=G2842;
			G117<=G2839;
			G121<=G2836;
			G125<=G2833;
			G129<=G24261;
			G130<=G24259;
			G131<=G24260;
			G132<=G24264;
			G133<=G24262;
			G134<=G24263;
			G135<=G138;
			G138<=G13405;
			G141<=G24267;
			G142<=G24265;
			G143<=G24266;
			G144<=G24270;
			G145<=G24268;
			G146<=G24269;
			G147<=G24273;
			G148<=G24271;
			G149<=G24272;
			G150<=G24276;
			G151<=G24274;
			G152<=G24275;
			G153<=G24279;
			G154<=G24277;
			G155<=G24278;
			G156<=G24282;
			G157<=G24280;
			G158<=G24281;
			G159<=G24285;
			G160<=G24283;
			G161<=G24284;
			G162<=G24288;
			G163<=G24286;
			G164<=G24287;
			G165<=G135;
			G168<=G26681;
			G169<=G26679;
			G170<=G26680;
			G171<=G26684;
			G172<=G26682;
			G173<=G26683;
			G174<=G26687;
			G175<=G26685;
			G176<=G26686;
			G177<=G26690;
			G178<=G26688;
			G179<=G26689;
			G180<=G20555;
			G181<=G182;
			G182<=G180;
			G185<=G29657;
			G186<=G30506;
			G189<=G30507;
			G192<=G30508;
			G195<=G30836;
			G198<=G30837;
			G201<=G30838;
			G204<=G30509;
			G207<=G30510;
			G210<=G30511;
			G213<=G30512;
			G216<=G30513;
			G219<=G30514;
			G222<=G30839;
			G225<=G30840;
			G228<=G30841;
			G231<=G30842;
			G234<=G30843;
			G237<=G30844;
			G240<=G30845;
			G243<=G30846;
			G246<=G30847;
			G249<=G30515;
			G252<=G30516;
			G255<=G30517;
			G258<=G30518;
			G261<=G30519;
			G264<=G30520;
			G267<=G30848;
			G270<=G30849;
			G273<=G30850;
			G276<=G13406;
			G279<=G454;
			G280<=G11491;
			G281<=G280;
			G282<=G11492;
			G283<=G282;
			G284<=G11493;
			G285<=G284;
			G286<=G11494;
			G287<=G286;
			G288<=G11495;
			G289<=G288;
			G290<=G13407;
			G291<=G290;
			G294<=G23153;
			G295<=G23152;
			G296<=G23151;
			G297<=G23150;
			G298<=G27190;
			G299<=G19012;
			G300<=G25130;
			G301<=G19013;
			G302<=G19014;
			G303<=G19015;
			G304<=G19016;
			G305<=G23148;
			G308<=G23149;
			G309<=G11496;
			G312<=G29795;
			G313<=G29796;
			G314<=G29797;
			G315<=G30851;
			G316<=G30852;
			G317<=G30853;
			G318<=G30710;
			G319<=G30711;
			G320<=G30712;
			G321<=G29630;
			G322<=G29628;
			G323<=G29629;
			G324<=G397;
			G325<=G13408;
			G331<=G325;
			G337<=G331;
			G342<=G11497;
			G343<=G28208;
			G346<=G28209;
			G349<=G342;
			G350<=G11498;
			G351<=G350;
			G352<=G11499;
			G353<=G352;
			G354<=G28207;
			G357<=G11500;
			G358<=G28211;
			G361<=G28212;
			G364<=G357;
			G365<=G11501;
			G366<=G365;
			G367<=G11502;
			G368<=G367;
			G369<=G28210;
			G372<=G11503;
			G373<=G28214;
			G376<=G28215;
			G379<=G372;
			G380<=G11504;
			G381<=G380;
			G382<=G11505;
			G383<=G382;
			G384<=G28213;
			G387<=G11506;
			G388<=G28217;
			G391<=G28218;
			G394<=G387;
			G395<=G11507;
			G396<=G395;
			G397<=G11508;
			G398<=G28216;
			G401<=G405;
			G402<=G27193;
			G403<=G27191;
			G404<=G27192;
			G405<=G276;
			G408<=G29414;
			G411<=G29415;
			G414<=G29416;
			G417<=G29631;
			G420<=G29632;
			G423<=G29633;
			G426<=G29419;
			G427<=G29417;
			G428<=G29418;
			G429<=G27684;
			G432<=G27685;
			G435<=G27686;
			G438<=G27687;
			G441<=G27688;
			G444<=G27689;
			G447<=G28676;
			G448<=G28674;
			G449<=G28675;
			G450<=G11509;
			G451<=G450;
			G452<=G11510;
			G453<=G452;
			G454<=G11511;
			G455<=G25139;
			G458<=G25131;
			G461<=G25132;
			G464<=G24291;
			G465<=G25133;
			G468<=G25134;
			G471<=G25135;
			G474<=G13409;
			G477<=G25136;
			G478<=G25137;
			G479<=G25138;
			G480<=G24289;
			G481<=G474;
			G484<=G24290;
			G485<=G481;
			G486<=G24292;
			G487<=G24293;
			G488<=G24294;
			G489<=G568;
			G490<=G27194;
			G493<=G27195;
			G496<=G27196;
			G499<=G549;
			G506<=G8284;
			G507<=G24295;
			G508<=G19017;
			G509<=G19018;
			G510<=G20557;
			G513<=G16467;
			G514<=G19019;
			G515<=G19020;
			G516<=G23158;
			G517<=G23157;
			G518<=G23156;
			G519<=G23155;
			G520<=G23154;
			G523<=G513;
			G524<=G523;
			G525<=G520;
			G528<=G16468;
			G529<=G13410;
			G530<=G13411;
			G531<=G13412;
			G532<=G13413;
			G533<=G13414;
			G534<=G13415;
			G535<=G528;
			G536<=G13416;
			G537<=G13417;
			G538<=G25984;
			G541<=G13418;
			G542<=G535;
			G543<=G19021;
			G544<=G543;
			G545<=G13419;
			G548<=G23159;
			G549<=G19022;
			G550<=G551;
			G551<=G545;
			G554<=G23160;
			G557<=G20556;
			G558<=G19023;
			G559<=G558;
			G564<=G11512;
			G565<=G574;
			G566<=G11513;
			G567<=G566;
			G568<=G11514;
			G569<=G564;
			G570<=G11515;
			G571<=G570;
			G572<=G11516;
			G573<=G572;
			G574<=G11517;
			G575<=G28221;
			G576<=G28219;
			G577<=G28220;
			G578<=G28224;
			G579<=G28222;
			G580<=G28223;
			G581<=G28227;
			G582<=G28225;
			G583<=G28226;
			G584<=G28230;
			G585<=G28228;
			G586<=G28229;
			G587<=G25985;
			G590<=G25986;
			G593<=G25987;
			G596<=G25988;
			G599<=G25989;
			G602<=G25990;
			G605<=G29132;
			G608<=G29133;
			G611<=G29134;
			G614<=G29135;
			G617<=G29136;
			G620<=G29137;
			G623<=G13420;
			G626<=G623;
			G629<=G626;
			G630<=G20558;
			G633<=G24296;
			G640<=G23161;
			G646<=G25991;
			G653<=G25140;
			G659<=G21943;
			G660<=G26691;
			G666<=G27690;
			G672<=G27197;
			G679<=G28231;
			G686<=G28677;
			G692<=G29138;
			G698<=G23164;
			G699<=G23162;
			G700<=G23163;
			G701<=G23167;
			G702<=G23165;
			G703<=G23166;
			G704<=G23170;
			G705<=G23168;
			G706<=G23169;
			G707<=G23173;
			G708<=G23171;
			G709<=G23172;
			G710<=G23176;
			G711<=G23174;
			G712<=G23175;
			G713<=G23179;
			G714<=G23177;
			G715<=G23178;
			G716<=G23182;
			G717<=G23180;
			G718<=G23181;
			G719<=G23185;
			G720<=G23183;
			G721<=G23184;
			G722<=G23188;
			G723<=G23186;
			G724<=G23187;
			G725<=G23191;
			G726<=G23189;
			G727<=G23190;
			G728<=G23194;
			G729<=G23192;
			G730<=G23193;
			G731<=G23197;
			G732<=G23195;
			G733<=G23196;
			G734<=G26694;
			G735<=G26692;
			G736<=G26693;
			G737<=G24299;
			G738<=G24297;
			G739<=G24298;
			G740<=G29798;
			G744<=G29634;
			G749<=G29420;
			G753<=G29139;
			G758<=G28678;
			G762<=G28232;
			G767<=G27691;
			G771<=G27198;
			G776<=G26695;
			G780<=G25992;
			G785<=G2827;
			G789<=G2824;
			G793<=G2821;
			G797<=G2818;
			G801<=G2870;
			G805<=G2867;
			G809<=G2864;
			G813<=G2861;
			G817<=G24302;
			G818<=G24300;
			G819<=G24301;
			G820<=G24305;
			G821<=G24303;
			G822<=G24304;
			G823<=G826;
			G826<=G13421;
			G829<=G24308;
			G830<=G24306;
			G831<=G24307;
			G832<=G24311;
			G833<=G24309;
			G834<=G24310;
			G835<=G24314;
			G836<=G24312;
			G837<=G24313;
			G838<=G24317;
			G839<=G24315;
			G840<=G24316;
			G841<=G24320;
			G842<=G24318;
			G843<=G24319;
			G844<=G24323;
			G845<=G24321;
			G846<=G24322;
			G847<=G24326;
			G848<=G24324;
			G849<=G24325;
			G850<=G24329;
			G851<=G24327;
			G852<=G24328;
			G853<=G823;
			G856<=G26698;
			G857<=G26696;
			G858<=G26697;
			G859<=G26701;
			G860<=G26699;
			G861<=G26700;
			G862<=G26704;
			G863<=G26702;
			G864<=G26703;
			G865<=G26707;
			G866<=G26705;
			G867<=G26706;
			G868<=G20559;
			G869<=G870;
			G870<=G868;
			G873<=G30521;
			G876<=G30522;
			G879<=G30523;
			G882<=G30854;
			G885<=G30855;
			G888<=G30856;
			G891<=G30524;
			G894<=G30525;
			G897<=G30526;
			G900<=G30527;
			G903<=G30528;
			G906<=G30529;
			G909<=G30857;
			G912<=G30858;
			G915<=G30859;
			G918<=G30860;
			G921<=G30861;
			G924<=G30862;
			G927<=G30863;
			G930<=G30864;
			G933<=G30865;
			G936<=G30530;
			G939<=G30531;
			G942<=G30532;
			G945<=G30533;
			G948<=G30534;
			G951<=G30535;
			G954<=G30866;
			G957<=G30867;
			G960<=G30868;
			G963<=G13422;
			G966<=G1141;
			G967<=G11518;
			G968<=G967;
			G969<=G11519;
			G970<=G969;
			G971<=G11520;
			G972<=G971;
			G973<=G11521;
			G974<=G973;
			G975<=G11522;
			G976<=G975;
			G977<=G13423;
			G978<=G977;
			G981<=G27205;
			G982<=G27204;
			G983<=G27203;
			G984<=G27202;
			G985<=G27199;
			G986<=G19024;
			G987<=G25141;
			G988<=G19025;
			G989<=G19026;
			G990<=G19027;
			G991<=G19028;
			G992<=G27200;
			G995<=G27201;
			G996<=G11523;
			G999<=G29799;
			G1000<=G29800;
			G1001<=G29801;
			G1002<=G30869;
			G1003<=G30870;
			G1004<=G30871;
			G1005<=G30713;
			G1006<=G30714;
			G1007<=G30715;
			G1008<=G29637;
			G1009<=G29635;
			G1010<=G29636;
			G1011<=G1084;
			G1012<=G13424;
			G1018<=G1012;
			G1024<=G1018;
			G1029<=G11524;
			G1030<=G28234;
			G1033<=G28235;
			G1036<=G1029;
			G1037<=G11525;
			G1038<=G1037;
			G1039<=G11526;
			G1040<=G1039;
			G1041<=G28233;
			G1044<=G11527;
			G1045<=G28237;
			G1048<=G28238;
			G1051<=G1044;
			G1052<=G11528;
			G1053<=G1052;
			G1054<=G11529;
			G1055<=G1054;
			G1056<=G28236;
			G1059<=G11530;
			G1060<=G28240;
			G1063<=G28241;
			G1066<=G1059;
			G1067<=G11531;
			G1068<=G1067;
			G1069<=G11532;
			G1070<=G1069;
			G1071<=G28239;
			G1074<=G11533;
			G1075<=G28243;
			G1078<=G28244;
			G1081<=G1074;
			G1082<=G11534;
			G1083<=G1082;
			G1084<=G11535;
			G1085<=G28242;
			G1088<=G1092;
			G1089<=G27208;
			G1090<=G27206;
			G1091<=G27207;
			G1092<=G963;
			G1095<=G29421;
			G1098<=G29422;
			G1101<=G29423;
			G1104<=G29638;
			G1107<=G29639;
			G1110<=G29640;
			G1113<=G29426;
			G1114<=G29424;
			G1115<=G29425;
			G1116<=G27692;
			G1119<=G27693;
			G1122<=G27694;
			G1125<=G27695;
			G1128<=G27696;
			G1131<=G27697;
			G1134<=G28681;
			G1135<=G28679;
			G1136<=G28680;
			G1137<=G11536;
			G1138<=G1137;
			G1139<=G11537;
			G1140<=G1139;
			G1141<=G11538;
			G1142<=G25150;
			G1145<=G25142;
			G1148<=G25143;
			G1151<=G24332;
			G1152<=G25144;
			G1155<=G25145;
			G1158<=G25146;
			G1161<=G13425;
			G1164<=G25147;
			G1165<=G25148;
			G1166<=G25149;
			G1167<=G24330;
			G1168<=G1161;
			G1171<=G24331;
			G1172<=G1168;
			G1173<=G24333;
			G1174<=G24334;
			G1175<=G24335;
			G1176<=G1254;
			G1177<=G27209;
			G1180<=G27210;
			G1183<=G27211;
			G1186<=G1235;
			G1192<=G8293;
			G1193<=G24336;
			G1194<=G19029;
			G1195<=G19030;
			G1196<=G20561;
			G1199<=G16469;
			G1200<=G19031;
			G1201<=G19032;
			G1202<=G27216;
			G1203<=G27215;
			G1204<=G27214;
			G1205<=G27213;
			G1206<=G27212;
			G1209<=G1199;
			G1210<=G1209;
			G1211<=G1206;
			G1214<=G16470;
			G1215<=G13426;
			G1216<=G13427;
			G1217<=G13428;
			G1218<=G13429;
			G1219<=G13430;
			G1220<=G13431;
			G1221<=G1214;
			G1222<=G13432;
			G1223<=G13433;
			G1224<=G25993;
			G1227<=G13434;
			G1228<=G1221;
			G1229<=G19033;
			G1230<=G1229;
			G1231<=G13435;
			G1234<=G27217;
			G1235<=G19034;
			G1236<=G1237;
			G1237<=G1231;
			G1240<=G23198;
			G1243<=G20560;
			G1244<=G19035;
			G1245<=G1244;
			G1250<=G11539;
			G1251<=G1260;
			G1252<=G11540;
			G1253<=G1252;
			G1254<=G11541;
			G1255<=G1250;
			G1256<=G11542;
			G1257<=G1256;
			G1258<=G11543;
			G1259<=G1258;
			G1260<=G11544;
			G1261<=G28247;
			G1262<=G28245;
			G1263<=G28246;
			G1264<=G28250;
			G1265<=G28248;
			G1266<=G28249;
			G1267<=G28253;
			G1268<=G28251;
			G1269<=G28252;
			G1270<=G28256;
			G1271<=G28254;
			G1272<=G28255;
			G1273<=G25994;
			G1276<=G25995;
			G1279<=G25996;
			G1282<=G25997;
			G1285<=G25998;
			G1288<=G25999;
			G1291<=G29140;
			G1294<=G29141;
			G1297<=G29142;
			G1300<=G29143;
			G1303<=G29144;
			G1306<=G29145;
			G1309<=G13436;
			G1312<=G1309;
			G1315<=G1312;
			G1316<=G20562;
			G1319<=G24337;
			G1326<=G23199;
			G1332<=G26000;
			G1339<=G25151;
			G1345<=G21944;
			G1346<=G26708;
			G1352<=G27698;
			G1358<=G27218;
			G1365<=G28257;
			G1372<=G28682;
			G1378<=G29146;
			G1384<=G23202;
			G1385<=G23200;
			G1386<=G23201;
			G1387<=G23205;
			G1388<=G23203;
			G1389<=G23204;
			G1390<=G23208;
			G1391<=G23206;
			G1392<=G23207;
			G1393<=G23211;
			G1394<=G23209;
			G1395<=G23210;
			G1396<=G23214;
			G1397<=G23212;
			G1398<=G23213;
			G1399<=G23217;
			G1400<=G23215;
			G1401<=G23216;
			G1402<=G23220;
			G1403<=G23218;
			G1404<=G23219;
			G1405<=G23223;
			G1406<=G23221;
			G1407<=G23222;
			G1408<=G23226;
			G1409<=G23224;
			G1410<=G23225;
			G1411<=G23229;
			G1412<=G23227;
			G1413<=G23228;
			G1414<=G23232;
			G1415<=G23230;
			G1416<=G23231;
			G1417<=G23235;
			G1418<=G23233;
			G1419<=G23234;
			G1420<=G26711;
			G1421<=G26709;
			G1422<=G26710;
			G1423<=G24340;
			G1424<=G24338;
			G1425<=G24339;
			G1426<=G29802;
			G1430<=G29641;
			G1435<=G29427;
			G1439<=G29147;
			G1444<=G28683;
			G1448<=G28258;
			G1453<=G27699;
			G1457<=G27219;
			G1462<=G26712;
			G1466<=G26001;
			G1471<=G20579;
			G1476<=G20578;
			G1481<=G20577;
			G1486<=G20576;
			G1491<=G20575;
			G1496<=G20574;
			G1501<=G20573;
			G1506<=G20572;
			G1511<=G24343;
			G1512<=G24341;
			G1513<=G24342;
			G1514<=G24346;
			G1515<=G24344;
			G1516<=G24345;
			G1517<=G1520;
			G1520<=G13437;
			G1523<=G24349;
			G1524<=G24347;
			G1525<=G24348;
			G1526<=G24352;
			G1527<=G24350;
			G1528<=G24351;
			G1529<=G24355;
			G1530<=G24353;
			G1531<=G24354;
			G1532<=G24358;
			G1533<=G24356;
			G1534<=G24357;
			G1535<=G24361;
			G1536<=G24359;
			G1537<=G24360;
			G1538<=G24364;
			G1539<=G24362;
			G1540<=G24363;
			G1541<=G24367;
			G1542<=G24365;
			G1543<=G24366;
			G1544<=G24370;
			G1545<=G24368;
			G1546<=G24369;
			G1547<=G1517;
			G1550<=G26715;
			G1551<=G26713;
			G1552<=G26714;
			G1553<=G26718;
			G1554<=G26716;
			G1555<=G26717;
			G1556<=G26721;
			G1557<=G26719;
			G1558<=G26720;
			G1559<=G26724;
			G1560<=G26722;
			G1561<=G26723;
			G1562<=G20563;
			G1563<=G1564;
			G1564<=G1562;
			G1567<=G30536;
			G1570<=G30537;
			G1573<=G30538;
			G1576<=G30872;
			G1579<=G30873;
			G1582<=G30874;
			G1585<=G30539;
			G1588<=G30540;
			G1591<=G30541;
			G1594<=G30542;
			G1597<=G30543;
			G1600<=G30544;
			G1603<=G30875;
			G1606<=G30876;
			G1609<=G30877;
			G1612<=G30878;
			G1615<=G30879;
			G1618<=G30880;
			G1621<=G30881;
			G1624<=G30882;
			G1627<=G30883;
			G1630<=G30545;
			G1633<=G30546;
			G1636<=G30547;
			G1639<=G30548;
			G1642<=G30549;
			G1645<=G30550;
			G1648<=G30884;
			G1651<=G30885;
			G1654<=G30886;
			G1657<=G13438;
			G1660<=G1835;
			G1661<=G11545;
			G1662<=G1661;
			G1663<=G11546;
			G1664<=G1663;
			G1665<=G11547;
			G1666<=G1665;
			G1667<=G11548;
			G1668<=G1667;
			G1669<=G11549;
			G1670<=G1669;
			G1671<=G13439;
			G1672<=G1671;
			G1675<=G29433;
			G1676<=G29432;
			G1677<=G29431;
			G1678<=G29430;
			G1679<=G27220;
			G1680<=G19036;
			G1681<=G25152;
			G1682<=G19037;
			G1683<=G19038;
			G1684<=G19039;
			G1685<=G19040;
			G1686<=G29428;
			G1689<=G29429;
			G1690<=G11550;
			G1693<=G29803;
			G1694<=G29804;
			G1695<=G29805;
			G1696<=G30887;
			G1697<=G30888;
			G1698<=G30889;
			G1699<=G30716;
			G1700<=G30717;
			G1701<=G30718;
			G1702<=G29644;
			G1703<=G29642;
			G1704<=G29643;
			G1705<=G1778;
			G1706<=G13440;
			G1712<=G1706;
			G1718<=G1712;
			G1723<=G11551;
			G1724<=G28260;
			G1727<=G28261;
			G1730<=G1723;
			G1731<=G11552;
			G1732<=G1731;
			G1733<=G11553;
			G1734<=G1733;
			G1735<=G28259;
			G1738<=G11554;
			G1739<=G28263;
			G1742<=G28264;
			G1745<=G1738;
			G1746<=G11555;
			G1747<=G1746;
			G1748<=G11556;
			G1749<=G1748;
			G1750<=G28262;
			G1753<=G11557;
			G1754<=G28266;
			G1757<=G28267;
			G1760<=G1753;
			G1761<=G11558;
			G1762<=G1761;
			G1763<=G11559;
			G1764<=G1763;
			G1765<=G28265;
			G1768<=G11560;
			G1769<=G28269;
			G1772<=G28270;
			G1775<=G1768;
			G1776<=G11561;
			G1777<=G1776;
			G1778<=G11562;
			G1779<=G28268;
			G1782<=G1786;
			G1783<=G27223;
			G1784<=G27221;
			G1785<=G27222;
			G1786<=G1657;
			G1789<=G29434;
			G1792<=G29435;
			G1795<=G29436;
			G1798<=G29645;
			G1801<=G29646;
			G1804<=G29647;
			G1807<=G29439;
			G1808<=G29437;
			G1809<=G29438;
			G1810<=G27700;
			G1813<=G27701;
			G1816<=G27702;
			G1819<=G27703;
			G1822<=G27704;
			G1825<=G27705;
			G1828<=G28686;
			G1829<=G28684;
			G1830<=G28685;
			G1831<=G11563;
			G1832<=G1831;
			G1833<=G11564;
			G1834<=G1833;
			G1835<=G11565;
			G1836<=G25161;
			G1839<=G25153;
			G1842<=G25154;
			G1845<=G24373;
			G1846<=G25155;
			G1849<=G25156;
			G1852<=G25157;
			G1855<=G13441;
			G1858<=G25158;
			G1859<=G25159;
			G1860<=G25160;
			G1861<=G24371;
			G1862<=G1855;
			G1865<=G24372;
			G1866<=G1862;
			G1867<=G24374;
			G1868<=G24375;
			G1869<=G24376;
			G1870<=G1948;
			G1871<=G27224;
			G1874<=G27225;
			G1877<=G27226;
			G1880<=G1929;
			G1886<=G8302;
			G1887<=G24377;
			G1888<=G19041;
			G1889<=G19042;
			G1890<=G20565;
			G1893<=G16471;
			G1894<=G19043;
			G1895<=G19044;
			G1896<=G29444;
			G1897<=G29443;
			G1898<=G29442;
			G1899<=G29441;
			G1900<=G29440;
			G1903<=G1893;
			G1904<=G1903;
			G1905<=G1900;
			G1908<=G16472;
			G1909<=G13442;
			G1910<=G13443;
			G1911<=G13444;
			G1912<=G13445;
			G1913<=G13446;
			G1914<=G13447;
			G1915<=G1908;
			G1916<=G13448;
			G1917<=G13449;
			G1918<=G26002;
			G1921<=G13450;
			G1922<=G1915;
			G1923<=G19045;
			G1924<=G1923;
			G1925<=G13451;
			G1928<=G29445;
			G1929<=G19046;
			G1930<=G1931;
			G1931<=G1925;
			G1934<=G23236;
			G1937<=G20564;
			G1938<=G19047;
			G1939<=G1938;
			G1944<=G11566;
			G1945<=G1954;
			G1946<=G11567;
			G1947<=G1946;
			G1948<=G11568;
			G1949<=G1944;
			G1950<=G11569;
			G1951<=G1950;
			G1952<=G11570;
			G1953<=G1952;
			G1954<=G11571;
			G1955<=G28273;
			G1956<=G28271;
			G1957<=G28272;
			G1958<=G28276;
			G1959<=G28274;
			G1960<=G28275;
			G1961<=G28279;
			G1962<=G28277;
			G1963<=G28278;
			G1964<=G28282;
			G1965<=G28280;
			G1966<=G28281;
			G1967<=G26003;
			G1970<=G26004;
			G1973<=G26005;
			G1976<=G26006;
			G1979<=G26007;
			G1982<=G26008;
			G1985<=G29148;
			G1988<=G29149;
			G1991<=G29150;
			G1994<=G29151;
			G1997<=G29152;
			G2000<=G29153;
			G2003<=G13452;
			G2006<=G2003;
			G2009<=G2006;
			G2010<=G20566;
			G2013<=G24378;
			G2020<=G23237;
			G2026<=G26009;
			G2033<=G25162;
			G2039<=G21945;
			G2040<=G26725;
			G2046<=G27706;
			G2052<=G27227;
			G2059<=G28283;
			G2066<=G28687;
			G2072<=G29154;
			G2078<=G23240;
			G2079<=G23238;
			G2080<=G23239;
			G2081<=G23243;
			G2082<=G23241;
			G2083<=G23242;
			G2084<=G23246;
			G2085<=G23244;
			G2086<=G23245;
			G2087<=G23249;
			G2088<=G23247;
			G2089<=G23248;
			G2090<=G23252;
			G2091<=G23250;
			G2092<=G23251;
			G2093<=G23255;
			G2094<=G23253;
			G2095<=G23254;
			G2096<=G23258;
			G2097<=G23256;
			G2098<=G23257;
			G2099<=G23261;
			G2100<=G23259;
			G2101<=G23260;
			G2102<=G23264;
			G2103<=G23262;
			G2104<=G23263;
			G2105<=G23267;
			G2106<=G23265;
			G2107<=G23266;
			G2108<=G23270;
			G2109<=G23268;
			G2110<=G23269;
			G2111<=G23273;
			G2112<=G23271;
			G2113<=G23272;
			G2114<=G26728;
			G2115<=G26726;
			G2116<=G26727;
			G2117<=G24381;
			G2118<=G24379;
			G2119<=G24380;
			G2120<=G29806;
			G2124<=G29648;
			G2129<=G29446;
			G2133<=G29155;
			G2138<=G28688;
			G2142<=G28284;
			G2147<=G27707;
			G2151<=G27228;
			G2156<=G26729;
			G2160<=G26010;
			G2165<=G20580;
			G2170<=G20581;
			G2175<=G20582;
			G2180<=G20583;
			G2185<=G20584;
			G2190<=G20586;
			G2195<=G20585;
			G2200<=G20587;
			G2205<=G24384;
			G2206<=G24382;
			G2207<=G24383;
			G2208<=G24387;
			G2209<=G24385;
			G2210<=G24386;
			G2211<=G2214;
			G2214<=G13453;
			G2217<=G24390;
			G2218<=G24388;
			G2219<=G24389;
			G2220<=G24393;
			G2221<=G24391;
			G2222<=G24392;
			G2223<=G24396;
			G2224<=G24394;
			G2225<=G24395;
			G2226<=G24399;
			G2227<=G24397;
			G2228<=G24398;
			G2229<=G24402;
			G2230<=G24400;
			G2231<=G24401;
			G2232<=G24405;
			G2233<=G24403;
			G2234<=G24404;
			G2235<=G24408;
			G2236<=G24406;
			G2237<=G24407;
			G2238<=G24411;
			G2239<=G24409;
			G2240<=G24410;
			G2241<=G2211;
			G2244<=G26732;
			G2245<=G26730;
			G2246<=G26731;
			G2247<=G26735;
			G2248<=G26733;
			G2249<=G26734;
			G2250<=G26738;
			G2251<=G26736;
			G2252<=G26737;
			G2253<=G26741;
			G2254<=G26739;
			G2255<=G26740;
			G2256<=G20567;
			G2257<=G2258;
			G2258<=G2256;
			G2261<=G30551;
			G2264<=G30552;
			G2267<=G30553;
			G2270<=G30890;
			G2273<=G30891;
			G2276<=G30892;
			G2279<=G30554;
			G2282<=G30555;
			G2285<=G30556;
			G2288<=G30557;
			G2291<=G30558;
			G2294<=G30559;
			G2297<=G30893;
			G2300<=G30894;
			G2303<=G30895;
			G2306<=G30896;
			G2309<=G30897;
			G2312<=G30898;
			G2315<=G30899;
			G2318<=G30900;
			G2321<=G30901;
			G2324<=G30560;
			G2327<=G30561;
			G2330<=G30562;
			G2333<=G30563;
			G2336<=G30564;
			G2339<=G30565;
			G2342<=G30902;
			G2345<=G30903;
			G2348<=G30904;
			G2351<=G13454;
			G2354<=G2529;
			G2355<=G11572;
			G2356<=G2355;
			G2357<=G11573;
			G2358<=G2357;
			G2359<=G11574;
			G2360<=G2359;
			G2361<=G11575;
			G2362<=G2361;
			G2363<=G11576;
			G2364<=G2363;
			G2365<=G13455;
			G2366<=G2365;
			G2369<=G30319;
			G2370<=G30318;
			G2371<=G30317;
			G2372<=G30316;
			G2373<=G27229;
			G2374<=G19048;
			G2375<=G25163;
			G2376<=G19049;
			G2377<=G19050;
			G2378<=G19051;
			G2379<=G19052;
			G2380<=G30314;
			G2383<=G30315;
			G2384<=G11577;
			G2387<=G29807;
			G2388<=G29808;
			G2389<=G29809;
			G2390<=G30905;
			G2391<=G30906;
			G2392<=G30907;
			G2393<=G30719;
			G2394<=G30720;
			G2395<=G30721;
			G2396<=G29651;
			G2397<=G29649;
			G2398<=G29650;
			G2399<=G2472;
			G2400<=G13456;
			G2406<=G2400;
			G2412<=G2406;
			G2417<=G11578;
			G2418<=G28286;
			G2421<=G28287;
			G2424<=G2417;
			G2425<=G11579;
			G2426<=G2425;
			G2427<=G11580;
			G2428<=G2427;
			G2429<=G28285;
			G2432<=G11581;
			G2433<=G28289;
			G2436<=G28290;
			G2439<=G2432;
			G2440<=G11582;
			G2441<=G2440;
			G2442<=G11583;
			G2443<=G2442;
			G2444<=G28288;
			G2447<=G11584;
			G2448<=G28292;
			G2451<=G28293;
			G2454<=G2447;
			G2455<=G11585;
			G2456<=G2455;
			G2457<=G11586;
			G2458<=G2457;
			G2459<=G28291;
			G2462<=G11587;
			G2463<=G28295;
			G2466<=G28296;
			G2469<=G2462;
			G2470<=G11588;
			G2471<=G2470;
			G2472<=G11589;
			G2473<=G28294;
			G2476<=G2480;
			G2477<=G27232;
			G2478<=G27230;
			G2479<=G27231;
			G2480<=G2351;
			G2483<=G29447;
			G2486<=G29448;
			G2489<=G29449;
			G2492<=G29652;
			G2495<=G29653;
			G2498<=G29654;
			G2501<=G29452;
			G2502<=G29450;
			G2503<=G29451;
			G2504<=G27708;
			G2507<=G27709;
			G2510<=G27710;
			G2513<=G27711;
			G2516<=G27712;
			G2519<=G27713;
			G2522<=G28691;
			G2523<=G28689;
			G2524<=G28690;
			G2525<=G11590;
			G2526<=G2525;
			G2527<=G11591;
			G2528<=G2527;
			G2529<=G11592;
			G2530<=G25172;
			G2533<=G25164;
			G2536<=G25165;
			G2539<=G24414;
			G2540<=G25166;
			G2543<=G25167;
			G2546<=G25168;
			G2549<=G13457;
			G2552<=G25169;
			G2553<=G25170;
			G2554<=G25171;
			G2555<=G24412;
			G2556<=G2549;
			G2559<=G24413;
			G2560<=G2556;
			G2561<=G24415;
			G2562<=G24416;
			G2563<=G24417;
			G2564<=G2642;
			G2565<=G27233;
			G2568<=G27234;
			G2571<=G27235;
			G2574<=G2623;
			G2580<=G8311;
			G2581<=G24418;
			G2582<=G19053;
			G2583<=G19054;
			G2584<=G20569;
			G2587<=G16473;
			G2588<=G19055;
			G2589<=G19056;
			G2590<=G30324;
			G2591<=G30323;
			G2592<=G30322;
			G2593<=G30321;
			G2594<=G30320;
			G2597<=G2587;
			G2598<=G2597;
			G2599<=G2594;
			G2602<=G16474;
			G2603<=G13458;
			G2604<=G13459;
			G2605<=G13460;
			G2606<=G13461;
			G2607<=G13462;
			G2608<=G13463;
			G2609<=G2602;
			G2610<=G13464;
			G2611<=G13465;
			G2612<=G26011;
			G2615<=G13466;
			G2616<=G2609;
			G2617<=G19057;
			G2618<=G2617;
			G2619<=G13467;
			G2622<=G30325;
			G2623<=G19058;
			G2624<=G2625;
			G2625<=G2619;
			G2628<=G23274;
			G2631<=G20568;
			G2632<=G19059;
			G2633<=G2632;
			G2638<=G11593;
			G2639<=G2648;
			G2640<=G11594;
			G2641<=G2640;
			G2642<=G11595;
			G2643<=G2638;
			G2644<=G11596;
			G2645<=G2644;
			G2646<=G11597;
			G2647<=G2646;
			G2648<=G11598;
			G2649<=G28299;
			G2650<=G28297;
			G2651<=G28298;
			G2652<=G28302;
			G2653<=G28300;
			G2654<=G28301;
			G2655<=G28305;
			G2656<=G28303;
			G2657<=G28304;
			G2658<=G28308;
			G2659<=G28306;
			G2660<=G28307;
			G2661<=G26012;
			G2664<=G26013;
			G2667<=G26014;
			G2670<=G26015;
			G2673<=G26016;
			G2676<=G26017;
			G2679<=G29156;
			G2682<=G29157;
			G2685<=G29158;
			G2688<=G29159;
			G2691<=G29160;
			G2694<=G29161;
			G2697<=G13468;
			G2700<=G2697;
			G2703<=G2700;
			G2704<=G20570;
			G2707<=G24419;
			G2714<=G23275;
			G2720<=G26018;
			G2727<=G25173;
			G2733<=G21946;
			G2734<=G26742;
			G2740<=G27714;
			G2746<=G27236;
			G2753<=G28309;
			G2760<=G28692;
			G2766<=G29162;
			G2772<=G23278;
			G2773<=G23276;
			G2774<=G23277;
			G2775<=G23281;
			G2776<=G23279;
			G2777<=G23280;
			G2778<=G23284;
			G2779<=G23282;
			G2780<=G23283;
			G2781<=G23287;
			G2782<=G23285;
			G2783<=G23286;
			G2784<=G23290;
			G2785<=G23288;
			G2786<=G23289;
			G2787<=G23293;
			G2788<=G23291;
			G2789<=G23292;
			G2790<=G23296;
			G2791<=G23294;
			G2792<=G23295;
			G2793<=G23299;
			G2794<=G23297;
			G2795<=G23298;
			G2796<=G23302;
			G2797<=G23300;
			G2798<=G23301;
			G2799<=G23305;
			G2800<=G23303;
			G2801<=G23304;
			G2802<=G23308;
			G2803<=G23306;
			G2804<=G23307;
			G2805<=G23311;
			G2806<=G23309;
			G2807<=G23310;
			G2808<=G26745;
			G2809<=G26743;
			G2810<=G26744;
			G2811<=G24422;
			G2812<=G24420;
			G2813<=G24421;
			G2814<=G16475;
			G2817<=G20571;
			G2818<=G21947;
			G2821<=G21948;
			G2824<=G21949;
			G2827<=G21950;
			G2830<=G23312;
			G2833<=G21952;
			G2836<=G21953;
			G2839<=G21954;
			G2842<=G21955;
			G2845<=G21956;
			G2848<=G21957;
			G2851<=G21958;
			G2854<=G21959;
			G2857<=G2858;
			G2858<=G23316;
			G2861<=G21960;
			G2864<=G21961;
			G2867<=G21962;
			G2870<=G21963;
			G2873<=G2830;
			G2874<=G16493;
			G2877<=G23313;
			G2878<=G23314;
			G2879<=G16494;
			G2883<=G23315;
			G2888<=G24423;
			G2892<=G26019;
			G2896<=G25175;
			G2900<=G27237;
			G2903<=G26747;
			G2908<=G27715;
			G2912<=G24424;
			G2917<=G25174;
			G2920<=G26746;
			G2924<=G26020;
			G2929<=G2930;
			G2930<=G19062;
			G2933<=G20588;
			G2934<=G16476;
			G2935<=G16477;
			G2938<=G16478;
			G2941<=G16479;
			G2944<=G16480;
			G2947<=G16481;
			G2950<=G21951;
			G2953<=G16482;
			G2956<=G16483;
			G2959<=G16484;
			G2962<=G16485;
			G2963<=G16486;
			G2966<=G16487;
			G2969<=G16488;
			G2972<=G16489;
			G2975<=G16490;
			G2978<=G16491;
			G2981<=G16492;
			G2984<=G19061;
			G2985<=G19060;
			G2986<=G3040;
			G2987<=G16495;
			G2990<=G20593;
			G2991<=G21964;
			G2992<=G21966;
			G2993<=G26748;
			G2997<=G30989;
			G2998<=G27238;
			G3002<=G26021;
			G3006<=G25177;
			G3010<=G27239;
			G3013<=G26750;
			G3018<=G24425;
			G3024<=G27716;
			G3028<=G25176;
			G3032<=G26749;
			G3036<=G26022;
			G3040<=G16497;
			G3043<=G29453;
			G3044<=G29454;
			G3045<=G29455;
			G3046<=G29456;
			G3047<=G29457;
			G3048<=G29458;
			G3049<=G29459;
			G3050<=G29460;
			G3051<=G29655;
			G3052<=G29972;
			G3053<=G29973;
			G3054<=G23317;
			G3055<=G29974;
			G3056<=G29975;
			G3057<=G29976;
			G3058<=G29977;
			G3059<=G29978;
			G3060<=G29979;
			G3061<=G30119;
			G3062<=G30908;
			G3063<=G30909;
			G3064<=G30910;
			G3065<=G30911;
			G3066<=G30912;
			G3067<=G30913;
			G3068<=G30914;
			G3069<=G30915;
			G3070<=G30940;
			G3071<=G30980;
			G3072<=G30981;
			G3073<=G30982;
			G3074<=G30983;
			G3075<=G30984;
			G3076<=G30985;
			G3077<=G30986;
			G3078<=G30987;
			G3079<=G23318;
			G3080<=G21965;
			G3083<=G20603;
			G3084<=G20632;
			G3085<=G20609;
			G3086<=G20610;
			G3087<=G20611;
			G3088<=G20629;
			G3091<=G20612;
			G3092<=G20613;
			G3093<=G20614;
			G3094<=G20615;
			G3095<=G20616;
			G3096<=G20617;
			G3097<=G26751;
			G3098<=G26752;
			G3099<=G26753;
			G3100<=G29163;
			G3101<=G29164;
			G3102<=G29165;
			G3103<=G30120;
			G3104<=G30121;
			G3105<=G30122;
			G3106<=G30941;
			G3107<=G30942;
			G3108<=G30943;
			G3109<=G3117;
			G3110<=G28311;
			G3111<=G28310;
			G3112<=G28312;
			G3113<=G28693;
			G3114<=G28694;
			G3117<=G3129;
			G3120<=G28695;
			G3123<=G28313;
			G3124<=G28314;
			G3125<=G28696;
			G3126<=G28315;
			G3127<=G28697;
			G3128<=G29166;
			G3129<=G13475;
			G3132<=G28698;
			G3133<=G29656;
			G3134<=G28700;
			G3135<=G28699;
			G3136<=G28701;
			G3139<=G29461;
			G3142<=G28703;
			G3147<=G28702;
			G3151<=G29462;
			G3155<=G20618;
			G3158<=G20619;
			G3161<=G20620;
			G3164<=G20621;
			G3167<=G20622;
			G3170<=G20623;
			G3173<=G20624;
			G3176<=G20625;
			G3179<=G20626;
			G3182<=G20627;
			G3185<=G20628;
			G3188<=G29463;
			G3191<=G27717;
			G3194<=G28316;
			G3197<=G28317;
			G3198<=G28318;
			G3201<=G28704;
			G3204<=G28705;
			G3207<=G28706;
			G3210<=G20630;
			G3211<=G20631;
		end if;
	end process;
	G562<= not I13089;
	G1248<= not I13092;
	G1942<= not I13095;
	G2636<= not I13098;
	G3235<= not I13101;
	G3236<= not I13104;
	G3237<= not I13107;
	G3238<= not I13110;
	G3239<= not I13113;
	G3240<= not I13116;
	G3241<= not I13119;
	G3242<= not I13122;
	G3243<= not I13125;
	G3244<= not I13128;
	G3245<= not I13131;
	G3246<= not I13134;
	G3247<= not I13137;
	G3248<= not I13140;
	G3249<= not I13143;
	G3250<= not I13146;
	G3251<= not I13149;
	G3252<= not I13152;
	G3253<= not I13155;
	G3254<= not I13158;
	G3304<= not I13161;
	G3305<= not G305;
	G3306<= not I13165;
	G3337<= not G309;
	G3338<= not I13169;
	G3365<= not G499;
	G3366<= not I13173;
	G3398<= not I13176;
	G3410<= not I13179;
	G3460<= not I13182;
	G3461<= not G992;
	G3462<= not I13186;
	G3493<= not G996;
	G3494<= not I13190;
	G3521<= not G1186;
	G3522<= not I13194;
	G3554<= not I13197;
	G3566<= not I13200;
	G3616<= not I13203;
	G3617<= not G1686;
	G3618<= not I13207;
	G3649<= not G1690;
	G3650<= not I13211;
	G3677<= not G1880;
	G3678<= not I13215;
	G3710<= not I13218;
	G3722<= not I13221;
	G3772<= not I13224;
	G3773<= not G2380;
	G3774<= not I13228;
	G3805<= not G2384;
	G3806<= not I13232;
	G3833<= not G2574;
	G3834<= not I13236;
	G3866<= not I13239;
	G3878<= not I13242;
	G3897<= not G2950;
	G3900<= not I13246;
	G3919<= not G3080;
	G3922<= not G150;
	G3925<= not G155;
	G3928<= not G157;
	G3931<= not G171;
	G3934<= not G176;
	G3937<= not G178;
	G3940<= not G408;
	G3941<= not G455;
	G3942<= not G699;
	G3945<= not G726;
	G3948<= not G835;
	G3951<= not G840;
	G3954<= not G842;
	G3957<= not G856;
	G3960<= not G861;
	G3963<= not G863;
	G3966<= not G1526;
	G3969<= not G1531;
	G3972<= not G1533;
	G3975<= not G1552;
	G3978<= not G1554;
	G3981<= not G2217;
	G3984<= not G2222;
	G3987<= not G2224;
	G3990<= not G2245;
	G3993<= not I13275;
	G3994<= not G2848;
	G3995<= not G3064;
	G3996<= not G3073;
	G3997<= not G45;
	G3998<= not G23;
	G3999<= not G3204;
	G4000<= not G153;
	G4003<= not G158;
	G4006<= not G160;
	G4009<= not G174;
	G4012<= not G179;
	G4015<= not G411;
	G4016<= not G417;
	G4017<= not G427;
	G4020<= not G700;
	G4023<= not G702;
	G4026<= not G727;
	G4029<= not G838;
	G4032<= not G843;
	G4035<= not G845;
	G4038<= not G859;
	G4041<= not G864;
	G4044<= not G866;
	G4047<= not G1095;
	G4048<= not G1142;
	G4049<= not G1385;
	G4052<= not G1412;
	G4055<= not G1529;
	G4058<= not G1534;
	G4061<= not G1536;
	G4064<= not G1550;
	G4067<= not G1555;
	G4070<= not G1557;
	G4073<= not G2220;
	G4076<= not G2225;
	G4079<= not G2227;
	G4082<= not G2246;
	G4085<= not G2248;
	G4088<= not I13316;
	G4089<= not G2836;
	G4090<= not I13320;
	G4091<= not G2864;
	G4092<= not G3074;
	G4093<= not G33;
	G4094<= not G3207;
	G4095<= not G130;
	G4098<= not G156;
	G4101<= not G161;
	G4104<= not G163;
	G4107<= not G177;
	G4110<= not G414;
	G4111<= not G420;
	G4112<= not G428;
	G4115<= not G698;
	G4118<= not G703;
	G4121<= not G705;
	G4124<= not G725;
	G4127<= not G841;
	G4130<= not G846;
	G4133<= not G848;
	G4136<= not G862;
	G4139<= not G867;
	G4142<= not G1098;
	G4143<= not G1104;
	G4144<= not G1114;
	G4147<= not G1386;
	G4150<= not G1388;
	G4153<= not G1413;
	G4156<= not G1532;
	G4159<= not G1537;
	G4162<= not G1539;
	G4165<= not G1553;
	G4168<= not G1558;
	G4171<= not G1560;
	G4174<= not G1789;
	G4175<= not G1836;
	G4176<= not G2079;
	G4179<= not G2106;
	G4182<= not G2223;
	G4185<= not G2228;
	G4188<= not G2230;
	G4191<= not G2244;
	G4194<= not G2249;
	G4197<= not G2251;
	G4200<= not I13366;
	G4201<= not G2851;
	G4202<= not G42;
	G4203<= not G20;
	G4204<= not G3188;
	G4205<= not G131;
	G4208<= not G133;
	G4211<= not G159;
	G4214<= not G164;
	G4217<= not G354;
	G4220<= not G423;
	G4221<= not G426;
	G4224<= not G429;
	G4225<= not G701;
	G4228<= not G706;
	G4231<= not G708;
	G4234<= not G818;
	G4237<= not G844;
	G4240<= not G849;
	G4243<= not G851;
	G4246<= not G865;
	G4249<= not G1101;
	G4250<= not G1107;
	G4251<= not G1115;
	G4254<= not G1384;
	G4257<= not G1389;
	G4260<= not G1391;
	G4263<= not G1411;
	G4266<= not G1535;
	G4269<= not G1540;
	G4272<= not G1542;
	G4275<= not G1556;
	G4278<= not G1561;
	G4281<= not G1792;
	G4282<= not G1798;
	G4283<= not G1808;
	G4286<= not G2080;
	G4289<= not G2082;
	G4292<= not G2107;
	G4295<= not G2226;
	G4298<= not G2231;
	G4301<= not G2233;
	G4304<= not G2247;
	G4307<= not G2252;
	G4310<= not G2254;
	G4313<= not G2483;
	G4314<= not G2530;
	G4315<= not G2773;
	G4318<= not G2800;
	G4321<= not I13417;
	G4322<= not G2839;
	G4323<= not I13421;
	G4324<= not G2867;
	G4325<= not G36;
	G4326<= not G181;
	G4329<= not G129;
	G4332<= not G134;
	G4335<= not G162;
	G4338<= not I13430;
	G4339<= not I13433;
	G4340<= not G343;
	G4343<= not G369;
	G4346<= not G432;
	G4347<= not G438;
	G4348<= not G704;
	G4351<= not G709;
	G4354<= not G711;
	G4357<= not G729;
	G4360<= not G819;
	G4363<= not G821;
	G4366<= not G847;
	G4369<= not G852;
	G4372<= not G1041;
	G4375<= not G1110;
	G4376<= not G1113;
	G4379<= not G1116;
	G4380<= not G1387;
	G4383<= not G1392;
	G4386<= not G1394;
	G4389<= not G1512;
	G4392<= not G1538;
	G4395<= not G1543;
	G4398<= not G1545;
	G4401<= not G1559;
	G4404<= not G1795;
	G4405<= not G1801;
	G4406<= not G1809;
	G4409<= not G2078;
	G4412<= not G2083;
	G4415<= not G2085;
	G4418<= not G2105;
	G4421<= not G2229;
	G4424<= not G2234;
	G4427<= not G2236;
	G4430<= not G2250;
	G4433<= not G2255;
	G4436<= not G2486;
	G4437<= not G2492;
	G4438<= not G2502;
	G4441<= not G2774;
	G4444<= not G2776;
	G4447<= not G2801;
	G4450<= not I13478;
	G4451<= not G2854;
	G4452<= not G17;
	G4453<= not G132;
	G4456<= not G309;
	G4465<= not G346;
	G4468<= not G358;
	G4471<= not G384;
	G4474<= not G435;
	G4475<= not G441;
	G4476<= not G576;
	G4479<= not G587;
	G4480<= not G707;
	G4483<= not G712;
	G4486<= not G714;
	G4489<= not G730;
	G4492<= not G732;
	G4495<= not G869;
	G4498<= not G817;
	G4501<= not G822;
	G4504<= not G850;
	G4507<= not I13501;
	G4508<= not I13504;
	G4509<= not G1030;
	G4512<= not G1056;
	G4515<= not G1119;
	G4516<= not G1125;
	G4517<= not G1390;
	G4520<= not G1395;
	G4523<= not G1397;
	G4526<= not G1415;
	G4529<= not G1513;
	G4532<= not G1515;
	G4535<= not G1541;
	G4538<= not G1546;
	G4541<= not G1735;
	G4544<= not G1804;
	G4545<= not G1807;
	G4548<= not G1810;
	G4549<= not G2081;
	G4552<= not G2086;
	G4555<= not G2088;
	G4558<= not G2206;
	G4561<= not G2232;
	G4564<= not G2237;
	G4567<= not G2239;
	G4570<= not G2253;
	G4573<= not G2489;
	G4574<= not G2495;
	G4575<= not G2503;
	G4578<= not G2772;
	G4581<= not G2777;
	G4584<= not G2779;
	G4587<= not G2799;
	G4590<= not I13538;
	G4591<= not G2870;
	G4592<= not G361;
	G4595<= not G373;
	G4598<= not G398;
	G4601<= not G444;
	G4602<= not G525;
	G4603<= not G577;
	G4606<= not G579;
	G4609<= not G590;
	G4610<= not G596;
	G4611<= not G710;
	G4614<= not G715;
	G4617<= not G717;
	G4620<= not G728;
	G4623<= not G733;
	G4626<= not G735;
	G4629<= not G820;
	G4632<= not G996;
	G4641<= not G1033;
	G4644<= not G1045;
	G4647<= not G1071;
	G4650<= not G1122;
	G4651<= not G1128;
	G4652<= not G1262;
	G4655<= not G1273;
	G4656<= not G1393;
	G4659<= not G1398;
	G4662<= not G1400;
	G4665<= not G1416;
	G4668<= not G1418;
	G4671<= not G1563;
	G4674<= not G1511;
	G4677<= not G1516;
	G4680<= not G1544;
	G4683<= not I13575;
	G4684<= not I13578;
	G4685<= not G1724;
	G4688<= not G1750;
	G4691<= not G1813;
	G4692<= not G1819;
	G4693<= not G2084;
	G4696<= not G2089;
	G4699<= not G2091;
	G4702<= not G2109;
	G4705<= not G2207;
	G4708<= not G2209;
	G4711<= not G2235;
	G4714<= not G2240;
	G4717<= not G2429;
	G4720<= not G2498;
	G4721<= not G2501;
	G4724<= not G2504;
	G4725<= not G2775;
	G4728<= not G2780;
	G4731<= not G2782;
	G4734<= not G11;
	G4735<= not I13601;
	G4736<= not I13604;
	G4737<= not G376;
	G4740<= not G388;
	G4743<= not G575;
	G4746<= not G580;
	G4749<= not G582;
	G4752<= not G593;
	G4753<= not G599;
	G4754<= not G713;
	G4757<= not G718;
	G4760<= not G720;
	G4763<= not G731;
	G4766<= not G736;
	G4769<= not G1048;
	G4772<= not G1060;
	G4775<= not G1085;
	G4778<= not G1131;
	G4779<= not G1211;
	G4780<= not G1263;
	G4783<= not G1265;
	G4786<= not G1276;
	G4787<= not G1282;
	G4788<= not G1396;
	G4791<= not G1401;
	G4794<= not G1403;
	G4797<= not G1414;
	G4800<= not G1419;
	G4803<= not G1421;
	G4806<= not G1514;
	G4809<= not G1690;
	G4818<= not G1727;
	G4821<= not G1739;
	G4824<= not G1765;
	G4827<= not G1816;
	G4828<= not G1822;
	G4829<= not G1956;
	G4832<= not G1967;
	G4833<= not G2087;
	G4836<= not G2092;
	G4839<= not G2094;
	G4842<= not G2110;
	G4845<= not G2112;
	G4848<= not G2257;
	G4851<= not G2205;
	G4854<= not G2210;
	G4857<= not G2238;
	G4860<= not I13652;
	G4861<= not I13655;
	G4862<= not G2418;
	G4865<= not G2444;
	G4868<= not G2507;
	G4869<= not G2513;
	G4870<= not G2778;
	G4873<= not G2783;
	G4876<= not G2785;
	G4879<= not G2803;
	G4882<= not G391;
	G4885<= not G448;
	G4888<= not G578;
	G4891<= not G583;
	G4894<= not G585;
	G4897<= not G602;
	G4898<= not G605;
	G4899<= not G716;
	G4902<= not G721;
	G4905<= not G723;
	G4908<= not G734;
	G4911<= not I13677;
	G4912<= not I13680;
	G4913<= not G1063;
	G4916<= not G1075;
	G4919<= not G1261;
	G4922<= not G1266;
	G4925<= not G1268;
	G4928<= not G1279;
	G4929<= not G1285;
	G4930<= not G1399;
	G4933<= not G1404;
	G4936<= not G1406;
	G4939<= not G1417;
	G4942<= not G1422;
	G4945<= not G1742;
	G4948<= not G1754;
	G4951<= not G1779;
	G4954<= not G1825;
	G4955<= not G1905;
	G4956<= not G1957;
	G4959<= not G1959;
	G4962<= not G1970;
	G4963<= not G1976;
	G4964<= not G2090;
	G4967<= not G2095;
	G4970<= not G2097;
	G4973<= not G2108;
	G4976<= not G2113;
	G4979<= not G2115;
	G4982<= not G2208;
	G4985<= not G2384;
	G4994<= not G2421;
	G4997<= not G2433;
	G5000<= not G2459;
	G5003<= not G2510;
	G5004<= not G2516;
	G5005<= not G2650;
	G5008<= not G2661;
	G5009<= not G2781;
	G5012<= not G2786;
	G5015<= not G2788;
	G5018<= not G2804;
	G5021<= not G2806;
	G5024<= not G449;
	G5027<= not G581;
	G5030<= not G586;
	G5033<= not G608;
	G5034<= not G614;
	G5035<= not G719;
	G5038<= not G724;
	G5041<= not G1078;
	G5044<= not G1135;
	G5047<= not G1264;
	G5050<= not G1269;
	G5053<= not G1271;
	G5056<= not G1288;
	G5057<= not G1291;
	G5058<= not G1402;
	G5061<= not G1407;
	G5064<= not G1409;
	G5067<= not G1420;
	G5070<= not I13742;
	G5071<= not I13745;
	G5072<= not G1757;
	G5075<= not G1769;
	G5078<= not G1955;
	G5081<= not G1960;
	G5084<= not G1962;
	G5087<= not G1973;
	G5088<= not G1979;
	G5089<= not G2093;
	G5092<= not G2098;
	G5095<= not G2100;
	G5098<= not G2111;
	G5101<= not G2116;
	G5104<= not G2436;
	G5107<= not G2448;
	G5110<= not G2473;
	G5113<= not G2519;
	G5114<= not G2599;
	G5115<= not G2651;
	G5118<= not G2653;
	G5121<= not G2664;
	G5122<= not G2670;
	G5123<= not G2784;
	G5126<= not G2789;
	G5129<= not G2791;
	G5132<= not G2802;
	G5135<= not G2807;
	G5138<= not G2809;
	G5141<= not I13775;
	G5142<= not G447;
	G5145<= not G584;
	G5148<= not G611;
	G5149<= not G617;
	G5150<= not G722;
	G5153<= not G1136;
	G5156<= not G1267;
	G5159<= not G1272;
	G5162<= not G1294;
	G5163<= not G1300;
	G5164<= not G1405;
	G5167<= not G1410;
	G5170<= not G1772;
	G5173<= not G1829;
	G5176<= not G1958;
	G5179<= not G1963;
	G5182<= not G1965;
	G5185<= not G1982;
	G5186<= not G1985;
	G5187<= not G2096;
	G5190<= not G2101;
	G5193<= not G2103;
	G5196<= not G2114;
	G5199<= not I13801;
	G5200<= not I13804;
	G5201<= not G2451;
	G5204<= not G2463;
	G5207<= not G2649;
	G5210<= not G2654;
	G5213<= not G2656;
	G5216<= not G2667;
	G5217<= not G2673;
	G5218<= not G2787;
	G5221<= not G2792;
	G5224<= not G2794;
	G5227<= not G2805;
	G5230<= not G2810;
	G5233<= not G620;
	G5234<= not I13820;
	G5235<= not G1134;
	G5238<= not G1270;
	G5241<= not G1297;
	G5242<= not G1303;
	G5243<= not G1408;
	G5246<= not G1830;
	G5249<= not G1961;
	G5252<= not G1966;
	G5255<= not G1988;
	G5256<= not G1994;
	G5257<= not G2099;
	G5260<= not G2104;
	G5263<= not G2466;
	G5266<= not G2523;
	G5269<= not G2652;
	G5272<= not G2657;
	G5275<= not G2659;
	G5278<= not G2676;
	G5279<= not G2679;
	G5280<= not G2790;
	G5283<= not G2795;
	G5286<= not G2797;
	G5289<= not G2808;
	G5292<= not G2857;
	G5293<= not G738;
	G5296<= not G1306;
	G5297<= not I13849;
	G5298<= not G1828;
	G5301<= not G1964;
	G5304<= not G1991;
	G5305<= not G1997;
	G5306<= not G2102;
	G5309<= not G2524;
	G5312<= not G2655;
	G5315<= not G2660;
	G5318<= not G2682;
	G5319<= not G2688;
	G5320<= not G2793;
	G5323<= not G2798;
	G5326<= not G2873;
	G5327<= not G739;
	G5330<= not G1424;
	G5333<= not G2000;
	G5334<= not I13868;
	G5335<= not G2522;
	G5338<= not G2658;
	G5341<= not G2685;
	G5342<= not G2691;
	G5343<= not G2796;
	G5346<= not G3106;
	G5349<= not G2877;
	G5352<= not G737;
	G5355<= not G1425;
	G5358<= not G2118;
	G5361<= not G2694;
	G5362<= not G2817;
	G5363<= not G3107;
	G5366<= not G2878;
	G5369<= not G1423;
	G5372<= not G2119;
	G5375<= not G2812;
	G5378<= not G2933;
	G5379<= not G3108;
	G5382<= not G2117;
	G5385<= not G2813;
	G5388<= not I13892;
	G5389<= not G3040;
	G5390<= not I13896;
	G5391<= not G2811;
	G5394<= not G3054;
	G5395<= not I13901;
	G5396<= not I13904;
	G5397<= not I13907;
	G5398<= not I13910;
	G5399<= not I13913;
	G5400<= not I13916;
	G5401<= not I13919;
	G5402<= not I13922;
	G5403<= not I13925;
	G5404<= not I13928;
	G5405<= not I13931;
	G5406<= not I13934;
	G5407<= not I13937;
	G5408<= not I13940;
	G5409<= not I13943;
	G5410<= not G3079;
	G5411<= not I13947;
	G5412<= not I13950;
	G5413<= not I13953;
	G5414<= not I13956;
	G5415<= not I13959;
	G5416<= not I13962;
	G5417<= not I13965;
	G5418<= not I13968;
	G5419<= not I13971;
	G5420<= not I13974;
	G5421<= not I13977;
	G5422<= not I13980;
	G5423<= not G2879;
	G5424<= not I13984;
	G5425<= not I13987;
	G5426<= not I13990;
	G5427<= not I13993;
	G5428<= not G3210;
	G5431<= not G3211;
	G5434<= not G3084;
	G5437<= not I13999;
	G5438<= not I14002;
	G5469<= not G3085;
	G5472<= not I14006;
	G5473<= not I14009;
	G5504<= not G3086;
	G5507<= not G3155;
	G5508<= not I14014;
	G5511<= not I14017;
	G5512<= not I14020;
	G5543<= not G3087;
	G5546<= not G3164;
	G5547<= not G101;
	G5548<= not G105;
	G5549<= not I14027;
	G5550<= not I14030;
	G5551<= not G514;
	G5552<= not I14034;
	G5555<= not I14037;
	G5556<= not I14040;
	G5587<= not G3091;
	G5590<= not G3158;
	G5591<= not G3173;
	G5592<= not G515;
	G5593<= not G789;
	G5594<= not G793;
	G5595<= not I14049;
	G5596<= not I14052;
	G5597<= not G1200;
	G5598<= not I14056;
	G5601<= not G3092;
	G5604<= not G3167;
	G5605<= not G3182;
	G5606<= not G79;
	G5609<= not G1201;
	G5610<= not G1476;
	G5611<= not G1481;
	G5612<= not I14066;
	G5613<= not I14069;
	G5614<= not G1894;
	G5615<= not I14073;
	G5618<= not G3093;
	G5621<= not G3161;
	G5622<= not G3176;
	G5623<= not G70;
	G5626<= not G121;
	G5627<= not G125;
	G5628<= not G300;
	G5629<= not I14083;
	G5631<= not G767;
	G5634<= not G1895;
	G5635<= not G2170;
	G5636<= not G2175;
	G5637<= not I14091;
	G5638<= not I14094;
	G5639<= not G2588;
	G5640<= not G3170;
	G5641<= not G3185;
	G5642<= not G61;
	G5645<= not G101;
	G5646<= not G213;
	G5647<= not G301;
	G5648<= not I14104;
	G5651<= not G758;
	G5654<= not G809;
	G5655<= not G813;
	G5656<= not G987;
	G5657<= not I14113;
	G5659<= not G1453;
	G5662<= not G2589;
	G5663<= not G3179;
	G5664<= not G65;
	G5665<= not G105;
	G5666<= not G216;
	G5667<= not G222;
	G5668<= not G299;
	G5675<= not G302;
	G5679<= not G506;
	G5680<= not G749;
	G5683<= not G789;
	G5684<= not G900;
	G5685<= not G988;
	G5686<= not I14134;
	G5689<= not G1444;
	G5692<= not G1501;
	G5693<= not G1506;
	G5694<= not G1681;
	G5695<= not I14143;
	G5697<= not G2147;
	G5700<= not G3088;
	G5701<= not I14149;
	G5702<= not G56;
	G5703<= not G109;
	G5704<= not G219;
	G5705<= not G225;
	G5706<= not G231;
	G5707<= not G109;
	G5708<= not G303;
	G5712<= not G305;
	G5713<= not I14163;
	G5714<= not G507;
	G5715<= not G541;
	G5716<= not G753;
	G5717<= not G793;
	G5718<= not G903;
	G5719<= not G909;
	G5720<= not G986;
	G5727<= not G989;
	G5731<= not G1192;
	G5732<= not G1435;
	G5735<= not G1476;
	G5736<= not G1594;
	G5737<= not G1682;
	G5738<= not I14182;
	G5741<= not G2138;
	G5744<= not G2195;
	G5745<= not G2200;
	G5746<= not G2375;
	G5747<= not I14191;
	G5749<= not I14195;
	G5750<= not G92;
	G5751<= not G52;
	G5752<= not G113;
	G5753<= not G228;
	G5754<= not G234;
	G5755<= not G240;
	G5756<= not G304;
	G5759<= not G508;
	G5760<= not G744;
	G5761<= not G797;
	G5762<= not G906;
	G5763<= not G912;
	G5764<= not G918;
	G5765<= not G797;
	G5766<= not G990;
	G5770<= not G992;
	G5771<= not I14219;
	G5772<= not G1193;
	G5773<= not G1227;
	G5774<= not G1439;
	G5775<= not G1481;
	G5776<= not G1597;
	G5777<= not G1603;
	G5778<= not G1680;
	G5785<= not G1683;
	G5789<= not G1886;
	G5790<= not G2129;
	G5793<= not G2170;
	G5794<= not G2288;
	G5795<= not G2376;
	G5796<= not I14238;
	G5799<= not I14243;
	G5800<= not I14246;
	G5801<= not I14249;
	G5802<= not G83;
	G5803<= not G117;
	G5804<= not G237;
	G5805<= not G243;
	G5806<= not G249;
	G5808<= not G509;
	G5809<= not G780;
	G5810<= not G740;
	G5811<= not G801;
	G5812<= not G915;
	G5813<= not G921;
	G5814<= not G927;
	G5815<= not G991;
	G5818<= not G1194;
	G5819<= not G1430;
	G5820<= not G1486;
	G5821<= not G1600;
	G5822<= not G1606;
	G5823<= not G1612;
	G5824<= not G1486;
	G5825<= not G1684;
	G5829<= not G1686;
	G5830<= not I14280;
	G5831<= not G1887;
	G5832<= not G1921;
	G5833<= not G2133;
	G5834<= not G2175;
	G5835<= not G2291;
	G5836<= not G2297;
	G5837<= not G2374;
	G5844<= not G2377;
	G5848<= not G2580;
	G5849<= not I14295;
	G5850<= not I14298;
	G5851<= not G74;
	G5852<= not G121;
	G5853<= not G246;
	G5854<= not G252;
	G5855<= not G258;
	G5856<= not I14306;
	G5857<= not G538;
	G5858<= not G771;
	G5859<= not G805;
	G5860<= not G924;
	G5861<= not G930;
	G5862<= not G936;
	G5864<= not G1195;
	G5865<= not G1466;
	G5866<= not G1426;
	G5867<= not G1491;
	G5868<= not G1609;
	G5869<= not G1615;
	G5870<= not G1621;
	G5871<= not G1685;
	G5874<= not G1888;
	G5875<= not G2124;
	G5876<= not G2180;
	G5877<= not G2294;
	G5878<= not G2300;
	G5879<= not G2306;
	G5880<= not G2180;
	G5881<= not G2378;
	G5885<= not G2380;
	G5886<= not I14338;
	G5887<= not G2581;
	G5888<= not G2615;
	G5889<= not I14343;
	G5890<= not G88;
	G5893<= not G125;
	G5894<= not G186;
	G5895<= not G255;
	G5896<= not G261;
	G5897<= not G267;
	G5898<= not G762;
	G5899<= not G809;
	G5900<= not G933;
	G5901<= not G939;
	G5902<= not G945;
	G5903<= not I14357;
	G5904<= not G1224;
	G5905<= not G1457;
	G5906<= not G1496;
	G5907<= not G1618;
	G5908<= not G1624;
	G5909<= not G1630;
	G5911<= not G1889;
	G5912<= not G2160;
	G5913<= not G2120;
	G5914<= not G2185;
	G5915<= not G2303;
	G5916<= not G2309;
	G5917<= not G2315;
	G5918<= not G2379;
	G5921<= not G2582;
	G5922<= not I14378;
	G5923<= not I14381;
	G5924<= not I14384;
	G5925<= not G189;
	G5926<= not G195;
	G5927<= not G264;
	G5928<= not G270;
	G5929<= not G776;
	G5932<= not G813;
	G5933<= not G873;
	G5934<= not G942;
	G5935<= not G948;
	G5936<= not G954;
	G5937<= not G1448;
	G5938<= not G1501;
	G5939<= not G1627;
	G5940<= not G1633;
	G5941<= not G1639;
	G5942<= not I14402;
	G5943<= not G1918;
	G5944<= not G2151;
	G5945<= not G2190;
	G5946<= not G2312;
	G5947<= not G2318;
	G5948<= not G2324;
	G5950<= not G2583;
	G5951<= not I14413;
	G5952<= not I14416;
	G5953<= not G97;
	G5954<= not G192;
	G5955<= not G198;
	G5956<= not G204;
	G5957<= not G273;
	G5958<= not I14424;
	G5959<= not G876;
	G5960<= not G882;
	G5961<= not G951;
	G5962<= not G957;
	G5963<= not G1462;
	G5966<= not G1506;
	G5967<= not G1567;
	G5968<= not G1636;
	G5969<= not G1642;
	G5970<= not G1648;
	G5971<= not G2142;
	G5972<= not G2195;
	G5973<= not G2321;
	G5974<= not G2327;
	G5975<= not G2333;
	G5976<= not I14442;
	G5977<= not G2612;
	G5978<= not I14446;
	G5979<= not I14449;
	G5980<= not G201;
	G5981<= not G207;
	G5982<= not G785;
	G5983<= not G879;
	G5984<= not G885;
	G5985<= not G891;
	G5986<= not G960;
	G5987<= not I14459;
	G5988<= not G1570;
	G5989<= not G1576;
	G5990<= not G1645;
	G5991<= not G1651;
	G5992<= not G2156;
	G5995<= not G2200;
	G5996<= not G2261;
	G5997<= not G2330;
	G5998<= not G2336;
	G5999<= not G2342;
	G6000<= not I14472;
	G6014<= not I14475;
	G6015<= not I14478;
	G6016<= not G210;
	G6017<= not G888;
	G6018<= not G894;
	G6019<= not G1471;
	G6020<= not G1573;
	G6021<= not G1579;
	G6022<= not G1585;
	G6023<= not G1654;
	G6024<= not I14489;
	G6025<= not G2264;
	G6026<= not G2270;
	G6027<= not G2339;
	G6028<= not G2345;
	G6029<= not I14496;
	G6030<= not I14499;
	G6031<= not I14502;
	G6032<= not G897;
	G6033<= not G1582;
	G6034<= not G1588;
	G6035<= not G2165;
	G6036<= not G2267;
	G6037<= not G2273;
	G6038<= not G2279;
	G6039<= not G2348;
	G6040<= not I14513;
	G6041<= not I14516;
	G6042<= not I14519;
	G6043<= not G1591;
	G6044<= not G2276;
	G6045<= not G2282;
	G6046<= not I14525;
	G6047<= not G2285;
	G6048<= not I14529;
	G6051<= not I14532;
	G6052<= not I14535;
	G6053<= not I14538;
	G6054<= not I14541;
	G6055<= not I14544;
	G6056<= not I14547;
	G6057<= not I14550;
	G6058<= not I14553;
	G6059<= not I14556;
	G6060<= not I14559;
	G6061<= not I14562;
	G6062<= not I14565;
	G6063<= not I14568;
	G6064<= not I14571;
	G6065<= not I14574;
	G6066<= not I14577;
	G6067<= not I14580;
	G6068<= not G499;
	G6079<= not I14584;
	G6080<= not I14587;
	G6081<= not I14590;
	G6082<= not I14593;
	G6083<= not I14596;
	G6084<= not I14599;
	G6085<= not I14602;
	G6086<= not I14605;
	G6087<= not G1186;
	G6098<= not I14609;
	G6099<= not I14612;
	G6100<= not I14615;
	G6101<= not I14618;
	G6102<= not I14621;
	G6103<= not I14624;
	G6104<= not G1880;
	G6115<= not I14628;
	G6116<= not I14631;
	G6117<= not I14634;
	G6118<= not I14637;
	G6119<= not G2574;
	G6130<= not I14641;
	G6131<= not I14644;
	G6134<= not I14647;
	G6135<= not I14650;
	G6136<= not G672;
	G6139<= not I14654;
	G6140<= not G524;
	G6141<= not G554;
	G6142<= not G679;
	G6145<= not I14660;
	G6146<= not G1358;
	G6149<= not G3097;
	G6153<= not I14665;
	G6156<= not I14668;
	G6157<= not G686;
	G6161<= not G1210;
	G6162<= not G1240;
	G6163<= not G1365;
	G6166<= not I14675;
	G6167<= not G2052;
	G6170<= not G3098;
	G6173<= not G557;
	G6177<= not G633;
	G6180<= not G692;
	G6183<= not G291;
	G6184<= not G1372;
	G6188<= not G1904;
	G6189<= not G1934;
	G6190<= not G2059;
	G6193<= not I14688;
	G6194<= not G2746;
	G6197<= not G3099;
	G6200<= not G542;
	G6201<= not G646;
	G6204<= not G289;
	G6205<= not G1243;
	G6209<= not G1319;
	G6212<= not G1378;
	G6215<= not G978;
	G6216<= not G2066;
	G6220<= not G2598;
	G6221<= not G2628;
	G6222<= not G2753;
	G6225<= not I14704;
	G6226<= not G2818;
	G6227<= not G3100;
	G6230<= not I14709;
	G6231<= not I14712;
	G6232<= not I14715;
	G6281<= not G510;
	G6284<= not G640;
	G6288<= not G287;
	G6289<= not G1228;
	G6290<= not G1332;
	G6293<= not G976;
	G6294<= not G1937;
	G6298<= not G2013;
	G6301<= not G2072;
	G6304<= not G1672;
	G6305<= not G2760;
	G6309<= not G14;
	G6310<= not G3101;
	G6313<= not I14731;
	G6314<= not I14734;
	G6363<= not G653;
	G6367<= not G285;
	G6368<= not I14739;
	G6369<= not I14742;
	G6418<= not G1196;
	G6421<= not G1326;
	G6425<= not G974;
	G6426<= not G1922;
	G6427<= not G2026;
	G6430<= not G1670;
	G6431<= not G2631;
	G6435<= not G2707;
	G6438<= not G2766;
	G6441<= not G2366;
	G6442<= not I14755;
	G6443<= not G2821;
	G6444<= not G3102;
	G6447<= not I14760;
	G6448<= not I14763;
	G6485<= not I14766;
	G6486<= not I14769;
	G6512<= not G544;
	G6513<= not G660;
	G6517<= not G283;
	G6518<= not I14775;
	G6519<= not I14778;
	G6568<= not G1339;
	G6572<= not G972;
	G6573<= not I14783;
	G6574<= not I14786;
	G6623<= not G1890;
	G6626<= not G2020;
	G6630<= not G1668;
	G6631<= not G2616;
	G6632<= not G2720;
	G6635<= not G2364;
	G6636<= not G1491;
	G6637<= not G5;
	G6638<= not G3103;
	G6641<= not G113;
	G6642<= not I14799;
	G6643<= not I14802;
	G6672<= not G464;
	G6675<= not G458;
	G6676<= not G559;
	G6677<= not I14808;
	G6678<= not I14811;
	G6707<= not G666;
	G6711<= not G281;
	G6712<= not I14816;
	G6713<= not I14819;
	G6750<= not I14822;
	G6751<= not I14825;
	G6776<= not G1230;
	G6777<= not G1346;
	G6781<= not G970;
	G6782<= not I14831;
	G6783<= not I14834;
	G6832<= not G2033;
	G6836<= not G1666;
	G6837<= not I14839;
	G6838<= not I14842;
	G6887<= not G2584;
	G6890<= not G2714;
	G6894<= not G2362;
	G6895<= not I14848;
	G6896<= not G2824;
	G6897<= not G1486;
	G6898<= not G2993;
	G6901<= not G3006;
	G6905<= not G3104;
	G6908<= not G484;
	G6911<= not I14857;
	G6912<= not I14860;
	G6942<= not G279;
	G6943<= not G801;
	G6944<= not I14865;
	G6945<= not I14868;
	G6974<= not G1151;
	G6977<= not G1145;
	G6978<= not G1245;
	G6979<= not I14874;
	G6980<= not I14877;
	G7009<= not G1352;
	G7013<= not G968;
	G7014<= not I14882;
	G7015<= not I14885;
	G7052<= not I14888;
	G7053<= not I14891;
	G7078<= not G1924;
	G7079<= not G2040;
	G7083<= not G1664;
	G7084<= not I14897;
	G7085<= not I14900;
	G7134<= not G2727;
	G7138<= not G2360;
	G7139<= not G1481;
	G7140<= not G2170;
	G7141<= not G2195;
	G7142<= not G8;
	G7143<= not G2998;
	G7146<= not G3013;
	G7149<= not G3105;
	G7152<= not G3136;
	G7153<= not G480;
	G7156<= not G461;
	G7157<= not G453;
	G7158<= not G1171;
	G7161<= not I14917;
	G7162<= not I14920;
	G7192<= not G966;
	G7193<= not G1491;
	G7194<= not I14925;
	G7195<= not I14928;
	G7224<= not G1845;
	G7227<= not G1839;
	G7228<= not G1939;
	G7229<= not I14934;
	G7230<= not I14937;
	G7259<= not G2046;
	G7263<= not G1662;
	G7264<= not I14942;
	G7265<= not I14945;
	G7302<= not I14948;
	G7303<= not I14951;
	G7328<= not G2618;
	G7329<= not G2734;
	G7333<= not G2358;
	G7334<= not I14957;
	G7335<= not G2827;
	G7336<= not G1476;
	G7337<= not G2190;
	G7338<= not G3002;
	G7342<= not G3024;
	G7345<= not G3139;
	G7346<= not G97;
	G7347<= not G490;
	G7348<= not G451;
	G7349<= not G1167;
	G7352<= not G1148;
	G7353<= not G1140;
	G7354<= not G1865;
	G7357<= not I14973;
	G7358<= not I14976;
	G7388<= not G1660;
	G7389<= not G2185;
	G7390<= not I14981;
	G7391<= not I14984;
	G7420<= not G2539;
	G7423<= not G2533;
	G7424<= not G2633;
	G7425<= not I14990;
	G7426<= not I14993;
	G7455<= not G2740;
	G7459<= not G2356;
	G7460<= not G1471;
	G7461<= not G2175;
	G7462<= not G2912;
	G7465<= not G2;
	G7466<= not G3010;
	G7471<= not G3036;
	G7475<= not G493;
	G7476<= not G785;
	G7477<= not G1177;
	G7478<= not G1138;
	G7479<= not G1861;
	G7482<= not G1842;
	G7483<= not G1834;
	G7484<= not G2559;
	G7487<= not I15012;
	G7488<= not I15015;
	G7518<= not G2354;
	G7519<= not I15019;
	G7520<= not G2830;
	G7521<= not G2200;
	G7522<= not G2917;
	G7527<= not G3018;
	G7529<= not G465;
	G7530<= not G496;
	G7531<= not G1180;
	G7532<= not G1471;
	G7533<= not G1871;
	G7534<= not G1832;
	G7535<= not G2555;
	G7538<= not G2536;
	G7539<= not G2528;
	G7540<= not G1506;
	G7541<= not G2180;
	G7542<= not G2883;
	G7545<= not G2920;
	G7548<= not G2990;
	G7549<= not G3028;
	G7553<= not G3114;
	G7554<= not G117;
	G7555<= not G1152;
	G7556<= not G1183;
	G7557<= not G1874;
	G7558<= not G2165;
	G7559<= not G2565;
	G7560<= not G2526;
	G7561<= not G1501;
	G7562<= not G2888;
	G7566<= not G2896;
	G7570<= not G3032;
	G7573<= not G3120;
	G7574<= not G3128;
	G7576<= not G468;
	G7577<= not G805;
	G7578<= not G1846;
	G7579<= not G1877;
	G7580<= not G2568;
	G7581<= not G1496;
	G7582<= not G2185;
	G7583<= not G2892;
	G7587<= not G2903;
	G7590<= not G1155;
	G7591<= not G1496;
	G7592<= not G2540;
	G7593<= not G2571;
	G7594<= not G2165;
	G7595<= not G2900;
	G7600<= not G2908;
	G7603<= not G3133;
	G7604<= not G471;
	G7605<= not G1849;
	G7606<= not G2190;
	G7607<= not G2924;
	G7610<= not G312;
	G7613<= not G1158;
	G7614<= not G2543;
	G7615<= not G3123;
	G7616<= not G313;
	G7619<= not G999;
	G7622<= not G1852;
	G7623<= not G314;
	G7626<= not G315;
	G7629<= not G403;
	G7632<= not G1000;
	G7635<= not G1693;
	G7638<= not G2546;
	G7639<= not G3094;
	G7642<= not G3125;
	G7643<= not G316;
	G7646<= not G318;
	G7649<= not G404;
	G7652<= not G1001;
	G7655<= not G1002;
	G7658<= not G1090;
	G7661<= not G1694;
	G7664<= not G2387;
	G7667<= not G3095;
	G7670<= not G317;
	G7673<= not G319;
	G7676<= not G402;
	G7679<= not G1003;
	G7682<= not G1005;
	G7685<= not G1091;
	G7688<= not G1695;
	G7691<= not G1696;
	G7694<= not G1784;
	G7697<= not G2388;
	G7700<= not G3096;
	G7703<= not G320;
	G7706<= not G1004;
	G7709<= not G1006;
	G7712<= not G1089;
	G7715<= not G1697;
	G7718<= not G1699;
	G7721<= not G1785;
	G7724<= not G2389;
	G7727<= not G2390;
	G7730<= not G2478;
	G7733<= not G1007;
	G7736<= not G1698;
	G7739<= not G1700;
	G7742<= not G1783;
	G7745<= not G2391;
	G7748<= not G2393;
	G7751<= not G2479;
	G7754<= not G322;
	G7757<= not G1701;
	G7760<= not G2392;
	G7763<= not G2394;
	G7766<= not G2477;
	G7769<= not G323;
	G7772<= not G659;
	G7776<= not G1009;
	G7779<= not G2395;
	G7782<= not G321;
	G7785<= not G1010;
	G7788<= not G1345;
	G7792<= not G1703;
	G7796<= not G1008;
	G7799<= not G1704;
	G7802<= not G2039;
	G7806<= not G2397;
	G7809<= not G1702;
	G7812<= not G2398;
	G7815<= not G2733;
	G7819<= not G479;
	G7822<= not G510;
	G7823<= not G2396;
	G7826<= not G2987;
	G7827<= not G478;
	G7830<= not G1166;
	G7833<= not G1196;
	G7834<= not G2953;
	G7837<= not G3044;
	G7838<= not G477;
	G7841<= not G630;
	G7842<= not G1165;
	G7845<= not G1860;
	G7848<= not G1890;
	G7849<= not G2956;
	G7852<= not G2981;
	G7856<= not G3045;
	G7857<= not G3055;
	G7858<= not G1164;
	G7861<= not G1316;
	G7862<= not G1859;
	G7865<= not G2554;
	G7868<= not G2584;
	G7869<= not G2959;
	G7872<= not G2874;
	G7877<= not G3046;
	G7878<= not G3056;
	G7879<= not G3065;
	G7880<= not G3201;
	G7888<= not G1858;
	G7891<= not G2010;
	G7892<= not G2553;
	G7897<= not G3047;
	G7898<= not G3057;
	G7899<= not G3066;
	G7900<= not G3075;
	G7901<= not I15222;
	G7906<= not G488;
	G7909<= not I15226;
	G7910<= not G474;
	G7911<= not I15230;
	G7912<= not G2552;
	G7915<= not G2704;
	G7916<= not G2935;
	G7919<= not G2963;
	G7924<= not G3048;
	G7925<= not G3058;
	G7926<= not G3067;
	G7927<= not G3076;
	G7928<= not G3204;
	G7936<= not I15256;
	G7949<= not G165;
	G7950<= not G142;
	G7953<= not G487;
	G7956<= not I15262;
	G7957<= not G481;
	G7958<= not G1175;
	G7961<= not I15267;
	G7962<= not G1161;
	G7963<= not I15271;
	G7964<= not G2938;
	G7967<= not G2966;
	G7971<= not G3049;
	G7972<= not G3059;
	G7973<= not G3068;
	G7974<= not G3077;
	G7975<= not G39;
	G7976<= not I15288;
	G7989<= not G3191;
	G7990<= not G143;
	G7993<= not G145;
	G7996<= not G486;
	G7999<= not G485;
	G8000<= not G853;
	G8001<= not G830;
	G8004<= not G1174;
	G8007<= not I15299;
	G8008<= not G1168;
	G8009<= not G1869;
	G8012<= not I15304;
	G8013<= not G1855;
	G8014<= not I15308;
	G8015<= not G2941;
	G8018<= not G2969;
	G8021<= not I15313;
	G8022<= not G2930;
	G8023<= not I15317;
	G8024<= not G2842;
	G8025<= not G3050;
	G8026<= not G3060;
	G8027<= not G3069;
	G8028<= not G3078;
	G8029<= not G3083;
	G8030<= not I15326;
	G8031<= not I15329;
	G8044<= not G3194;
	G8045<= not G3207;
	G8053<= not G141;
	G8056<= not G146;
	G8059<= not G148;
	G8062<= not G169;
	G8065<= not G831;
	G8068<= not G833;
	G8071<= not G1173;
	G8074<= not G1172;
	G8075<= not G1547;
	G8076<= not G1524;
	G8079<= not G1868;
	G8082<= not I15345;
	G8083<= not G1862;
	G8084<= not G2563;
	G8087<= not I15350;
	G8088<= not G2549;
	G8089<= not I15354;
	G8090<= not G2944;
	G8093<= not G2972;
	G8096<= not I15359;
	G8097<= not G2858;
	G8098<= not G3051;
	G8099<= not G3061;
	G8100<= not G3070;
	G8101<= not G2997;
	G8102<= not G27;
	G8103<= not G185;
	G8106<= not I15369;
	G8107<= not I15372;
	G8120<= not G3197;
	G8123<= not G144;
	G8126<= not G149;
	G8129<= not G151;
	G8132<= not G170;
	G8135<= not G172;
	G8138<= not G829;
	G8141<= not G834;
	G8144<= not G836;
	G8147<= not G857;
	G8150<= not G1525;
	G8153<= not G1527;
	G8156<= not G1867;
	G8159<= not G1866;
	G8160<= not G2241;
	G8161<= not G2218;
	G8164<= not G2562;
	G8167<= not I15392;
	G8168<= not G2556;
	G8169<= not G2947;
	G8172<= not G2975;
	G8175<= not I15398;
	G8176<= not G2845;
	G8177<= not G3043;
	G8178<= not G3052;
	G8179<= not G3062;
	G8180<= not G3071;
	G8181<= not G48;
	G8182<= not G3198;
	G8183<= not G3188;
	G8191<= not G147;
	G8194<= not G152;
	G8197<= not G154;
	G8200<= not G168;
	G8203<= not G173;
	G8206<= not G175;
	G8209<= not G832;
	G8212<= not G837;
	G8215<= not G839;
	G8218<= not G858;
	G8221<= not G860;
	G8224<= not G1523;
	G8227<= not G1528;
	G8230<= not G1530;
	G8233<= not G1551;
	G8236<= not G2219;
	G8239<= not G2221;
	G8242<= not G2561;
	G8245<= not G2560;
	G8246<= not G2978;
	G8249<= not I15429;
	G8250<= not G2833;
	G8251<= not I15433;
	G8252<= not G2861;
	G8253<= not G3053;
	G8254<= not G3063;
	G8255<= not G3072;
	G8256<= not G30;
	G8257<= not G3201;
	G8258<= not I15442;
	G8259<= not I15445;
	G8260<= not I15448;
	G8261<= not I15451;
	G8262<= not I15454;
	G8263<= not I15457;
	G8264<= not I15460;
	G8265<= not I15463;
	G8266<= not I15466;
	G8267<= not I15469;
	G8268<= not I15472;
	G8269<= not I15475;
	G8270<= not I15478;
	G8271<= not I15481;
	G8272<= not I15484;
	G8273<= not I15487;
	G8274<= not I15490;
	G8275<= not I15493;
	G8276<= not G3253;
	G8277<= not G3305;
	G8278<= not G3337;
	G8284<= not I15499;
	G8285<= not G3365;
	G8286<= not G3461;
	G8287<= not G3493;
	G8293<= not I15505;
	G8294<= not G3521;
	G8295<= not G3617;
	G8296<= not G3649;
	G8302<= not I15511;
	G8303<= not G3677;
	G8304<= not G3773;
	G8305<= not G3805;
	G8311<= not I15517;
	G8312<= not G3833;
	G8313<= not G3897;
	G8317<= not G3919;
	G8321<= not I15523;
	G8324<= not I15526;
	G8330<= not I15532;
	G8333<= not I15535;
	G8336<= not I15538;
	G8341<= not I15543;
	G8344<= not I15546;
	G8347<= not I15549;
	G8351<= not I15553;
	G8354<= not I15556;
	G8357<= not I15559;
	G8360<= not I15562;
	G8363<= not I15565;
	G8366<= not I15568;
	G8369<= not I15571;
	G8372<= not I15574;
	G8375<= not I15577;
	G8378<= not I15580;
	G8382<= not I15584;
	G8388<= not I15590;
	G8391<= not I15593;
	G8397<= not I15599;
	G8400<= not I15602;
	G8403<= not I15605;
	G8408<= not I15610;
	G8411<= not I15613;
	G8414<= not I15616;
	G8418<= not I15620;
	G8421<= not I15623;
	G8424<= not I15626;
	G8427<= not I15629;
	G8434<= not I15636;
	G8440<= not I15642;
	G8443<= not I15645;
	G8449<= not I15651;
	G8452<= not I15654;
	G8455<= not I15657;
	G8460<= not I15662;
	G8469<= not I15671;
	G8475<= not I15677;
	G8478<= not I15680;
	G8494<= not I15696;
	G8514<= not G6139;
	G8530<= not G6156;
	G8568<= not G6230;
	G8569<= not I15771;
	G8575<= not I15779;
	G8578<= not I15784;
	G8579<= not I15787;
	G8580<= not G6281;
	G8587<= not G6418;
	G8594<= not G6623;
	G8602<= not I15794;
	G8605<= not G6887;
	G8614<= not I15800;
	G8617<= not I15803;
	G8620<= not I15806;
	G8622<= not I15810;
	G8627<= not I15815;
	G8630<= not I15818;
	G8632<= not I15822;
	G8637<= not I15827;
	G8640<= not I15830;
	G8643<= not I15833;
	G8646<= not I15836;
	G8649<= not I15839;
	G8651<= not I15843;
	G8655<= not I15847;
	G8658<= not I15850;
	G8659<= not I15853;
	G8662<= not I15856;
	G8665<= not I15859;
	G8667<= not I15863;
	G8670<= not I15866;
	G8673<= not I15869;
	G8677<= not I15873;
	G8678<= not I15876;
	G8681<= not I15879;
	G8684<= not I15882;
	G8689<= not I15887;
	G8690<= not I15890;
	G8693<= not I15893;
	G8696<= not I15896;
	G8699<= not I15899;
	G8700<= not I15902;
	G8707<= not I15909;
	G8708<= not I15912;
	G8711<= not I15915;
	G8714<= not I15918;
	G8718<= not I15922;
	G8719<= not I15925;
	G8726<= not I15932;
	G8745<= not I15935;
	G8748<= not I15938;
	G8752<= not I15942;
	G8756<= not I15946;
	G8757<= not I15949;
	G8763<= not I15955;
	G8766<= not I15958;
	G8769<= not I15961;
	G8770<= not I15964;
	G8771<= not I15967;
	G8775<= not I15971;
	G8779<= not I15975;
	G8780<= not I15978;
	G8785<= not I15983;
	G8788<= not I15986;
	G8791<= not I15989;
	G8792<= not I15992;
	G8793<= not I15995;
	G8794<= not I15998;
	G8798<= not I16002;
	G8802<= not I16006;
	G8805<= not I16009;
	G8808<= not I16012;
	G8809<= not I16015;
	G8810<= not I16018;
	G8811<= not I16021;
	G8812<= not I16024;
	G8813<= not I16027;
	G8817<= not I16031;
	G8820<= not I16034;
	G8821<= not I16037;
	G8822<= not G4602;
	G8823<= not I16041;
	G8824<= not I16044;
	G8825<= not I16047;
	G8826<= not I16050;
	G8827<= not I16053;
	G8828<= not I16056;
	G8829<= not I16059;
	G8832<= not I16062;
	G8835<= not I16065;
	G8836<= not I16068;
	G8839<= not I16071;
	G8840<= not I16074;
	G8843<= not I16079;
	G8844<= not I16082;
	G8845<= not I16085;
	G8846<= not G4779;
	G8847<= not I16089;
	G8850<= not I16092;
	G8851<= not I16095;
	G8852<= not I16098;
	G8853<= not I16101;
	G8856<= not I16104;
	G8859<= not I16107;
	G8860<= not I16110;
	G8862<= not I16114;
	G8863<= not I16117;
	G8866<= not I16120;
	G8867<= not I16123;
	G8870<= not I16128;
	G8871<= not I16131;
	G8872<= not I16134;
	G8873<= not G4955;
	G8874<= not I16138;
	G8877<= not I16141;
	G8878<= not I16144;
	G8879<= not I16147;
	G8882<= not I16150;
	G8885<= not I16153;
	G8888<= not I16156;
	G8891<= not I16159;
	G8893<= not I16163;
	G8894<= not I16166;
	G8897<= not I16169;
	G8898<= not I16172;
	G8900<= not I16176;
	G8901<= not I16179;
	G8904<= not I16182;
	G8905<= not I16185;
	G8908<= not I16190;
	G8909<= not I16193;
	G8910<= not I16196;
	G8911<= not G5114;
	G8912<= not I16200;
	G8915<= not I16203;
	G8918<= not I16206;
	G8921<= not I16209;
	G8924<= not I16212;
	G8925<= not I16215;
	G8928<= not I16218;
	G8931<= not I16221;
	G8933<= not I16225;
	G8934<= not I16228;
	G8937<= not I16231;
	G8938<= not I16234;
	G8940<= not I16238;
	G8941<= not I16241;
	G8944<= not I16244;
	G8945<= not I16247;
	G8948<= not I16252;
	G8949<= not I16255;
	G8952<= not I16258;
	G8955<= not I16261;
	G8958<= not I16264;
	G8961<= not I16267;
	G8964<= not I16270;
	G8965<= not I16273;
	G8968<= not I16276;
	G8971<= not I16279;
	G8973<= not I16283;
	G8974<= not I16286;
	G8977<= not I16289;
	G8978<= not I16292;
	G8980<= not I16296;
	G8983<= not G6486;
	G8984<= not I16300;
	G8987<= not I16303;
	G8990<= not I16306;
	G8993<= not I16309;
	G8996<= not I16312;
	G8997<= not I16315;
	G9000<= not I16318;
	G9003<= not I16321;
	G9005<= not I16325;
	G9006<= not I16328;
	G9010<= not I16332;
	G9013<= not I16335;
	G9016<= not I16338;
	G9019<= not I16341;
	G9022<= not I16344;
	G9025<= not I16347;
	G9027<= not G5679;
	G9035<= not I16354;
	G9038<= not I16357;
	G9041<= not I16360;
	G9044<= not I16363;
	G9050<= not G5731;
	G9058<= not I16372;
	G9067<= not G5789;
	G9084<= not G5848;
	G9128<= not I16432;
	G9134<= not I16438;
	G9140<= not I16444;
	G9146<= not I16450;
	G9149<= not I16453;
	G9150<= not G5893;
	G9159<= not I16457;
	G9160<= not G6170;
	G9161<= not G5852;
	G9170<= not I16462;
	G9173<= not I16465;
	G9174<= not G5932;
	G9183<= not I16469;
	G9184<= not I16472;
	G9187<= not G5803;
	G9196<= not I16476;
	G9199<= not I16479;
	G9202<= not I16482;
	G9203<= not G5899;
	G9212<= not I16486;
	G9215<= not I16489;
	G9216<= not G5966;
	G9225<= not I16493;
	G9226<= not G5434;
	G9227<= not G5587;
	G9228<= not G7667;
	G9229<= not I16499;
	G9232<= not G5752;
	G9242<= not I16504;
	G9245<= not I16507;
	G9248<= not G5859;
	G9257<= not I16511;
	G9260<= not I16514;
	G9263<= not I16517;
	G9264<= not G5938;
	G9273<= not I16521;
	G9276<= not I16524;
	G9277<= not G5995;
	G9286<= not G6197;
	G9287<= not G6638;
	G9288<= not G5363;
	G9289<= not G5379;
	G9290<= not I16532;
	G9293<= not G5703;
	G9303<= not I16538;
	G9306<= not I16541;
	G9309<= not I16544;
	G9310<= not G5811;
	G9320<= not I16549;
	G9323<= not I16552;
	G9326<= not G5906;
	G9335<= not I16556;
	G9338<= not I16559;
	G9341<= not I16562;
	G9342<= not G5972;
	G9351<= not I16566;
	G9354<= not I16569;
	G9355<= not G7639;
	G9356<= not G5665;
	G9368<= not I16578;
	G9371<= not I16581;
	G9374<= not G5761;
	G9384<= not I16587;
	G9387<= not I16590;
	G9390<= not I16593;
	G9391<= not G5867;
	G9401<= not I16598;
	G9404<= not I16601;
	G9407<= not G5945;
	G9416<= not I16605;
	G9419<= not I16608;
	G9422<= not I16611;
	G9423<= not G5428;
	G9424<= not G5469;
	G9425<= not G5346;
	G9426<= not G5543;
	G9427<= not G5645;
	G9443<= not I16624;
	G9446<= not I16627;
	G9449<= not I16630;
	G9450<= not I16633;
	G9453<= not G5717;
	G9465<= not I16641;
	G9468<= not I16644;
	G9471<= not G5820;
	G9481<= not I16650;
	G9484<= not I16653;
	G9487<= not I16656;
	G9488<= not G5914;
	G9498<= not I16661;
	G9501<= not I16664;
	G9504<= not G6149;
	G9505<= not G6227;
	G9506<= not G6444;
	G9507<= not G5953;
	G9524<= not I16677;
	G9527<= not G5508;
	G9528<= not I16681;
	G9531<= not I16684;
	G9569<= not G5683;
	G9585<= not I16694;
	G9588<= not I16697;
	G9591<= not I16700;
	G9592<= not I16703;
	G9595<= not G5775;
	G9607<= not I16711;
	G9610<= not I16714;
	G9613<= not G5876;
	G9623<= not I16720;
	G9626<= not I16723;
	G9629<= not I16726;
	G9640<= not I16741;
	G9641<= not I16744;
	G9644<= not I16747;
	G9649<= not G5982;
	G9666<= not I16759;
	G9669<= not G5552;
	G9670<= not I16763;
	G9673<= not I16766;
	G9711<= not G5735;
	G9727<= not I16776;
	G9730<= not I16779;
	G9733<= not I16782;
	G9734<= not I16785;
	G9737<= not G5834;
	G9749<= not I16793;
	G9752<= not I16796;
	G9755<= not G5431;
	G9756<= not G5504;
	G9757<= not G5601;
	G9758<= not G5618;
	G9767<= not I16811;
	G9770<= not I16814;
	G9786<= not I16832;
	G9787<= not I16835;
	G9790<= not I16838;
	G9795<= not G6019;
	G9812<= not I16850;
	G9815<= not G5598;
	G9816<= not I16854;
	G9819<= not I16857;
	G9857<= not G5793;
	G9873<= not I16867;
	G9876<= not I16870;
	G9879<= not I16873;
	G9880<= not I16876;
	G9884<= not G6310;
	G9885<= not G6905;
	G9886<= not G7149;
	G9895<= not I16897;
	G9898<= not I16900;
	G9913<= not I16915;
	G9916<= not I16918;
	G9932<= not I16936;
	G9933<= not I16939;
	G9936<= not I16942;
	G9941<= not G6035;
	G9958<= not I16954;
	G9961<= not G5615;
	G9962<= not I16958;
	G9965<= not I16961;
	G10004<= not I16972;
	G10015<= not G5292;
	G10016<= not I16984;
	G10017<= not I16987;
	G10018<= not I16990;
	G10021<= not I16993;
	G10049<= not I17009;
	G10052<= not I17012;
	G10067<= not I17027;
	G10070<= not I17030;
	G10086<= not I17048;
	G10087<= not I17051;
	G10090<= not I17054;
	G10096<= not I17066;
	G10099<= not G7700;
	G10100<= not I17070;
	G10109<= not I17081;
	G10124<= not G5326;
	G10125<= not I17097;
	G10126<= not I17100;
	G10127<= not I17103;
	G10130<= not I17106;
	G10158<= not I17122;
	G10161<= not I17125;
	G10176<= not I17140;
	G10179<= not I17143;
	G10189<= not I17159;
	G10214<= not I17184;
	G10229<= not G5349;
	G10230<= not I17200;
	G10231<= not I17203;
	G10232<= not I17206;
	G10235<= not I17209;
	G10263<= not I17225;
	G10266<= not I17228;
	G10273<= not I17235;
	G10276<= not I17238;
	G10316<= not I17278;
	G10331<= not G5366;
	G10332<= not I17294;
	G10333<= not I17297;
	G10334<= not I17300;
	G10337<= not I17303;
	G10357<= not I17311;
	G10409<= not I17363;
	G10416<= not I17370;
	G10419<= not I17373;
	G10424<= not G7910;
	G10481<= not G7826;
	G10482<= not I17433;
	G10486<= not G7957;
	G10500<= not G7962;
	G10542<= not I17483;
	G10545<= not I17486;
	G10549<= not G7999;
	G10560<= not G8008;
	G10574<= not G8013;
	G10601<= not I17527;
	G10606<= not G8074;
	G10617<= not G8083;
	G10631<= not G8088;
	G10646<= not I17557;
	G10653<= not G8159;
	G10664<= not G8168;
	G10683<= not G8245;
	G10694<= not G4326;
	G10714<= not G4495;
	G10730<= not G6173;
	G10735<= not G4671;
	G10749<= not G6205;
	G10754<= not G4848;
	G10765<= not G6048;
	G10766<= not G6676;
	G10767<= not G6294;
	G10772<= not G6978;
	G10773<= not G6431;
	G10779<= not I17627;
	G10783<= not G7228;
	G10787<= not I17632;
	G10788<= not G7424;
	G10792<= not I17637;
	G10796<= not I17641;
	G10800<= not I17645;
	G10804<= not I17649;
	G10808<= not I17653;
	G10809<= not G5701;
	G10813<= not I17658;
	G10817<= not I17662;
	G10821<= not I17666;
	G10825<= not I17670;
	G10826<= not I17673;
	G10829<= not G5749;
	G10830<= not I17677;
	G10834<= not I17681;
	G10838<= not I17685;
	G10842<= not I17689;
	G10843<= not I17692;
	G10846<= not G5799;
	G10847<= not G5800;
	G10848<= not G5801;
	G10849<= not I17698;
	G10850<= not I17701;
	G10854<= not I17705;
	G10858<= not I17709;
	G10859<= not I17712;
	G10862<= not I17715;
	G10865<= not G6131;
	G10866<= not G5849;
	G10867<= not G5850;
	G10868<= not I17721;
	G10869<= not I17724;
	G10870<= not I17727;
	G10871<= not I17730;
	G10875<= not I17734;
	G10876<= not I17737;
	G10877<= not I17740;
	G10880<= not I17743;
	G10883<= not I17746;
	G10886<= not G5889;
	G10887<= not I17750;
	G10888<= not I17753;
	G10889<= not I17756;
	G10890<= not I17759;
	G10891<= not I17762;
	G10892<= not I17765;
	G10895<= not I17768;
	G10898<= not I17771;
	G10901<= not I17774;
	G10904<= not G5922;
	G10905<= not G5923;
	G10906<= not G5924;
	G10907<= not I17780;
	G10908<= not I17783;
	G10909<= not I17786;
	G10910<= not I17789;
	G10911<= not I17792;
	G10912<= not I17795;
	G10915<= not I17798;
	G10918<= not I17801;
	G10921<= not I17804;
	G10924<= not I17807;
	G10927<= not G6153;
	G10928<= not G5951;
	G10929<= not G5952;
	G10930<= not I17813;
	G10931<= not I17816;
	G10932<= not I17819;
	G10933<= not I17822;
	G10934<= not I17825;
	G10935<= not I17828;
	G10936<= not I17831;
	G10937<= not I17834;
	G10940<= not I17837;
	G10943<= not I17840;
	G10946<= not I17843;
	G10949<= not I17846;
	G10952<= not I17849;
	G10961<= not G5978;
	G10962<= not G5979;
	G10963<= not I17854;
	G10966<= not I17857;
	G10967<= not I17860;
	G10968<= not I17863;
	G10969<= not I17866;
	G10972<= not I17869;
	G10973<= not I17872;
	G10974<= not I17875;
	G10977<= not I17878;
	G10980<= not I17881;
	G10983<= not I17884;
	G10986<= not G6014;
	G10987<= not G6015;
	G10988<= not I17889;
	G10991<= not I17892;
	G10994<= not I17895;
	G10995<= not I17898;
	G10996<= not I17901;
	G10999<= not I17904;
	G11002<= not I17907;
	G11003<= not I17910;
	G11004<= not I17913;
	G11007<= not I17916;
	G11008<= not I17919;
	G11011<= not I17922;
	G11014<= not I17925;
	G11017<= not I17928;
	G11020<= not G6029;
	G11021<= not G6030;
	G11022<= not I17933;
	G11025<= not I17936;
	G11028<= not I17939;
	G11031<= not I17942;
	G11032<= not I17945;
	G11035<= not I17948;
	G11036<= not I17951;
	G11039<= not I17954;
	G11042<= not I17957;
	G11045<= not I17960;
	G11048<= not I17963;
	G11051<= not I17966;
	G11054<= not I17969;
	G11055<= not I17972;
	G11056<= not I17975;
	G11059<= not I17978;
	G11063<= not I17981;
	G11066<= not I17984;
	G11069<= not G8257;
	G11078<= not G6041;
	G11079<= not I17989;
	G11082<= not I17992;
	G11085<= not I17995;
	G11088<= not I17998;
	G11091<= not I18001;
	G11092<= not I18004;
	G11095<= not I18007;
	G11098<= not I18010;
	G11101<= not I18013;
	G11102<= not I18016;
	G11105<= not I18019;
	G11108<= not I18022;
	G11111<= not I18025;
	G11114<= not I18028;
	G11117<= not I18031;
	G11120<= not I18034;
	G11123<= not I18037;
	G11126<= not I18040;
	G11129<= not I18043;
	G11132<= not I18046;
	G11135<= not I18049;
	G11138<= not I18052;
	G11141<= not I18055;
	G11144<= not I18058;
	G11145<= not I18061;
	G11148<= not I18064;
	G11151<= not I18067;
	G11154<= not I18070;
	G11157<= not I18073;
	G11160<= not I18076;
	G11163<= not I18079;
	G11166<= not I18082;
	G11169<= not I18085;
	G11170<= not I18088;
	G11173<= not I18091;
	G11176<= not I18094;
	G11179<= not I18097;
	G11182<= not I18100;
	G11185<= not I18103;
	G11190<= not G3999;
	G11199<= not I18121;
	G11202<= not I18124;
	G11205<= not I18127;
	G11208<= not I18130;
	G11209<= not I18133;
	G11210<= not I18136;
	G11213<= not I18139;
	G11216<= not I18142;
	G11219<= not I18145;
	G11222<= not I18148;
	G11225<= not I18151;
	G11228<= not I18154;
	G11231<= not I18157;
	G11234<= not I18160;
	G11237<= not I18163;
	G11240<= not I18166;
	G11243<= not I18169;
	G11246<= not I18172;
	G11249<= not I18175;
	G11252<= not I18178;
	G11255<= not I18181;
	G11256<= not I18184;
	G11259<= not I18187;
	G11265<= not I18211;
	G11268<= not I18214;
	G11271<= not I18217;
	G11274<= not I18220;
	G11277<= not I18223;
	G11278<= not I18226;
	G11281<= not I18229;
	G11284<= not I18232;
	G11287<= not I18235;
	G11290<= not I18238;
	G11291<= not I18241;
	G11294<= not I18244;
	G11297<= not I18247;
	G11300<= not I18250;
	G11303<= not I18253;
	G11306<= not I18256;
	G11309<= not I18259;
	G11312<= not I18262;
	G11315<= not I18265;
	G11318<= not I18268;
	G11321<= not I18271;
	G11324<= not I18274;
	G11327<= not I18277;
	G11332<= not G4094;
	G11341<= not I18295;
	G11344<= not I18298;
	G11348<= not I18302;
	G11351<= not I18305;
	G11354<= not I18308;
	G11355<= not I18311;
	G11358<= not I18314;
	G11361<= not I18317;
	G11364<= not I18320;
	G11367<= not I18323;
	G11370<= not I18326;
	G11373<= not I18329;
	G11376<= not I18332;
	G11379<= not I18335;
	G11382<= not I18338;
	G11385<= not I18341;
	G11386<= not I18344;
	G11389<= not I18347;
	G11392<= not I18350;
	G11395<= not I18353;
	G11398<= not I18356;
	G11401<= not I18359;
	G11404<= not I18362;
	G11407<= not I18365;
	G11411<= not I18375;
	G11414<= not I18378;
	G11417<= not I18381;
	G11422<= not I18386;
	G11425<= not I18389;
	G11428<= not I18392;
	G11432<= not I18396;
	G11435<= not I18399;
	G11438<= not I18402;
	G11441<= not I18405;
	G11444<= not I18408;
	G11447<= not I18411;
	G11450<= not I18414;
	G11453<= not I18417;
	G11456<= not I18420;
	G11459<= not I18423;
	G11462<= not I18426;
	G11465<= not I18429;
	G11468<= not I18432;
	G11471<= not I18435;
	G11472<= not I18438;
	G11475<= not I18441;
	G11478<= not I18444;
	G11481<= not G4204;
	G11490<= not G8276;
	G11491<= not I18449;
	G11492<= not I18452;
	G11493<= not I18455;
	G11494<= not I18458;
	G11495<= not I18461;
	G11496<= not I18464;
	G11497<= not I18467;
	G11498<= not I18470;
	G11499<= not I18473;
	G11500<= not I18476;
	G11501<= not I18479;
	G11502<= not I18482;
	G11503<= not I18485;
	G11504<= not I18488;
	G11505<= not I18491;
	G11506<= not I18494;
	G11507<= not I18497;
	G11508<= not I18500;
	G11509<= not I18503;
	G11510<= not I18506;
	G11511<= not I18509;
	G11512<= not I18512;
	G11513<= not I18515;
	G11514<= not I18518;
	G11515<= not I18521;
	G11516<= not I18524;
	G11517<= not I18527;
	G11518<= not I18530;
	G11519<= not I18533;
	G11520<= not I18536;
	G11521<= not I18539;
	G11522<= not I18542;
	G11523<= not I18545;
	G11524<= not I18548;
	G11525<= not I18551;
	G11526<= not I18554;
	G11527<= not I18557;
	G11528<= not I18560;
	G11529<= not I18563;
	G11530<= not I18566;
	G11531<= not I18569;
	G11532<= not I18572;
	G11533<= not I18575;
	G11534<= not I18578;
	G11535<= not I18581;
	G11536<= not I18584;
	G11537<= not I18587;
	G11538<= not I18590;
	G11539<= not I18593;
	G11540<= not I18596;
	G11541<= not I18599;
	G11542<= not I18602;
	G11543<= not I18605;
	G11544<= not I18608;
	G11545<= not I18611;
	G11546<= not I18614;
	G11547<= not I18617;
	G11548<= not I18620;
	G11549<= not I18623;
	G11550<= not I18626;
	G11551<= not I18629;
	G11552<= not I18632;
	G11553<= not I18635;
	G11554<= not I18638;
	G11555<= not I18641;
	G11556<= not I18644;
	G11557<= not I18647;
	G11558<= not I18650;
	G11559<= not I18653;
	G11560<= not I18656;
	G11561<= not I18659;
	G11562<= not I18662;
	G11563<= not I18665;
	G11564<= not I18668;
	G11565<= not I18671;
	G11566<= not I18674;
	G11567<= not I18677;
	G11568<= not I18680;
	G11569<= not I18683;
	G11570<= not I18686;
	G11571<= not I18689;
	G11572<= not I18692;
	G11573<= not I18695;
	G11574<= not I18698;
	G11575<= not I18701;
	G11576<= not I18704;
	G11577<= not I18707;
	G11578<= not I18710;
	G11579<= not I18713;
	G11580<= not I18716;
	G11581<= not I18719;
	G11582<= not I18722;
	G11583<= not I18725;
	G11584<= not I18728;
	G11585<= not I18731;
	G11586<= not I18734;
	G11587<= not I18737;
	G11588<= not I18740;
	G11589<= not I18743;
	G11590<= not I18746;
	G11591<= not I18749;
	G11592<= not I18752;
	G11593<= not I18755;
	G11594<= not I18758;
	G11595<= not I18761;
	G11596<= not I18764;
	G11597<= not I18767;
	G11598<= not I18770;
	G11599<= not I18773;
	G11603<= not I18777;
	G11606<= not I18780;
	G11608<= not I18784;
	G11611<= not I18787;
	G11613<= not I18791;
	G11616<= not I18794;
	G11620<= not G10601;
	G11623<= not G10961;
	G11628<= not I18810;
	G11629<= not I18813;
	G11633<= not I18817;
	G11636<= not I18820;
	G11638<= not I18824;
	G11641<= not I18827;
	G11642<= not G10646;
	G11651<= not I18835;
	G11652<= not I18838;
	G11656<= not I18842;
	G11659<= not I18845;
	G11670<= not I18854;
	G11671<= not I18857;
	G11682<= not I18866;
	G11706<= not G10928;
	G11732<= not G10826;
	G11734<= not G10843;
	G11735<= not G10859;
	G11736<= not G10862;
	G11737<= not G10809;
	G11740<= not G10877;
	G11741<= not G10880;
	G11742<= not G10883;
	G11743<= not G8530;
	G11745<= not G10892;
	G11746<= not G10895;
	G11747<= not G10898;
	G11748<= not G10901;
	G11749<= not I18929;
	G11758<= not G8514;
	G11761<= not G10912;
	G11762<= not G10915;
	G11763<= not G10918;
	G11764<= not G10921;
	G11765<= not G10924;
	G11766<= not G10886;
	G11769<= not I18943;
	G11770<= not G10932;
	G11774<= not G10937;
	G11775<= not G10940;
	G11776<= not G10943;
	G11777<= not G10946;
	G11778<= not G10949;
	G11779<= not G10906;
	G11782<= not G10963;
	G11783<= not G10966;
	G11786<= not I18962;
	G11787<= not G10969;
	G11791<= not I18969;
	G11794<= not G10974;
	G11795<= not G10977;
	G11796<= not G10980;
	G11797<= not G10983;
	G11798<= not G10867;
	G11801<= not G10988;
	G11802<= not G10991;
	G11803<= not G10994;
	G11804<= not G10995;
	G11808<= not G10996;
	G11809<= not G10999;
	G11812<= not I18990;
	G11813<= not G11004;
	G11817<= not G11008;
	G11818<= not G11011;
	G11819<= not G11014;
	G11820<= not G11017;
	G11821<= not G10848;
	G11824<= not G11022;
	G11825<= not G11025;
	G11826<= not G11028;
	G11827<= not G11032;
	G11829<= not G11035;
	G11834<= not G11036;
	G11835<= not G11039;
	G11836<= not G11042;
	G11837<= not G11045;
	G11841<= not G11048;
	G11842<= not G11051;
	G11845<= not I19025;
	G11846<= not G11056;
	G11848<= not I19030;
	G11852<= not G11063;
	G11853<= not G11066;
	G11854<= not G11078;
	G11856<= not G11079;
	G11857<= not G11082;
	G11858<= not G11085;
	G11859<= not G11088;
	G11862<= not G11091;
	G11866<= not G11092;
	G11867<= not G11095;
	G11868<= not G11098;
	G11869<= not G11102;
	G11871<= not G11105;
	G11876<= not G11108;
	G11877<= not G11111;
	G11878<= not G11114;
	G11879<= not G11117;
	G11883<= not G11120;
	G11884<= not G11123;
	G11886<= not G11126;
	G11887<= not G11129;
	G11888<= not G11021;
	G11891<= not G11132;
	G11892<= not G11135;
	G11893<= not G11138;
	G11894<= not G11141;
	G11895<= not G11144;
	G11898<= not G11145;
	G11899<= not G11148;
	G11900<= not G11151;
	G11901<= not G11154;
	G11904<= not G11157;
	G11908<= not G11160;
	G11909<= not G11163;
	G11910<= not G11166;
	G11911<= not G11170;
	G11913<= not G11173;
	G11918<= not G11176;
	G11919<= not G11179;
	G11920<= not G11182;
	G11921<= not G11185;
	G11923<= not I19105;
	G11927<= not G10987;
	G11929<= not G11199;
	G11930<= not G11202;
	G11931<= not G11205;
	G11932<= not G11209;
	G11933<= not G11210;
	G11936<= not G11213;
	G11937<= not I19119;
	G11941<= not G11216;
	G11942<= not G11219;
	G11943<= not G11222;
	G11944<= not G11225;
	G11945<= not G11228;
	G11948<= not G11231;
	G11949<= not G11234;
	G11950<= not G11237;
	G11951<= not G11240;
	G11954<= not G11243;
	G11958<= not G11246;
	G11959<= not G11249;
	G11960<= not G11252;
	G11961<= not G11256;
	G11963<= not G11259;
	G11968<= not G11265;
	G11969<= not G11268;
	G11970<= not G11271;
	G11971<= not G11274;
	G11972<= not G11277;
	G11973<= not G11278;
	G11976<= not I19160;
	G11982<= not G11281;
	G11983<= not G11284;
	G11984<= not G11287;
	G11985<= not G11291;
	G11986<= not G11294;
	G11989<= not G11297;
	G11990<= not I19174;
	G11994<= not G11300;
	G11995<= not G11303;
	G11996<= not G11306;
	G11997<= not G11309;
	G11998<= not G11312;
	G12001<= not G11315;
	G12002<= not G11318;
	G12003<= not G11321;
	G12004<= not G11324;
	G12007<= not G11327;
	G12009<= not I19195;
	G12013<= not G10772;
	G12017<= not G10100;
	G12020<= not G11341;
	G12021<= not G11344;
	G12022<= not G11348;
	G12023<= not G11351;
	G12024<= not G11354;
	G12025<= not G11355;
	G12027<= not I19208;
	G12030<= not I19211;
	G12037<= not G11358;
	G12038<= not G11361;
	G12039<= not G11364;
	G12040<= not G11367;
	G12041<= not G11370;
	G12042<= not G11373;
	G12045<= not I19226;
	G12051<= not G11376;
	G12052<= not G11379;
	G12053<= not G11382;
	G12054<= not G11386;
	G12055<= not G11389;
	G12058<= not G11392;
	G12059<= not I19240;
	G12063<= not G11395;
	G12064<= not G11398;
	G12065<= not G11401;
	G12066<= not G11404;
	G12067<= not G11407;
	G12071<= not G10783;
	G12075<= not G11411;
	G12076<= not G11414;
	G12077<= not G11417;
	G12078<= not G11422;
	G12084<= not G11425;
	G12085<= not G11428;
	G12086<= not G11432;
	G12087<= not G11435;
	G12088<= not G11438;
	G12089<= not G11441;
	G12091<= not I19271;
	G12094<= not I19274;
	G12101<= not G11444;
	G12102<= not G11447;
	G12103<= not G11450;
	G12104<= not G11453;
	G12105<= not G11456;
	G12106<= not G11459;
	G12109<= not I19289;
	G12115<= not G11462;
	G12116<= not G11465;
	G12117<= not G11468;
	G12118<= not G11472;
	G12119<= not G11475;
	G12122<= not G11478;
	G12123<= not I19303;
	G12125<= not I19307;
	G12130<= not G10788;
	G12134<= not G8321;
	G12135<= not G8324;
	G12136<= not I19315;
	G12139<= not I19318;
	G12142<= not I19321;
	G12147<= not G8330;
	G12148<= not G8333;
	G12149<= not G8336;
	G12150<= not G8341;
	G12156<= not G8344;
	G12157<= not G8347;
	G12158<= not G8351;
	G12159<= not G8354;
	G12160<= not G8357;
	G12161<= not G8360;
	G12163<= not I19342;
	G12166<= not I19345;
	G12173<= not G8363;
	G12174<= not G8366;
	G12175<= not G8369;
	G12176<= not G8372;
	G12177<= not G8375;
	G12178<= not G8378;
	G12181<= not I19360;
	G12187<= not G8285;
	G12191<= not G8382;
	G12196<= not G8388;
	G12197<= not G8391;
	G12198<= not I19374;
	G12201<= not I19377;
	G12204<= not I19380;
	G12209<= not G8397;
	G12210<= not G8400;
	G12211<= not G8403;
	G12212<= not G8408;
	G12218<= not G8411;
	G12219<= not G8414;
	G12220<= not G8418;
	G12221<= not G8421;
	G12222<= not G8424;
	G12223<= not G8427;
	G12225<= not I19401;
	G12228<= not I19404;
	G12235<= not G8294;
	G12239<= not I19412;
	G12242<= not I19415;
	G12246<= not G8434;
	G12251<= not G8440;
	G12252<= not G8443;
	G12253<= not I19426;
	G12256<= not I19429;
	G12259<= not I19432;
	G12264<= not G8449;
	G12265<= not G8452;
	G12266<= not G8455;
	G12267<= not G8460;
	G12275<= not G8303;
	G12279<= not I19449;
	G12282<= not I19452;
	G12285<= not I19455;
	G12289<= not G8469;
	G12294<= not G8475;
	G12295<= not G8478;
	G12296<= not I19466;
	G12299<= not I19469;
	G12302<= not I19472;
	G12308<= not G8312;
	G12312<= not I19479;
	G12315<= not I19482;
	G12318<= not I19485;
	G12321<= not I19488;
	G12325<= not G8494;
	G12332<= not G10829;
	G12333<= not I19500;
	G12336<= not I19503;
	G12340<= not I19507;
	G12343<= not I19510;
	G12346<= not I19513;
	G12349<= not I19516;
	G12354<= not G8381;
	G12362<= not G10866;
	G12363<= not I19523;
	G12366<= not I19526;
	G12370<= not I19530;
	G12373<= not I19533;
	G12378<= not G10847;
	G12379<= not I19539;
	G12382<= not I19542;
	G12385<= not I19545;
	G12389<= not I19549;
	G12392<= not I19552;
	G12408<= not G11020;
	G12409<= not I19557;
	G12412<= not I19560;
	G12415<= not I19563;
	G12420<= not G10986;
	G12421<= not I19569;
	G12424<= not G10962;
	G12425<= not I19573;
	G12426<= not I19576;
	G12430<= not G10905;
	G12432<= not I19582;
	G12434<= not G10929;
	G12435<= not I19587;
	G12437<= not I19591;
	G12438<= not G10846;
	G12439<= not I19595;
	G12440<= not I19598;
	G12442<= not I19602;
	G12443<= not I19605;
	G12444<= not I19608;
	G12445<= not I19611;
	G12447<= not I19615;
	G12448<= not I19618;
	G12449<= not I19621;
	G12450<= not I19624;
	G12452<= not I19628;
	G12453<= not I19631;
	G12454<= not I19634;
	G12455<= not I19637;
	G12456<= not G8602;
	G12460<= not I19642;
	G12461<= not I19645;
	G12462<= not I19648;
	G12463<= not G10730;
	G12466<= not G8614;
	G12470<= not I19654;
	G12471<= not I19657;
	G12472<= not G8617;
	G12473<= not G8580;
	G12476<= not G8622;
	G12478<= not G10749;
	G12481<= not G8627;
	G12485<= not I19667;
	G12490<= not G8587;
	G12493<= not G8632;
	G12495<= not G10767;
	G12498<= not G8637;
	G12502<= not G8640;
	G12504<= not G8643;
	G12505<= not G8646;
	G12510<= not G8594;
	G12513<= not G8651;
	G12515<= not G10773;
	G12518<= not G8655;
	G12519<= not I19689;
	G12521<= not G8659;
	G12522<= not G8662;
	G12527<= not G8605;
	G12530<= not G8667;
	G12532<= not G8670;
	G12533<= not G8673;
	G12534<= not I19702;
	G12536<= not G8678;
	G12537<= not G8681;
	G12542<= not G8684;
	G12543<= not I19711;
	G12545<= not G8690;
	G12546<= not G8693;
	G12547<= not G8696;
	G12548<= not I19718;
	G12551<= not G8700;
	G12552<= not I19722;
	G12553<= not G8708;
	G12554<= not G8711;
	G12555<= not I19727;
	G12558<= not G8714;
	G12559<= not G8719;
	G12560<= not G8745;
	G12561<= not I19733;
	G12564<= not I19736;
	G12565<= not I19739;
	G12596<= not G8748;
	G12597<= not G8752;
	G12598<= not G8757;
	G12599<= not G8763;
	G12600<= not G8766;
	G12601<= not I19747;
	G12604<= not I19750;
	G12607<= not I19753;
	G12608<= not I19756;
	G12611<= not I19759;
	G12642<= not G8771;
	G12643<= not G8775;
	G12644<= not G8780;
	G12645<= not G8785;
	G12646<= not G8788;
	G12647<= not I19767;
	G12651<= not I19771;
	G12654<= not I19774;
	G12657<= not I19777;
	G12688<= not G8794;
	G12689<= not G8798;
	G12690<= not G8802;
	G12691<= not G8805;
	G12692<= not I19784;
	G12695<= not I19787;
	G12699<= not I19791;
	G12702<= not I19794;
	G12705<= not I19797;
	G12708<= not I19800;
	G12711<= not I19803;
	G12742<= not G8813;
	G12743<= not G8817;
	G12744<= not I19808;
	G12748<= not G8823;
	G12749<= not I19813;
	G12752<= not I19816;
	G12756<= not I19820;
	G12759<= not I19823;
	G12762<= not I19826;
	G12765<= not I19829;
	G12768<= not G8829;
	G12769<= not I19833;
	G12772<= not I19836;
	G12775<= not G8832;
	G12776<= not G10766;
	G12782<= not G8836;
	G12783<= not I19844;
	G12786<= not I19847;
	G12790<= not G8847;
	G12791<= not I19852;
	G12794<= not I19855;
	G12798<= not I19859;
	G12801<= not I19862;
	G12804<= not I19865;
	G12807<= not G8853;
	G12808<= not I19869;
	G12811<= not I19872;
	G12815<= not G8856;
	G12816<= not I19877;
	G12821<= not G8863;
	G12822<= not I19883;
	G12825<= not I19886;
	G12829<= not G8874;
	G12830<= not I19891;
	G12833<= not I19894;
	G12837<= not I19898;
	G12840<= not I19901;
	G12843<= not G8879;
	G12844<= not I19905;
	G12847<= not G8882;
	G12848<= not G11059;
	G12850<= not G8885;
	G12851<= not G8888;
	G12853<= not G8894;
	G12854<= not I19915;
	G12859<= not G8901;
	G12860<= not I19921;
	G12863<= not I19924;
	G12867<= not G8912;
	G12868<= not I19929;
	G12871<= not I19932;
	G12874<= not G8915;
	G12875<= not G10779;
	G12881<= not G8918;
	G12882<= not G8921;
	G12891<= not G8925;
	G12892<= not G8928;
	G12894<= not G8934;
	G12895<= not I19952;
	G12900<= not G8941;
	G12901<= not I19958;
	G12904<= not I19961;
	G12907<= not G8949;
	G12909<= not G10904;
	G12914<= not G8952;
	G12915<= not G8955;
	G12921<= not G8958;
	G12922<= not G8961;
	G12931<= not G8965;
	G12932<= not G8968;
	G12934<= not G8974;
	G12935<= not I19986;
	G12940<= not G8980;
	G12943<= not G8984;
	G12944<= not G8987;
	G12950<= not G8990;
	G12951<= not G8993;
	G12960<= not G8997;
	G12961<= not G9000;
	G12962<= not I20009;
	G12965<= not G9006;
	G12969<= not G9010;
	G12972<= not G9013;
	G12973<= not G9016;
	G12979<= not G9019;
	G12980<= not G9022;
	G12993<= not G9035;
	G12996<= not G9038;
	G12997<= not G9041;
	G12998<= not G9044;
	G13003<= not G9058;
	G13011<= not I20062;
	G13025<= not G10810;
	G13033<= not G10797;
	G13036<= not G10831;
	G13043<= not G10789;
	G13046<= not G10814;
	G13049<= not G10851;
	G13057<= not G10784;
	G13060<= not G10801;
	G13063<= not G10835;
	G13066<= not G10872;
	G13070<= not I20117;
	G13073<= not G10793;
	G13076<= not G10818;
	G13079<= not G10855;
	G13092<= not G10805;
	G13095<= not G10839;
	G13101<= not G9128;
	G13107<= not G10822;
	G13117<= not G9134;
	G13130<= not G9140;
	G13141<= not G9146;
	G13148<= not G9170;
	G13151<= not G9184;
	G13152<= not G9196;
	G13153<= not G9199;
	G13154<= not G9212;
	G13157<= not G9229;
	G13158<= not G9242;
	G13159<= not G9245;
	G13161<= not G9257;
	G13162<= not G9260;
	G13163<= not G9273;
	G13166<= not G9290;
	G13167<= not G9303;
	G13168<= not G9306;
	G13169<= not G9320;
	G13170<= not G9323;
	G13172<= not G9335;
	G13173<= not G9338;
	G13174<= not G9351;
	G13176<= not G9368;
	G13177<= not G9371;
	G13178<= not G9384;
	G13179<= not G9387;
	G13180<= not G9401;
	G13181<= not G9404;
	G13183<= not G9416;
	G13184<= not G9419;
	G13185<= not G9443;
	G13186<= not G9446;
	G13187<= not G9450;
	G13188<= not G9465;
	G13189<= not G9468;
	G13190<= not G9481;
	G13191<= not G9484;
	G13192<= not G9498;
	G13193<= not G9501;
	G13195<= not G9524;
	G13196<= not G9528;
	G13197<= not G9531;
	G13198<= not G9585;
	G13199<= not G9588;
	G13200<= not G9592;
	G13201<= not G9607;
	G13202<= not G9610;
	G13203<= not G9623;
	G13204<= not G9626;
	G13205<= not G9641;
	G13206<= not G9644;
	G13207<= not G9666;
	G13208<= not G9670;
	G13209<= not G9673;
	G13210<= not G9727;
	G13211<= not G9730;
	G13212<= not G9734;
	G13213<= not G9749;
	G13214<= not G9752;
	G13215<= not I20264;
	G13218<= not G9767;
	G13219<= not G9770;
	G13220<= not G9787;
	G13221<= not G9790;
	G13222<= not G9812;
	G13223<= not G9816;
	G13224<= not G9819;
	G13225<= not G9873;
	G13226<= not G9876;
	G13227<= not G9880;
	G13229<= not I20278;
	G13232<= not G9895;
	G13233<= not G9898;
	G13234<= not I20283;
	G13237<= not G9913;
	G13238<= not G9916;
	G13239<= not G9933;
	G13240<= not G9936;
	G13241<= not G9958;
	G13242<= not G9962;
	G13243<= not G9965;
	G13244<= not G10004;
	G13246<= not I20295;
	G13248<= not I20299;
	G13249<= not G10018;
	G13250<= not G10021;
	G13252<= not I20305;
	G13255<= not G10049;
	G13256<= not G10052;
	G13257<= not I20310;
	G13260<= not G10067;
	G13261<= not G10070;
	G13262<= not G10087;
	G13263<= not G10090;
	G13264<= not G10096;
	G13265<= not G8568;
	G13267<= not I20320;
	G13268<= not G10109;
	G13269<= not I20324;
	G13271<= not I20328;
	G13272<= not G10127;
	G13273<= not G10130;
	G13275<= not I20334;
	G13278<= not G10158;
	G13279<= not G10161;
	G13280<= not I20339;
	G13283<= not G10176;
	G13284<= not G10179;
	G13285<= not G10189;
	G13290<= not I20347;
	G13292<= not I20351;
	G13293<= not G10214;
	G13294<= not I20355;
	G13296<= not I20359;
	G13297<= not G10232;
	G13298<= not G10235;
	G13300<= not I20365;
	G13303<= not G10263;
	G13304<= not G10266;
	G13308<= not G10273;
	G13309<= not G10276;
	G13317<= not I20376;
	G13318<= not I20379;
	G13319<= not I20382;
	G13321<= not I20386;
	G13323<= not I20390;
	G13324<= not G10316;
	G13325<= not I20394;
	G13327<= not I20398;
	G13328<= not G10334;
	G13329<= not G10337;
	G13330<= not G10357;
	G13336<= not I20407;
	G13339<= not I20410;
	G13341<= not I20414;
	G13342<= not I20417;
	G13344<= not I20421;
	G13346<= not I20425;
	G13347<= not G10409;
	G13351<= not G10416;
	G13352<= not G10419;
	G13356<= not I20441;
	G13359<= not I20444;
	G13361<= not I20448;
	G13364<= not I20451;
	G13366<= not I20455;
	G13367<= not I20458;
	G13369<= not I20462;
	G13373<= not G10482;
	G13381<= not I20476;
	G13384<= not I20479;
	G13386<= not I20483;
	G13389<= not I20486;
	G13391<= not I20490;
	G13394<= not I20493;
	G13396<= not I20497;
	G13397<= not I20500;
	G13398<= not G10542;
	G13400<= not G10545;
	G13405<= not I20514;
	G13406<= not I20517;
	G13407<= not I20520;
	G13408<= not I20523;
	G13409<= not I20526;
	G13410<= not I20529;
	G13411<= not I20532;
	G13412<= not I20535;
	G13413<= not I20538;
	G13414<= not I20541;
	G13415<= not I20544;
	G13416<= not I20547;
	G13417<= not I20550;
	G13418<= not I20553;
	G13419<= not I20556;
	G13420<= not I20559;
	G13421<= not I20562;
	G13422<= not I20565;
	G13423<= not I20568;
	G13424<= not I20571;
	G13425<= not I20574;
	G13426<= not I20577;
	G13427<= not I20580;
	G13428<= not I20583;
	G13429<= not I20586;
	G13430<= not I20589;
	G13431<= not I20592;
	G13432<= not I20595;
	G13433<= not I20598;
	G13434<= not I20601;
	G13435<= not I20604;
	G13436<= not I20607;
	G13437<= not I20610;
	G13438<= not I20613;
	G13439<= not I20616;
	G13440<= not I20619;
	G13441<= not I20622;
	G13442<= not I20625;
	G13443<= not I20628;
	G13444<= not I20631;
	G13445<= not I20634;
	G13446<= not I20637;
	G13447<= not I20640;
	G13448<= not I20643;
	G13449<= not I20646;
	G13450<= not I20649;
	G13451<= not I20652;
	G13452<= not I20655;
	G13453<= not I20658;
	G13454<= not I20661;
	G13455<= not I20664;
	G13456<= not I20667;
	G13457<= not I20670;
	G13458<= not I20673;
	G13459<= not I20676;
	G13460<= not I20679;
	G13461<= not I20682;
	G13462<= not I20685;
	G13463<= not I20688;
	G13464<= not I20691;
	G13465<= not I20694;
	G13466<= not I20697;
	G13467<= not I20700;
	G13468<= not I20703;
	G13469<= not I20706;
	G13475<= not I20709;
	G13519<= not G13228;
	G13530<= not G13251;
	G13541<= not G13274;
	G13552<= not G13299;
	G13565<= not G12192;
	G13568<= not G11627;
	G13571<= not I20791;
	G13572<= not I20794;
	G13573<= not G12247;
	G13576<= not G11650;
	G13579<= not I20799;
	G13580<= not I20802;
	G13581<= not I20805;
	G13582<= not G12290;
	G13585<= not G11669;
	G13588<= not I20810;
	G13589<= not I20813;
	G13598<= not I20816;
	G13600<= not I20820;
	G13601<= not I20823;
	G13602<= not G12326;
	G13605<= not G11681;
	G13608<= not I20828;
	G13610<= not I20832;
	G13612<= not I20836;
	G13613<= not I20839;
	G13614<= not G11690;
	G13620<= not I20844;
	G13622<= not I20848;
	G13624<= not I20852;
	G13626<= not G11697;
	G13632<= not I20858;
	G13635<= not I20863;
	G13637<= not G11703;
	G13644<= not G13215;
	G13647<= not I20873;
	G13649<= not G11711;
	G13657<= not G12452;
	G13669<= not G13229;
	G13670<= not G13234;
	G13673<= not I20886;
	G13677<= not G12447;
	G13687<= not G12460;
	G13699<= not G13252;
	G13700<= not G13257;
	G13706<= not G12443;
	G13714<= not G12453;
	G13724<= not G12470;
	G13736<= not G13275;
	G13737<= not G13280;
	G13741<= not I20909;
	G13750<= not G12439;
	G13756<= not G12448;
	G13764<= not G12461;
	G13774<= not G12485;
	G13786<= not G13300;
	G13791<= not G12444;
	G13797<= not G12454;
	G13805<= not G12471;
	G13817<= not G13336;
	G13819<= not G12449;
	G13825<= not G12462;
	G13836<= not G13356;
	G13838<= not G13361;
	G13840<= not G12455;
	G13848<= not G11744;
	G13849<= not G13381;
	G13850<= not G13386;
	G13852<= not G13391;
	G13856<= not G11759;
	G13857<= not G11760;
	G13858<= not G11603;
	G13859<= not G11608;
	G13861<= not G11613;
	G13863<= not I20959;
	G13864<= not G11767;
	G13866<= not G11772;
	G13867<= not G11773;
	G13868<= not G11633;
	G13869<= not G11638;
	G13872<= not G11780;
	G13873<= not G12698;
	G13879<= not G11784;
	G13881<= not G11789;
	G13882<= not G11790;
	G13883<= not G11656;
	G13885<= not G11799;
	G13886<= not G12747;
	G13894<= not G11806;
	G13895<= not G12755;
	G13901<= not G11810;
	G13903<= not G11815;
	G13906<= not G11822;
	G13907<= not G12781;
	G13918<= not G11830;
	G13922<= not G11831;
	G13926<= not G11832;
	G13927<= not G12789;
	G13935<= not G11839;
	G13936<= not G12797;
	G13942<= not G11843;
	G13945<= not G11855;
	G13946<= not G12814;
	G13954<= not I21012;
	G13958<= not G11863;
	G13962<= not G11864;
	G13963<= not G12820;
	G13974<= not G11872;
	G13978<= not G11873;
	G13982<= not G11874;
	G13983<= not G12828;
	G13991<= not G11881;
	G13992<= not G12836;
	G13999<= not G11889;
	G14000<= not G11890;
	G14001<= not G12849;
	G14008<= not I21037;
	G14011<= not G11896;
	G14015<= not G11897;
	G14016<= not G12852;
	G14024<= not I21045;
	G14028<= not G11905;
	G14032<= not G11906;
	G14033<= not G12858;
	G14044<= not G11914;
	G14048<= not G11915;
	G14052<= not G11916;
	G14053<= not G12866;
	G14061<= not G11928;
	G14062<= not G12880;
	G14068<= not I21064;
	G14071<= not G11934;
	G14079<= not G11935;
	G14086<= not G11938;
	G14090<= not G11939;
	G14091<= not G11940;
	G14092<= not G12890;
	G14099<= not I21075;
	G14102<= not G11946;
	G14106<= not G11947;
	G14107<= not G12893;
	G14115<= not I21083;
	G14119<= not G11955;
	G14123<= not G11956;
	G14124<= not G12899;
	G14135<= not G11964;
	G14139<= not G11965;
	G14144<= not I21096;
	G14148<= not G12912;
	G14153<= not G12913;
	G14158<= not G11974;
	G14165<= not G11975;
	G14171<= not G11979;
	G14175<= not G11980;
	G14176<= not G11981;
	G14177<= not G12920;
	G14183<= not I21108;
	G14186<= not G11987;
	G14194<= not G11988;
	G14201<= not G11991;
	G14205<= not G11992;
	G14206<= not G11993;
	G14207<= not G12930;
	G14214<= not I21119;
	G14217<= not G11999;
	G14221<= not G12000;
	G14222<= not G12933;
	G14230<= not I21127;
	G14234<= not G12008;
	G14238<= not G12939;
	G14244<= not G12026;
	G14249<= not G12034;
	G14252<= not G12035;
	G14256<= not G12036;
	G14259<= not I21137;
	G14263<= not G12941;
	G14268<= not G12942;
	G14273<= not G12043;
	G14280<= not G12044;
	G14286<= not G12048;
	G14290<= not G12049;
	G14291<= not G12050;
	G14292<= not G12949;
	G14298<= not I21149;
	G14301<= not G12056;
	G14309<= not G12057;
	G14316<= not G12060;
	G14320<= not G12061;
	G14321<= not G12062;
	G14322<= not G12959;
	G14329<= not I21160;
	G14332<= not G12068;
	G14337<= not I21165;
	G14342<= not G12967;
	G14347<= not G12079;
	G14352<= not G12081;
	G14355<= not G12082;
	G14359<= not G12083;
	G14360<= not G12968;
	G14366<= not G12090;
	G14371<= not G12098;
	G14374<= not G12099;
	G14378<= not G12100;
	G14381<= not I21178;
	G14385<= not G12970;
	G14390<= not G12971;
	G14395<= not G12107;
	G14402<= not G12108;
	G14408<= not G12112;
	G14412<= not G12113;
	G14413<= not G12114;
	G14414<= not G12978;
	G14420<= not I21190;
	G14423<= not G12120;
	G14431<= not G12121;
	G14438<= not G12124;
	G14442<= not G11768;
	G14450<= not G12146;
	G14454<= not G12991;
	G14459<= not G12151;
	G14464<= not G12153;
	G14467<= not G12154;
	G14471<= not G12155;
	G14472<= not G12992;
	G14478<= not G12162;
	G14483<= not G12170;
	G14486<= not G12171;
	G14490<= not G12172;
	G14493<= not I21208;
	G14497<= not G12994;
	G14502<= not G12995;
	G14507<= not G12179;
	G14514<= not G12180;
	G14520<= not G12184;
	G14524<= not G12185;
	G14525<= not G12195;
	G14529<= not G11785;
	G14537<= not G12208;
	G14541<= not G13001;
	G14546<= not G12213;
	G14551<= not G12215;
	G14554<= not G12216;
	G14558<= not G12217;
	G14559<= not G13002;
	G14565<= not G12224;
	G14570<= not G12232;
	G14573<= not G12233;
	G14577<= not G12234;
	G14580<= not G12250;
	G14584<= not G11811;
	G14592<= not G12263;
	G14596<= not G13022;
	G14601<= not G12268;
	G14606<= not G12270;
	G14609<= not G12271;
	G14613<= not G12272;
	G14614<= not G12293;
	G14618<= not G11844;
	G14626<= not G12306;
	G14630<= not I21241;
	G14637<= not G12329;
	G14641<= not G11823;
	G14642<= not I21246;
	G14650<= not I21249;
	G14657<= not I21252;
	G14668<= not G11865;
	G14669<= not I21256;
	G14677<= not I21259;
	G14684<= not I21262;
	G14685<= not G12245;
	G14691<= not I21267;
	G14702<= not G11907;
	G14703<= not I21271;
	G14711<= not I21274;
	G14718<= not I21277;
	G14719<= not G12288;
	G14725<= not I21282;
	G14736<= not G11957;
	G14737<= not I21286;
	G14745<= not I21289;
	G14746<= not I21292;
	G14747<= not G12324;
	G14753<= not I21297;
	G14764<= not G11791;
	G14765<= not I21301;
	G14766<= not I21304;
	G14768<= not G12352;
	G14774<= not I21310;
	G14775<= not I21313;
	G14776<= not G12033;
	G14794<= not G11848;
	G14795<= not I21318;
	G14796<= not I21321;
	G14797<= not G12080;
	G14811<= not G12097;
	G14829<= not I21326;
	G14830<= not I21329;
	G14831<= not G11828;
	G14837<= not G12145;
	G14849<= not G12152;
	G14863<= not G12169;
	G14881<= not G11923;
	G14882<= not I21337;
	G14883<= not I21340;
	G14885<= not G11860;
	G14895<= not G12193;
	G14904<= not G11870;
	G14910<= not G12207;
	G14922<= not G12214;
	G14936<= not G12231;
	G14954<= not I21351;
	G14955<= not I21354;
	G14959<= not G11976;
	G14960<= not I21361;
	G14963<= not I21364;
	G14966<= not G11902;
	G14976<= not G12248;
	G14985<= not G11912;
	G14991<= not G12262;
	G15003<= not G12269;
	G15017<= not G12009;
	G15018<= not I21374;
	G15019<= not I21377;
	G15021<= not I21381;
	G15022<= not G11781;
	G15032<= not G12027;
	G15033<= not G12030;
	G15034<= not I21389;
	G15037<= not I21392;
	G15040<= not I21395;
	G15043<= not I21398;
	G15048<= not G12045;
	G15049<= not I21404;
	G15052<= not I21407;
	G15055<= not G11952;
	G15065<= not G12291;
	G15074<= not G11962;
	G15080<= not G12305;
	G15092<= not I21415;
	G15095<= not I21420;
	G15096<= not G11800;
	G15106<= not I21426;
	G15109<= not I21429;
	G15112<= not I21432;
	G15115<= not I21435;
	G15118<= not G11807;
	G15128<= not G12091;
	G15129<= not G12094;
	G15130<= not I21443;
	G15133<= not I21446;
	G15136<= not I21449;
	G15139<= not I21452;
	G15144<= not G12109;
	G15145<= not I21458;
	G15148<= not I21461;
	G15151<= not G12005;
	G15161<= not G12327;
	G15170<= not G12125;
	G15174<= not G12136;
	G15175<= not G12139;
	G15176<= not G12142;
	G15177<= not G12339;
	G15179<= not I21476;
	G15182<= not I21479;
	G15185<= not I21482;
	G15188<= not G11833;
	G15198<= not I21488;
	G15201<= not I21491;
	G15204<= not I21494;
	G15207<= not I21497;
	G15210<= not G11840;
	G15220<= not G12163;
	G15221<= not G12166;
	G15222<= not I21505;
	G15225<= not I21508;
	G15228<= not I21511;
	G15231<= not I21514;
	G15236<= not G12181;
	G15237<= not I21520;
	G15240<= not I21523;
	G15248<= not I21531;
	G15251<= not I21534;
	G15254<= not I21537;
	G15260<= not G12198;
	G15261<= not G12201;
	G15262<= not G12204;
	G15263<= not G12369;
	G15265<= not I21548;
	G15268<= not I21551;
	G15271<= not I21554;
	G15274<= not G11875;
	G15284<= not I21560;
	G15287<= not I21563;
	G15290<= not I21566;
	G15293<= not I21569;
	G15296<= not G11882;
	G15306<= not G12225;
	G15307<= not G12228;
	G15308<= not I21577;
	G15311<= not I21580;
	G15314<= not I21583;
	G15317<= not I21586;
	G15322<= not G12239;
	G15323<= not G12242;
	G15326<= not I21595;
	G15329<= not I21598;
	G15332<= not I21601;
	G15340<= not I21609;
	G15343<= not I21612;
	G15346<= not I21615;
	G15352<= not G12253;
	G15353<= not G12256;
	G15354<= not G12259;
	G15355<= not G12388;
	G15357<= not I21626;
	G15360<= not I21629;
	G15363<= not I21632;
	G15366<= not G11917;
	G15376<= not I21638;
	G15379<= not I21641;
	G15382<= not I21644;
	G15385<= not I21647;
	G15390<= not G12279;
	G15393<= not I21655;
	G15396<= not I21658;
	G15399<= not I21661;
	G15404<= not I21666;
	G15408<= not G12282;
	G15409<= not G12285;
	G15412<= not I21674;
	G15415<= not I21677;
	G15418<= not I21680;
	G15426<= not I21688;
	G15429<= not I21691;
	G15432<= not I21694;
	G15438<= not G12296;
	G15439<= not G12299;
	G15440<= not G12302;
	G15441<= not G12418;
	G15443<= not I21705;
	G15446<= not I21708;
	G15449<= not I21711;
	G15458<= not G12312;
	G15461<= not I21720;
	G15464<= not I21723;
	G15467<= not I21726;
	G15471<= not I21730;
	G15474<= not G12315;
	G15477<= not I21736;
	G15480<= not I21739;
	G15483<= not I21742;
	G15488<= not I21747;
	G15492<= not G12318;
	G15493<= not G12321;
	G15496<= not I21755;
	G15499<= not I21758;
	G15502<= not I21761;
	G15510<= not I21769;
	G15513<= not I21772;
	G15516<= not I21775;
	G15521<= not I21780;
	G15524<= not G12333;
	G15525<= not G12336;
	G15528<= not I21787;
	G15531<= not I21790;
	G15534<= not I21793;
	G15537<= not I21796;
	G15544<= not G12340;
	G15547<= not I21803;
	G15550<= not I21806;
	G15553<= not I21809;
	G15557<= not I21813;
	G15560<= not G12343;
	G15563<= not I21819;
	G15566<= not I21822;
	G15569<= not I21825;
	G15574<= not I21830;
	G15578<= not G12346;
	G15579<= not G12349;
	G15582<= not I21838;
	G15585<= not I21841;
	G15588<= not I21844;
	G15596<= not I21852;
	G15599<= not I21855;
	G15602<= not G12363;
	G15603<= not G12366;
	G15606<= not I21862;
	G15609<= not I21865;
	G15612<= not I21868;
	G15615<= not I21871;
	G15622<= not G12370;
	G15625<= not I21878;
	G15628<= not I21881;
	G15631<= not I21884;
	G15635<= not I21888;
	G15638<= not G12373;
	G15641<= not I21894;
	G15644<= not I21897;
	G15647<= not I21900;
	G15652<= not I21905;
	G15655<= not I21908;
	G15659<= not G11706;
	G15665<= not G12379;
	G15667<= not I21918;
	G15672<= not I21923;
	G15675<= not I21926;
	G15678<= not G12382;
	G15679<= not G12385;
	G15682<= not I21933;
	G15685<= not I21936;
	G15688<= not I21939;
	G15691<= not I21942;
	G15698<= not G12389;
	G15701<= not I21949;
	G15704<= not I21952;
	G15707<= not I21955;
	G15711<= not I21959;
	G15714<= not I21962;
	G15722<= not G13011;
	G15724<= not G12409;
	G15726<= not I21974;
	G15731<= not I21979;
	G15734<= not I21982;
	G15737<= not G12412;
	G15738<= not G12415;
	G15741<= not I21989;
	G15744<= not I21992;
	G15747<= not I21995;
	G15750<= not I21998;
	G15762<= not G13011;
	G15764<= not G12421;
	G15766<= not I22014;
	G15771<= not I22019;
	G15774<= not I22022;
	G15777<= not I22025;
	G15790<= not G13011;
	G15792<= not G12426;
	G15794<= not I22044;
	G15800<= not G12909;
	G15813<= not G13011;
	G15859<= not G13378;
	G15876<= not I22120;
	G15880<= not G11624;
	G15890<= not G11600;
	G15904<= not G11644;
	G15913<= not G11647;
	G15923<= not G11630;
	G15933<= not G11663;
	G15942<= not G11666;
	G15952<= not G11653;
	G15962<= not G11675;
	G15971<= not G11678;
	G15981<= not G11687;
	G15989<= not I22163;
	G15991<= not G12548;
	G15994<= not G12555;
	G15997<= not G12561;
	G16001<= not G12601;
	G16002<= not G12604;
	G16005<= not G12608;
	G16007<= not G12647;
	G16011<= not G12651;
	G16012<= not G12654;
	G16013<= not G12692;
	G16014<= not G12695;
	G16023<= not G12699;
	G16024<= not G12702;
	G16025<= not G12705;
	G16026<= not G12708;
	G16027<= not G12744;
	G16034<= not G12749;
	G16035<= not G12752;
	G16039<= not G12756;
	G16040<= not G12759;
	G16041<= not G12762;
	G16042<= not G12765;
	G16043<= not G12769;
	G16044<= not G12772;
	G16054<= not G12783;
	G16055<= not G12786;
	G16056<= not G12791;
	G16057<= not G12794;
	G16061<= not G12798;
	G16062<= not G12801;
	G16063<= not G12804;
	G16064<= not G12808;
	G16065<= not G12811;
	G16075<= not G11861;
	G16088<= not G12816;
	G16090<= not G12822;
	G16091<= not G12825;
	G16092<= not G12830;
	G16093<= not G12833;
	G16097<= not G12837;
	G16098<= not G12840;
	G16099<= not G12844;
	G16113<= not G11903;
	G16126<= not G12854;
	G16128<= not G12860;
	G16129<= not G12863;
	G16130<= not G12868;
	G16131<= not G12871;
	G16142<= not G13057;
	G16154<= not G12194;
	G16164<= not G11953;
	G16177<= not G12895;
	G16179<= not G12901;
	G16180<= not G12904;
	G16189<= not G13043;
	G16201<= not G13073;
	G16213<= not G12249;
	G16223<= not G12006;
	G16236<= not G12935;
	G16243<= not G13033;
	G16254<= not G13060;
	G16266<= not G13092;
	G16278<= not G12292;
	G16287<= not G12962;
	G16293<= not G13025;
	G16297<= not I22382;
	G16302<= not G13046;
	G16313<= not G13076;
	G16325<= not G13107;
	G16337<= not G12328;
	G16351<= not G13036;
	G16355<= not I22414;
	G16360<= not G13063;
	G16371<= not G13095;
	G16395<= not G13049;
	G16399<= not I22444;
	G16404<= not G13079;
	G16433<= not G13066;
	G16437<= not I22475;
	G16466<= not G12017;
	G16467<= not I22503;
	G16468<= not I22506;
	G16469<= not I22509;
	G16470<= not I22512;
	G16471<= not I22515;
	G16472<= not I22518;
	G16473<= not I22521;
	G16474<= not I22524;
	G16475<= not I22527;
	G16476<= not I22530;
	G16477<= not I22533;
	G16478<= not I22536;
	G16479<= not I22539;
	G16480<= not I22542;
	G16481<= not I22545;
	G16482<= not I22548;
	G16483<= not I22551;
	G16484<= not I22554;
	G16485<= not I22557;
	G16486<= not I22560;
	G16487<= not I22563;
	G16488<= not I22566;
	G16489<= not I22569;
	G16490<= not I22572;
	G16491<= not I22575;
	G16492<= not I22578;
	G16493<= not I22581;
	G16494<= not I22584;
	G16495<= not I22587;
	G16496<= not I22590;
	G16497<= not I22593;
	G16501<= not G14158;
	G16506<= not I22599;
	G16507<= not G14186;
	G16514<= not I22604;
	G16515<= not G14244;
	G16523<= not G14273;
	G16528<= not I22611;
	G16529<= not G14301;
	G16540<= not I22618;
	G16543<= not G14347;
	G16546<= not G14366;
	G16554<= not G14395;
	G16559<= not I22626;
	G16560<= not G14423;
	G16572<= not I22640;
	G16575<= not G14459;
	G16578<= not G14478;
	G16586<= not G14507;
	G16596<= not I22651;
	G16599<= not G14546;
	G16602<= not G14565;
	G16608<= not I22657;
	G16616<= not I22663;
	G16619<= not G14601;
	G16622<= not I22667;
	G16626<= not I22671;
	G16633<= not I22676;
	G16636<= not I22679;
	G16640<= not I22683;
	G16644<= not I22687;
	G16647<= not I22690;
	G16651<= not I22694;
	G16656<= not I22699;
	G16659<= not I22702;
	G16665<= not G14776;
	G16673<= not I22715;
	G16676<= not I22718;
	G16682<= not G14797;
	G16686<= not G14811;
	G16694<= not I22726;
	G16697<= not G14837;
	G16702<= not I22730;
	G16708<= not G14849;
	G16712<= not G14863;
	G16719<= not I22737;
	G16722<= not G14895;
	G16725<= not I22741;
	G16728<= not G14910;
	G16733<= not I22745;
	G16739<= not G14922;
	G16743<= not G14936;
	G16749<= not G15782;
	G16758<= not I22752;
	G16761<= not I22755;
	G16764<= not G14976;
	G16767<= not I22759;
	G16770<= not G14991;
	G16775<= not I22763;
	G16781<= not G15003;
	G16785<= not I22768;
	G16788<= not I22771;
	G16791<= not G15065;
	G16794<= not I22775;
	G16797<= not G15080;
	G16804<= not G15803;
	G16809<= not G15842;
	G16813<= not I22783;
	G16814<= not I22786;
	G16817<= not I22789;
	G16820<= not G15161;
	G16825<= not G15855;
	G16830<= not I22797;
	G16831<= not I22800;
	G16832<= not I22803;
	G16836<= not G15818;
	G16840<= not G15878;
	G16842<= not I22810;
	G16843<= not I22813;
	G16846<= not G15903;
	G16848<= not I22820;
	G16849<= not I22823;
	G16852<= not I22828;
	G16858<= not I22836;
	G16862<= not I22842;
	G16863<= not I22845;
	G16867<= not G13589;
	G16877<= not I22852;
	G16878<= not I22855;
	G16881<= not I22860;
	G16884<= not G13589;
	G16895<= not G13589;
	G16905<= not I22866;
	G16906<= not I22869;
	G16910<= not I22875;
	G16913<= not G13589;
	G16924<= not G13589;
	G16934<= not I22881;
	G16940<= not I22893;
	G16943<= not G13589;
	G16954<= not G13589;
	G16971<= not I22912;
	G16974<= not G13589;
	G17029<= not G14685;
	G17057<= not G13519;
	G17063<= not G14719;
	G17092<= not G13530;
	G17098<= not G14747;
	G17130<= not G13541;
	G17136<= not G14768;
	G17157<= not G13552;
	G17189<= not I23253;
	G17200<= not I23274;
	G17203<= not G13568;
	G17207<= not I23287;
	G17208<= not G13576;
	G17212<= not I23292;
	G17214<= not G13585;
	G17217<= not G13605;
	G17227<= not I23309;
	G17230<= not I23314;
	G17233<= not I23317;
	G17237<= not I23323;
	G17240<= not I23326;
	G17243<= not I23329;
	G17249<= not I23335;
	G17252<= not I23338;
	G17255<= not I23341;
	G17258<= not G16053;
	G17259<= not I23345;
	G17262<= not I23348;
	G17265<= not I23351;
	G17272<= not I23358;
	G17275<= not I23361;
	G17278<= not I23364;
	G17281<= not G16081;
	G17282<= not I23368;
	G17285<= not I23371;
	G17288<= not I23374;
	G17291<= not I23377;
	G17294<= not I23380;
	G17297<= not I23383;
	G17300<= not I23386;
	G17304<= not I23392;
	G17307<= not I23395;
	G17310<= not I23398;
	G17313<= not G16109;
	G17314<= not G16110;
	G17315<= not I23403;
	G17318<= not I23406;
	G17321<= not I23409;
	G17324<= not I23412;
	G17327<= not I23415;
	G17330<= not I23418;
	G17333<= not I23421;
	G17336<= not I23424;
	G17342<= not I23430;
	G17345<= not I23433;
	G17348<= not I23436;
	G17351<= not G16152;
	G17354<= not I23442;
	G17357<= not I23445;
	G17360<= not I23448;
	G17363<= not I23451;
	G17366<= not I23454;
	G17369<= not I23457;
	G17372<= not I23460;
	G17375<= not I23463;
	G17378<= not I23466;
	G17384<= not I23472;
	G17387<= not I23475;
	G17390<= not I23478;
	G17394<= not G16197;
	G17399<= not I23487;
	G17402<= not I23490;
	G17405<= not I23493;
	G17410<= not I23498;
	G17413<= not I23501;
	G17416<= not I23504;
	G17419<= not I23507;
	G17422<= not I23510;
	G17425<= not I23513;
	G17430<= not I23518;
	G17433<= not I23521;
	G17436<= not I23524;
	G17439<= not I23527;
	G17442<= not I23530;
	G17445<= not G16250;
	G17451<= not I23539;
	G17454<= not I23542;
	G17457<= not I23545;
	G17465<= not I23553;
	G17468<= not I23556;
	G17471<= not I23559;
	G17476<= not I23564;
	G17479<= not I23567;
	G17482<= not I23570;
	G17487<= not I23575;
	G17490<= not I23578;
	G17493<= not I23581;
	G17496<= not I23584;
	G17499<= not G16292;
	G17500<= not I23588;
	G17503<= not I23591;
	G17511<= not I23599;
	G17514<= not I23602;
	G17517<= not I23605;
	G17520<= not I23608;
	G17523<= not I23611;
	G17531<= not I23619;
	G17534<= not I23622;
	G17537<= not I23625;
	G17545<= not I23633;
	G17548<= not I23636;
	G17551<= not I23639;
	G17557<= not I23645;
	G17560<= not I23648;
	G17563<= not I23651;
	G17566<= not G16346;
	G17567<= not I23655;
	G17570<= not I23658;
	G17573<= not I23661;
	G17579<= not I23667;
	G17582<= not I23670;
	G17585<= not I23673;
	G17588<= not I23676;
	G17591<= not I23679;
	G17594<= not I23682;
	G17601<= not I23689;
	G17604<= not I23692;
	G17607<= not I23695;
	G17610<= not I23698;
	G17613<= not I23701;
	G17621<= not I23709;
	G17624<= not I23712;
	G17627<= not I23715;
	G17637<= not I23725;
	G17640<= not G13873;
	G17645<= not I23729;
	G17648<= not G16384;
	G17649<= not I23733;
	G17655<= not I23739;
	G17658<= not I23742;
	G17661<= not I23745;
	G17664<= not I23748;
	G17667<= not I23751;
	G17670<= not I23754;
	G17676<= not I23760;
	G17679<= not I23763;
	G17682<= not I23766;
	G17685<= not I23769;
	G17688<= not I23772;
	G17691<= not I23775;
	G17698<= not I23782;
	G17701<= not I23785;
	G17704<= not I23788;
	G17707<= not I23791;
	G17710<= not I23794;
	G17720<= not G15853;
	G17724<= not G13886;
	G17738<= not I23817;
	G17741<= not G13895;
	G17746<= not I23821;
	G17749<= not I23824;
	G17755<= not I23830;
	G17758<= not I23833;
	G17761<= not I23836;
	G17764<= not I23839;
	G17767<= not I23842;
	G17770<= not I23845;
	G17776<= not I23851;
	G17779<= not I23854;
	G17782<= not I23857;
	G17785<= not I23860;
	G17788<= not I23863;
	G17791<= not I23866;
	G17799<= not I23874;
	G17802<= not G13907;
	G17815<= not I23888;
	G17825<= not G13927;
	G17839<= not I23904;
	G17842<= not G13936;
	G17847<= not I23908;
	G17850<= not I23911;
	G17856<= not I23917;
	G17859<= not I23920;
	G17862<= not I23923;
	G17865<= not I23926;
	G17868<= not I23929;
	G17871<= not I23932;
	G17878<= not G15830;
	G17882<= not G13946;
	G17892<= not G13954;
	G17893<= not G14165;
	G17903<= not I23954;
	G17914<= not G13963;
	G17927<= not I23976;
	G17937<= not G13983;
	G17951<= not I23992;
	G17954<= not G13992;
	G17959<= not I23996;
	G17962<= not I23999;
	G17969<= not G15841;
	G17974<= not G14001;
	G17984<= not G14008;
	G17988<= not G14685;
	G17991<= not G14450;
	G17993<= not G14016;
	G18003<= not G14024;
	G18004<= not G14280;
	G18014<= not I24049;
	G18025<= not G14033;
	G18038<= not I24071;
	G18048<= not G14053;
	G18063<= not G15660;
	G18070<= not G15854;
	G18074<= not G14062;
	G18084<= not G14068;
	G18089<= not G14355;
	G18091<= not G14092;
	G18101<= not G14099;
	G18105<= not G14719;
	G18108<= not G14537;
	G18110<= not G14107;
	G18120<= not G14115;
	G18121<= not G14402;
	G18131<= not I24144;
	G18142<= not G14124;
	G18155<= not I24166;
	G18166<= not I24171;
	G18170<= not G15877;
	G18174<= not G14148;
	G18179<= not G14153;
	G18188<= not G14252;
	G18190<= not G14177;
	G18200<= not G14183;
	G18205<= not G14467;
	G18207<= not G14207;
	G18217<= not G14214;
	G18221<= not G14747;
	G18224<= not G14592;
	G18226<= not G14222;
	G18236<= not G14230;
	G18237<= not G14514;
	G18247<= not I24247;
	G18258<= not I24258;
	G18261<= not G15719;
	G18265<= not G14238;
	G18275<= not G14171;
	G18278<= not I24285;
	G18281<= not G14263;
	G18286<= not G14268;
	G18295<= not G14374;
	G18297<= not G14292;
	G18307<= not G14298;
	G18312<= not G14554;
	G18314<= not G14322;
	G18324<= not G14329;
	G18328<= not G14768;
	G18331<= not G14626;
	G18334<= not I24346;
	G18337<= not G15757;
	G18341<= not G14342;
	G18351<= not G13741;
	G18353<= not G13918;
	G18355<= not I24368;
	G18358<= not G14360;
	G18368<= not G14286;
	G18371<= not I24394;
	G18374<= not G14385;
	G18379<= not G14390;
	G18388<= not G14486;
	G18390<= not G14414;
	G18400<= not G14420;
	G18405<= not G14609;
	G18407<= not G15959;
	G18414<= not G15718;
	G18415<= not G15783;
	G18429<= not G14831;
	G18432<= not I24459;
	G18435<= not G14359;
	G18436<= not G14454;
	G18446<= not G13741;
	G18448<= not G13974;
	G18450<= not I24481;
	G18453<= not G14472;
	G18463<= not G14408;
	G18466<= not I24507;
	G18469<= not G14497;
	G18474<= not G14502;
	G18483<= not G14573;
	G18485<= not G15756;
	G18486<= not G15804;
	G18490<= not G13565;
	G18502<= not G14904;
	G18505<= not I24560;
	G18508<= not G14471;
	G18509<= not G14541;
	G18519<= not G13741;
	G18521<= not G14044;
	G18523<= not I24582;
	G18526<= not G14559;
	G18536<= not G14520;
	G18539<= not I24608;
	G18543<= not G15819;
	G18552<= not G16154;
	G18554<= not G13573;
	G18566<= not G14985;
	G18569<= not I24662;
	G18572<= not G14558;
	G18573<= not G14596;
	G18583<= not G13741;
	G18585<= not G14135;
	G18587<= not I24684;
	G18593<= not G15831;
	G18602<= not G16213;
	G18604<= not G13582;
	G18616<= not G15074;
	G18619<= not I24732;
	G18622<= not G14613;
	G18634<= not G16278;
	G18636<= not G13602;
	G18643<= not G16337;
	G18646<= not G16341;
	G18656<= not G14776;
	G18670<= not G14797;
	G18679<= not G14811;
	G18691<= not G14885;
	G18692<= not G14837;
	G18699<= not G14849;
	G18708<= not G14863;
	G18720<= not G14895;
	G18725<= not G13865;
	G18727<= not G14966;
	G18728<= not G14910;
	G18735<= not G14922;
	G18744<= not G14936;
	G18756<= not G14960;
	G18757<= not G14963;
	G18758<= not G14976;
	G18764<= not G15055;
	G18765<= not G14991;
	G18772<= not G15003;
	G18783<= not G15034;
	G18784<= not G15037;
	G18785<= not G15040;
	G18786<= not G15043;
	G18787<= not G15049;
	G18788<= not G15052;
	G18789<= not G15065;
	G18795<= not G15151;
	G18796<= not G15080;
	G18805<= not G15106;
	G18806<= not G15109;
	G18807<= not G15112;
	G18808<= not G15115;
	G18809<= not G15130;
	G18810<= not G15133;
	G18811<= not G15136;
	G18812<= not G15139;
	G18813<= not G15145;
	G18814<= not G15148;
	G18815<= not G15161;
	G18822<= not G15179;
	G18823<= not G15182;
	G18824<= not G15185;
	G18825<= not G15198;
	G18826<= not G15201;
	G18827<= not G15204;
	G18828<= not G15207;
	G18829<= not G15222;
	G18830<= not G15225;
	G18831<= not G15228;
	G18832<= not G15231;
	G18833<= not G15237;
	G18834<= not G15240;
	G18838<= not G15248;
	G18839<= not G15251;
	G18840<= not G15254;
	G18841<= not G15265;
	G18842<= not G15268;
	G18843<= not G15271;
	G18844<= not G15284;
	G18845<= not G15287;
	G18846<= not G15290;
	G18847<= not G15293;
	G18848<= not G15308;
	G18849<= not G15311;
	G18850<= not G15314;
	G18851<= not G15317;
	G18853<= not G15326;
	G18854<= not G15329;
	G18855<= not G15332;
	G18856<= not G15340;
	G18857<= not G15343;
	G18858<= not G15346;
	G18859<= not G15357;
	G18860<= not G15360;
	G18861<= not G15363;
	G18862<= not G15376;
	G18863<= not G15379;
	G18864<= not G15382;
	G18865<= not G15385;
	G18869<= not I24894;
	G18870<= not G15393;
	G18871<= not G15396;
	G18872<= not G15399;
	G18873<= not G15404;
	G18874<= not G15412;
	G18875<= not G15415;
	G18876<= not G15418;
	G18877<= not G15426;
	G18878<= not G15429;
	G18879<= not G15432;
	G18880<= not G15443;
	G18881<= not G15446;
	G18882<= not G15449;
	G18884<= not G13469;
	G18886<= not I24913;
	G18890<= not I24916;
	G18891<= not G15461;
	G18892<= not G15464;
	G18893<= not G15467;
	G18894<= not G15471;
	G18895<= not I24923;
	G18896<= not G15477;
	G18897<= not G15480;
	G18898<= not G15483;
	G18899<= not G15488;
	G18900<= not G15496;
	G18901<= not G15499;
	G18902<= not G15502;
	G18903<= not G15510;
	G18904<= not G15513;
	G18905<= not G15516;
	G18908<= not G15521;
	G18909<= not G15528;
	G18910<= not G15531;
	G18911<= not G15534;
	G18912<= not G15537;
	G18913<= not I24943;
	G18914<= not G15547;
	G18915<= not G15550;
	G18916<= not G15553;
	G18917<= not G15557;
	G18918<= not I24950;
	G18919<= not G15563;
	G18920<= not G15566;
	G18921<= not G15569;
	G18922<= not G15574;
	G18923<= not G15582;
	G18924<= not G15585;
	G18925<= not G15588;
	G18926<= not G15596;
	G18927<= not G15599;
	G18928<= not G15606;
	G18929<= not G15609;
	G18930<= not G15612;
	G18931<= not G15615;
	G18932<= not I24966;
	G18933<= not G15625;
	G18934<= not G15628;
	G18935<= not G15631;
	G18936<= not G15635;
	G18937<= not I24973;
	G18938<= not G15641;
	G18939<= not G15644;
	G18940<= not G15647;
	G18941<= not G15652;
	G18943<= not G15655;
	G18944<= not I24982;
	G18945<= not G15667;
	G18946<= not G15672;
	G18947<= not G15675;
	G18948<= not G15682;
	G18949<= not G15685;
	G18950<= not G15688;
	G18951<= not G15691;
	G18952<= not I24992;
	G18953<= not G15701;
	G18954<= not G15704;
	G18955<= not G15707;
	G18956<= not G15711;
	G18958<= not G15714;
	G18959<= not I25001;
	G18960<= not I25004;
	G18961<= not G15726;
	G18962<= not G15731;
	G18963<= not G15734;
	G18964<= not G15741;
	G18965<= not G15744;
	G18966<= not G15747;
	G18967<= not G15750;
	G18969<= not I25015;
	G18970<= not I25018;
	G18971<= not I25021;
	G18972<= not G15766;
	G18973<= not G15771;
	G18974<= not G15774;
	G18976<= not G15777;
	G18981<= not I25037;
	G18983<= not I25041;
	G18984<= not I25044;
	G18985<= not I25047;
	G18986<= not I25050;
	G18987<= not G15794;
	G18988<= not I25054;
	G18989<= not I25057;
	G18991<= not I25061;
	G18992<= not I25064;
	G18993<= not I25067;
	G18995<= not I25071;
	G18996<= not I25074;
	G18998<= not I25078;
	G18999<= not I25081;
	G19000<= not I25084;
	G19001<= not G14071;
	G19008<= not I25089;
	G19009<= not I25092;
	G19011<= not I25096;
	G19012<= not I25099;
	G19013<= not I25102;
	G19014<= not I25105;
	G19015<= not I25108;
	G19016<= not I25111;
	G19017<= not I25114;
	G19018<= not I25117;
	G19019<= not I25120;
	G19020<= not I25123;
	G19021<= not I25126;
	G19022<= not I25129;
	G19023<= not I25132;
	G19024<= not I25135;
	G19025<= not I25138;
	G19026<= not I25141;
	G19027<= not I25144;
	G19028<= not I25147;
	G19029<= not I25150;
	G19030<= not I25153;
	G19031<= not I25156;
	G19032<= not I25159;
	G19033<= not I25162;
	G19034<= not I25165;
	G19035<= not I25168;
	G19036<= not I25171;
	G19037<= not I25174;
	G19038<= not I25177;
	G19039<= not I25180;
	G19040<= not I25183;
	G19041<= not I25186;
	G19042<= not I25189;
	G19043<= not I25192;
	G19044<= not I25195;
	G19045<= not I25198;
	G19046<= not I25201;
	G19047<= not I25204;
	G19048<= not I25207;
	G19049<= not I25210;
	G19050<= not I25213;
	G19051<= not I25216;
	G19052<= not I25219;
	G19053<= not I25222;
	G19054<= not I25225;
	G19055<= not I25228;
	G19056<= not I25231;
	G19057<= not I25234;
	G19058<= not I25237;
	G19059<= not I25240;
	G19060<= not I25243;
	G19061<= not I25246;
	G19062<= not I25249;
	G19064<= not I25253;
	G19070<= not G18583;
	G19075<= not I25258;
	G19078<= not G18619;
	G19081<= not I25264;
	G19091<= not I25272;
	G19096<= not G18980;
	G19098<= not I25283;
	G19105<= not I25294;
	G19110<= not I25303;
	G19113<= not I25308;
	G19118<= not I25315;
	G19125<= not I25320;
	G19132<= not I25325;
	G19145<= not I25334;
	G19147<= not I25338;
	G19151<= not I25344;
	G19156<= not I25351;
	G19158<= not I25355;
	G19159<= not I25358;
	G19164<= not I25365;
	G19168<= not I25371;
	G19169<= not I25374;
	G19170<= not I25377;
	G19174<= not I25383;
	G19175<= not I25386;
	G19176<= not I25389;
	G19180<= not I25395;
	G19182<= not I25399;
	G19183<= not I25402;
	G19185<= not I25406;
	G19189<= not I25412;
	G19190<= not I25415;
	G19196<= not I25423;
	G19197<= not I25426;
	G19198<= not I25429;
	G19199<= not I25432;
	G19207<= not I25442;
	G19208<= not I25445;
	G19217<= not I25456;
	G19218<= not I25459;
	G19220<= not I25463;
	G19229<= not I25474;
	G19237<= not I25486;
	G19238<= not I25489;
	G19239<= not I25492;
	G19247<= not I25506;
	G19249<= not I25510;
	G19251<= not G16540;
	G19258<= not I25525;
	G19259<= not I25528;
	G19265<= not G16572;
	G19270<= not I25557;
	G19272<= not I25567;
	G19280<= not G16596;
	G19287<= not G16608;
	G19291<= not I25612;
	G19299<= not G16616;
	G19301<= not G16622;
	G19302<= not G17025;
	G19305<= not G16626;
	G19309<= not I25660;
	G19319<= not G16633;
	G19322<= not G16636;
	G19323<= not G17059;
	G19326<= not G16640;
	G19330<= not I25717;
	G19335<= not I25728;
	G19346<= not G16644;
	G19349<= not G16647;
	G19350<= not G17094;
	G19353<= not G16651;
	G19358<= not I25768;
	G19369<= not I25778;
	G19380<= not G16656;
	G19383<= not G16659;
	G19384<= not G17132;
	G19387<= not G16567;
	G19388<= not G17139;
	G19390<= not I25816;
	G19401<= not I25826;
	G19412<= not G16673;
	G19415<= not G16676;
	G19417<= not G16591;
	G19418<= not G17162;
	G19420<= not I25862;
	G19431<= not I25872;
	G19441<= not G17213;
	G19444<= not G17985;
	G19448<= not G16694;
	G19452<= not G16702;
	G19454<= not G16611;
	G19455<= not G17177;
	G19457<= not I25904;
	G19467<= not G16719;
	G19468<= not G17216;
	G19471<= not G18102;
	G19475<= not G16725;
	G19479<= not G16733;
	G19481<= not G16629;
	G19482<= not G17194;
	G19483<= not G16758;
	G19484<= not G16867;
	G19490<= not G16761;
	G19491<= not G17219;
	G19494<= not G18218;
	G19498<= not G16767;
	G19502<= not G16775;
	G19504<= not G16785;
	G19505<= not G16895;
	G19511<= not G16788;
	G19512<= not G17221;
	G19515<= not G18325;
	G19519<= not G16794;
	G19523<= not G16814;
	G19524<= not G16924;
	G19530<= not G16817;
	G19533<= not G16832;
	G19534<= not G16954;
	G19543<= not I25966;
	G19546<= not I25971;
	G19550<= not I25977;
	G19556<= not I25985;
	G19563<= not I25994;
	G19573<= not I26006;
	G19577<= not G16881;
	G19578<= not G16884;
	G19595<= not I26025;
	G19596<= not I26028;
	G19607<= not G16910;
	G19608<= not G16913;
	G19622<= not I26051;
	G19640<= not G16940;
	G19641<= not G16943;
	G19652<= not I26078;
	G19657<= not I26085;
	G19680<= not G16971;
	G19681<= not G16974;
	G19689<= not I26112;
	G19690<= not I26115;
	G19696<= not I26123;
	G19705<= not I26134;
	G19725<= not I26154;
	G19740<= not I26171;
	G19749<= not I26182;
	G19762<= not I26195;
	G19763<= not I26198;
	G19783<= not I26220;
	G19792<= not I26231;
	G19798<= not I26237;
	G19825<= not I26266;
	G19830<= not G18886;
	G19838<= not I26276;
	G19890<= not I26334;
	G19893<= not I26337;
	G19894<= not I26340;
	G19915<= not I26365;
	G19918<= not G18646;
	G19919<= not I26369;
	G19933<= not G18548;
	G19934<= not I26388;
	G19945<= not I26401;
	G19948<= not G17896;
	G19950<= not G18598;
	G19951<= not I26407;
	G19957<= not I26413;
	G19972<= not I26420;
	G19975<= not G18007;
	G19977<= not G18630;
	G19978<= not I26426;
	G19987<= not I26437;
	G20002<= not I26444;
	G20005<= not G18124;
	G20007<= not G18639;
	G20016<= not I26458;
	G20025<= not I26469;
	G20040<= not I26476;
	G20043<= not G18240;
	G20045<= not I26481;
	G20058<= not I26494;
	G20067<= not I26505;
	G20082<= not I26512;
	G20083<= not G17968;
	G20099<= not I26535;
	G20105<= not I26545;
	G20124<= not I26574;
	G20127<= not G18623;
	G20140<= not G16830;
	G20163<= not G17973;
	G20164<= not I26612;
	G20178<= not G16842;
	G20193<= not G18691;
	G20198<= not I26642;
	G20212<= not G16848;
	G20223<= not G18727;
	G20228<= not I26664;
	G20242<= not G16852;
	G20250<= not G18764;
	G20255<= not I26679;
	G20269<= not G17230;
	G20273<= not G18795;
	G20278<= not G17237;
	G20279<= not G17240;
	G20281<= not G17243;
	G20286<= not G17249;
	G20287<= not G17252;
	G20288<= not G17255;
	G20289<= not G17259;
	G20290<= not G17262;
	G20292<= not G17265;
	G20295<= not I26714;
	G20296<= not G17272;
	G20297<= not G17275;
	G20298<= not G17278;
	G20302<= not G17282;
	G20303<= not G17285;
	G20304<= not G17288;
	G20305<= not G17291;
	G20306<= not G17294;
	G20308<= not G17297;
	G20311<= not G17304;
	G20312<= not G17307;
	G20313<= not G17310;
	G20315<= not G17315;
	G20316<= not G17318;
	G20317<= not G17321;
	G20321<= not G17324;
	G20322<= not G17327;
	G20323<= not G17330;
	G20324<= not G17333;
	G20325<= not G17336;
	G20327<= not G17342;
	G20328<= not G17345;
	G20329<= not G17348;
	G20330<= not G17354;
	G20331<= not G17357;
	G20332<= not G17360;
	G20334<= not G17363;
	G20335<= not G17366;
	G20336<= not G17369;
	G20340<= not G17372;
	G20341<= not G17375;
	G20342<= not G17378;
	G20344<= not G17384;
	G20345<= not G17387;
	G20346<= not G17390;
	G20347<= not G17399;
	G20348<= not G17402;
	G20349<= not G17405;
	G20350<= not G17410;
	G20351<= not G17413;
	G20352<= not G17416;
	G20354<= not G17419;
	G20355<= not G17422;
	G20356<= not G17425;
	G20360<= not I26777;
	G20361<= not G17430;
	G20362<= not G17433;
	G20363<= not G17436;
	G20364<= not G17439;
	G20365<= not G17442;
	G20366<= not G17451;
	G20367<= not G17454;
	G20368<= not G17457;
	G20369<= not G17465;
	G20370<= not G17468;
	G20371<= not G17471;
	G20372<= not G17476;
	G20373<= not G17479;
	G20374<= not G17482;
	G20377<= not I26796;
	G20378<= not G17487;
	G20379<= not G17490;
	G20380<= not G17493;
	G20381<= not G17496;
	G20382<= not G17500;
	G20383<= not G17503;
	G20384<= not G17511;
	G20385<= not G17514;
	G20386<= not G17517;
	G20387<= not G17520;
	G20388<= not G17523;
	G20389<= not G17531;
	G20390<= not G17534;
	G20391<= not G17537;
	G20392<= not G17545;
	G20393<= not G17548;
	G20394<= not G17551;
	G20395<= not I26816;
	G20396<= not I26819;
	G20397<= not G17557;
	G20398<= not G17560;
	G20399<= not G17563;
	G20400<= not G17567;
	G20401<= not G17570;
	G20402<= not G17573;
	G20403<= not G17579;
	G20404<= not G17582;
	G20405<= not G17585;
	G20406<= not G17588;
	G20407<= not G17591;
	G20408<= not G17594;
	G20409<= not G17601;
	G20410<= not G17604;
	G20411<= not G17607;
	G20412<= not G17610;
	G20413<= not G17613;
	G20414<= not G17621;
	G20415<= not G17624;
	G20416<= not G17627;
	G20418<= not I26843;
	G20419<= not I26846;
	G20420<= not G17637;
	G20421<= not G17649;
	G20422<= not G17655;
	G20423<= not G17658;
	G20424<= not G17661;
	G20425<= not G17664;
	G20426<= not G17667;
	G20427<= not G17670;
	G20428<= not G17676;
	G20429<= not G17679;
	G20430<= not G17682;
	G20431<= not G17685;
	G20432<= not G17688;
	G20433<= not G17691;
	G20434<= not G17698;
	G20435<= not G17701;
	G20436<= not G17704;
	G20437<= not G17707;
	G20438<= not G17710;
	G20439<= not I26868;
	G20440<= not I26871;
	G20441<= not I26874;
	G20442<= not G17738;
	G20443<= not G17749;
	G20444<= not G17755;
	G20445<= not G17758;
	G20446<= not G17761;
	G20447<= not G17764;
	G20448<= not G17767;
	G20449<= not G17770;
	G20450<= not G17776;
	G20451<= not G17779;
	G20452<= not G17782;
	G20453<= not G17785;
	G20454<= not G17788;
	G20455<= not G17791;
	G20456<= not G17799;
	G20457<= not I26892;
	G20458<= not I26895;
	G20459<= not I26898;
	G20461<= not G17839;
	G20462<= not G17850;
	G20463<= not G17856;
	G20464<= not G17859;
	G20465<= not G17862;
	G20466<= not G17865;
	G20467<= not G17868;
	G20468<= not G17871;
	G20469<= not I26910;
	G20470<= not I26913;
	G20471<= not I26916;
	G20476<= not G17951;
	G20477<= not G17962;
	G20478<= not I26923;
	G20479<= not I26926;
	G20484<= not I26931;
	G20485<= not I26934;
	G20490<= not G18166;
	G20491<= not I26940;
	G20496<= not G18258;
	G20498<= not I26947;
	G20500<= not G18278;
	G20501<= not G18334;
	G20504<= not G18355;
	G20505<= not G18371;
	G20507<= not G18351;
	G20513<= not I26960;
	G20516<= not G18432;
	G20517<= not G18450;
	G20518<= not G18466;
	G20519<= not I26966;
	G20526<= not G18446;
	G20531<= not I26972;
	G20534<= not G18505;
	G20535<= not G18523;
	G20536<= not G18539;
	G20539<= not I26980;
	G20545<= not G18519;
	G20550<= not I26985;
	G20553<= not G18569;
	G20554<= not G18587;
	G20555<= not I26990;
	G20556<= not I26993;
	G20557<= not I26996;
	G20558<= not I26999;
	G20559<= not I27002;
	G20560<= not I27005;
	G20561<= not I27008;
	G20562<= not I27011;
	G20563<= not I27014;
	G20564<= not I27017;
	G20565<= not I27020;
	G20566<= not I27023;
	G20567<= not I27026;
	G20568<= not I27029;
	G20569<= not I27032;
	G20570<= not I27035;
	G20571<= not I27038;
	G20572<= not I27041;
	G20573<= not I27044;
	G20574<= not I27047;
	G20575<= not I27050;
	G20576<= not I27053;
	G20577<= not I27056;
	G20578<= not I27059;
	G20579<= not I27062;
	G20580<= not I27065;
	G20581<= not I27068;
	G20582<= not I27071;
	G20583<= not I27074;
	G20584<= not I27077;
	G20585<= not I27080;
	G20586<= not I27083;
	G20587<= not I27086;
	G20588<= not I27089;
	G20589<= not I27092;
	G20590<= not I27095;
	G20591<= not I27098;
	G20592<= not I27101;
	G20593<= not I27104;
	G20594<= not I27107;
	G20595<= not I27110;
	G20596<= not I27113;
	G20597<= not I27116;
	G20598<= not I27119;
	G20599<= not I27122;
	G20600<= not I27125;
	G20601<= not I27128;
	G20602<= not I27131;
	G20603<= not I27134;
	G20604<= not I27137;
	G20605<= not I27140;
	G20606<= not I27143;
	G20607<= not I27146;
	G20608<= not I27149;
	G20609<= not I27152;
	G20610<= not I27155;
	G20611<= not I27158;
	G20612<= not I27161;
	G20613<= not I27164;
	G20614<= not I27167;
	G20615<= not I27170;
	G20616<= not I27173;
	G20617<= not I27176;
	G20618<= not I27179;
	G20619<= not I27182;
	G20620<= not I27185;
	G20621<= not I27188;
	G20622<= not I27191;
	G20623<= not I27194;
	G20624<= not I27197;
	G20625<= not I27200;
	G20626<= not I27203;
	G20627<= not I27206;
	G20628<= not I27209;
	G20629<= not I27212;
	G20630<= not I27215;
	G20631<= not I27218;
	G20632<= not I27221;
	G20634<= not I27225;
	G20637<= not I27228;
	G20641<= not I27232;
	G20644<= not I27235;
	G20649<= not I27240;
	G20652<= not I27243;
	G20655<= not I27246;
	G20659<= not I27250;
	G20662<= not I27253;
	G20666<= not I27257;
	G20669<= not I27260;
	G20673<= not I27264;
	G20676<= not I27267;
	G20679<= not I27270;
	G20684<= not I27275;
	G20687<= not I27278;
	G20690<= not I27281;
	G20694<= not I27285;
	G20697<= not I27288;
	G20704<= not I27293;
	G20708<= not I27297;
	G20711<= not I27300;
	G20714<= not I27303;
	G20719<= not I27308;
	G20722<= not I27311;
	G20725<= not I27314;
	G20729<= not I27318;
	G20732<= not I27321;
	G20735<= not I27324;
	G20739<= not I27328;
	G20743<= not I27332;
	G20746<= not I27335;
	G20749<= not I27338;
	G20754<= not I27343;
	G20757<= not I27346;
	G20760<= not I27349;
	G20763<= not I27352;
	G20766<= not I27355;
	G20769<= not I27358;
	G20772<= not I27361;
	G20776<= not I27365;
	G20780<= not I27369;
	G20783<= not I27372;
	G20786<= not I27375;
	G20790<= not I27379;
	G20793<= not I27382;
	G20796<= not I27385;
	G20799<= not I27388;
	G20802<= not I27391;
	G20806<= not I27395;
	G20810<= not I27399;
	G20813<= not I27402;
	G20816<= not I27405;
	G20819<= not I27408;
	G20822<= not I27411;
	G20827<= not I27416;
	G20830<= not I27419;
	G20833<= not I27422;
	G20837<= not I27426;
	G20842<= not G19441;
	G20850<= not G19468;
	G20858<= not G19491;
	G20866<= not G19512;
	G20885<= not G19865;
	G20904<= not G19896;
	G20928<= not G19921;
	G20942<= not I27488;
	G20943<= not I27491;
	G20956<= not G19936;
	G20971<= not I27516;
	G20984<= not I27531;
	G20985<= not I27534;
	G20986<= not I27537;
	G20998<= not I27549;
	G21012<= not I27565;
	G21024<= not I27577;
	G21030<= not I27585;
	G21036<= not I27593;
	G21050<= not G20513;
	G21057<= not I27614;
	G21064<= not I27621;
	G21066<= not G20519;
	G21069<= not G20531;
	G21076<= not G20539;
	G21079<= not G20550;
	G21087<= not I27646;
	G21090<= not G19064;
	G21093<= not G19075;
	G21099<= not I27658;
	G21102<= not G19081;
	G21108<= not I27667;
	G21113<= not I27672;
	G21125<= not I27684;
	G21130<= not I27689;
	G21144<= not I27705;
	G21164<= not I27727;
	G21184<= not I27749;
	G21187<= not G19113;
	G21199<= not I27766;
	G21202<= not G19118;
	G21214<= not I27779;
	G21217<= not G19125;
	G21222<= not I27785;
	G21225<= not G19132;
	G21241<= not G19945;
	G21249<= not G19972;
	G21258<= not G20002;
	G21266<= not G20040;
	G21271<= not I27822;
	G21278<= not I27827;
	G21285<= not I27832;
	G21293<= not I27838;
	G21327<= not I27868;
	G21358<= not I27897;
	G21359<= not I27900;
	G21376<= not I27917;
	G21377<= not I27920;
	G21382<= not I27927;
	G21399<= not I27942;
	G21400<= not G19918;
	G21404<= not I27949;
	G21415<= not I27958;
	G21426<= not I27969;
	G21427<= not I27972;
	G21429<= not I27976;
	G21441<= not I27984;
	G21449<= not I27992;
	G21457<= not I28000;
	G21458<= not I28003;
	G21461<= not G19957;
	G21473<= not I28009;
	G21477<= not I28013;
	G21483<= not I28019;
	G21491<= not I28027;
	G21495<= not I28031;
	G21496<= not I28034;
	G21498<= not I28038;
	G21505<= not I28043;
	G21508<= not G19987;
	G21514<= not I28047;
	G21518<= not I28051;
	G21524<= not I28057;
	G21528<= not I28061;
	G21529<= not G19272;
	G21530<= not I28065;
	G21537<= not I28072;
	G21541<= not I28076;
	G21544<= not G20025;
	G21550<= not I28080;
	G21554<= not I28084;
	G21557<= not I28087;
	G21558<= not I28090;
	G21561<= not I28093;
	G21565<= not G19291;
	G21566<= not I28100;
	G21573<= not I28107;
	G21577<= not I28111;
	G21580<= not G20067;
	G21586<= not I28115;
	G21590<= not I28119;
	G21594<= not I28123;
	G21598<= not G19309;
	G21599<= not I28130;
	G21606<= not I28137;
	G21612<= not I28143;
	G21619<= not I28148;
	G21623<= not I28152;
	G21627<= not G19330;
	G21628<= not I28159;
	G21640<= not I28169;
	G21647<= not I28174;
	G21651<= not I28178;
	G21655<= not I28184;
	G21661<= not G19091;
	G21671<= not I28201;
	G21678<= not I28206;
	G21682<= not I28210;
	G21690<= not G19098;
	G21700<= not I28229;
	G21708<= not I28235;
	G21716<= not G19894;
	G21726<= not G19105;
	G21742<= not G19919;
	G21752<= not G19110;
	G21766<= not G19934;
	G21782<= not G19951;
	G21795<= not I28314;
	G21824<= not I28357;
	G21825<= not I28360;
	G21861<= not G19657;
	G21867<= not G19705;
	G21872<= not G19749;
	G21876<= not G19792;
	G21883<= not G19890;
	G21886<= not G19915;
	G21895<= not G19945;
	G21902<= not G19978;
	G21907<= not G19972;
	G21914<= not I28432;
	G21917<= not I28435;
	G21921<= not G20002;
	G21927<= not G20045;
	G21928<= not I28443;
	G21932<= not I28447;
	G21935<= not I28450;
	G21939<= not G20040;
	G21943<= not I28455;
	G21944<= not I28458;
	G21945<= not I28461;
	G21946<= not I28464;
	G21947<= not I28467;
	G21948<= not I28470;
	G21949<= not I28473;
	G21950<= not I28476;
	G21951<= not I28479;
	G21952<= not I28482;
	G21953<= not I28485;
	G21954<= not I28488;
	G21955<= not I28491;
	G21956<= not I28494;
	G21957<= not I28497;
	G21958<= not I28500;
	G21959<= not I28503;
	G21960<= not I28506;
	G21961<= not I28509;
	G21962<= not I28512;
	G21963<= not I28515;
	G21964<= not I28518;
	G21965<= not I28521;
	G21966<= not I28524;
	G21967<= not I28527;
	G21982<= not I28541;
	G21995<= not I28550;
	G22003<= not I28557;
	G22014<= not I28564;
	G22082<= not I28628;
	G22107<= not I28649;
	G22133<= not I28671;
	G22156<= not I28693;
	G22176<= not I28712;
	G22212<= not G21914;
	G22213<= not G21917;
	G22217<= not G21928;
	G22219<= not I28781;
	G22221<= not G21932;
	G22222<= not G21935;
	G22225<= not I28789;
	G22226<= not I28792;
	G22230<= not G20634;
	G22232<= not I28800;
	G22233<= not G20637;
	G22236<= not G20641;
	G22237<= not G20644;
	G22239<= not G20649;
	G22240<= not G20652;
	G22241<= not G20655;
	G22243<= not I28813;
	G22246<= not G20659;
	G22248<= not G20662;
	G22251<= not G20666;
	G22252<= not G20669;
	G22253<= not I28825;
	G22256<= not G20673;
	G22257<= not G20676;
	G22258<= not G20679;
	G22259<= not I28833;
	G22260<= not G20684;
	G22261<= not G20687;
	G22262<= not G20690;
	G22266<= not G20694;
	G22268<= not G20697;
	G22271<= not G20704;
	G22274<= not G20708;
	G22275<= not G20711;
	G22276<= not G20714;
	G22277<= not G20719;
	G22278<= not G20722;
	G22279<= not G20725;
	G22283<= not G20729;
	G22286<= not G20732;
	G22287<= not G20735;
	G22290<= not G20739;
	G22293<= not G20743;
	G22294<= not G20746;
	G22295<= not G20749;
	G22296<= not G20754;
	G22297<= not G20757;
	G22298<= not G20760;
	G22300<= not I28876;
	G22303<= not G20763;
	G22304<= not G20766;
	G22306<= not G20769;
	G22307<= not G20772;
	G22310<= not G20776;
	G22313<= not G20780;
	G22314<= not G20783;
	G22315<= not G20786;
	G22316<= not G21149;
	G22318<= not G20790;
	G22319<= not G21228;
	G22328<= not I28896;
	G22331<= not G20793;
	G22332<= not G20796;
	G22334<= not G20799;
	G22335<= not G20802;
	G22338<= not G20806;
	G22341<= not G21169;
	G22343<= not G20810;
	G22344<= not G21233;
	G22353<= not I28913;
	G22356<= not G20813;
	G22357<= not G20816;
	G22359<= not G20819;
	G22360<= not G20822;
	G22364<= not G21189;
	G22366<= not G20827;
	G22367<= not G21242;
	G22376<= not I28928;
	G22379<= not G20830;
	G22380<= not G20833;
	G22384<= not G21204;
	G22386<= not G20837;
	G22387<= not G21250;
	G22401<= not G21533;
	G22402<= not G21569;
	G22403<= not G21602;
	G22404<= not G21631;
	G22405<= not I28949;
	G22408<= not G20986;
	G22409<= not I28953;
	G22412<= not I28956;
	G22415<= not I28959;
	G22418<= not I28962;
	G22421<= not G21012;
	G22422<= not I28966;
	G22425<= not I28969;
	G22428<= not I28972;
	G22431<= not I28975;
	G22434<= not I28978;
	G22437<= not I28981;
	G22440<= not I28984;
	G22443<= not G21036;
	G22444<= not I28988;
	G22445<= not I28991;
	G22448<= not I28994;
	G22451<= not I28997;
	G22455<= not I29001;
	G22458<= not I29004;
	G22461<= not I29007;
	G22464<= not I29010;
	G22467<= not I29013;
	G22470<= not I29016;
	G22473<= not I29019;
	G22476<= not G21057;
	G22477<= not I29023;
	G22480<= not I29026;
	G22484<= not I29030;
	G22487<= not I29033;
	G22490<= not I29036;
	G22494<= not I29040;
	G22497<= not I29043;
	G22500<= not I29046;
	G22503<= not I29049;
	G22506<= not I29052;
	G22509<= not I29055;
	G22512<= not I29058;
	G22518<= not I29064;
	G22519<= not I29067;
	G22520<= not I29070;
	G22523<= not I29073;
	G22527<= not I29077;
	G22530<= not I29080;
	G22533<= not I29083;
	G22537<= not I29087;
	G22540<= not I29090;
	G22543<= not I29093;
	G22547<= not G21087;
	G22548<= not I29098;
	G22549<= not I29101;
	G22550<= not I29104;
	G22551<= not I29107;
	G22552<= not I29110;
	G22558<= not I29116;
	G22559<= not I29119;
	G22560<= not I29122;
	G22563<= not I29125;
	G22567<= not I29129;
	G22570<= not I29132;
	G22573<= not I29135;
	G22582<= not I29142;
	G22583<= not I29145;
	G22584<= not I29148;
	G22585<= not I29151;
	G22586<= not I29154;
	G22588<= not G21099;
	G22589<= not I29159;
	G22590<= not I29162;
	G22591<= not I29165;
	G22592<= not I29168;
	G22598<= not I29174;
	G22599<= not I29177;
	G22600<= not I29180;
	G22603<= not I29183;
	G22609<= not G21108;
	G22611<= not I29191;
	G22612<= not I29194;
	G22613<= not I29197;
	G22619<= not I29203;
	G22620<= not I29206;
	G22621<= not I29209;
	G22622<= not I29212;
	G22623<= not I29215;
	G22625<= not G21113;
	G22626<= not I29220;
	G22627<= not I29223;
	G22628<= not I29226;
	G22629<= not I29229;
	G22635<= not I29235;
	G22636<= not I29238;
	G22639<= not I29243;
	G22640<= not I29246;
	G22641<= not I29249;
	G22642<= not I29252;
	G22645<= not G21125;
	G22647<= not I29259;
	G22648<= not I29262;
	G22649<= not I29265;
	G22655<= not I29271;
	G22656<= not I29274;
	G22657<= not I29277;
	G22658<= not I29280;
	G22659<= not I29283;
	G22661<= not G21130;
	G22662<= not I29288;
	G22663<= not I29291;
	G22664<= not I29294;
	G22669<= not I29301;
	G22670<= not I29304;
	G22671<= not I29307;
	G22672<= not I29310;
	G22673<= not I29313;
	G22675<= not I29317;
	G22676<= not I29320;
	G22677<= not I29323;
	G22678<= not I29326;
	G22681<= not G21144;
	G22683<= not I29333;
	G22684<= not I29336;
	G22685<= not I29339;
	G22691<= not I29345;
	G22692<= not I29348;
	G22693<= not I29351;
	G22694<= not I29354;
	G22695<= not I29357;
	G22696<= not I29360;
	G22702<= not I29366;
	G22703<= not I29369;
	G22704<= not I29372;
	G22705<= not I29375;
	G22706<= not I29378;
	G22709<= not I29383;
	G22710<= not I29386;
	G22711<= not I29389;
	G22712<= not I29392;
	G22713<= not I29395;
	G22715<= not I29399;
	G22716<= not I29402;
	G22717<= not I29405;
	G22718<= not I29408;
	G22721<= not G21164;
	G22723<= not I29415;
	G22724<= not I29418;
	G22725<= not I29421;
	G22728<= not I29426;
	G22729<= not I29429;
	G22730<= not I29432;
	G22731<= not I29435;
	G22733<= not I29439;
	G22734<= not I29442;
	G22735<= not I29445;
	G22736<= not I29448;
	G22737<= not I29451;
	G22740<= not I29456;
	G22741<= not I29459;
	G22742<= not I29462;
	G22743<= not I29465;
	G22744<= not I29468;
	G22746<= not I29472;
	G22747<= not I29475;
	G22748<= not I29478;
	G22749<= not I29481;
	G22750<= not I29484;
	G22753<= not G21184;
	G22756<= not I29490;
	G22757<= not I29493;
	G22758<= not I29496;
	G22760<= not I29500;
	G22761<= not I29503;
	G22762<= not I29506;
	G22763<= not I29509;
	G22765<= not I29513;
	G22766<= not I29516;
	G22767<= not I29519;
	G22768<= not I29522;
	G22769<= not I29525;
	G22772<= not I29530;
	G22773<= not I29533;
	G22774<= not I29536;
	G22775<= not I29539;
	G22776<= not I29542;
	G22777<= not G21796;
	G22785<= not I29547;
	G22786<= not I29550;
	G22787<= not G21199;
	G22790<= not I29556;
	G22791<= not I29559;
	G22792<= not I29562;
	G22794<= not I29566;
	G22795<= not I29569;
	G22796<= not I29572;
	G22797<= not I29575;
	G22799<= not I29579;
	G22800<= not I29582;
	G22801<= not I29585;
	G22802<= not I29588;
	G22803<= not I29591;
	G22805<= not G21894;
	G22806<= not G21615;
	G22812<= not I29600;
	G22824<= not I29603;
	G22825<= not I29606;
	G22827<= not I29610;
	G22828<= not I29613;
	G22829<= not G21214;
	G22832<= not I29619;
	G22833<= not I29622;
	G22834<= not I29625;
	G22836<= not I29629;
	G22837<= not I29632;
	G22838<= not I29635;
	G22839<= not I29638;
	G22840<= not I29641;
	G22843<= not G21889;
	G22847<= not G21643;
	G22852<= not I29653;
	G22864<= not I29656;
	G22866<= not I29660;
	G22867<= not I29663;
	G22868<= not G21222;
	G22871<= not I29669;
	G22872<= not I29672;
	G22873<= not I29675;
	G22875<= not G21884;
	G22882<= not G21674;
	G22887<= not I29687;
	G22899<= not I29690;
	G22901<= not I29694;
	G22902<= not I29697;
	G22903<= not I29700;
	G22907<= not G21711;
	G22917<= not G21703;
	G22922<= not I29712;
	G22934<= not I29715;
	G22945<= not I29724;
	G22948<= not I29727;
	G22949<= not G21665;
	G22954<= not G21739;
	G22958<= not G21694;
	G22962<= not G21763;
	G22966<= not G21730;
	G22970<= not I29736;
	G22971<= not G21779;
	G22975<= not G21756;
	G22979<= not I29741;
	G22980<= not G21794;
	G22986<= not G21382;
	G22988<= not G21404;
	G22989<= not G21415;
	G22991<= not G21429;
	G22995<= not G21441;
	G22996<= not G21449;
	G22998<= not G21458;
	G23001<= not G21473;
	G23002<= not G21477;
	G23006<= not G21483;
	G23007<= not G21491;
	G23008<= not G21498;
	G23012<= not G21505;
	G23015<= not G21514;
	G23016<= not G21518;
	G23020<= not G21524;
	G23021<= not G21530;
	G23024<= not G21537;
	G23028<= not G21541;
	G23031<= not G21550;
	G23032<= not G21554;
	G23036<= not G21558;
	G23037<= not G21561;
	G23038<= not G21566;
	G23041<= not G21573;
	G23045<= not G21577;
	G23048<= not G21586;
	G23049<= not G21590;
	G23050<= not I29797;
	G23055<= not I29802;
	G23056<= not G21594;
	G23057<= not G21599;
	G23060<= not G21606;
	G23064<= not G21612;
	G23065<= not I29812;
	G23068<= not I29817;
	G23069<= not G21619;
	G23074<= not G21623;
	G23075<= not G21628;
	G23078<= not I29827;
	G23079<= not G21640;
	G23082<= not G21647;
	G23087<= not G21651;
	G23088<= not G21655;
	G23094<= not I29841;
	G23095<= not G21671;
	G23098<= not G21678;
	G23103<= not G21682;
	G23105<= not I29852;
	G23112<= not G21700;
	G23115<= not G21708;
	G23116<= not I29863;
	G23125<= not I29872;
	G23134<= not I29881;
	G23140<= not G21825;
	G23141<= not G21825;
	G23142<= not G21825;
	G23143<= not G21825;
	G23144<= not G21825;
	G23145<= not G21825;
	G23146<= not G21825;
	G23147<= not G21825;
	G23148<= not I29897;
	G23149<= not I29900;
	G23150<= not I29903;
	G23151<= not I29906;
	G23152<= not I29909;
	G23153<= not I29912;
	G23154<= not I29915;
	G23155<= not I29918;
	G23156<= not I29921;
	G23157<= not I29924;
	G23158<= not I29927;
	G23159<= not I29930;
	G23160<= not I29933;
	G23161<= not I29936;
	G23162<= not I29939;
	G23163<= not I29942;
	G23164<= not I29945;
	G23165<= not I29948;
	G23166<= not I29951;
	G23167<= not I29954;
	G23168<= not I29957;
	G23169<= not I29960;
	G23170<= not I29963;
	G23171<= not I29966;
	G23172<= not I29969;
	G23173<= not I29972;
	G23174<= not I29975;
	G23175<= not I29978;
	G23176<= not I29981;
	G23177<= not I29984;
	G23178<= not I29987;
	G23179<= not I29990;
	G23180<= not I29993;
	G23181<= not I29996;
	G23182<= not I29999;
	G23183<= not I30002;
	G23184<= not I30005;
	G23185<= not I30008;
	G23186<= not I30011;
	G23187<= not I30014;
	G23188<= not I30017;
	G23189<= not I30020;
	G23190<= not I30023;
	G23191<= not I30026;
	G23192<= not I30029;
	G23193<= not I30032;
	G23194<= not I30035;
	G23195<= not I30038;
	G23196<= not I30041;
	G23197<= not I30044;
	G23198<= not I30047;
	G23199<= not I30050;
	G23200<= not I30053;
	G23201<= not I30056;
	G23202<= not I30059;
	G23203<= not I30062;
	G23204<= not I30065;
	G23205<= not I30068;
	G23206<= not I30071;
	G23207<= not I30074;
	G23208<= not I30077;
	G23209<= not I30080;
	G23210<= not I30083;
	G23211<= not I30086;
	G23212<= not I30089;
	G23213<= not I30092;
	G23214<= not I30095;
	G23215<= not I30098;
	G23216<= not I30101;
	G23217<= not I30104;
	G23218<= not I30107;
	G23219<= not I30110;
	G23220<= not I30113;
	G23221<= not I30116;
	G23222<= not I30119;
	G23223<= not I30122;
	G23224<= not I30125;
	G23225<= not I30128;
	G23226<= not I30131;
	G23227<= not I30134;
	G23228<= not I30137;
	G23229<= not I30140;
	G23230<= not I30143;
	G23231<= not I30146;
	G23232<= not I30149;
	G23233<= not I30152;
	G23234<= not I30155;
	G23235<= not I30158;
	G23236<= not I30161;
	G23237<= not I30164;
	G23238<= not I30167;
	G23239<= not I30170;
	G23240<= not I30173;
	G23241<= not I30176;
	G23242<= not I30179;
	G23243<= not I30182;
	G23244<= not I30185;
	G23245<= not I30188;
	G23246<= not I30191;
	G23247<= not I30194;
	G23248<= not I30197;
	G23249<= not I30200;
	G23250<= not I30203;
	G23251<= not I30206;
	G23252<= not I30209;
	G23253<= not I30212;
	G23254<= not I30215;
	G23255<= not I30218;
	G23256<= not I30221;
	G23257<= not I30224;
	G23258<= not I30227;
	G23259<= not I30230;
	G23260<= not I30233;
	G23261<= not I30236;
	G23262<= not I30239;
	G23263<= not I30242;
	G23264<= not I30245;
	G23265<= not I30248;
	G23266<= not I30251;
	G23267<= not I30254;
	G23268<= not I30257;
	G23269<= not I30260;
	G23270<= not I30263;
	G23271<= not I30266;
	G23272<= not I30269;
	G23273<= not I30272;
	G23274<= not I30275;
	G23275<= not I30278;
	G23276<= not I30281;
	G23277<= not I30284;
	G23278<= not I30287;
	G23279<= not I30290;
	G23280<= not I30293;
	G23281<= not I30296;
	G23282<= not I30299;
	G23283<= not I30302;
	G23284<= not I30305;
	G23285<= not I30308;
	G23286<= not I30311;
	G23287<= not I30314;
	G23288<= not I30317;
	G23289<= not I30320;
	G23290<= not I30323;
	G23291<= not I30326;
	G23292<= not I30329;
	G23293<= not I30332;
	G23294<= not I30335;
	G23295<= not I30338;
	G23296<= not I30341;
	G23297<= not I30344;
	G23298<= not I30347;
	G23299<= not I30350;
	G23300<= not I30353;
	G23301<= not I30356;
	G23302<= not I30359;
	G23303<= not I30362;
	G23304<= not I30365;
	G23305<= not I30368;
	G23306<= not I30371;
	G23307<= not I30374;
	G23308<= not I30377;
	G23309<= not I30380;
	G23310<= not I30383;
	G23311<= not I30386;
	G23312<= not I30389;
	G23313<= not I30392;
	G23314<= not I30395;
	G23315<= not I30398;
	G23316<= not I30401;
	G23317<= not I30404;
	G23318<= not I30407;
	G23403<= not G23052;
	G23410<= not G23071;
	G23415<= not G23084;
	G23420<= not G23089;
	G23424<= not G23100;
	G23429<= not G23107;
	G23435<= not G23120;
	G23438<= not I30467;
	G23439<= not I30470;
	G23441<= not G23129;
	G23444<= not G22945;
	G23448<= not I30476;
	G23452<= not I30480;
	G23453<= not I30483;
	G23454<= not I30486;
	G23455<= not I30489;
	G23459<= not I30493;
	G23460<= not I30496;
	G23463<= not I30501;
	G23464<= not I30504;
	G23468<= not I30508;
	G23469<= not I30511;
	G23470<= not G22188;
	G23472<= not I30516;
	G23473<= not I30519;
	G23481<= not I30525;
	G23482<= not G22197;
	G23485<= not I30531;
	G23492<= not I30536;
	G23493<= not G22203;
	G23500<= not I30544;
	G23501<= not I30547;
	G23508<= not I30552;
	G23509<= not G22209;
	G23516<= not I30560;
	G23517<= not I30563;
	G23524<= not I30568;
	G23531<= not I30575;
	G23532<= not I30578;
	G23542<= not I30586;
	G23543<= not I30589;
	G23546<= not I30594;
	G23548<= not I30598;
	G23549<= not I30601;
	G23553<= not I30607;
	G23555<= not I30611;
	G23556<= not I30614;
	G23557<= not I30617;
	G23561<= not I30623;
	G23562<= not I30626;
	G23566<= not I30632;
	G23568<= not I30636;
	G23569<= not I30639;
	G23570<= not I30642;
	G23574<= not I30648;
	G23575<= not I30651;
	G23576<= not I30654;
	G23580<= not I30660;
	G23581<= not I30663;
	G23585<= not I30669;
	G23587<= not I30673;
	G23588<= not I30676;
	G23589<= not I30679;
	G23594<= not I30686;
	G23595<= not I30689;
	G23596<= not I30692;
	G23597<= not I30695;
	G23601<= not I30701;
	G23602<= not I30704;
	G23603<= not I30707;
	G23607<= not I30713;
	G23608<= not I30716;
	G23612<= not I30722;
	G23613<= not I30725;
	G23614<= not I30728;
	G23619<= not I30735;
	G23620<= not I30738;
	G23621<= not I30741;
	G23626<= not I30748;
	G23627<= not I30751;
	G23628<= not I30754;
	G23629<= not I30757;
	G23633<= not I30763;
	G23634<= not I30766;
	G23635<= not I30769;
	G23640<= not I30776;
	G23641<= not I30779;
	G23642<= not I30782;
	G23644<= not I30786;
	G23661<= not I30797;
	G23662<= not I30800;
	G23663<= not I30803;
	G23668<= not I30810;
	G23669<= not I30813;
	G23670<= not I30816;
	G23675<= not I30823;
	G23676<= not I30826;
	G23677<= not I30829;
	G23678<= not I30832;
	G23682<= not I30838;
	G23683<= not I30841;
	G23684<= not I30844;
	G23685<= not I30847;
	G23690<= not I30854;
	G23691<= not I30857;
	G23692<= not I30860;
	G23694<= not I30864;
	G23711<= not I30875;
	G23712<= not I30878;
	G23713<= not I30881;
	G23718<= not I30888;
	G23719<= not I30891;
	G23720<= not I30894;
	G23725<= not I30901;
	G23727<= not I30905;
	G23728<= not I30908;
	G23729<= not I30911;
	G23730<= not I30914;
	G23731<= not I30917;
	G23736<= not I30922;
	G23737<= not I30925;
	G23738<= not I30928;
	G23739<= not I30931;
	G23744<= not I30938;
	G23745<= not I30941;
	G23746<= not I30944;
	G23748<= not I30948;
	G23765<= not I30959;
	G23766<= not I30962;
	G23767<= not I30965;
	G23773<= not I30973;
	G23774<= not I30976;
	G23775<= not I30979;
	G23779<= not I30985;
	G23782<= not I30988;
	G23783<= not I30991;
	G23784<= not I30994;
	G23785<= not I30997;
	G23786<= not I31000;
	G23791<= not I31005;
	G23792<= not I31008;
	G23793<= not I31011;
	G23794<= not I31014;
	G23799<= not I31021;
	G23800<= not I31024;
	G23801<= not I31027;
	G23803<= not I31031;
	G23821<= not I31043;
	G23826<= not I31050;
	G23827<= not I31053;
	G23828<= not I31056;
	G23832<= not I31062;
	G23835<= not I31065;
	G23836<= not I31068;
	G23837<= not I31071;
	G23838<= not I31074;
	G23839<= not I31077;
	G23844<= not I31082;
	G23845<= not I31085;
	G23846<= not I31088;
	G23847<= not I31091;
	G23853<= not G22300;
	G23856<= not I31102;
	G23861<= not I31109;
	G23862<= not I31112;
	G23863<= not I31115;
	G23867<= not I31121;
	G23870<= not I31124;
	G23871<= not I31127;
	G23872<= not I31130;
	G23873<= not I31133;
	G23874<= not I31136;
	G23879<= not I31141;
	G23882<= not I31144;
	G23885<= not G22062;
	G23887<= not G22328;
	G23890<= not I31152;
	G23895<= not I31159;
	G23896<= not I31162;
	G23897<= not I31165;
	G23901<= not I31171;
	G23905<= not G22046;
	G23908<= not G22353;
	G23911<= not I31181;
	G23916<= not I31188;
	G23918<= not G22036;
	G23923<= not I31195;
	G23940<= not G22376;
	G23943<= not I31205;
	G23955<= not I31213;
	G23984<= not I31226;
	G24000<= not I31232;
	G24001<= not I31235;
	G24014<= not I31244;
	G24030<= not I31250;
	G24033<= not I31253;
	G24035<= not I31257;
	G24047<= not G23023;
	G24051<= not I31266;
	G24053<= not I31270;
	G24055<= not I31274;
	G24060<= not G23040;
	G24064<= not I31282;
	G24066<= not I31286;
	G24068<= not I31290;
	G24073<= not G23059;
	G24077<= not I31298;
	G24079<= not I31302;
	G24084<= not G23077;
	G24088<= not I31310;
	G24094<= not G22339;
	G24095<= not G22362;
	G24096<= not G22405;
	G24097<= not G22382;
	G24098<= not G22409;
	G24099<= not G22412;
	G24101<= not G22415;
	G24102<= not G22418;
	G24103<= not G22397;
	G24104<= not G22422;
	G24105<= not G22425;
	G24106<= not G22428;
	G24107<= not G22431;
	G24108<= not G22434;
	G24110<= not G22437;
	G24111<= not G22440;
	G24112<= not G22445;
	G24113<= not G22448;
	G24114<= not G22451;
	G24115<= not G22381;
	G24121<= not G22455;
	G24122<= not G22458;
	G24123<= not G22461;
	G24124<= not G22464;
	G24125<= not G22467;
	G24127<= not G22470;
	G24128<= not G22473;
	G24129<= not G22477;
	G24130<= not G22480;
	G24131<= not G22484;
	G24132<= not G22487;
	G24133<= not G22490;
	G24134<= not G22396;
	G24140<= not G22494;
	G24141<= not G22497;
	G24142<= not G22500;
	G24143<= not G22503;
	G24144<= not G22506;
	G24146<= not G22509;
	G24147<= not G22512;
	G24148<= not G22520;
	G24149<= not G22523;
	G24150<= not G22527;
	G24151<= not G22530;
	G24152<= not G22533;
	G24153<= not G22399;
	G24159<= not G22537;
	G24160<= not G22540;
	G24161<= not G22543;
	G24162<= not G22552;
	G24163<= not G22560;
	G24164<= not G22563;
	G24165<= not G22567;
	G24166<= not G22570;
	G24167<= not G22573;
	G24168<= not G22400;
	G24175<= not G22592;
	G24176<= not G22600;
	G24177<= not G22603;
	G24180<= not G22629;
	G24183<= not I31387;
	G24210<= not G22696;
	G24220<= not G22750;
	G24233<= not I31417;
	G24240<= not I31426;
	G24248<= not I31436;
	G24251<= not G22903;
	G24255<= not I31445;
	G24259<= not I31451;
	G24260<= not I31454;
	G24261<= not I31457;
	G24262<= not I31460;
	G24263<= not I31463;
	G24264<= not I31466;
	G24265<= not I31469;
	G24266<= not I31472;
	G24267<= not I31475;
	G24268<= not I31478;
	G24269<= not I31481;
	G24270<= not I31484;
	G24271<= not I31487;
	G24272<= not I31490;
	G24273<= not I31493;
	G24274<= not I31496;
	G24275<= not I31499;
	G24276<= not I31502;
	G24277<= not I31505;
	G24278<= not I31508;
	G24279<= not I31511;
	G24280<= not I31514;
	G24281<= not I31517;
	G24282<= not I31520;
	G24283<= not I31523;
	G24284<= not I31526;
	G24285<= not I31529;
	G24286<= not I31532;
	G24287<= not I31535;
	G24288<= not I31538;
	G24289<= not I31541;
	G24290<= not I31544;
	G24291<= not I31547;
	G24292<= not I31550;
	G24293<= not I31553;
	G24294<= not I31556;
	G24295<= not I31559;
	G24296<= not I31562;
	G24297<= not I31565;
	G24298<= not I31568;
	G24299<= not I31571;
	G24300<= not I31574;
	G24301<= not I31577;
	G24302<= not I31580;
	G24303<= not I31583;
	G24304<= not I31586;
	G24305<= not I31589;
	G24306<= not I31592;
	G24307<= not I31595;
	G24308<= not I31598;
	G24309<= not I31601;
	G24310<= not I31604;
	G24311<= not I31607;
	G24312<= not I31610;
	G24313<= not I31613;
	G24314<= not I31616;
	G24315<= not I31619;
	G24316<= not I31622;
	G24317<= not I31625;
	G24318<= not I31628;
	G24319<= not I31631;
	G24320<= not I31634;
	G24321<= not I31637;
	G24322<= not I31640;
	G24323<= not I31643;
	G24324<= not I31646;
	G24325<= not I31649;
	G24326<= not I31652;
	G24327<= not I31655;
	G24328<= not I31658;
	G24329<= not I31661;
	G24330<= not I31664;
	G24331<= not I31667;
	G24332<= not I31670;
	G24333<= not I31673;
	G24334<= not I31676;
	G24335<= not I31679;
	G24336<= not I31682;
	G24337<= not I31685;
	G24338<= not I31688;
	G24339<= not I31691;
	G24340<= not I31694;
	G24341<= not I31697;
	G24342<= not I31700;
	G24343<= not I31703;
	G24344<= not I31706;
	G24345<= not I31709;
	G24346<= not I31712;
	G24347<= not I31715;
	G24348<= not I31718;
	G24349<= not I31721;
	G24350<= not I31724;
	G24351<= not I31727;
	G24352<= not I31730;
	G24353<= not I31733;
	G24354<= not I31736;
	G24355<= not I31739;
	G24356<= not I31742;
	G24357<= not I31745;
	G24358<= not I31748;
	G24359<= not I31751;
	G24360<= not I31754;
	G24361<= not I31757;
	G24362<= not I31760;
	G24363<= not I31763;
	G24364<= not I31766;
	G24365<= not I31769;
	G24366<= not I31772;
	G24367<= not I31775;
	G24368<= not I31778;
	G24369<= not I31781;
	G24370<= not I31784;
	G24371<= not I31787;
	G24372<= not I31790;
	G24373<= not I31793;
	G24374<= not I31796;
	G24375<= not I31799;
	G24376<= not I31802;
	G24377<= not I31805;
	G24378<= not I31808;
	G24379<= not I31811;
	G24380<= not I31814;
	G24381<= not I31817;
	G24382<= not I31820;
	G24383<= not I31823;
	G24384<= not I31826;
	G24385<= not I31829;
	G24386<= not I31832;
	G24387<= not I31835;
	G24388<= not I31838;
	G24389<= not I31841;
	G24390<= not I31844;
	G24391<= not I31847;
	G24392<= not I31850;
	G24393<= not I31853;
	G24394<= not I31856;
	G24395<= not I31859;
	G24396<= not I31862;
	G24397<= not I31865;
	G24398<= not I31868;
	G24399<= not I31871;
	G24400<= not I31874;
	G24401<= not I31877;
	G24402<= not I31880;
	G24403<= not I31883;
	G24404<= not I31886;
	G24405<= not I31889;
	G24406<= not I31892;
	G24407<= not I31895;
	G24408<= not I31898;
	G24409<= not I31901;
	G24410<= not I31904;
	G24411<= not I31907;
	G24412<= not I31910;
	G24413<= not I31913;
	G24414<= not I31916;
	G24415<= not I31919;
	G24416<= not I31922;
	G24417<= not I31925;
	G24418<= not I31928;
	G24419<= not I31931;
	G24420<= not I31934;
	G24421<= not I31937;
	G24422<= not I31940;
	G24423<= not I31943;
	G24424<= not I31946;
	G24425<= not I31949;
	G24482<= not G24183;
	G24518<= not I32042;
	G24531<= not I32057;
	G24539<= not I32067;
	G24544<= not I32074;
	G24549<= not I32081;
	G24551<= not I32085;
	G24556<= not I32092;
	G24560<= not I32098;
	G24562<= not I32102;
	G24567<= not I32109;
	G24568<= not I32112;
	G24570<= not I32116;
	G24572<= not I32120;
	G24576<= not I32126;
	G24577<= not I32129;
	G24579<= not I32133;
	G24581<= not I32137;
	G24582<= not I32140;
	G24583<= not I32143;
	G24584<= not I32146;
	G24586<= not I32150;
	G24587<= not I32153;
	G24588<= not I32156;
	G24589<= not I32159;
	G24592<= not I32164;
	G24593<= not I32167;
	G24594<= not I32170;
	G24597<= not I32175;
	G24598<= not I32178;
	G24599<= not I32181;
	G24600<= not I32184;
	G24605<= not I32189;
	G24607<= not I32193;
	G24612<= not I32198;
	G24619<= not I32203;
	G24630<= not I32210;
	G24648<= not G23470;
	G24668<= not G23482;
	G24687<= not G23493;
	G24704<= not G23509;
	G24734<= not I32248;
	G24735<= not I32251;
	G24763<= not I32281;
	G24784<= not I32320;
	G24805<= not I32365;
	G24815<= not G23448;
	G24816<= not I32388;
	G24827<= not I32419;
	G24834<= not G23455;
	G24835<= not I32439;
	G24850<= not G23464;
	G24851<= not I32487;
	G24856<= not I32506;
	G24864<= not G23473;
	G24865<= not I32535;
	G24872<= not I32556;
	G24879<= not I32583;
	G24886<= not I32604;
	G24893<= not G23486;
	G24903<= not I32642;
	G24912<= not G23495;
	G24916<= not G23502;
	G24929<= not G23511;
	G24933<= not G23518;
	G24939<= not G23660;
	G24941<= not G23526;
	G24945<= not G23533;
	G24949<= not I32704;
	G24950<= not G23710;
	G24952<= not G23537;
	G24956<= not I32716;
	G24957<= not I32719;
	G24958<= not G23478;
	G24962<= not G23764;
	G24969<= not G23489;
	G24973<= not G23819;
	G24982<= not G23505;
	G24993<= not G23521;
	G25087<= not G23731;
	G25094<= not G23779;
	G25095<= not G23786;
	G25103<= not I32829;
	G25104<= not G23832;
	G25105<= not G23839;
	G25109<= not I32835;
	G25110<= not G23867;
	G25111<= not G23874;
	G25115<= not G23879;
	G25116<= not G23882;
	G25118<= not I32844;
	G25119<= not I32847;
	G25120<= not G23901;
	G25121<= not I32851;
	G25122<= not I32854;
	G25123<= not I32857;
	G25124<= not I32860;
	G25126<= not G24030;
	G25130<= not I32868;
	G25131<= not I32871;
	G25132<= not I32874;
	G25133<= not I32877;
	G25134<= not I32880;
	G25135<= not I32883;
	G25136<= not I32886;
	G25137<= not I32889;
	G25138<= not I32892;
	G25139<= not I32895;
	G25140<= not I32898;
	G25141<= not I32901;
	G25142<= not I32904;
	G25143<= not I32907;
	G25144<= not I32910;
	G25145<= not I32913;
	G25146<= not I32916;
	G25147<= not I32919;
	G25148<= not I32922;
	G25149<= not I32925;
	G25150<= not I32928;
	G25151<= not I32931;
	G25152<= not I32934;
	G25153<= not I32937;
	G25154<= not I32940;
	G25155<= not I32943;
	G25156<= not I32946;
	G25157<= not I32949;
	G25158<= not I32952;
	G25159<= not I32955;
	G25160<= not I32958;
	G25161<= not I32961;
	G25162<= not I32964;
	G25163<= not I32967;
	G25164<= not I32970;
	G25165<= not I32973;
	G25166<= not I32976;
	G25167<= not I32979;
	G25168<= not I32982;
	G25169<= not I32985;
	G25170<= not I32988;
	G25171<= not I32991;
	G25172<= not I32994;
	G25173<= not I32997;
	G25174<= not I33000;
	G25175<= not I33003;
	G25176<= not I33006;
	G25177<= not I33009;
	G25179<= not I33013;
	G25180<= not I33016;
	G25274<= not G24912;
	G25283<= not G24929;
	G25291<= not G24941;
	G25296<= not I33128;
	G25301<= not G24952;
	G25305<= not G24880;
	G25306<= not I33136;
	G25313<= not G24868;
	G25314<= not G24897;
	G25315<= not I33145;
	G25319<= not G24857;
	G25322<= not G24883;
	G25323<= not G24920;
	G25324<= not I33154;
	G25327<= not I33157;
	G25329<= not G24844;
	G25330<= not G24873;
	G25332<= not G24900;
	G25333<= not G24937;
	G25335<= not G24832;
	G25336<= not I33168;
	G25338<= not G24860;
	G25339<= not G24887;
	G25341<= not G24923;
	G25347<= not G24817;
	G25349<= not G24848;
	G25350<= not I33182;
	G25352<= not G24875;
	G25353<= not G24904;
	G25354<= not I33188;
	G25355<= not G24797;
	G25361<= not G24837;
	G25363<= not G24862;
	G25364<= not I33198;
	G25366<= not G24889;
	G25367<= not G24676;
	G25368<= not G24778;
	G25369<= not I33205;
	G25370<= not G24820;
	G25376<= not G24852;
	G25378<= not G24877;
	G25379<= not G24893;
	G25383<= not G24766;
	G25384<= not G24695;
	G25385<= not G24801;
	G25386<= not I33219;
	G25387<= not G24839;
	G25393<= not G24866;
	G25394<= not G24753;
	G25395<= not G24916;
	G25399<= not G24787;
	G25400<= not G24712;
	G25401<= not G24823;
	G25402<= not I33232;
	G25403<= not G24854;
	G25404<= not G24771;
	G25405<= not G24933;
	G25409<= not G24808;
	G25410<= not G24723;
	G25411<= not G24842;
	G25412<= not G24791;
	G25413<= not G24945;
	G25417<= not G24830;
	G25419<= not G24812;
	G25420<= not I33246;
	G25421<= not I33249;
	G25422<= not G24958;
	G25430<= not G24616;
	G25431<= not G24969;
	G25435<= not I33257;
	G25436<= not I33260;
	G25437<= not G24627;
	G25438<= not G24982;
	G25442<= not I33265;
	G25443<= not I33268;
	G25444<= not G24641;
	G25445<= not G24993;
	G25449<= not G24660;
	G25454<= not I33278;
	G25458<= not I33282;
	G25462<= not I33286;
	G25463<= not I33289;
	G25467<= not I33293;
	G25471<= not I33297;
	G25472<= not I33300;
	G25476<= not I33304;
	G25479<= not I33307;
	G25484<= not I33312;
	G25488<= not I33316;
	G25493<= not I33321;
	G25496<= not I33324;
	G25499<= not I33327;
	G25502<= not I33330;
	G25507<= not I33335;
	G25510<= not I33338;
	G25515<= not I33343;
	G25519<= not I33347;
	G25524<= not I33352;
	G25527<= not I33355;
	G25530<= not I33358;
	G25533<= not I33361;
	G25536<= not I33364;
	G25540<= not I33368;
	G25543<= not I33371;
	G25546<= not I33374;
	G25549<= not I33377;
	G25554<= not I33382;
	G25557<= not I33385;
	G25562<= not I33390;
	G25573<= not I33396;
	G25576<= not I33399;
	G25579<= not I33402;
	G25582<= not I33405;
	G25585<= not I33408;
	G25588<= not I33411;
	G25590<= not I33415;
	G25593<= not I33418;
	G25596<= not I33421;
	G25599<= not I33424;
	G25602<= not I33427;
	G25606<= not I33431;
	G25609<= not I33434;
	G25612<= not I33437;
	G25615<= not I33440;
	G25620<= not I33445;
	G25623<= not I33448;
	G25630<= not G24478;
	G25634<= not I33457;
	G25637<= not I33460;
	G25640<= not I33463;
	G25643<= not I33466;
	G25646<= not I33469;
	G25647<= not I33472;
	G25652<= not I33476;
	G25655<= not I33479;
	G25658<= not I33482;
	G25661<= not I33485;
	G25664<= not I33488;
	G25667<= not I33491;
	G25669<= not I33495;
	G25672<= not I33498;
	G25675<= not I33501;
	G25678<= not I33504;
	G25681<= not I33507;
	G25685<= not I33511;
	G25688<= not I33514;
	G25691<= not I33517;
	G25694<= not I33520;
	G25698<= not G24600;
	G25700<= not I33526;
	G25703<= not I33529;
	G25706<= not I33532;
	G25707<= not I33535;
	G25711<= not I33539;
	G25714<= not I33542;
	G25717<= not I33545;
	G25720<= not I33548;
	G25723<= not I33551;
	G25724<= not I33554;
	G25729<= not I33558;
	G25732<= not I33561;
	G25735<= not I33564;
	G25738<= not I33567;
	G25741<= not I33570;
	G25744<= not I33573;
	G25746<= not I33577;
	G25749<= not I33580;
	G25752<= not I33583;
	G25755<= not I33586;
	G25758<= not I33589;
	G25762<= not I33593;
	G25763<= not I33596;
	G25767<= not I33600;
	G25770<= not I33603;
	G25771<= not G24607;
	G25773<= not I33608;
	G25776<= not I33611;
	G25779<= not I33614;
	G25780<= not I33617;
	G25784<= not I33621;
	G25787<= not I33624;
	G25790<= not I33627;
	G25793<= not I33630;
	G25796<= not I33633;
	G25797<= not I33636;
	G25802<= not I33640;
	G25805<= not I33643;
	G25808<= not I33646;
	G25811<= not I33649;
	G25814<= not I33652;
	G25817<= not I33655;
	G25821<= not I33659;
	G25824<= not I33662;
	G25825<= not G24619;
	G25827<= not I33667;
	G25830<= not I33670;
	G25833<= not I33673;
	G25834<= not I33676;
	G25838<= not I33680;
	G25841<= not I33683;
	G25844<= not I33686;
	G25847<= not I33689;
	G25850<= not I33692;
	G25851<= not I33695;
	G25856<= not I33700;
	G25859<= not I33703;
	G25860<= not G24630;
	G25862<= not I33708;
	G25865<= not I33711;
	G25868<= not I33714;
	G25869<= not I33717;
	G25877<= not I33723;
	G25880<= not I33726;
	G25886<= not I33732;
	G25891<= not I33737;
	G25895<= not G24939;
	G25899<= not G24928;
	G25903<= not G24950;
	G25907<= not G24940;
	G25911<= not G24962;
	G25915<= not G24951;
	G25919<= not G24973;
	G25923<= not G24963;
	G25937<= not G24763;
	G25939<= not G24784;
	G25942<= not G24805;
	G25945<= not G24827;
	G25952<= not G24735;
	G25976<= not I33790;
	G25982<= not I33798;
	G25983<= not I33801;
	G25984<= not I33804;
	G25985<= not I33807;
	G25986<= not I33810;
	G25987<= not I33813;
	G25988<= not I33816;
	G25989<= not I33819;
	G25990<= not I33822;
	G25991<= not I33825;
	G25992<= not I33828;
	G25993<= not I33831;
	G25994<= not I33834;
	G25995<= not I33837;
	G25996<= not I33840;
	G25997<= not I33843;
	G25998<= not I33846;
	G25999<= not I33849;
	G26000<= not I33852;
	G26001<= not I33855;
	G26002<= not I33858;
	G26003<= not I33861;
	G26004<= not I33864;
	G26005<= not I33867;
	G26006<= not I33870;
	G26007<= not I33873;
	G26008<= not I33876;
	G26009<= not I33879;
	G26010<= not I33882;
	G26011<= not I33885;
	G26012<= not I33888;
	G26013<= not I33891;
	G26014<= not I33894;
	G26015<= not I33897;
	G26016<= not I33900;
	G26017<= not I33903;
	G26018<= not I33906;
	G26019<= not I33909;
	G26020<= not I33912;
	G26021<= not I33915;
	G26022<= not I33918;
	G26056<= not I33954;
	G26063<= not I33961;
	G26070<= not I33968;
	G26076<= not I33974;
	G26086<= not I33984;
	G26092<= not I33990;
	G26102<= not I33995;
	G26104<= not I33999;
	G26105<= not I34002;
	G26114<= not I34009;
	G26118<= not I34012;
	G26121<= not I34017;
	G26125<= not I34020;
	G26131<= not I34026;
	G26135<= not I34029;
	G26136<= not I34032;
	G26149<= not I34041;
	G26150<= not I34044;
	G26159<= not I34051;
	G26164<= not I34056;
	G26165<= not I34059;
	G26167<= not I34063;
	G26172<= not I34068;
	G26173<= not I34071;
	G26174<= not I34074;
	G26175<= not I34077;
	G26178<= not I34080;
	G26181<= not I34083;
	G26182<= not I34086;
	G26187<= not I34091;
	G26189<= not G25952;
	G26190<= not I34096;
	G26191<= not I34099;
	G26192<= not I34102;
	G26193<= not I34105;
	G26194<= not I34108;
	G26195<= not I34111;
	G26196<= not I34114;
	G26202<= not I34118;
	G26205<= not I34121;
	G26206<= not I34124;
	G26208<= not I34128;
	G26209<= not G25296;
	G26210<= not I34132;
	G26211<= not I34135;
	G26214<= not I34140;
	G26215<= not I34143;
	G26216<= not I34146;
	G26220<= not I34150;
	G26221<= not I34153;
	G26222<= not I34156;
	G26223<= not I34159;
	G26226<= not I34162;
	G26229<= not I34165;
	G26230<= not I34168;
	G26232<= not I34172;
	G26237<= not G25306;
	G26238<= not I34180;
	G26239<= not I34183;
	G26245<= not I34189;
	G26246<= not I34192;
	G26247<= not I34195;
	G26248<= not I34198;
	G26249<= not I34201;
	G26250<= not I34204;
	G26251<= not I34207;
	G26254<= not I34210;
	G26264<= not I34220;
	G26275<= not G25315;
	G26276<= not I34230;
	G26277<= not I34233;
	G26280<= not I34238;
	G26281<= not I34241;
	G26282<= not I34244;
	G26294<= not I34254;
	G26308<= not I34266;
	G26313<= not G25324;
	G26314<= not I34274;
	G26315<= not I34277;
	G26341<= not I34296;
	G26349<= not I34306;
	G26354<= not I34313;
	G26355<= not I34316;
	G26358<= not I34321;
	G26364<= not I34327;
	G26385<= not I34343;
	G26393<= not I34353;
	G26398<= not I34358;
	G26401<= not I34363;
	G26407<= not I34369;
	G26428<= not I34385;
	G26429<= not I34388;
	G26433<= not I34392;
	G26434<= not I34395;
	G26439<= not I34400;
	G26442<= not I34405;
	G26448<= not I34411;
	G26461<= not I34421;
	G26465<= not I34425;
	G26466<= not I34428;
	G26471<= not I34433;
	G26474<= not I34438;
	G26480<= not I34444;
	G26481<= not G25764;
	G26485<= not I34449;
	G26489<= not I34453;
	G26490<= not I34456;
	G26495<= not I34461;
	G26496<= not I34464;
	G26497<= not G25818;
	G26501<= not I34469;
	G26505<= not I34473;
	G26506<= not I34476;
	G26507<= not I34479;
	G26508<= not G25312;
	G26512<= not G25853;
	G26516<= not G25320;
	G26520<= not G25874;
	G26521<= not G25331;
	G26525<= not G25340;
	G26533<= not G25454;
	G26538<= not G25458;
	G26539<= not G25463;
	G26540<= not G25467;
	G26542<= not G25472;
	G26543<= not G25476;
	G26544<= not G25479;
	G26546<= not G25484;
	G26548<= not I34505;
	G26549<= not G25421;
	G26550<= not G25493;
	G26551<= not G25496;
	G26552<= not G25499;
	G26554<= not G25502;
	G26555<= not G25507;
	G26556<= not G25510;
	G26558<= not G25515;
	G26561<= not G25524;
	G26562<= not G25527;
	G26563<= not G25530;
	G26564<= not G25533;
	G26565<= not G25536;
	G26566<= not G25540;
	G26567<= not G25543;
	G26568<= not G25546;
	G26570<= not G25549;
	G26571<= not G25554;
	G26572<= not G25557;
	G26574<= not G25562;
	G26576<= not I34535;
	G26577<= not G25436;
	G26578<= not G25573;
	G26579<= not G25576;
	G26580<= not G25579;
	G26581<= not G25582;
	G26582<= not G25585;
	G26584<= not G25590;
	G26585<= not G25593;
	G26586<= not G25596;
	G26587<= not G25599;
	G26588<= not G25602;
	G26589<= not G25606;
	G26590<= not G25609;
	G26591<= not G25612;
	G26593<= not G25615;
	G26594<= not G25620;
	G26595<= not G25623;
	G26597<= not G25443;
	G26598<= not G25634;
	G26599<= not G25637;
	G26600<= not G25640;
	G26601<= not G25643;
	G26602<= not G25652;
	G26603<= not G25655;
	G26604<= not G25658;
	G26605<= not G25661;
	G26606<= not G25664;
	G26608<= not G25669;
	G26609<= not G25672;
	G26610<= not G25675;
	G26611<= not G25678;
	G26612<= not G25681;
	G26613<= not G25685;
	G26614<= not G25688;
	G26615<= not G25691;
	G26617<= not G25694;
	G26618<= not I34579;
	G26619<= not G25700;
	G26620<= not G25703;
	G26621<= not G25711;
	G26622<= not G25714;
	G26623<= not G25717;
	G26624<= not G25720;
	G26625<= not G25729;
	G26626<= not G25732;
	G26627<= not G25735;
	G26628<= not G25738;
	G26629<= not G25741;
	G26631<= not G25746;
	G26632<= not G25749;
	G26633<= not G25752;
	G26634<= not G25755;
	G26635<= not G25758;
	G26636<= not G25767;
	G26637<= not G25773;
	G26638<= not G25776;
	G26639<= not G25784;
	G26640<= not G25787;
	G26641<= not G25790;
	G26642<= not G25793;
	G26643<= not G25802;
	G26644<= not G25805;
	G26645<= not G25808;
	G26646<= not G25811;
	G26647<= not G25814;
	G26648<= not G25821;
	G26649<= not G25827;
	G26650<= not G25830;
	G26651<= not G25838;
	G26652<= not G25841;
	G26653<= not G25844;
	G26654<= not G25847;
	G26656<= not G25856;
	G26657<= not G25862;
	G26658<= not G25865;
	G26662<= not G25877;
	G26678<= not I34641;
	G26679<= not I34644;
	G26680<= not I34647;
	G26681<= not I34650;
	G26682<= not I34653;
	G26683<= not I34656;
	G26684<= not I34659;
	G26685<= not I34662;
	G26686<= not I34665;
	G26687<= not I34668;
	G26688<= not I34671;
	G26689<= not I34674;
	G26690<= not I34677;
	G26691<= not I34680;
	G26692<= not I34683;
	G26693<= not I34686;
	G26694<= not I34689;
	G26695<= not I34692;
	G26696<= not I34695;
	G26697<= not I34698;
	G26698<= not I34701;
	G26699<= not I34704;
	G26700<= not I34707;
	G26701<= not I34710;
	G26702<= not I34713;
	G26703<= not I34716;
	G26704<= not I34719;
	G26705<= not I34722;
	G26706<= not I34725;
	G26707<= not I34728;
	G26708<= not I34731;
	G26709<= not I34734;
	G26710<= not I34737;
	G26711<= not I34740;
	G26712<= not I34743;
	G26713<= not I34746;
	G26714<= not I34749;
	G26715<= not I34752;
	G26716<= not I34755;
	G26717<= not I34758;
	G26718<= not I34761;
	G26719<= not I34764;
	G26720<= not I34767;
	G26721<= not I34770;
	G26722<= not I34773;
	G26723<= not I34776;
	G26724<= not I34779;
	G26725<= not I34782;
	G26726<= not I34785;
	G26727<= not I34788;
	G26728<= not I34791;
	G26729<= not I34794;
	G26730<= not I34797;
	G26731<= not I34800;
	G26732<= not I34803;
	G26733<= not I34806;
	G26734<= not I34809;
	G26735<= not I34812;
	G26736<= not I34815;
	G26737<= not I34818;
	G26738<= not I34821;
	G26739<= not I34824;
	G26740<= not I34827;
	G26741<= not I34830;
	G26742<= not I34833;
	G26743<= not I34836;
	G26744<= not I34839;
	G26745<= not I34842;
	G26746<= not I34845;
	G26747<= not I34848;
	G26748<= not I34851;
	G26749<= not I34854;
	G26750<= not I34857;
	G26751<= not I34860;
	G26752<= not I34863;
	G26753<= not I34866;
	G26757<= not I34872;
	G26762<= not I34879;
	G26782<= not I34901;
	G26788<= not I34909;
	G26793<= not I34916;
	G26796<= not I34921;
	G26819<= not I34946;
	G26828<= not I34957;
	G26830<= not I34961;
	G26831<= not I34964;
	G26832<= not I34967;
	G26834<= not I34971;
	G26835<= not I34974;
	G26836<= not I34977;
	G26837<= not I34980;
	G26840<= not I34983;
	G26841<= not I34986;
	G26843<= not I34990;
	G26844<= not I34993;
	G26846<= not I34997;
	G26849<= not I35000;
	G26850<= not I35003;
	G26852<= not I35007;
	G26854<= not I35011;
	G26855<= not I35014;
	G26858<= not I35017;
	G26861<= not I35028;
	G26864<= not I35031;
	G26868<= not I35049;
	G26872<= not I35053;
	G26875<= not I35064;
	G26876<= not I35067;
	G26881<= not I35072;
	G26883<= not I35076;
	G26884<= not I35079;
	G26886<= not I35083;
	G26890<= not I35087;
	G26895<= not I35092;
	G26896<= not I35095;
	G26900<= not I35099;
	G26909<= not I35106;
	G26910<= not I35109;
	G26921<= not I35116;
	G26922<= not G26283;
	G26935<= not G26327;
	G26944<= not G26374;
	G26950<= not G26417;
	G26953<= not I35136;
	G26954<= not G26549;
	G26956<= not I35141;
	G26957<= not G26577;
	G26959<= not I35146;
	G26960<= not G26597;
	G26964<= not I35153;
	G26983<= not I35172;
	G26987<= not G26056;
	G27010<= not G26063;
	G27036<= not G26070;
	G27064<= not G26076;
	G27075<= not I35254;
	G27102<= not I35283;
	G27114<= not I35297;
	G27116<= not I35301;
	G27126<= not I35313;
	G27132<= not I35319;
	G27133<= not G26105;
	G27134<= not G26175;
	G27135<= not G26178;
	G27136<= not G26196;
	G27137<= not G26202;
	G27138<= not G26223;
	G27139<= not G26226;
	G27140<= not G26136;
	G27141<= not G26251;
	G27142<= not G26254;
	G27143<= not G26150;
	G27145<= not I35334;
	G27146<= not G26358;
	G27148<= not G26393;
	G27150<= not I35341;
	G27151<= not G26401;
	G27153<= not G26429;
	G27154<= not I35347;
	G27155<= not G26434;
	G27156<= not I35351;
	G27158<= not I35355;
	G27159<= not G26442;
	G27161<= not I35360;
	G27162<= not G26461;
	G27163<= not I35364;
	G27164<= not G26466;
	G27166<= not I35369;
	G27167<= not G26474;
	G27168<= not I35373;
	G27171<= not I35376;
	G27172<= not G26485;
	G27173<= not G26490;
	G27176<= not I35383;
	G27177<= not G26501;
	G27180<= not I35389;
	G27183<= not I35394;
	G27186<= not I35399;
	G27189<= not I35404;
	G27190<= not I35407;
	G27191<= not I35410;
	G27192<= not I35413;
	G27193<= not I35416;
	G27194<= not I35419;
	G27195<= not I35422;
	G27196<= not I35425;
	G27197<= not I35428;
	G27198<= not I35431;
	G27199<= not I35434;
	G27200<= not I35437;
	G27201<= not I35440;
	G27202<= not I35443;
	G27203<= not I35446;
	G27204<= not I35449;
	G27205<= not I35452;
	G27206<= not I35455;
	G27207<= not I35458;
	G27208<= not I35461;
	G27209<= not I35464;
	G27210<= not I35467;
	G27211<= not I35470;
	G27212<= not I35473;
	G27213<= not I35476;
	G27214<= not I35479;
	G27215<= not I35482;
	G27216<= not I35485;
	G27217<= not I35488;
	G27218<= not I35491;
	G27219<= not I35494;
	G27220<= not I35497;
	G27221<= not I35500;
	G27222<= not I35503;
	G27223<= not I35506;
	G27224<= not I35509;
	G27225<= not I35512;
	G27226<= not I35515;
	G27227<= not I35518;
	G27228<= not I35521;
	G27229<= not I35524;
	G27230<= not I35527;
	G27231<= not I35530;
	G27232<= not I35533;
	G27233<= not I35536;
	G27234<= not I35539;
	G27235<= not I35542;
	G27236<= not I35545;
	G27237<= not I35548;
	G27238<= not I35551;
	G27239<= not I35554;
	G27349<= not G27126;
	G27353<= not I35667;
	G27357<= not I35673;
	G27360<= not I35678;
	G27361<= not I35681;
	G27366<= not I35686;
	G27367<= not I35689;
	G27373<= not I35695;
	G27376<= not I35698;
	G27380<= not I35708;
	G27381<= not I35711;
	G27383<= not G27133;
	G27384<= not G27140;
	G27385<= not I35723;
	G27386<= not G27143;
	G27387<= not I35727;
	G27391<= not I35731;
	G27397<= not I35737;
	G27401<= not I35741;
	G27404<= not I35744;
	G27410<= not I35750;
	G27416<= not I35756;
	G27419<= not I35759;
	G27422<= not I35762;
	G27428<= not I35768;
	G27432<= not I35772;
	G27437<= not I35777;
	G27440<= not I35780;
	G27443<= not I35783;
	G27449<= not G26837;
	G27451<= not I35791;
	G27456<= not I35796;
	G27459<= not I35799;
	G27463<= not I35803;
	G27465<= not G26846;
	G27467<= not I35809;
	G27472<= not I35814;
	G27475<= not I35817;
	G27479<= not I35821;
	G27480<= not I35824;
	G27483<= not I35829;
	G27484<= not G26855;
	G27486<= not I35834;
	G27489<= not I35837;
	G27493<= not I35841;
	G27494<= not I35844;
	G27497<= not I35849;
	G27498<= not I35852;
	G27502<= not I35856;
	G27503<= not I35859;
	G27505<= not I35863;
	G27506<= not G26861;
	G27508<= not I35868;
	G27510<= not I35872;
	G27514<= not I35876;
	G27515<= not I35879;
	G27517<= not I35883;
	G27518<= not I35886;
	G27522<= not I35890;
	G27523<= not I35893;
	G27525<= not I35897;
	G27526<= not I35900;
	G27533<= not I35915;
	G27535<= not I35919;
	G27539<= not I35923;
	G27540<= not I35926;
	G27542<= not I35930;
	G27543<= not I35933;
	G27547<= not I35937;
	G27548<= not I35940;
	G27553<= not I35953;
	G27555<= not I35957;
	G27559<= not I35961;
	G27560<= not I35964;
	G27562<= not I35968;
	G27569<= not I35983;
	G27586<= not I36008;
	G27589<= not G27168;
	G27590<= not G27144;
	G27595<= not G27149;
	G27599<= not G27147;
	G27604<= not G27157;
	G27608<= not G27152;
	G27613<= not G27165;
	G27617<= not G27160;
	G27622<= not G27174;
	G27632<= not I36032;
	G27662<= not I36042;
	G27667<= not I36046;
	G27674<= not I36052;
	G27683<= not I36060;
	G27684<= not I36063;
	G27685<= not I36066;
	G27686<= not I36069;
	G27687<= not I36072;
	G27688<= not I36075;
	G27689<= not I36078;
	G27690<= not I36081;
	G27691<= not I36084;
	G27692<= not I36087;
	G27693<= not I36090;
	G27694<= not I36093;
	G27695<= not I36096;
	G27696<= not I36099;
	G27697<= not I36102;
	G27698<= not I36105;
	G27699<= not I36108;
	G27700<= not I36111;
	G27701<= not I36114;
	G27702<= not I36117;
	G27703<= not I36120;
	G27704<= not I36123;
	G27705<= not I36126;
	G27706<= not I36129;
	G27707<= not I36132;
	G27708<= not I36135;
	G27709<= not I36138;
	G27710<= not I36141;
	G27711<= not I36144;
	G27712<= not I36147;
	G27713<= not I36150;
	G27714<= not I36153;
	G27715<= not I36156;
	G27716<= not I36159;
	G27717<= not I36162;
	G27748<= not G27632;
	G27776<= not I36213;
	G27780<= not I36217;
	G27784<= not I36221;
	G27785<= not I36224;
	G27786<= not I36227;
	G27787<= not I36230;
	G27791<= not I36234;
	G27792<= not I36237;
	G27793<= not I36240;
	G27794<= not I36243;
	G27797<= not I36246;
	G27799<= not I36250;
	G27800<= not I36253;
	G27805<= not I36264;
	G27806<= not I36267;
	G27817<= not I36280;
	G27820<= not I36283;
	G27831<= not I36296;
	G27839<= not I36307;
	G27843<= not I36311;
	G27847<= not I36321;
	G27858<= not I36327;
	G27861<= not I36330;
	G27872<= not I36337;
	G27879<= not I36341;
	G27889<= not I36347;
	G27903<= not I36354;
	G27905<= not I36358;
	G27907<= not I36362;
	G27910<= not I36367;
	G27912<= not I36371;
	G27918<= not I36379;
	G27919<= not I36382;
	G27927<= not I36390;
	G27928<= not I36393;
	G27932<= not I36397;
	G27939<= not I36404;
	G27942<= not I36407;
	G27946<= not I36411;
	G27952<= not I36417;
	G27955<= not I36420;
	G27956<= not I36423;
	G27959<= not I36426;
	G27965<= not I36432;
	G27969<= not G27361;
	G27971<= not I36438;
	G27972<= not I36441;
	G27973<= not I36444;
	G27976<= not I36447;
	G27977<= not I36450;
	G27981<= not I36454;
	G27986<= not I36459;
	G27987<= not I36462;
	G27988<= not I36465;
	G27989<= not I36468;
	G27990<= not G27367;
	G27992<= not I36473;
	G27993<= not I36476;
	G27994<= not I36479;
	G27998<= not I36483;
	G27999<= not I36486;
	G28003<= not I36490;
	G28004<= not I36493;
	G28005<= not I36496;
	G28006<= not I36499;
	G28007<= not I36502;
	G28010<= not I36507;
	G28011<= not I36510;
	G28012<= not I36513;
	G28013<= not I36516;
	G28014<= not G27373;
	G28016<= not I36521;
	G28017<= not I36524;
	G28018<= not I36527;
	G28021<= not I36530;
	G28022<= not I36533;
	G28023<= not I36536;
	G28024<= not I36539;
	G28025<= not I36542;
	G28026<= not I36545;
	G28030<= not I36551;
	G28031<= not I36554;
	G28032<= not I36557;
	G28033<= not I36560;
	G28034<= not I36563;
	G28037<= not I36568;
	G28038<= not I36571;
	G28039<= not I36574;
	G28040<= not I36577;
	G28041<= not G27376;
	G28043<= not I36582;
	G28044<= not I36585;
	G28045<= not I36588;
	G28047<= not I36598;
	G28048<= not I36601;
	G28049<= not I36604;
	G28052<= not I36609;
	G28053<= not I36612;
	G28054<= not I36615;
	G28055<= not I36618;
	G28056<= not I36621;
	G28060<= not I36627;
	G28061<= not I36630;
	G28062<= not I36633;
	G28063<= not I36636;
	G28064<= not I36639;
	G28067<= not I36644;
	G28068<= not I36647;
	G28069<= not I36650;
	G28070<= not I36653;
	G28071<= not I36656;
	G28072<= not I36659;
	G28074<= not I36663;
	G28076<= not I36673;
	G28077<= not I36676;
	G28078<= not I36679;
	G28081<= not I36684;
	G28082<= not I36687;
	G28083<= not I36690;
	G28084<= not I36693;
	G28085<= not I36696;
	G28089<= not I36702;
	G28090<= not I36705;
	G28091<= not I36708;
	G28092<= not I36711;
	G28093<= not I36714;
	G28095<= not I36718;
	G28096<= not I36721;
	G28097<= not I36724;
	G28099<= not I36728;
	G28101<= not I36738;
	G28102<= not I36741;
	G28103<= not I36744;
	G28106<= not I36749;
	G28107<= not I36752;
	G28108<= not I36755;
	G28109<= not I36758;
	G28110<= not I36761;
	G28113<= not I36766;
	G28114<= not I36769;
	G28115<= not I36772;
	G28117<= not I36776;
	G28119<= not I36786;
	G28120<= not I36789;
	G28121<= not I36792;
	G28124<= not I36797;
	G28125<= not I36800;
	G28126<= not I36803;
	G28128<= not G27528;
	G28132<= not I36808;
	G28133<= not G27550;
	G28137<= not G27566;
	G28141<= not G27576;
	G28149<= not G27667;
	G28150<= not G27387;
	G28151<= not G27381;
	G28152<= not G27391;
	G28153<= not G27397;
	G28154<= not G27401;
	G28155<= not G27404;
	G28156<= not G27410;
	G28158<= not G27416;
	G28159<= not G27419;
	G28160<= not G27422;
	G28161<= not G27428;
	G28162<= not G27432;
	G28163<= not G27437;
	G28164<= not G27440;
	G28165<= not G27443;
	G28166<= not G27451;
	G28167<= not G27456;
	G28168<= not G27459;
	G28169<= not G27467;
	G28170<= not G27472;
	G28172<= not G27475;
	G28173<= not G27486;
	G28174<= not G27489;
	G28175<= not G27498;
	G28177<= not G27510;
	G28178<= not G27518;
	G28179<= not I36848;
	G28186<= not G27535;
	G28187<= not G27543;
	G28190<= not G27555;
	G28194<= not I36860;
	G28200<= not I36864;
	G28206<= not I36867;
	G28207<= not I36870;
	G28208<= not I36873;
	G28209<= not I36876;
	G28210<= not I36879;
	G28211<= not I36882;
	G28212<= not I36885;
	G28213<= not I36888;
	G28214<= not I36891;
	G28215<= not I36894;
	G28216<= not I36897;
	G28217<= not I36900;
	G28218<= not I36903;
	G28219<= not I36906;
	G28220<= not I36909;
	G28221<= not I36912;
	G28222<= not I36915;
	G28223<= not I36918;
	G28224<= not I36921;
	G28225<= not I36924;
	G28226<= not I36927;
	G28227<= not I36930;
	G28228<= not I36933;
	G28229<= not I36936;
	G28230<= not I36939;
	G28231<= not I36942;
	G28232<= not I36945;
	G28233<= not I36948;
	G28234<= not I36951;
	G28235<= not I36954;
	G28236<= not I36957;
	G28237<= not I36960;
	G28238<= not I36963;
	G28239<= not I36966;
	G28240<= not I36969;
	G28241<= not I36972;
	G28242<= not I36975;
	G28243<= not I36978;
	G28244<= not I36981;
	G28245<= not I36984;
	G28246<= not I36987;
	G28247<= not I36990;
	G28248<= not I36993;
	G28249<= not I36996;
	G28250<= not I36999;
	G28251<= not I37002;
	G28252<= not I37005;
	G28253<= not I37008;
	G28254<= not I37011;
	G28255<= not I37014;
	G28256<= not I37017;
	G28257<= not I37020;
	G28258<= not I37023;
	G28259<= not I37026;
	G28260<= not I37029;
	G28261<= not I37032;
	G28262<= not I37035;
	G28263<= not I37038;
	G28264<= not I37041;
	G28265<= not I37044;
	G28266<= not I37047;
	G28267<= not I37050;
	G28268<= not I37053;
	G28269<= not I37056;
	G28270<= not I37059;
	G28271<= not I37062;
	G28272<= not I37065;
	G28273<= not I37068;
	G28274<= not I37071;
	G28275<= not I37074;
	G28276<= not I37077;
	G28277<= not I37080;
	G28278<= not I37083;
	G28279<= not I37086;
	G28280<= not I37089;
	G28281<= not I37092;
	G28282<= not I37095;
	G28283<= not I37098;
	G28284<= not I37101;
	G28285<= not I37104;
	G28286<= not I37107;
	G28287<= not I37110;
	G28288<= not I37113;
	G28289<= not I37116;
	G28290<= not I37119;
	G28291<= not I37122;
	G28292<= not I37125;
	G28293<= not I37128;
	G28294<= not I37131;
	G28295<= not I37134;
	G28296<= not I37137;
	G28297<= not I37140;
	G28298<= not I37143;
	G28299<= not I37146;
	G28300<= not I37149;
	G28301<= not I37152;
	G28302<= not I37155;
	G28303<= not I37158;
	G28304<= not I37161;
	G28305<= not I37164;
	G28306<= not I37167;
	G28307<= not I37170;
	G28308<= not I37173;
	G28309<= not I37176;
	G28310<= not I37179;
	G28311<= not I37182;
	G28312<= not I37185;
	G28313<= not I37188;
	G28314<= not I37191;
	G28315<= not I37194;
	G28316<= not I37197;
	G28317<= not I37200;
	G28318<= not I37203;
	G28341<= not I37228;
	G28343<= not I37232;
	G28347<= not I37238;
	G28359<= not I37252;
	G28365<= not I37260;
	G28369<= not I37266;
	G28370<= not I37269;
	G28372<= not I37273;
	G28374<= not I37277;
	G28375<= not I37280;
	G28377<= not I37284;
	G28382<= not I37291;
	G28390<= not I37319;
	G28393<= not I37330;
	G28395<= not I37334;
	G28419<= not G28151;
	G28432<= not I37379;
	G28437<= not I37386;
	G28443<= not I37394;
	G28447<= not I37400;
	G28455<= not I37410;
	G28458<= not I37415;
	G28467<= not I37426;
	G28483<= not G27776;
	G28491<= not G27780;
	G28496<= not G27787;
	G28498<= not I37459;
	G28500<= not G27794;
	G28524<= not I37467;
	G28526<= not I37471;
	G28527<= not I37474;
	G28552<= not I37481;
	G28553<= not I37484;
	G28554<= not G27806;
	G28555<= not I37488;
	G28579<= not I37494;
	G28580<= not I37497;
	G28581<= not G27817;
	G28582<= not G27820;
	G28583<= not I37502;
	G28607<= not I37508;
	G28608<= not G27831;
	G28609<= not G27839;
	G28610<= not G27843;
	G28611<= not I37514;
	G28612<= not G28046;
	G28616<= not G27847;
	G28617<= not G27858;
	G28618<= not G27861;
	G28619<= not G28075;
	G28623<= not G27872;
	G28624<= not G27879;
	G28625<= not G28100;
	G28629<= not G27889;
	G28630<= not G28118;
	G28638<= not G28200;
	G28639<= not G27919;
	G28640<= not G27928;
	G28641<= not G27932;
	G28642<= not G27939;
	G28643<= not G27942;
	G28644<= not G27946;
	G28645<= not G27952;
	G28646<= not G27956;
	G28647<= not G27959;
	G28648<= not G27965;
	G28649<= not G27973;
	G28650<= not G27977;
	G28651<= not G27981;
	G28652<= not G27994;
	G28653<= not G27999;
	G28655<= not G28018;
	G28673<= not I37566;
	G28674<= not I37569;
	G28675<= not I37572;
	G28676<= not I37575;
	G28677<= not I37578;
	G28678<= not I37581;
	G28679<= not I37584;
	G28680<= not I37587;
	G28681<= not I37590;
	G28682<= not I37593;
	G28683<= not I37596;
	G28684<= not I37599;
	G28685<= not I37602;
	G28686<= not I37605;
	G28687<= not I37608;
	G28688<= not I37611;
	G28689<= not I37614;
	G28690<= not I37617;
	G28691<= not I37620;
	G28692<= not I37623;
	G28693<= not I37626;
	G28694<= not I37629;
	G28695<= not I37632;
	G28696<= not I37635;
	G28697<= not I37638;
	G28698<= not I37641;
	G28699<= not I37644;
	G28700<= not I37647;
	G28701<= not I37650;
	G28702<= not I37653;
	G28703<= not I37656;
	G28704<= not I37659;
	G28705<= not I37662;
	G28706<= not I37665;
	G28720<= not G28495;
	G28721<= not G28490;
	G28723<= not G28528;
	G28725<= not G28499;
	G28727<= not G28489;
	G28730<= not G28470;
	G28734<= not G28525;
	G28740<= not G28488;
	G28741<= not I37702;
	G28751<= not I37712;
	G28755<= not I37716;
	G28764<= not I37725;
	G28768<= not I37729;
	G28775<= not I37736;
	G28779<= not I37740;
	G28785<= not I37746;
	G28791<= not I37752;
	G28796<= not I37757;
	G28799<= not I37760;
	G28804<= not I37765;
	G28807<= not I37768;
	G28810<= not I37771;
	G28814<= not I37775;
	G28817<= not I37778;
	G28820<= not I37781;
	G28823<= not I37784;
	G28826<= not I37787;
	G28829<= not I37790;
	G28832<= not I37793;
	G28833<= not I37796;
	G28835<= not I37800;
	G28837<= not I37804;
	G28839<= not I37808;
	G28855<= not G28409;
	G28859<= not G28413;
	G28863<= not G28417;
	G28867<= not G28418;
	G28871<= not I37842;
	G28877<= not I37846;
	G28882<= not I37851;
	G28883<= not I37854;
	G28889<= not I37858;
	G28894<= not I37863;
	G28899<= not I37868;
	G28900<= not I37871;
	G28906<= not I37875;
	G28911<= not I37880;
	G28916<= not I37885;
	G28924<= not I37891;
	G28925<= not I37894;
	G28928<= not I37897;
	G28932<= not I37901;
	G28937<= not I37906;
	G28945<= not I37912;
	G28950<= not I37917;
	G28951<= not I37920;
	G28955<= not I37924;
	G28959<= not I37928;
	G28967<= not I37934;
	G28972<= not I37939;
	G28975<= not I37942;
	G28979<= not I37946;
	G28983<= not I37950;
	G28993<= not I37956;
	G28998<= not I37961;
	G29002<= not I37965;
	G29005<= not I37968;
	G29010<= not I37973;
	G29019<= not I37978;
	G29023<= not I37982;
	G29027<= not I37986;
	G29032<= not I37991;
	G29035<= not I37994;
	G29042<= not I37999;
	G29046<= not I38003;
	G29050<= not I38007;
	G29054<= not I38011;
	G29057<= not I38014;
	G29061<= not I38018;
	G29065<= not I38024;
	G29069<= not I38028;
	G29073<= not I38032;
	G29074<= not I38035;
	G29075<= not I38038;
	G29077<= not I38042;
	G29081<= not I38046;
	G29082<= not I38049;
	G29084<= not I38053;
	G29085<= not I38056;
	G29086<= not I38059;
	G29089<= not I38064;
	G29091<= not I38068;
	G29092<= not I38071;
	G29093<= not I38074;
	G29094<= not I38077;
	G29095<= not I38080;
	G29098<= not I38085;
	G29099<= not I38088;
	G29100<= not I38091;
	G29101<= not I38094;
	G29102<= not I38097;
	G29104<= not I38101;
	G29105<= not I38104;
	G29106<= not I38107;
	G29108<= not I38111;
	G29117<= not I38119;
	G29118<= not I38122;
	G29119<= not I38125;
	G29120<= not I38128;
	G29131<= not I38136;
	G29132<= not I38139;
	G29133<= not I38142;
	G29134<= not I38145;
	G29135<= not I38148;
	G29136<= not I38151;
	G29137<= not I38154;
	G29138<= not I38157;
	G29139<= not I38160;
	G29140<= not I38163;
	G29141<= not I38166;
	G29142<= not I38169;
	G29143<= not I38172;
	G29144<= not I38175;
	G29145<= not I38178;
	G29146<= not I38181;
	G29147<= not I38184;
	G29148<= not I38187;
	G29149<= not I38190;
	G29150<= not I38193;
	G29151<= not I38196;
	G29152<= not I38199;
	G29153<= not I38202;
	G29154<= not I38205;
	G29155<= not I38208;
	G29156<= not I38211;
	G29157<= not I38214;
	G29158<= not I38217;
	G29159<= not I38220;
	G29160<= not I38223;
	G29161<= not I38226;
	G29162<= not I38229;
	G29163<= not I38232;
	G29164<= not I38235;
	G29165<= not I38238;
	G29166<= not I38241;
	G29168<= not I38245;
	G29171<= not I38250;
	G29177<= not I38258;
	G29189<= not I38272;
	G29190<= not I38275;
	G29191<= not I38278;
	G29192<= not G28954;
	G29193<= not I38282;
	G29230<= not I38321;
	G29237<= not I38330;
	G29244<= not I38339;
	G29245<= not I38342;
	G29246<= not I38345;
	G29247<= not I38348;
	G29249<= not I38352;
	G29250<= not I38355;
	G29253<= not I38360;
	G29254<= not I38363;
	G29258<= not I38369;
	G29266<= not G28741;
	G29267<= not I38386;
	G29268<= not G28751;
	G29269<= not G28755;
	G29270<= not I38391;
	G29271<= not G28764;
	G29272<= not G28768;
	G29273<= not I38396;
	G29274<= not G28775;
	G29275<= not G28779;
	G29276<= not I38401;
	G29277<= not G28785;
	G29278<= not I38405;
	G29279<= not I38408;
	G29280<= not G28791;
	G29281<= not I38412;
	G29282<= not G28796;
	G29283<= not G28799;
	G29285<= not G28804;
	G29286<= not G28807;
	G29287<= not G28810;
	G29288<= not I38421;
	G29290<= not G28814;
	G29291<= not G28817;
	G29292<= not G28820;
	G29293<= not I38428;
	G29295<= not G28823;
	G29296<= not G28826;
	G29297<= not I38434;
	G29298<= not I38437;
	G29299<= not I38440;
	G29301<= not G28829;
	G29304<= not I38447;
	G29305<= not I38450;
	G29306<= not I38453;
	G29307<= not I38456;
	G29308<= not I38459;
	G29309<= not I38462;
	G29311<= not I38466;
	G29314<= not I38471;
	G29315<= not I38474;
	G29316<= not I38477;
	G29317<= not I38480;
	G29318<= not I38483;
	G29319<= not I38486;
	G29322<= not I38491;
	G29325<= not I38496;
	G29326<= not I38499;
	G29327<= not I38502;
	G29328<= not I38505;
	G29331<= not I38510;
	G29334<= not I38515;
	G29335<= not I38518;
	G29339<= not I38524;
	G29349<= not I38536;
	G29350<= not I38539;
	G29356<= not G29120;
	G29358<= not G29120;
	G29359<= not I38548;
	G29360<= not G28871;
	G29361<= not G28877;
	G29362<= not G28883;
	G29363<= not G28889;
	G29364<= not G28894;
	G29365<= not G28900;
	G29366<= not G28906;
	G29367<= not G28911;
	G29368<= not G28916;
	G29369<= not G28925;
	G29370<= not G28928;
	G29371<= not G28932;
	G29372<= not G28937;
	G29373<= not G28945;
	G29374<= not G28951;
	G29375<= not G28955;
	G29376<= not G28959;
	G29377<= not G28967;
	G29378<= not G28972;
	G29379<= not G28975;
	G29380<= not G28979;
	G29381<= not G28983;
	G29382<= not G28993;
	G29383<= not G28998;
	G29384<= not G29002;
	G29385<= not G29005;
	G29386<= not G29010;
	G29387<= not G29019;
	G29388<= not G29023;
	G29389<= not G29027;
	G29390<= not G29032;
	G29391<= not G29035;
	G29392<= not G29042;
	G29393<= not G29046;
	G29394<= not G29050;
	G29395<= not G29054;
	G29396<= not G29057;
	G29397<= not G29065;
	G29398<= not G29069;
	G29400<= not I38591;
	G29401<= not I38594;
	G29402<= not G29077;
	G29404<= not I38599;
	G29405<= not I38602;
	G29407<= not I38606;
	G29408<= not I38609;
	G29410<= not I38613;
	G29412<= not I38617;
	G29413<= not I38620;
	G29414<= not I38623;
	G29415<= not I38626;
	G29416<= not I38629;
	G29417<= not I38632;
	G29418<= not I38635;
	G29419<= not I38638;
	G29420<= not I38641;
	G29421<= not I38644;
	G29422<= not I38647;
	G29423<= not I38650;
	G29424<= not I38653;
	G29425<= not I38656;
	G29426<= not I38659;
	G29427<= not I38662;
	G29428<= not I38665;
	G29429<= not I38668;
	G29430<= not I38671;
	G29431<= not I38674;
	G29432<= not I38677;
	G29433<= not I38680;
	G29434<= not I38683;
	G29435<= not I38686;
	G29436<= not I38689;
	G29437<= not I38692;
	G29438<= not I38695;
	G29439<= not I38698;
	G29440<= not I38701;
	G29441<= not I38704;
	G29442<= not I38707;
	G29443<= not I38710;
	G29444<= not I38713;
	G29445<= not I38716;
	G29446<= not I38719;
	G29447<= not I38722;
	G29448<= not I38725;
	G29449<= not I38728;
	G29450<= not I38731;
	G29451<= not I38734;
	G29452<= not I38737;
	G29453<= not I38740;
	G29454<= not I38743;
	G29455<= not I38746;
	G29456<= not I38749;
	G29457<= not I38752;
	G29458<= not I38755;
	G29459<= not I38758;
	G29460<= not I38761;
	G29461<= not I38764;
	G29462<= not I38767;
	G29463<= not I38770;
	G29491<= not G29350;
	G29495<= not I38801;
	G29496<= not I38804;
	G29497<= not I38807;
	G29499<= not I38817;
	G29501<= not I38827;
	G29504<= not I38838;
	G29506<= not I38848;
	G29507<= not I38851;
	G29508<= not I38854;
	G29509<= not I38857;
	G29510<= not I38860;
	G29511<= not I38863;
	G29512<= not I38866;
	G29513<= not I38869;
	G29514<= not I38872;
	G29515<= not I38875;
	G29516<= not I38878;
	G29517<= not I38881;
	G29519<= not I38885;
	G29530<= not I38898;
	G29535<= not I38905;
	G29537<= not I38909;
	G29542<= not I38916;
	G29544<= not I38920;
	G29546<= not I38924;
	G29551<= not I38931;
	G29554<= not I38936;
	G29556<= not I38940;
	G29561<= not I38947;
	G29563<= not I38951;
	G29568<= not I38958;
	G29583<= not I38975;
	G29627<= not I38999;
	G29628<= not I39002;
	G29629<= not I39005;
	G29630<= not I39008;
	G29631<= not I39011;
	G29632<= not I39014;
	G29633<= not I39017;
	G29634<= not I39020;
	G29635<= not I39023;
	G29636<= not I39026;
	G29637<= not I39029;
	G29638<= not I39032;
	G29639<= not I39035;
	G29640<= not I39038;
	G29641<= not I39041;
	G29642<= not I39044;
	G29643<= not I39047;
	G29644<= not I39050;
	G29645<= not I39053;
	G29646<= not I39056;
	G29647<= not I39059;
	G29648<= not I39062;
	G29649<= not I39065;
	G29650<= not I39068;
	G29651<= not I39071;
	G29652<= not I39074;
	G29653<= not I39077;
	G29654<= not I39080;
	G29655<= not I39083;
	G29656<= not I39086;
	G29657<= not I39089;
	G29658<= not G29574;
	G29659<= not G29571;
	G29660<= not G29578;
	G29661<= not G29576;
	G29662<= not G29570;
	G29664<= not G29552;
	G29666<= not G29577;
	G29668<= not G29569;
	G29673<= not G29583;
	G29689<= not I39121;
	G29690<= not I39124;
	G29691<= not I39127;
	G29692<= not I39130;
	G29693<= not I39133;
	G29694<= not I39136;
	G29695<= not I39139;
	G29696<= not I39142;
	G29697<= not I39145;
	G29698<= not I39148;
	G29699<= not I39151;
	G29700<= not I39154;
	G29701<= not I39157;
	G29702<= not I39160;
	G29704<= not I39164;
	G29708<= not I39168;
	G29716<= not G29498;
	G29724<= not G29500;
	G29726<= not G29503;
	G29739<= not G29505;
	G29794<= not I39234;
	G29795<= not I39237;
	G29796<= not I39240;
	G29797<= not I39243;
	G29798<= not I39246;
	G29799<= not I39249;
	G29800<= not I39252;
	G29801<= not I39255;
	G29802<= not I39258;
	G29803<= not I39261;
	G29804<= not I39264;
	G29805<= not I39267;
	G29806<= not I39270;
	G29807<= not I39273;
	G29808<= not I39276;
	G29809<= not I39279;
	G29823<= not G29663;
	G29829<= not G29665;
	G29835<= not G29667;
	G29840<= not G29669;
	G29844<= not G29670;
	G29848<= not G29761;
	G29849<= not G29671;
	G29853<= not G29672;
	G29857<= not G29676;
	G29861<= not G29677;
	G29865<= not G29678;
	G29869<= not G29679;
	G29873<= not G29680;
	G29877<= not G29681;
	G29881<= not G29682;
	G29885<= not G29683;
	G29889<= not G29684;
	G29893<= not G29685;
	G29897<= not G29686;
	G29901<= not G29687;
	G29905<= not G29688;
	G29932<= not I39398;
	G29933<= not I39401;
	G29934<= not I39404;
	G29935<= not I39407;
	G29937<= not I39411;
	G29938<= not I39414;
	G29940<= not I39418;
	G29943<= not I39423;
	G29972<= not I39454;
	G29973<= not I39457;
	G29974<= not I39460;
	G29975<= not I39463;
	G29976<= not I39466;
	G29977<= not I39469;
	G29978<= not I39472;
	G29979<= not I39475;
	G30036<= not G29912;
	G30040<= not G29914;
	G30044<= not G29916;
	G30048<= not G29920;
	G30052<= not I39550;
	G30076<= not I39573;
	G30078<= not I39577;
	G30084<= not I39585;
	G30119<= not I39622;
	G30120<= not I39625;
	G30121<= not I39628;
	G30122<= not I39631;
	G30124<= not I39635;
	G30125<= not I39638;
	G30126<= not I39641;
	G30130<= not I39647;
	G30134<= not G30010;
	G30139<= not G30011;
	G30143<= not G30012;
	G30147<= not G30013;
	G30151<= not G30014;
	G30155<= not G30015;
	G30159<= not G30016;
	G30163<= not G30017;
	G30167<= not G30018;
	G30171<= not G30019;
	G30175<= not G30020;
	G30179<= not G30021;
	G30183<= not G30022;
	G30187<= not G30023;
	G30191<= not G30024;
	G30195<= not G30025;
	G30199<= not G30026;
	G30203<= not G30027;
	G30207<= not G30028;
	G30211<= not G30029;
	G30215<= not I39674;
	G30229<= not G30030;
	G30233<= not G30031;
	G30237<= not G30032;
	G30241<= not G30033;
	G30306<= not I39761;
	G30307<= not I39764;
	G30308<= not I39767;
	G30309<= not I39770;
	G30310<= not I39773;
	G30311<= not I39776;
	G30312<= not I39779;
	G30313<= not I39782;
	G30314<= not I39785;
	G30315<= not I39788;
	G30316<= not I39791;
	G30317<= not I39794;
	G30318<= not I39797;
	G30319<= not I39800;
	G30320<= not I39803;
	G30321<= not I39806;
	G30322<= not I39809;
	G30323<= not I39812;
	G30324<= not I39815;
	G30325<= not I39818;
	G30326<= not I39821;
	G30328<= not I39825;
	G30329<= not I39828;
	G30331<= not I39832;
	G30332<= not I39835;
	G30335<= not I39840;
	G30336<= not I39843;
	G30339<= not I39848;
	G30342<= not I39853;
	G30343<= not I39856;
	G30344<= not I39859;
	G30346<= not I39863;
	G30347<= not I39866;
	G30349<= not I39870;
	G30350<= not I39873;
	G30353<= not I39878;
	G30354<= not I39881;
	G30357<= not I39886;
	G30358<= not I39889;
	G30359<= not I39892;
	G30360<= not I39895;
	G30362<= not I39899;
	G30363<= not I39902;
	G30365<= not I39906;
	G30366<= not I39909;
	G30368<= not I39913;
	G30369<= not I39916;
	G30370<= not I39919;
	G30371<= not I39922;
	G30373<= not I39926;
	G30375<= not I39930;
	G30376<= not I39933;
	G30377<= not I39936;
	G30378<= not I39939;
	G30379<= not I39942;
	G30380<= not I39945;
	G30381<= not I39948;
	G30382<= not I39951;
	G30383<= not G30306;
	G30408<= not I39976;
	G30412<= not I39982;
	G30435<= not I39985;
	G30439<= not I39991;
	G30443<= not I39997;
	G30446<= not I40002;
	G30450<= not I40008;
	G30456<= not I40016;
	G30459<= not I40021;
	G30463<= not I40027;
	G30466<= not I40032;
	G30471<= not I40039;
	G30474<= not I40044;
	G30479<= not I40051;
	G30480<= not I40054;
	G30483<= not I40059;
	G30488<= not I40066;
	G30491<= not I40071;
	G30493<= not I40075;
	G30494<= not I40078;
	G30497<= not I40083;
	G30498<= not I40086;
	G30501<= not I40091;
	G30506<= not I40098;
	G30507<= not I40101;
	G30508<= not I40104;
	G30509<= not I40107;
	G30510<= not I40110;
	G30511<= not I40113;
	G30512<= not I40116;
	G30513<= not I40119;
	G30514<= not I40122;
	G30515<= not I40125;
	G30516<= not I40128;
	G30517<= not I40131;
	G30518<= not I40134;
	G30519<= not I40137;
	G30520<= not I40140;
	G30521<= not I40143;
	G30522<= not I40146;
	G30523<= not I40149;
	G30524<= not I40152;
	G30525<= not I40155;
	G30526<= not I40158;
	G30527<= not I40161;
	G30528<= not I40164;
	G30529<= not I40167;
	G30530<= not I40170;
	G30531<= not I40173;
	G30532<= not I40176;
	G30533<= not I40179;
	G30534<= not I40182;
	G30535<= not I40185;
	G30536<= not I40188;
	G30537<= not I40191;
	G30538<= not I40194;
	G30539<= not I40197;
	G30540<= not I40200;
	G30541<= not I40203;
	G30542<= not I40206;
	G30543<= not I40209;
	G30544<= not I40212;
	G30545<= not I40215;
	G30546<= not I40218;
	G30547<= not I40221;
	G30548<= not I40224;
	G30549<= not I40227;
	G30550<= not I40230;
	G30551<= not I40233;
	G30552<= not I40236;
	G30553<= not I40239;
	G30554<= not I40242;
	G30555<= not I40245;
	G30556<= not I40248;
	G30557<= not I40251;
	G30558<= not I40254;
	G30559<= not I40257;
	G30560<= not I40260;
	G30561<= not I40263;
	G30562<= not I40266;
	G30563<= not I40269;
	G30564<= not I40272;
	G30565<= not I40275;
	G30567<= not G30403;
	G30568<= not G30402;
	G30569<= not G30406;
	G30570<= not G30404;
	G30571<= not G30401;
	G30572<= not G30399;
	G30573<= not G30405;
	G30574<= not G30400;
	G30575<= not G30412;
	G30578<= not I40288;
	G30579<= not I40291;
	G30580<= not I40294;
	G30581<= not I40297;
	G30582<= not I40300;
	G30583<= not I40303;
	G30585<= not I40307;
	G30586<= not I40310;
	G30587<= not I40313;
	G30591<= not I40317;
	G30592<= not I40320;
	G30600<= not I40326;
	G30710<= not I40420;
	G30711<= not I40423;
	G30712<= not I40426;
	G30713<= not I40429;
	G30714<= not I40432;
	G30715<= not I40435;
	G30716<= not I40438;
	G30717<= not I40441;
	G30718<= not I40444;
	G30719<= not I40447;
	G30720<= not I40450;
	G30721<= not I40453;
	G30722<= not I40456;
	G30723<= not I40459;
	G30724<= not I40462;
	G30725<= not I40465;
	G30726<= not I40468;
	G30727<= not I40471;
	G30729<= not I40475;
	G30730<= not I40478;
	G30731<= not I40481;
	G30732<= not I40484;
	G30733<= not I40487;
	G30734<= not I40490;
	G30737<= not I40495;
	G30738<= not I40498;
	G30739<= not I40501;
	G30740<= not I40504;
	G30741<= not I40507;
	G30742<= not I40510;
	G30745<= not I40515;
	G30746<= not I40518;
	G30747<= not I40521;
	G30748<= not I40524;
	G30749<= not I40527;
	G30751<= not I40531;
	G30752<= not I40534;
	G30753<= not I40537;
	G30756<= not I40542;
	G30765<= not G30685;
	G30767<= not I40555;
	G30769<= not I40565;
	G30770<= not I40568;
	G30772<= not I40578;
	G30773<= not I40581;
	G30774<= not I40584;
	G30776<= not I40594;
	G30777<= not I40597;
	G30778<= not I40600;
	G30781<= not I40611;
	G30782<= not I40614;
	G30784<= not I40618;
	G30792<= not I40634;
	G30793<= not I40637;
	G30794<= not I40640;
	G30795<= not I40643;
	G30797<= not I40647;
	G30799<= not I40651;
	G30800<= not I40654;
	G30802<= not I40658;
	G30803<= not I40661;
	G30804<= not I40664;
	G30805<= not I40667;
	G30806<= not I40670;
	G30807<= not I40673;
	G30808<= not I40676;
	G30809<= not I40679;
	G30810<= not I40682;
	G30811<= not I40685;
	G30812<= not I40688;
	G30813<= not I40691;
	G30814<= not I40694;
	G30815<= not I40697;
	G30816<= not I40700;
	G30817<= not I40703;
	G30818<= not I40706;
	G30819<= not I40709;
	G30820<= not I40712;
	G30821<= not I40715;
	G30822<= not I40718;
	G30823<= not I40721;
	G30824<= not I40724;
	G30825<= not I40727;
	G30826<= not I40730;
	G30827<= not I40733;
	G30828<= not I40736;
	G30829<= not I40739;
	G30830<= not I40742;
	G30831<= not I40745;
	G30832<= not I40748;
	G30833<= not I40751;
	G30834<= not I40754;
	G30835<= not I40757;
	G30836<= not I40760;
	G30837<= not I40763;
	G30838<= not I40766;
	G30839<= not I40769;
	G30840<= not I40772;
	G30841<= not I40775;
	G30842<= not I40778;
	G30843<= not I40781;
	G30844<= not I40784;
	G30845<= not I40787;
	G30846<= not I40790;
	G30847<= not I40793;
	G30848<= not I40796;
	G30849<= not I40799;
	G30850<= not I40802;
	G30851<= not I40805;
	G30852<= not I40808;
	G30853<= not I40811;
	G30854<= not I40814;
	G30855<= not I40817;
	G30856<= not I40820;
	G30857<= not I40823;
	G30858<= not I40826;
	G30859<= not I40829;
	G30860<= not I40832;
	G30861<= not I40835;
	G30862<= not I40838;
	G30863<= not I40841;
	G30864<= not I40844;
	G30865<= not I40847;
	G30866<= not I40850;
	G30867<= not I40853;
	G30868<= not I40856;
	G30869<= not I40859;
	G30870<= not I40862;
	G30871<= not I40865;
	G30872<= not I40868;
	G30873<= not I40871;
	G30874<= not I40874;
	G30875<= not I40877;
	G30876<= not I40880;
	G30877<= not I40883;
	G30878<= not I40886;
	G30879<= not I40889;
	G30880<= not I40892;
	G30881<= not I40895;
	G30882<= not I40898;
	G30883<= not I40901;
	G30884<= not I40904;
	G30885<= not I40907;
	G30886<= not I40910;
	G30887<= not I40913;
	G30888<= not I40916;
	G30889<= not I40919;
	G30890<= not I40922;
	G30891<= not I40925;
	G30892<= not I40928;
	G30893<= not I40931;
	G30894<= not I40934;
	G30895<= not I40937;
	G30896<= not I40940;
	G30897<= not I40943;
	G30898<= not I40946;
	G30899<= not I40949;
	G30900<= not I40952;
	G30901<= not I40955;
	G30902<= not I40958;
	G30903<= not I40961;
	G30904<= not I40964;
	G30905<= not I40967;
	G30906<= not I40970;
	G30907<= not I40973;
	G30908<= not I40976;
	G30909<= not I40979;
	G30910<= not I40982;
	G30911<= not I40985;
	G30912<= not I40988;
	G30913<= not I40991;
	G30914<= not I40994;
	G30915<= not I40997;
	G30928<= not I41024;
	G30937<= not I41035;
	G30938<= not I41038;
	G30939<= not I41041;
	G30940<= not I41044;
	G30941<= not I41047;
	G30942<= not I41050;
	G30943<= not I41053;
	G30962<= not G30958;
	G30963<= not G30957;
	G30964<= not G30961;
	G30965<= not G30959;
	G30966<= not G30956;
	G30967<= not G30954;
	G30968<= not G30960;
	G30969<= not G30955;
	G30971<= not G30970;
	G30972<= not I41090;
	G30973<= not I41093;
	G30974<= not I41096;
	G30975<= not I41099;
	G30976<= not I41102;
	G30977<= not I41105;
	G30978<= not I41108;
	G30979<= not I41111;
	G30980<= not I41114;
	G30981<= not I41117;
	G30982<= not I41120;
	G30983<= not I41123;
	G30984<= not I41126;
	G30985<= not I41129;
	G30986<= not I41132;
	G30987<= not I41135;
	G30988<= not I41138;
	G30989<= not I41141;
	I13089<= not G563;
	I13092<= not G1249;
	I13095<= not G1943;
	I13098<= not G2637;
	I13101<= not G1;
	I13104<= not G2;
	I13107<= not G5;
	I13110<= not G8;
	I13113<= not G11;
	I13116<= not G14;
	I13119<= not G17;
	I13122<= not G20;
	I13125<= not G23;
	I13128<= not G26;
	I13131<= not G27;
	I13134<= not G30;
	I13137<= not G33;
	I13140<= not G36;
	I13143<= not G39;
	I13146<= not G42;
	I13149<= not G45;
	I13152<= not G48;
	I13155<= not G51;
	I13158<= not G165;
	I13161<= not G308;
	I13165<= not G401;
	I13169<= not G550;
	I13173<= not G629;
	I13176<= not G630;
	I13179<= not G853;
	I13182<= not G995;
	I13186<= not G1088;
	I13190<= not G1236;
	I13194<= not G1315;
	I13197<= not G1316;
	I13200<= not G1547;
	I13203<= not G1689;
	I13207<= not G1782;
	I13211<= not G1930;
	I13215<= not G2009;
	I13218<= not G2010;
	I13221<= not G2241;
	I13224<= not G2383;
	I13228<= not G2476;
	I13232<= not G2624;
	I13236<= not G2703;
	I13239<= not G2704;
	I13242<= not G2879;
	I13246<= not G2987;
	I13275<= not G2848;
	I13316<= not G2836;
	I13320<= not G2864;
	I13366<= not G2851;
	I13417<= not G2839;
	I13421<= not G2867;
	I13430<= not G101;
	I13433<= not G105;
	I13478<= not G2854;
	I13501<= not G789;
	I13504<= not G793;
	I13538<= not G2870;
	I13575<= not G1476;
	I13578<= not G1481;
	I13601<= not G121;
	I13604<= not G125;
	I13652<= not G2170;
	I13655<= not G2175;
	I13677<= not G809;
	I13680<= not G813;
	I13742<= not G1501;
	I13745<= not G1506;
	I13775<= not G109;
	I13801<= not G2195;
	I13804<= not G2200;
	I13820<= not G797;
	I13849<= not G1486;
	I13868<= not G2180;
	I13892<= not G3040;
	I13896<= not G343;
	I13901<= not G346;
	I13904<= not G358;
	I13907<= not G1030;
	I13910<= not G361;
	I13913<= not G373;
	I13916<= not G1033;
	I13919<= not G1045;
	I13922<= not G1724;
	I13925<= not G376;
	I13928<= not G388;
	I13931<= not G1048;
	I13934<= not G1060;
	I13937<= not G1727;
	I13940<= not G1739;
	I13943<= not G2418;
	I13947<= not G391;
	I13950<= not G1063;
	I13953<= not G1075;
	I13956<= not G1742;
	I13959<= not G1754;
	I13962<= not G2421;
	I13965<= not G2433;
	I13968<= not G1078;
	I13971<= not G1757;
	I13974<= not G1769;
	I13977<= not G2436;
	I13980<= not G2448;
	I13984<= not G1772;
	I13987<= not G2451;
	I13990<= not G2463;
	I13993<= not G2466;
	I13999<= not G276;
	I14002<= not G276;
	I14006<= not G963;
	I14009<= not G963;
	I14014<= not G499;
	I14017<= not G1657;
	I14020<= not G1657;
	I14027<= not G182;
	I14030<= not G182;
	I14034<= not G1186;
	I14037<= not G2351;
	I14040<= not G2351;
	I14049<= not G870;
	I14052<= not G870;
	I14056<= not G1880;
	I14066<= not G1564;
	I14069<= not G1564;
	I14073<= not G2574;
	I14083<= not G325;
	I14091<= not G2258;
	I14094<= not G2258;
	I14104<= not G331;
	I14113<= not G1012;
	I14134<= not G1018;
	I14143<= not G1706;
	I14149<= not G3231;
	I14163<= not G113;
	I14182<= not G1712;
	I14191<= not G2400;
	I14195<= not G3212;
	I14219<= not G801;
	I14238<= not G2406;
	I14243<= not G3221;
	I14246<= not G3227;
	I14249<= not G3216;
	I14280<= not G1491;
	I14295<= not G3228;
	I14298<= not G3217;
	I14306<= not G97;
	I14338<= not G2185;
	I14343<= not G3219;
	I14357<= not G785;
	I14378<= not G3234;
	I14381<= not G3223;
	I14384<= not G3218;
	I14402<= not G1471;
	I14413<= not G3233;
	I14416<= not G3222;
	I14424<= not G117;
	I14442<= not G2165;
	I14446<= not G3230;
	I14449<= not G3224;
	I14459<= not G805;
	I14472<= not G3080;
	I14475<= not G3225;
	I14478<= not G3213;
	I14489<= not G1496;
	I14496<= not G3226;
	I14499<= not G3214;
	I14502<= not G471;
	I14513<= not G2190;
	I14516<= not G3215;
	I14519<= not G1158;
	I14525<= not G1852;
	I14529<= not G3142;
	I14532<= not G354;
	I14535<= not G2546;
	I14538<= not G369;
	I14541<= not G455;
	I14544<= not G1041;
	I14547<= not G384;
	I14550<= not G458;
	I14553<= not G1056;
	I14556<= not G1142;
	I14559<= not G1735;
	I14562<= not G398;
	I14565<= not G461;
	I14568<= not G1071;
	I14571<= not G1145;
	I14574<= not G1750;
	I14577<= not G1836;
	I14580<= not G2429;
	I14584<= not G465;
	I14587<= not G1085;
	I14590<= not G1148;
	I14593<= not G1765;
	I14596<= not G1839;
	I14599<= not G2444;
	I14602<= not G2530;
	I14605<= not G468;
	I14609<= not G1152;
	I14612<= not G1779;
	I14615<= not G1842;
	I14618<= not G2459;
	I14621<= not G2533;
	I14624<= not G1155;
	I14628<= not G1846;
	I14631<= not G2473;
	I14634<= not G2536;
	I14637<= not G1849;
	I14641<= not G2540;
	I14644<= not G3142;
	I14647<= not G2543;
	I14650<= not G525;
	I14654<= not G3220;
	I14660<= not G1211;
	I14665<= not G3147;
	I14668<= not G3232;
	I14675<= not G1905;
	I14688<= not G2599;
	I14704<= not G2818;
	I14709<= not G3229;
	I14712<= not G138;
	I14715<= not G138;
	I14731<= not G135;
	I14734<= not G135;
	I14739<= not G826;
	I14742<= not G826;
	I14755<= not G2821;
	I14760<= not G405;
	I14763<= not G405;
	I14766<= not G545;
	I14769<= not G545;
	I14775<= not G823;
	I14778<= not G823;
	I14783<= not G1520;
	I14786<= not G1520;
	I14799<= not G551;
	I14802<= not G551;
	I14808<= not G623;
	I14811<= not G623;
	I14816<= not G1092;
	I14819<= not G1092;
	I14822<= not G1231;
	I14825<= not G1231;
	I14831<= not G1517;
	I14834<= not G1517;
	I14839<= not G2214;
	I14842<= not G2214;
	I14848<= not G2824;
	I14857<= not G626;
	I14860<= not G626;
	I14865<= not G1237;
	I14868<= not G1237;
	I14874<= not G1309;
	I14877<= not G1309;
	I14882<= not G1786;
	I14885<= not G1786;
	I14888<= not G1925;
	I14891<= not G1925;
	I14897<= not G2211;
	I14900<= not G2211;
	I14917<= not G1312;
	I14920<= not G1312;
	I14925<= not G1931;
	I14928<= not G1931;
	I14934<= not G2003;
	I14937<= not G2003;
	I14942<= not G2480;
	I14945<= not G2480;
	I14948<= not G2619;
	I14951<= not G2619;
	I14957<= not G2827;
	I14973<= not G2006;
	I14976<= not G2006;
	I14981<= not G2625;
	I14984<= not G2625;
	I14990<= not G2697;
	I14993<= not G2697;
	I15012<= not G2700;
	I15015<= not G2700;
	I15019<= not G2830;
	I15222<= not G3151;
	I15226<= not G474;
	I15230<= not G499;
	I15256<= not G2950;
	I15262<= not G481;
	I15267<= not G1161;
	I15271<= not G1186;
	I15288<= not G3109;
	I15299<= not G1168;
	I15304<= not G1855;
	I15308<= not G1880;
	I15313<= not G2930;
	I15317<= not G2842;
	I15326<= not G3117;
	I15329<= not G3117;
	I15345<= not G1862;
	I15350<= not G2549;
	I15354<= not G2574;
	I15359<= not G2858;
	I15369<= not G3129;
	I15372<= not G3129;
	I15392<= not G2556;
	I15398<= not G2845;
	I15429<= not G2833;
	I15433<= not G2861;
	I15442<= not G3235;
	I15445<= not G3236;
	I15448<= not G3237;
	I15451<= not G3238;
	I15454<= not G3239;
	I15457<= not G3240;
	I15460<= not G3241;
	I15463<= not G3242;
	I15466<= not G3243;
	I15469<= not G3244;
	I15472<= not G3245;
	I15475<= not G3246;
	I15478<= not G3247;
	I15481<= not G3248;
	I15484<= not G3249;
	I15487<= not G3250;
	I15490<= not G3251;
	I15493<= not G3252;
	I15499<= not G7911;
	I15505<= not G7963;
	I15511<= not G8014;
	I15517<= not G8089;
	I15523<= not G3254;
	I15526<= not G6314;
	I15532<= not G3410;
	I15535<= not G6519;
	I15538<= not G6369;
	I15543<= not G3410;
	I15546<= not G6783;
	I15549<= not G6574;
	I15553<= not G3566;
	I15556<= not G6783;
	I15559<= not G7015;
	I15562<= not G5778;
	I15565<= not G6838;
	I15568<= not G3722;
	I15571<= not G7085;
	I15574<= not G6838;
	I15577<= not G7265;
	I15580<= not G5837;
	I15584<= not G3254;
	I15590<= not G3410;
	I15593<= not G6519;
	I15599<= not G3566;
	I15602<= not G6783;
	I15605<= not G6574;
	I15610<= not G3566;
	I15613<= not G7085;
	I15616<= not G6838;
	I15620<= not G3722;
	I15623<= not G7085;
	I15626<= not G7265;
	I15629<= not G5837;
	I15636<= not G3410;
	I15642<= not G3566;
	I15645<= not G6783;
	I15651<= not G3722;
	I15654<= not G7085;
	I15657<= not G6838;
	I15662<= not G3722;
	I15671<= not G3566;
	I15677<= not G3722;
	I15680<= not G7085;
	I15696<= not G3722;
	I15771<= not G6000;
	I15779<= not G6000;
	I15784<= not G6000;
	I15787<= not G6000;
	I15794<= not G3338;
	I15800<= not G3494;
	I15803<= not G8107;
	I15806<= not G5550;
	I15810<= not G3338;
	I15815<= not G3650;
	I15818<= not G5596;
	I15822<= not G3494;
	I15827<= not G3806;
	I15830<= not G8031;
	I15833<= not G3338;
	I15836<= not G3366;
	I15839<= not G5613;
	I15843<= not G3650;
	I15847<= not G3878;
	I15850<= not G5627;
	I15853<= not G3494;
	I15856<= not G3522;
	I15859<= not G5638;
	I15863<= not G3806;
	I15866<= not G3878;
	I15869<= not G7976;
	I15873<= not G5655;
	I15876<= not G3650;
	I15879<= not G3678;
	I15882<= not G3878;
	I15887<= not G5693;
	I15890<= not G3806;
	I15893<= not G3834;
	I15896<= not G3878;
	I15899<= not G5626;
	I15902<= not G6486;
	I15909<= not G5745;
	I15912<= not G3878;
	I15915<= not G3878;
	I15918<= not G6643;
	I15922<= not G5654;
	I15925<= not G6751;
	I15932<= not G5423;
	I15935<= not G3878;
	I15938<= not G3338;
	I15942<= not G6945;
	I15946<= not G5692;
	I15949<= not G7053;
	I15955<= not G3878;
	I15958<= not G3878;
	I15961<= not G6051;
	I15964<= not G7554;
	I15967<= not G3494;
	I15971<= not G7195;
	I15975<= not G5744;
	I15978<= not G7303;
	I15983<= not G3878;
	I15986<= not G3878;
	I15989<= not G6053;
	I15992<= not G6055;
	I15995<= not G7577;
	I15998<= not G3650;
	I16002<= not G7391;
	I16006<= not G3878;
	I16009<= not G3878;
	I16012<= not G5390;
	I16015<= not G6056;
	I16018<= not G6058;
	I16021<= not G6060;
	I16024<= not G7591;
	I16027<= not G3806;
	I16031<= not G3878;
	I16034<= not G5396;
	I16037<= not G6061;
	I16041<= not G6486;
	I16044<= not G5397;
	I16047<= not G6063;
	I16050<= not G6065;
	I16053<= not G6067;
	I16056<= not G7606;
	I16059<= not G3878;
	I16062<= not G3900;
	I16065<= not G7936;
	I16068<= not G5438;
	I16071<= not G5395;
	I16074<= not G5399;
	I16079<= not G6086;
	I16082<= not G5401;
	I16085<= not G6080;
	I16089<= not G6751;
	I16092<= not G5402;
	I16095<= not G6082;
	I16098<= not G6084;
	I16101<= not G3878;
	I16104<= not G6448;
	I16107<= not G5398;
	I16110<= not G5404;
	I16114<= not G7936;
	I16117<= not G5473;
	I16120<= not G5400;
	I16123<= not G5406;
	I16128<= not G6103;
	I16131<= not G5408;
	I16134<= not G6099;
	I16138<= not G7053;
	I16141<= not G5409;
	I16144<= not G6101;
	I16147<= not G3878;
	I16150<= not G3900;
	I16153<= not G3306;
	I16156<= not G5438;
	I16159<= not G5403;
	I16163<= not G6031;
	I16166<= not G6713;
	I16169<= not G5405;
	I16172<= not G5413;
	I16176<= not G7936;
	I16179<= not G5512;
	I16182<= not G5407;
	I16185<= not G5415;
	I16190<= not G6118;
	I16193<= not G5417;
	I16196<= not G6116;
	I16200<= not G7303;
	I16203<= not G3878;
	I16206<= not G6448;
	I16209<= not G5438;
	I16212<= not G5411;
	I16215<= not G3462;
	I16218<= not G5473;
	I16221<= not G5412;
	I16225<= not G6042;
	I16228<= not G7015;
	I16231<= not G5414;
	I16234<= not G5420;
	I16238<= not G7936;
	I16241<= not G5556;
	I16244<= not G5416;
	I16247<= not G5422;
	I16252<= not G6134;
	I16255<= not G3900;
	I16258<= not G3306;
	I16261<= not G6448;
	I16264<= not G6713;
	I16267<= not G5473;
	I16270<= not G5418;
	I16273<= not G3618;
	I16276<= not G5512;
	I16279<= not G5419;
	I16283<= not G6046;
	I16286<= not G7265;
	I16289<= not G5421;
	I16292<= not G5426;
	I16296<= not G3306;
	I16300<= not G3462;
	I16303<= not G6713;
	I16306<= not G7015;
	I16309<= not G5512;
	I16312<= not G5424;
	I16315<= not G3774;
	I16318<= not G5556;
	I16321<= not G5425;
	I16325<= not G6052;
	I16328<= not G3900;
	I16332<= not G3462;
	I16335<= not G3618;
	I16338<= not G7015;
	I16341<= not G7265;
	I16344<= not G5556;
	I16347<= not G5427;
	I16354<= not G3618;
	I16357<= not G3774;
	I16360<= not G7265;
	I16363<= not G3900;
	I16372<= not G3774;
	I16432<= not G3366;
	I16438<= not G3522;
	I16444<= not G3678;
	I16450<= not G3834;
	I16453<= not G7936;
	I16457<= not G7936;
	I16462<= not G5438;
	I16465<= not G6000;
	I16469<= not G7936;
	I16472<= not G7901;
	I16476<= not G6448;
	I16479<= not G5438;
	I16482<= not G6000;
	I16486<= not G5473;
	I16489<= not G6000;
	I16493<= not G7936;
	I16499<= not G7901;
	I16504<= not G3306;
	I16507<= not G6448;
	I16511<= not G6713;
	I16514<= not G5473;
	I16517<= not G6000;
	I16521<= not G5512;
	I16524<= not G6000;
	I16532<= not G7901;
	I16538<= not G3306;
	I16541<= not G5438;
	I16544<= not G6054;
	I16549<= not G3462;
	I16552<= not G6713;
	I16556<= not G7015;
	I16559<= not G5512;
	I16562<= not G6000;
	I16566<= not G5556;
	I16569<= not G6000;
	I16578<= not G6448;
	I16581<= not G5438;
	I16587<= not G3462;
	I16590<= not G5473;
	I16593<= not G6059;
	I16598<= not G3618;
	I16601<= not G7015;
	I16605<= not G7265;
	I16608<= not G5556;
	I16611<= not G6000;
	I16624<= not G3306;
	I16627<= not G6448;
	I16630<= not G6057;
	I16633<= not G6486;
	I16641<= not G6713;
	I16644<= not G5473;
	I16650<= not G3618;
	I16653<= not G5512;
	I16656<= not G6066;
	I16661<= not G3774;
	I16664<= not G7265;
	I16677<= not G3306;
	I16681<= not G6643;
	I16684<= not G6486;
	I16694<= not G3462;
	I16697<= not G6713;
	I16700<= not G6064;
	I16703<= not G6751;
	I16711<= not G7015;
	I16714<= not G5512;
	I16720<= not G3774;
	I16723<= not G5556;
	I16726<= not G6085;
	I16741<= not G6062;
	I16744<= not G3338;
	I16747<= not G6643;
	I16759<= not G3462;
	I16763<= not G6945;
	I16766<= not G6751;
	I16776<= not G3618;
	I16779<= not G7015;
	I16782<= not G6083;
	I16785<= not G7053;
	I16793<= not G7265;
	I16796<= not G5556;
	I16811<= not G3338;
	I16814<= not G6486;
	I16832<= not G6081;
	I16835<= not G3494;
	I16838<= not G6945;
	I16850<= not G3618;
	I16854<= not G7195;
	I16857<= not G7053;
	I16867<= not G3774;
	I16870<= not G7265;
	I16873<= not G6102;
	I16876<= not G7303;
	I16897<= not G6643;
	I16900<= not G6486;
	I16915<= not G3494;
	I16918<= not G6751;
	I16936<= not G6100;
	I16939<= not G3650;
	I16942<= not G7195;
	I16954<= not G3774;
	I16958<= not G7391;
	I16961<= not G7303;
	I16972<= not G3900;
	I16984<= not G7936;
	I16987<= not G6079;
	I16990<= not G3338;
	I16993<= not G6643;
	I17009<= not G6945;
	I17012<= not G6751;
	I17027<= not G3650;
	I17030<= not G7053;
	I17048<= not G6117;
	I17051<= not G3806;
	I17054<= not G7391;
	I17066<= not G3900;
	I17070<= not G7528;
	I17081<= not G3338;
	I17097<= not G7936;
	I17100<= not G6098;
	I17103<= not G3494;
	I17106<= not G6945;
	I17122<= not G7195;
	I17125<= not G7053;
	I17140<= not G3806;
	I17143<= not G7303;
	I17159<= not G3900;
	I17184<= not G3494;
	I17200<= not G7936;
	I17203<= not G6115;
	I17206<= not G3650;
	I17209<= not G7195;
	I17225<= not G7391;
	I17228<= not G7303;
	I17235<= not G3900;
	I17238<= not G3900;
	I17278<= not G3650;
	I17294<= not G7936;
	I17297<= not G6130;
	I17300<= not G3806;
	I17303<= not G7391;
	I17311<= not G3900;
	I17363<= not G3806;
	I17370<= not G3900;
	I17373<= not G3900;
	I17433<= not G3900;
	I17483<= not G3900;
	I17486<= not G3900;
	I17527<= not G3900;
	I17557<= not G3900;
	I17627<= not G7575;
	I17632<= not G6183;
	I17637<= not G6204;
	I17641<= not G6215;
	I17645<= not G6288;
	I17649<= not G6293;
	I17653<= not G6304;
	I17658<= not G6367;
	I17662<= not G6425;
	I17666<= not G6430;
	I17670<= not G6441;
	I17673<= not G8107;
	I17677<= not G6517;
	I17681<= not G6572;
	I17685<= not G6630;
	I17689<= not G6635;
	I17692<= not G8107;
	I17698<= not G6711;
	I17701<= not G6781;
	I17705<= not G6836;
	I17709<= not G6894;
	I17712<= not G8031;
	I17715<= not G8107;
	I17721<= not G6641;
	I17724<= not G6942;
	I17727<= not G7013;
	I17730<= not G7083;
	I17734<= not G7138;
	I17737<= not G6000;
	I17740<= not G8031;
	I17743<= not G8107;
	I17746<= not G8107;
	I17750<= not G7157;
	I17753<= not G6943;
	I17756<= not G7192;
	I17759<= not G7263;
	I17762<= not G7333;
	I17765<= not G7976;
	I17768<= not G8031;
	I17771<= not G8107;
	I17774<= not G8107;
	I17780<= not G7348;
	I17783<= not G7353;
	I17786<= not G7193;
	I17789<= not G7388;
	I17792<= not G7459;
	I17795<= not G7976;
	I17798<= not G8031;
	I17801<= not G8107;
	I17804<= not G8031;
	I17807<= not G8107;
	I17813<= not G5707;
	I17816<= not G7346;
	I17819<= not G6448;
	I17822<= not G7478;
	I17825<= not G7483;
	I17828<= not G7389;
	I17831<= not G7518;
	I17834<= not G7976;
	I17837<= not G8031;
	I17840<= not G8107;
	I17843<= not G8031;
	I17846<= not G8107;
	I17849<= not G8103;
	I17854<= not G6232;
	I17857<= not G6448;
	I17860<= not G5765;
	I17863<= not G7476;
	I17866<= not G6713;
	I17869<= not G7534;
	I17872<= not G7539;
	I17875<= not G7976;
	I17878<= not G8031;
	I17881<= not G7976;
	I17884<= not G8031;
	I17889<= not G6314;
	I17892<= not G6232;
	I17895<= not G6448;
	I17898<= not G6643;
	I17901<= not G6369;
	I17904<= not G6713;
	I17907<= not G5824;
	I17910<= not G7532;
	I17913<= not G7015;
	I17916<= not G7560;
	I17919<= not G7976;
	I17922<= not G8031;
	I17925<= not G7976;
	I17928<= not G8031;
	I17933<= not G3254;
	I17936<= not G6314;
	I17939<= not G6232;
	I17942<= not G5548;
	I17945<= not G5668;
	I17948<= not G6643;
	I17951<= not G6519;
	I17954<= not G6369;
	I17957<= not G6713;
	I17960<= not G6945;
	I17963<= not G6574;
	I17966<= not G7015;
	I17969<= not G5880;
	I17972<= not G7558;
	I17975<= not G7265;
	I17978<= not G7795;
	I17981<= not G7976;
	I17984<= not G7976;
	I17989<= not G3254;
	I17992<= not G6314;
	I17995<= not G6232;
	I17998<= not G5668;
	I18001<= not G6643;
	I18004<= not G3410;
	I18007<= not G6519;
	I18010<= not G6369;
	I18013<= not G5594;
	I18016<= not G5720;
	I18019<= not G6945;
	I18022<= not G6783;
	I18025<= not G6574;
	I18028<= not G7015;
	I18031<= not G7195;
	I18034<= not G6838;
	I18037<= not G7265;
	I18040<= not G7976;
	I18043<= not G7976;
	I18046<= not G3254;
	I18049<= not G6314;
	I18052<= not G6232;
	I18055<= not G5668;
	I18058<= not G6643;
	I18061<= not G3410;
	I18064<= not G6519;
	I18067<= not G6369;
	I18070<= not G5720;
	I18073<= not G6945;
	I18076<= not G3566;
	I18079<= not G6783;
	I18082<= not G6574;
	I18085<= not G5611;
	I18088<= not G5778;
	I18091<= not G7195;
	I18094<= not G7085;
	I18097<= not G6838;
	I18100<= not G7265;
	I18103<= not G7391;
	I18121<= not G3254;
	I18124<= not G6314;
	I18127<= not G6232;
	I18130<= not G5547;
	I18133<= not G6448;
	I18136<= not G5668;
	I18139<= not G6643;
	I18142<= not G3410;
	I18145<= not G6519;
	I18148<= not G6369;
	I18151<= not G5720;
	I18154<= not G6945;
	I18157<= not G3566;
	I18160<= not G6783;
	I18163<= not G6574;
	I18166<= not G5778;
	I18169<= not G7195;
	I18172<= not G3722;
	I18175<= not G7085;
	I18178<= not G6838;
	I18181<= not G5636;
	I18184<= not G5837;
	I18187<= not G7391;
	I18211<= not G6232;
	I18214<= not G3254;
	I18217<= not G6314;
	I18220<= not G6232;
	I18223<= not G6448;
	I18226<= not G5668;
	I18229<= not G3410;
	I18232<= not G6519;
	I18235<= not G6369;
	I18238<= not G5593;
	I18241<= not G6713;
	I18244<= not G5720;
	I18247<= not G6945;
	I18250<= not G3566;
	I18253<= not G6783;
	I18256<= not G6574;
	I18259<= not G5778;
	I18262<= not G7195;
	I18265<= not G3722;
	I18268<= not G7085;
	I18271<= not G6838;
	I18274<= not G5837;
	I18277<= not G7391;
	I18295<= not G6314;
	I18298<= not G6232;
	I18302<= not G3254;
	I18305<= not G6314;
	I18308<= not G6448;
	I18311<= not G5668;
	I18314<= not G6369;
	I18317<= not G3410;
	I18320<= not G6519;
	I18323<= not G6369;
	I18326<= not G6713;
	I18329<= not G5720;
	I18332<= not G3566;
	I18335<= not G6783;
	I18338<= not G6574;
	I18341<= not G5610;
	I18344<= not G7015;
	I18347<= not G5778;
	I18350<= not G7195;
	I18353<= not G3722;
	I18356<= not G7085;
	I18359<= not G6838;
	I18362<= not G5837;
	I18365<= not G7391;
	I18375<= not G3254;
	I18378<= not G6314;
	I18381<= not G6232;
	I18386<= not G3254;
	I18389<= not G6519;
	I18392<= not G6369;
	I18396<= not G3410;
	I18399<= not G6519;
	I18402<= not G6713;
	I18405<= not G5720;
	I18408<= not G6574;
	I18411<= not G3566;
	I18414<= not G6783;
	I18417<= not G6574;
	I18420<= not G7015;
	I18423<= not G5778;
	I18426<= not G3722;
	I18429<= not G7085;
	I18432<= not G6838;
	I18435<= not G5635;
	I18438<= not G7265;
	I18441<= not G5837;
	I18444<= not G7391;
	I18449<= not G10868;
	I18452<= not G10930;
	I18455<= not G11031;
	I18458<= not G11208;
	I18461<= not G10931;
	I18464<= not G8620;
	I18467<= not G8769;
	I18470<= not G8808;
	I18473<= not G8839;
	I18476<= not G8791;
	I18479<= not G8820;
	I18482<= not G8859;
	I18485<= not G8809;
	I18488<= not G8840;
	I18491<= not G8891;
	I18494<= not G8821;
	I18497<= not G8860;
	I18500<= not G8924;
	I18503<= not G8658;
	I18506<= not G8699;
	I18509<= not G8770;
	I18512<= not G9309;
	I18515<= not G8843;
	I18518<= not G8893;
	I18521<= not G9449;
	I18524<= not G9640;
	I18527<= not G10017;
	I18530<= not G10888;
	I18533<= not G10967;
	I18536<= not G11101;
	I18539<= not G11290;
	I18542<= not G10968;
	I18545<= not G8630;
	I18548<= not G8792;
	I18551<= not G8824;
	I18554<= not G8866;
	I18557<= not G8810;
	I18560<= not G8844;
	I18563<= not G8897;
	I18566<= not G8825;
	I18569<= not G8867;
	I18572<= not G8931;
	I18575<= not G8845;
	I18578<= not G8898;
	I18581<= not G8964;
	I18584<= not G8677;
	I18587<= not G8718;
	I18590<= not G8793;
	I18593<= not G9390;
	I18596<= not G8870;
	I18599<= not G8933;
	I18602<= not G9591;
	I18605<= not G9786;
	I18608<= not G10126;
	I18611<= not G10909;
	I18614<= not G11002;
	I18617<= not G11169;
	I18620<= not G11385;
	I18623<= not G11003;
	I18626<= not G8649;
	I18629<= not G8811;
	I18632<= not G8850;
	I18635<= not G8904;
	I18638<= not G8826;
	I18641<= not G8871;
	I18644<= not G8937;
	I18647<= not G8851;
	I18650<= not G8905;
	I18653<= not G8971;
	I18656<= not G8872;
	I18659<= not G8938;
	I18662<= not G8996;
	I18665<= not G8689;
	I18668<= not G8756;
	I18671<= not G8812;
	I18674<= not G9487;
	I18677<= not G8908;
	I18680<= not G8973;
	I18683<= not G9733;
	I18686<= not G9932;
	I18689<= not G10231;
	I18692<= not G10935;
	I18695<= not G11054;
	I18698<= not G11255;
	I18701<= not G11471;
	I18704<= not G11055;
	I18707<= not G8665;
	I18710<= not G8827;
	I18713<= not G8877;
	I18716<= not G8944;
	I18719<= not G8852;
	I18722<= not G8909;
	I18725<= not G8977;
	I18728<= not G8878;
	I18731<= not G8945;
	I18734<= not G9003;
	I18737<= not G8910;
	I18740<= not G8978;
	I18743<= not G9025;
	I18746<= not G8707;
	I18749<= not G8779;
	I18752<= not G8828;
	I18755<= not G9629;
	I18758<= not G8948;
	I18761<= not G9005;
	I18764<= not G9879;
	I18767<= not G10086;
	I18770<= not G10333;
	I18773<= not G10830;
	I18777<= not G9050;
	I18780<= not G10870;
	I18784<= not G9067;
	I18787<= not G10910;
	I18791<= not G9084;
	I18794<= not G10973;
	I18810<= not G10813;
	I18813<= not G10850;
	I18817<= not G9067;
	I18820<= not G10890;
	I18824<= not G9084;
	I18827<= not G10936;
	I18835<= not G10834;
	I18838<= not G10871;
	I18842<= not G9084;
	I18845<= not G10911;
	I18854<= not G10854;
	I18857<= not G10891;
	I18866<= not G10875;
	I18929<= not G10711;
	I18943<= not G9149;
	I18962<= not G9159;
	I18969<= not G8726;
	I18990<= not G9183;
	I19025<= not G9225;
	I19030<= not G8726;
	I19105<= not G8726;
	I19119<= not G9202;
	I19160<= not G10549;
	I19174<= not G9263;
	I19195<= not G8726;
	I19208<= not G10424;
	I19211<= not G10486;
	I19226<= not G10606;
	I19240<= not G9341;
	I19271<= not G10500;
	I19274<= not G10560;
	I19289<= not G10653;
	I19303<= not G9422;
	I19307<= not G8726;
	I19315<= not G10424;
	I19318<= not G10486;
	I19321<= not G10549;
	I19342<= not G10574;
	I19345<= not G10617;
	I19360<= not G10683;
	I19374<= not G10500;
	I19377<= not G10560;
	I19380<= not G10606;
	I19401<= not G10631;
	I19404<= not G10664;
	I19412<= not G10486;
	I19415<= not G10549;
	I19426<= not G10574;
	I19429<= not G10617;
	I19432<= not G10653;
	I19449<= not G10424;
	I19452<= not G10560;
	I19455<= not G10606;
	I19466<= not G10631;
	I19469<= not G10664;
	I19472<= not G10683;
	I19479<= not G10549;
	I19482<= not G10500;
	I19485<= not G10617;
	I19488<= not G10653;
	I19500<= not G10424;
	I19503<= not G10486;
	I19507<= not G10606;
	I19510<= not G10574;
	I19513<= not G10664;
	I19516<= not G10683;
	I19523<= not G10500;
	I19526<= not G10560;
	I19530<= not G10653;
	I19533<= not G10631;
	I19539<= not G10549;
	I19542<= not G10574;
	I19545<= not G10617;
	I19549<= not G10683;
	I19552<= not G8430;
	I19557<= not G10606;
	I19560<= not G10631;
	I19563<= not G10664;
	I19569<= not G10653;
	I19573<= not G8835;
	I19576<= not G10683;
	I19582<= not G8862;
	I19587<= not G9173;
	I19591<= not G8900;
	I19595<= not G10810;
	I19598<= not G9215;
	I19602<= not G8940;
	I19605<= not G10797;
	I19608<= not G10831;
	I19611<= not G9276;
	I19615<= not G10789;
	I19618<= not G10814;
	I19621<= not G10851;
	I19624<= not G9354;
	I19628<= not G10784;
	I19631<= not G10801;
	I19634<= not G10835;
	I19637<= not G10872;
	I19642<= not G10793;
	I19645<= not G10818;
	I19648<= not G10855;
	I19654<= not G10805;
	I19657<= not G10839;
	I19667<= not G10822;
	I19689<= not G10016;
	I19702<= not G10125;
	I19711<= not G10230;
	I19718<= not G8726;
	I19722<= not G10332;
	I19727<= not G8726;
	I19733<= not G8726;
	I19736<= not G9184;
	I19739<= not G10694;
	I19747<= not G8726;
	I19750<= not G8726;
	I19753<= not G9229;
	I19756<= not G10424;
	I19759<= not G10714;
	I19767<= not G8726;
	I19771<= not G10038;
	I19774<= not G10500;
	I19777<= not G10735;
	I19784<= not G8726;
	I19787<= not G8726;
	I19791<= not G10486;
	I19794<= not G10676;
	I19797<= not G10147;
	I19800<= not G10574;
	I19803<= not G10754;
	I19808<= not G8726;
	I19813<= not G10649;
	I19816<= not G10703;
	I19820<= not G10560;
	I19823<= not G10705;
	I19826<= not G10252;
	I19829<= not G10631;
	I19833<= not G8726;
	I19836<= not G8726;
	I19844<= not G8533;
	I19847<= not G10677;
	I19852<= not G10679;
	I19855<= not G10723;
	I19859<= not G10617;
	I19862<= not G10725;
	I19865<= not G10354;
	I19869<= not G8726;
	I19872<= not G8317;
	I19877<= not G8547;
	I19883<= not G8550;
	I19886<= not G10706;
	I19891<= not G10708;
	I19894<= not G10744;
	I19898<= not G10664;
	I19901<= not G10746;
	I19905<= not G8726;
	I19915<= not G8560;
	I19921<= not G8563;
	I19924<= not G10726;
	I19929<= not G10728;
	I19932<= not G10763;
	I19952<= not G8571;
	I19958<= not G8574;
	I19961<= not G10747;
	I19986<= not G8577;
	I20009<= not G8313;
	I20062<= not G10480;
	I20117<= not G10876;
	I20264<= not G9027;
	I20278<= not G9027;
	I20283<= not G9050;
	I20295<= not G10015;
	I20299<= not G10800;
	I20305<= not G9050;
	I20310<= not G9067;
	I20320<= not G10792;
	I20324<= not G10124;
	I20328<= not G10817;
	I20334<= not G9067;
	I20339<= not G9084;
	I20347<= not G10787;
	I20351<= not G10804;
	I20355<= not G10229;
	I20359<= not G10838;
	I20365<= not G9084;
	I20376<= not G8569;
	I20379<= not G11213;
	I20382<= not G10907;
	I20386<= not G10796;
	I20390<= not G10821;
	I20394<= not G10331;
	I20398<= not G10858;
	I20407<= not G9027;
	I20410<= not G10887;
	I20414<= not G8575;
	I20417<= not G10933;
	I20421<= not G10808;
	I20425<= not G10842;
	I20441<= not G9027;
	I20444<= not G10869;
	I20448<= not G9050;
	I20451<= not G10908;
	I20455<= not G8578;
	I20458<= not G10972;
	I20462<= not G10825;
	I20476<= not G9027;
	I20479<= not G10849;
	I20483<= not G9050;
	I20486<= not G10889;
	I20490<= not G9067;
	I20493<= not G10934;
	I20497<= not G8579;
	I20500<= not G11007;
	I20514<= not G11769;
	I20517<= not G12425;
	I20520<= not G13246;
	I20523<= not G13317;
	I20526<= not G12519;
	I20529<= not G13319;
	I20532<= not G13339;
	I20535<= not G13359;
	I20538<= not G13384;
	I20541<= not G11599;
	I20544<= not G11628;
	I20547<= not G13248;
	I20550<= not G13267;
	I20553<= not G13290;
	I20556<= not G12435;
	I20559<= not G11937;
	I20562<= not G11786;
	I20565<= not G12432;
	I20568<= not G13269;
	I20571<= not G13341;
	I20574<= not G12534;
	I20577<= not G13342;
	I20580<= not G13364;
	I20583<= not G13389;
	I20586<= not G11606;
	I20589<= not G11629;
	I20592<= not G11651;
	I20595<= not G13271;
	I20598<= not G13292;
	I20601<= not G13321;
	I20604<= not G12440;
	I20607<= not G11990;
	I20610<= not G11812;
	I20613<= not G12437;
	I20616<= not G13294;
	I20619<= not G13366;
	I20622<= not G12543;
	I20625<= not G13367;
	I20628<= not G13394;
	I20631<= not G11611;
	I20634<= not G11636;
	I20637<= not G11652;
	I20640<= not G11670;
	I20643<= not G13296;
	I20646<= not G13323;
	I20649<= not G13344;
	I20652<= not G12445;
	I20655<= not G12059;
	I20658<= not G11845;
	I20661<= not G12442;
	I20664<= not G13325;
	I20667<= not G13396;
	I20670<= not G12552;
	I20673<= not G13397;
	I20676<= not G11616;
	I20679<= not G11641;
	I20682<= not G11659;
	I20685<= not G11671;
	I20688<= not G11682;
	I20691<= not G13327;
	I20694<= not G13346;
	I20697<= not G13369;
	I20700<= not G12450;
	I20703<= not G12123;
	I20706<= not G11490;
	I20709<= not G13070;
	I20791<= not G13149;
	I20794<= not G13111;
	I20799<= not G13155;
	I20802<= not G13160;
	I20805<= not G13124;
	I20810<= not G13164;
	I20813<= not G13265;
	I20816<= not G12487;
	I20820<= not G13171;
	I20823<= not G13135;
	I20828<= not G13175;
	I20832<= not G12507;
	I20836<= not G13182;
	I20839<= not G13143;
	I20844<= not G12524;
	I20848<= not G13194;
	I20852<= not G12457;
	I20858<= not G12539;
	I20863<= not G12467;
	I20873<= not G12482;
	I20886<= not G12499;
	I20909<= not G13055;
	I20959<= not G11713;
	I21012<= not G12503;
	I21037<= not G12486;
	I21045<= not G12520;
	I21064<= not G13147;
	I21075<= not G12506;
	I21083<= not G12535;
	I21096<= not G11749;
	I21108<= not G13150;
	I21119<= not G12523;
	I21127<= not G12544;
	I21137<= not G11749;
	I21149<= not G13156;
	I21160<= not G12538;
	I21165<= not G13110;
	I21178<= not G11749;
	I21190<= not G13165;
	I21208<= not G11749;
	I21241<= not G13378;
	I21246<= not G11624;
	I21249<= not G11600;
	I21252<= not G11644;
	I21256<= not G11647;
	I21259<= not G11630;
	I21262<= not G11713;
	I21267<= not G11663;
	I21271<= not G11666;
	I21274<= not G11653;
	I21277<= not G12430;
	I21282<= not G11675;
	I21286<= not G11678;
	I21289<= not G12434;
	I21292<= not G11888;
	I21297<= not G11687;
	I21301<= not G12438;
	I21304<= not G11927;
	I21310<= not G12332;
	I21313<= not G11743;
	I21318<= not G12362;
	I21321<= not G11758;
	I21326<= not G12378;
	I21329<= not G11766;
	I21337<= not G12408;
	I21340<= not G11779;
	I21351<= not G12420;
	I21354<= not G11798;
	I21361<= not G13026;
	I21364<= not G13028;
	I21374<= not G12424;
	I21377<= not G11821;
	I21381<= not G13157;
	I21389<= not G12883;
	I21392<= not G13020;
	I21395<= not G13034;
	I21398<= not G13021;
	I21404<= not G13037;
	I21407<= not G13039;
	I21415<= not G11854;
	I21420<= not G13166;
	I21426<= not G11661;
	I21429<= not G13027;
	I21432<= not G13044;
	I21435<= not G11662;
	I21443<= not G12923;
	I21446<= not G13029;
	I21449<= not G13047;
	I21452<= not G13030;
	I21458<= not G13050;
	I21461<= not G13052;
	I21476<= not G11672;
	I21479<= not G13035;
	I21482<= not G13058;
	I21488<= not G11673;
	I21491<= not G13038;
	I21494<= not G13061;
	I21497<= not G11674;
	I21505<= not G12952;
	I21508<= not G13040;
	I21511<= not G13064;
	I21514<= not G13041;
	I21520<= not G13067;
	I21523<= not G13069;
	I21531<= not G11683;
	I21534<= not G13045;
	I21537<= not G13071;
	I21548<= not G11684;
	I21551<= not G13048;
	I21554<= not G13074;
	I21560<= not G11685;
	I21563<= not G13051;
	I21566<= not G13077;
	I21569<= not G11686;
	I21577<= not G12981;
	I21580<= not G13053;
	I21583<= not G13080;
	I21586<= not G13054;
	I21595<= not G11691;
	I21598<= not G13059;
	I21601<= not G13087;
	I21609<= not G11692;
	I21612<= not G13062;
	I21615<= not G13090;
	I21626<= not G11693;
	I21629<= not G13065;
	I21632<= not G13093;
	I21638<= not G11694;
	I21641<= not G13068;
	I21644<= not G13096;
	I21647<= not G11695;
	I21655<= not G11696;
	I21658<= not G13072;
	I21661<= not G13098;
	I21666<= not G13100;
	I21674<= not G11698;
	I21677<= not G13075;
	I21680<= not G13102;
	I21688<= not G11699;
	I21691<= not G13078;
	I21694<= not G13105;
	I21705<= not G11700;
	I21708<= not G13081;
	I21711<= not G13108;
	I21720<= not G11701;
	I21723<= not G13088;
	I21726<= not G13112;
	I21730<= not G13089;
	I21736<= not G11702;
	I21739<= not G13091;
	I21742<= not G13114;
	I21747<= not G13116;
	I21755<= not G11704;
	I21758<= not G13094;
	I21761<= not G13118;
	I21769<= not G11705;
	I21772<= not G13097;
	I21775<= not G13121;
	I21780<= not G13305;
	I21787<= not G11707;
	I21790<= not G13099;
	I21793<= not G13123;
	I21796<= not G11708;
	I21803<= not G11709;
	I21806<= not G13103;
	I21809<= not G13125;
	I21813<= not G13104;
	I21819<= not G11710;
	I21822<= not G13106;
	I21825<= not G13127;
	I21830<= not G13129;
	I21838<= not G11712;
	I21841<= not G13109;
	I21844<= not G13131;
	I21852<= not G11716;
	I21855<= not G13113;
	I21862<= not G11717;
	I21865<= not G13115;
	I21868<= not G13134;
	I21871<= not G11718;
	I21878<= not G11719;
	I21881<= not G13119;
	I21884<= not G13136;
	I21888<= not G13120;
	I21894<= not G11720;
	I21897<= not G13122;
	I21900<= not G13138;
	I21905<= not G13140;
	I21908<= not G13082;
	I21918<= not G11721;
	I21923<= not G11722;
	I21926<= not G13126;
	I21933<= not G11723;
	I21936<= not G13128;
	I21939<= not G13142;
	I21942<= not G11724;
	I21949<= not G11725;
	I21952<= not G13132;
	I21955<= not G13144;
	I21959<= not G13133;
	I21962<= not G13004;
	I21974<= not G11726;
	I21979<= not G11727;
	I21982<= not G13137;
	I21989<= not G11728;
	I21992<= not G13139;
	I21995<= not G13146;
	I21998<= not G11729;
	I22014<= not G11730;
	I22019<= not G11731;
	I22022<= not G13145;
	I22025<= not G11617;
	I22044<= not G11733;
	I22120<= not G12909;
	I22163<= not G12433;
	I22382<= not G520;
	I22414<= not G1206;
	I22444<= not G1900;
	I22475<= not G2594;
	I22503<= not G13598;
	I22506<= not G13624;
	I22509<= not G13610;
	I22512<= not G13635;
	I22515<= not G13620;
	I22518<= not G13647;
	I22521<= not G13632;
	I22524<= not G13673;
	I22527<= not G13469;
	I22530<= not G14774;
	I22533<= not G14795;
	I22536<= not G14829;
	I22539<= not G14882;
	I22542<= not G14954;
	I22545<= not G15018;
	I22548<= not G14718;
	I22551<= not G14745;
	I22554<= not G14765;
	I22557<= not G14775;
	I22560<= not G14796;
	I22563<= not G14830;
	I22566<= not G14883;
	I22569<= not G14955;
	I22572<= not G15019;
	I22575<= not G15092;
	I22578<= not G14746;
	I22581<= not G14766;
	I22584<= not G15989;
	I22587<= not G14684;
	I22590<= not G13863;
	I22593<= not G15876;
	I22599<= not G14966;
	I22604<= not G15080;
	I22611<= not G15055;
	I22618<= not G14630;
	I22626<= not G15151;
	I22640<= not G14650;
	I22651<= not G14677;
	I22657<= not G14657;
	I22663<= not G14711;
	I22667<= not G14642;
	I22671<= not G14691;
	I22676<= not G14630;
	I22679<= not G14669;
	I22683<= not G14725;
	I22687<= not G14650;
	I22690<= not G14703;
	I22694<= not G14753;
	I22699<= not G14677;
	I22702<= not G14737;
	I22715<= not G14711;
	I22718<= not G14657;
	I22726<= not G14642;
	I22730<= not G14691;
	I22737<= not G14630;
	I22741<= not G14669;
	I22745<= not G14725;
	I22752<= not G14657;
	I22755<= not G14650;
	I22759<= not G14703;
	I22763<= not G14753;
	I22768<= not G14691;
	I22771<= not G14677;
	I22775<= not G14737;
	I22783<= not G13572;
	I22786<= not G14725;
	I22789<= not G14711;
	I22797<= not G14165;
	I22800<= not G13581;
	I22803<= not G14753;
	I22810<= not G14280;
	I22813<= not G13601;
	I22820<= not G14402;
	I22823<= not G13613;
	I22828<= not G14514;
	I22836<= not G13571;
	I22842<= not G13580;
	I22845<= not G13579;
	I22852<= not G13600;
	I22855<= not G13588;
	I22860<= not G14885;
	I22866<= not G13612;
	I22869<= not G13608;
	I22875<= not G14966;
	I22881<= not G13622;
	I22893<= not G15055;
	I22912<= not G15151;
	I23253<= not G13741;
	I23274<= not G13741;
	I23287<= not G13741;
	I23292<= not G13741;
	I23309<= not G16132;
	I23314<= not G15720;
	I23317<= not G16181;
	I23323<= not G15664;
	I23326<= not G15758;
	I23329<= not G15760;
	I23335<= not G16412;
	I23338<= not G15721;
	I23341<= not G15784;
	I23345<= not G15723;
	I23348<= not G15786;
	I23351<= not G15788;
	I23358<= not G16442;
	I23361<= not G15759;
	I23364<= not G15805;
	I23368<= not G16446;
	I23371<= not G15761;
	I23374<= not G15807;
	I23377<= not G15763;
	I23380<= not G15809;
	I23383<= not G15811;
	I23386<= not G13469;
	I23392<= not G13476;
	I23395<= not G15785;
	I23398<= not G15820;
	I23403<= not G13478;
	I23406<= not G15787;
	I23409<= not G15822;
	I23412<= not G13482;
	I23415<= not G15789;
	I23418<= not G15824;
	I23421<= not G15791;
	I23424<= not G15826;
	I23430<= not G13494;
	I23433<= not G15806;
	I23436<= not G15832;
	I23442<= not G13495;
	I23445<= not G15808;
	I23448<= not G15834;
	I23451<= not G13497;
	I23454<= not G15810;
	I23457<= not G15836;
	I23460<= not G13501;
	I23463<= not G15812;
	I23466<= not G15838;
	I23472<= not G13510;
	I23475<= not G15821;
	I23478<= not G15844;
	I23487<= not G13511;
	I23490<= not G15823;
	I23493<= not G15846;
	I23498<= not G13512;
	I23501<= not G15825;
	I23504<= not G15848;
	I23507<= not G13514;
	I23510<= not G15827;
	I23513<= not G15850;
	I23518<= not G15856;
	I23521<= not G13518;
	I23524<= not G15833;
	I23527<= not G15858;
	I23530<= not G14885;
	I23539<= not G13524;
	I23542<= not G15835;
	I23545<= not G15867;
	I23553<= not G13525;
	I23556<= not G15837;
	I23559<= not G15869;
	I23564<= not G13526;
	I23567<= not G15839;
	I23570<= not G15871;
	I23575<= not G15843;
	I23578<= not G15879;
	I23581<= not G13528;
	I23584<= not G15845;
	I23588<= not G14885;
	I23591<= not G14885;
	I23599<= not G15887;
	I23602<= not G13529;
	I23605<= not G15847;
	I23608<= not G15889;
	I23611<= not G14966;
	I23619<= not G13535;
	I23622<= not G15849;
	I23625<= not G15898;
	I23633<= not G13536;
	I23636<= not G15851;
	I23639<= not G15900;
	I23645<= not G13537;
	I23648<= not G15857;
	I23651<= not G13538;
	I23655<= not G14831;
	I23658<= not G14885;
	I23661<= not G16085;
	I23667<= not G15866;
	I23670<= not G15912;
	I23673<= not G13539;
	I23676<= not G15868;
	I23679<= not G14966;
	I23682<= not G14966;
	I23689<= not G15920;
	I23692<= not G13540;
	I23695<= not G15870;
	I23698<= not G15922;
	I23701<= not G15055;
	I23709<= not G13546;
	I23712<= not G15872;
	I23715<= not G15931;
	I23725<= not G13547;
	I23729<= not G14337;
	I23733<= not G14831;
	I23739<= not G13548;
	I23742<= not G15888;
	I23745<= not G13549;
	I23748<= not G14904;
	I23751<= not G14966;
	I23754<= not G16123;
	I23760<= not G15897;
	I23763<= not G15941;
	I23766<= not G13550;
	I23769<= not G15899;
	I23772<= not G15055;
	I23775<= not G15055;
	I23782<= not G15949;
	I23785<= not G13551;
	I23788<= not G15901;
	I23791<= not G15951;
	I23794<= not G15151;
	I23817<= not G13557;
	I23821<= not G14337;
	I23824<= not G14904;
	I23830<= not G13558;
	I23833<= not G15921;
	I23836<= not G13559;
	I23839<= not G14985;
	I23842<= not G15055;
	I23845<= not G16174;
	I23851<= not G15930;
	I23854<= not G15970;
	I23857<= not G13560;
	I23860<= not G15932;
	I23863<= not G15151;
	I23866<= not G15151;
	I23874<= not G15797;
	I23888<= not G14685;
	I23904<= not G13561;
	I23908<= not G14337;
	I23911<= not G14985;
	I23917<= not G13562;
	I23920<= not G15950;
	I23923<= not G13563;
	I23926<= not G15074;
	I23929<= not G15151;
	I23932<= not G16233;
	I23954<= not G16154;
	I23976<= not G14719;
	I23992<= not G13564;
	I23996<= not G14337;
	I23999<= not G15074;
	I24049<= not G16213;
	I24071<= not G14747;
	I24144<= not G16278;
	I24166<= not G14768;
	I24171<= not G16439;
	I24247<= not G16337;
	I24258<= not G16463;
	I24285<= not G15992;
	I24346<= not G15873;
	I24368<= not G15990;
	I24394<= not G15995;
	I24459<= not G13599;
	I24481<= not G15993;
	I24507<= not G15999;
	I24560<= not G13611;
	I24582<= not G15996;
	I24608<= not G16006;
	I24662<= not G13621;
	I24684<= not G16000;
	I24732<= not G13633;
	I24894<= not G14797;
	I24913<= not G15800;
	I24916<= not G14776;
	I24923<= not G14849;
	I24943<= not G14811;
	I24950<= not G14922;
	I24966<= not G14863;
	I24973<= not G15003;
	I24982<= not G14347;
	I24992<= not G14936;
	I25001<= not G14244;
	I25004<= not G14459;
	I25015<= not G14158;
	I25018<= not G14366;
	I25021<= not G14546;
	I25037<= not G14071;
	I25041<= not G14895;
	I25044<= not G14273;
	I25047<= not G14478;
	I25050<= not G14601;
	I25054<= not G14837;
	I25057<= not G14186;
	I25061<= not G14976;
	I25064<= not G14395;
	I25067<= not G14565;
	I25071<= not G14910;
	I25074<= not G14301;
	I25078<= not G15065;
	I25081<= not G14507;
	I25084<= not G14885;
	I25089<= not G14991;
	I25092<= not G14423;
	I25096<= not G15161;
	I25099<= not G19000;
	I25102<= not G18944;
	I25105<= not G18959;
	I25108<= not G18969;
	I25111<= not G18981;
	I25114<= not G18983;
	I25117<= not G18988;
	I25120<= not G18869;
	I25123<= not G18890;
	I25126<= not G16858;
	I25129<= not G16813;
	I25132<= not G16862;
	I25135<= not G16506;
	I25138<= not G18960;
	I25141<= not G18970;
	I25144<= not G18984;
	I25147<= not G18989;
	I25150<= not G18991;
	I25153<= not G18995;
	I25156<= not G18895;
	I25159<= not G18913;
	I25162<= not G16863;
	I25165<= not G16831;
	I25168<= not G16877;
	I25171<= not G16528;
	I25174<= not G18971;
	I25177<= not G18985;
	I25180<= not G18992;
	I25183<= not G18996;
	I25186<= not G18998;
	I25189<= not G19008;
	I25192<= not G18918;
	I25195<= not G18932;
	I25198<= not G16878;
	I25201<= not G16843;
	I25204<= not G16905;
	I25207<= not G16559;
	I25210<= not G18986;
	I25213<= not G18993;
	I25216<= not G18999;
	I25219<= not G19009;
	I25222<= not G19011;
	I25225<= not G16514;
	I25228<= not G18937;
	I25231<= not G18952;
	I25234<= not G16906;
	I25237<= not G16849;
	I25240<= not G16934;
	I25243<= not G17227;
	I25246<= not G17233;
	I25249<= not G17300;
	I25253<= not G17124;
	I25258<= not G16974;
	I25264<= not G17151;
	I25272<= not G17051;
	I25283<= not G17086;
	I25294<= not G17124;
	I25303<= not G17151;
	I25308<= not G16867;
	I25315<= not G16895;
	I25320<= not G16924;
	I25325<= not G16954;
	I25334<= not G17645;
	I25338<= not G17746;
	I25344<= not G17847;
	I25351<= not G17959;
	I25355<= not G18669;
	I25358<= not G18678;
	I25365<= not G18707;
	I25371<= not G18719;
	I25374<= not G18726;
	I25377<= not G18743;
	I25383<= not G18755;
	I25386<= not G18763;
	I25389<= not G18780;
	I25395<= not G18782;
	I25399<= not G18794;
	I25402<= not G18821;
	I25406<= not G18804;
	I25412<= not G18820;
	I25415<= not G18835;
	I25423<= not G18852;
	I25426<= not G18836;
	I25429<= not G18975;
	I25432<= not G18837;
	I25442<= not G18866;
	I25445<= not G18968;
	I25456<= not G18883;
	I25459<= not G18867;
	I25463<= not G18868;
	I25474<= not G18885;
	I25486<= not G18754;
	I25489<= not G18906;
	I25492<= not G18907;
	I25506<= not G18781;
	I25510<= not G18542;
	I25525<= not G18803;
	I25528<= not G18942;
	I25557<= not G18957;
	I25567<= not G17186;
	I25612<= not G17197;
	I25660<= not G17204;
	I25717<= not G17209;
	I25728<= not G17118;
	I25768<= not G17139;
	I25778<= not G17145;
	I25816<= not G17162;
	I25826<= not G17168;
	I25862<= not G17177;
	I25872<= not G17183;
	I25904<= not G17194;
	I25966<= not G16654;
	I25971<= not G16671;
	I25977<= not G16692;
	I25985<= not G16718;
	I25994<= not G16860;
	I26006<= not G16866;
	I26025<= not G16803;
	I26028<= not G16566;
	I26051<= not G16824;
	I26078<= not G16835;
	I26085<= not G18085;
	I26112<= not G16844;
	I26115<= not G16845;
	I26123<= not G17503;
	I26134<= not G18201;
	I26154<= not G16851;
	I26171<= not G17594;
	I26182<= not G18308;
	I26195<= not G16853;
	I26198<= not G16854;
	I26220<= not G17691;
	I26231<= not G18401;
	I26237<= not G16857;
	I26266<= not G17791;
	I26276<= not G16861;
	I26334<= not G18977;
	I26337<= not G16880;
	I26340<= not G17025;
	I26365<= not G18626;
	I26369<= not G17059;
	I26388<= not G17094;
	I26401<= not G17012;
	I26407<= not G17132;
	I26413<= not G16643;
	I26420<= not G17042;
	I26426<= not G16536;
	I26437<= not G16655;
	I26444<= not G17076;
	I26458<= not G17985;
	I26469<= not G16672;
	I26476<= not G17111;
	I26481<= not G18590;
	I26494<= not G18102;
	I26505<= not G16693;
	I26512<= not G16802;
	I26535<= not G18218;
	I26545<= not G16823;
	I26574<= not G18325;
	I26612<= not G17645;
	I26642<= not G17746;
	I26664<= not G17847;
	I26679<= not G17959;
	I26714<= not G17720;
	I26777<= not G17222;
	I26796<= not G17224;
	I26816<= not G17225;
	I26819<= not G17226;
	I26843<= not G17228;
	I26846<= not G17229;
	I26868<= not G17234;
	I26871<= not G17235;
	I26874<= not G17236;
	I26892<= not G17246;
	I26895<= not G17247;
	I26898<= not G17248;
	I26910<= not G17269;
	I26913<= not G17270;
	I26916<= not G17271;
	I26923<= not G17302;
	I26926<= not G17303;
	I26931<= not G17340;
	I26934<= not G17341;
	I26940<= not G17383;
	I26947<= not G17429;
	I26960<= not G16884;
	I26966<= not G17051;
	I26972<= not G16913;
	I26980<= not G17086;
	I26985<= not G16943;
	I26990<= not G19145;
	I26993<= not G19159;
	I26996<= not G19169;
	I26999<= not G19543;
	I27002<= not G19147;
	I27005<= not G19164;
	I27008<= not G19175;
	I27011<= not G19546;
	I27014<= not G19151;
	I27017<= not G19170;
	I27020<= not G19182;
	I27023<= not G19550;
	I27026<= not G19156;
	I27029<= not G19176;
	I27032<= not G19189;
	I27035<= not G19556;
	I27038<= not G20082;
	I27041<= not G19237;
	I27044<= not G19247;
	I27047<= not G19258;
	I27050<= not G19183;
	I27053<= not G19190;
	I27056<= not G19196;
	I27059<= not G19207;
	I27062<= not G19217;
	I27065<= not G19270;
	I27068<= not G19197;
	I27071<= not G19218;
	I27074<= not G19238;
	I27077<= not G19259;
	I27080<= not G19198;
	I27083<= not G19208;
	I27086<= not G19229;
	I27089<= not G20105;
	I27092<= not G19174;
	I27095<= not G19185;
	I27098<= not G19199;
	I27101<= not G19220;
	I27104<= not G19239;
	I27107<= not G19249;
	I27110<= not G19622;
	I27113<= not G19689;
	I27116<= not G19762;
	I27119<= not G19563;
	I27122<= not G19595;
	I27125<= not G19652;
	I27128<= not G19725;
	I27131<= not G19798;
	I27134<= not G19573;
	I27137<= not G19596;
	I27140<= not G19690;
	I27143<= not G19763;
	I27146<= not G19838;
	I27149<= not G19893;
	I27152<= not G20360;
	I27155<= not G20395;
	I27158<= not G20439;
	I27161<= not G20377;
	I27164<= not G20418;
	I27167<= not G20457;
	I27170<= not G20396;
	I27173<= not G20440;
	I27176<= not G20469;
	I27179<= not G20419;
	I27182<= not G20458;
	I27185<= not G20478;
	I27188<= not G20441;
	I27191<= not G20470;
	I27194<= not G20484;
	I27197<= not G20459;
	I27200<= not G20479;
	I27203<= not G20491;
	I27206<= not G20471;
	I27209<= not G20485;
	I27212<= not G20498;
	I27215<= not G19158;
	I27218<= not G19168;
	I27221<= not G19180;
	I27225<= not G19358;
	I27228<= not G19390;
	I27232<= not G19401;
	I27235<= not G19420;
	I27240<= not G19335;
	I27243<= not G19335;
	I27246<= not G19335;
	I27250<= not G19390;
	I27253<= not G19420;
	I27257<= not G19431;
	I27260<= not G19457;
	I27264<= not G19358;
	I27267<= not G19358;
	I27270<= not G19335;
	I27275<= not G19369;
	I27278<= not G19369;
	I27281<= not G19369;
	I27285<= not G19420;
	I27288<= not G19457;
	I27293<= not G19335;
	I27297<= not G19390;
	I27300<= not G19390;
	I27303<= not G19369;
	I27308<= not G19401;
	I27311<= not G19401;
	I27314<= not G19401;
	I27318<= not G19457;
	I27321<= not G19335;
	I27324<= not G19358;
	I27328<= not G19369;
	I27332<= not G19420;
	I27335<= not G19420;
	I27338<= not G19401;
	I27343<= not G19431;
	I27346<= not G19431;
	I27349<= not G19431;
	I27352<= not G19358;
	I27355<= not G19335;
	I27358<= not G19369;
	I27361<= not G19390;
	I27365<= not G19401;
	I27369<= not G19457;
	I27372<= not G19457;
	I27375<= not G19431;
	I27379<= not G19358;
	I27382<= not G19390;
	I27385<= not G19369;
	I27388<= not G19401;
	I27391<= not G19420;
	I27395<= not G19431;
	I27399<= not G19390;
	I27402<= not G19420;
	I27405<= not G19401;
	I27408<= not G19431;
	I27411<= not G19457;
	I27416<= not G19420;
	I27419<= not G19457;
	I27422<= not G19431;
	I27426<= not G19457;
	I27488<= not G20310;
	I27491<= not G20314;
	I27516<= not G20333;
	I27531<= not G20343;
	I27534<= not G20083;
	I27537<= not G19957;
	I27549<= not G20353;
	I27565<= not G19987;
	I27577<= not G20375;
	I27585<= not G20376;
	I27593<= not G20025;
	I27614<= not G20067;
	I27621<= not G20417;
	I27646<= not G20507;
	I27658<= not G20526;
	I27667<= not G20507;
	I27672<= not G20545;
	I27684<= not G20526;
	I27689<= not G19070;
	I27705<= not G20545;
	I27727<= not G19070;
	I27749<= not G19954;
	I27766<= not G19984;
	I27779<= not G20022;
	I27785<= not G20064;
	I27822<= not G19865;
	I27827<= not G19896;
	I27832<= not G19921;
	I27838<= not G19936;
	I27868<= not G19144;
	I27897<= not G19149;
	I27900<= not G19096;
	I27917<= not G19153;
	I27920<= not G19154;
	I27927<= not G19957;
	I27942<= not G19157;
	I27949<= not G19957;
	I27958<= not G19987;
	I27969<= not G19162;
	I27972<= not G19163;
	I27976<= not G19957;
	I27984<= not G19987;
	I27992<= not G20025;
	I28000<= not G19167;
	I28003<= not G19957;
	I28009<= not G20473;
	I28013<= not G19987;
	I28019<= not G20025;
	I28027<= not G20067;
	I28031<= not G19172;
	I28034<= not G19173;
	I28038<= not G19957;
	I28043<= not G19987;
	I28047<= not G20481;
	I28051<= not G20025;
	I28057<= not G20067;
	I28061<= not G19178;
	I28065<= not G19957;
	I28072<= not G19987;
	I28076<= not G20025;
	I28080<= not G20487;
	I28084<= not G20067;
	I28087<= not G19184;
	I28090<= not G20008;
	I28093<= not G19957;
	I28100<= not G19987;
	I28107<= not G20025;
	I28111<= not G20067;
	I28115<= not G20493;
	I28119<= not G19957;
	I28123<= not G19987;
	I28130<= not G20025;
	I28137<= not G20067;
	I28143<= not G19957;
	I28148<= not G19987;
	I28152<= not G20025;
	I28159<= not G20067;
	I28169<= not G19987;
	I28174<= not G20025;
	I28178<= not G20067;
	I28184<= not G19103;
	I28201<= not G20025;
	I28206<= not G20067;
	I28210<= not G20537;
	I28229<= not G20067;
	I28235<= not G20153;
	I28314<= not G19152;
	I28357<= not G20497;
	I28360<= not G20163;
	I28432<= not G19335;
	I28435<= not G19358;
	I28443<= not G19358;
	I28447<= not G19369;
	I28450<= not G19390;
	I28455<= not G20943;
	I28458<= not G20971;
	I28461<= not G20998;
	I28464<= not G21024;
	I28467<= not G20942;
	I28470<= not G20984;
	I28473<= not G21030;
	I28476<= not G21064;
	I28479<= not G21795;
	I28482<= not G21376;
	I28485<= not G21426;
	I28488<= not G21495;
	I28491<= not G21327;
	I28494<= not G21358;
	I28497<= not G21399;
	I28500<= not G21457;
	I28503<= not G21528;
	I28506<= not G21377;
	I28509<= not G21427;
	I28512<= not G21496;
	I28515<= not G21557;
	I28518<= not G20985;
	I28521<= not G21824;
	I28524<= not G21359;
	I28527<= not G21407;
	I28541<= not G21467;
	I28550<= not G21432;
	I28557<= not G21407;
	I28564<= not G21385;
	I28628<= not G21842;
	I28649<= not G21843;
	I28671<= not G21845;
	I28693<= not G21847;
	I28712<= not G21851;
	I28781<= not G21331;
	I28789<= not G21878;
	I28792<= not G21880;
	I28800<= not G21316;
	I28813<= not G21502;
	I28825<= not G21882;
	I28833<= not G21470;
	I28876<= not G21238;
	I28896<= not G21246;
	I28913<= not G21255;
	I28928<= not G21263;
	I28949<= not G21685;
	I28953<= not G21659;
	I28956<= not G21714;
	I28959<= not G21636;
	I28962<= not G21721;
	I28966<= not G20633;
	I28969<= not G21686;
	I28972<= not G21736;
	I28975<= not G21688;
	I28978<= not G21740;
	I28981<= not G21667;
	I28984<= not G21747;
	I28988<= not G20874;
	I28991<= not G20648;
	I28994<= not G21715;
	I28997<= not G21759;
	I29001<= not G20658;
	I29004<= not G21722;
	I29007<= not G21760;
	I29010<= not G21724;
	I29013<= not G21764;
	I29016<= not G21696;
	I29019<= not G21771;
	I29023<= not G20672;
	I29026<= not G21737;
	I29030<= not G20683;
	I29033<= not G21741;
	I29036<= not G21775;
	I29040<= not G20693;
	I29043<= not G21748;
	I29046<= not G21776;
	I29049<= not G21750;
	I29052<= not G21780;
	I29055<= not G21732;
	I29058<= not G20703;
	I29064<= not G20875;
	I29067<= not G20876;
	I29070<= not G20707;
	I29073<= not G21761;
	I29077<= not G20718;
	I29080<= not G21765;
	I29083<= not G21790;
	I29087<= not G20728;
	I29090<= not G21772;
	I29093<= not G21791;
	I29098<= not G20879;
	I29101<= not G20880;
	I29104<= not G20881;
	I29107<= not G21435;
	I29110<= not G20738;
	I29116<= not G20882;
	I29119<= not G20883;
	I29122<= not G20742;
	I29125<= not G21777;
	I29129<= not G20753;
	I29132<= not G21781;
	I29135<= not G21804;
	I29142<= not G20682;
	I29145<= not G20891;
	I29148<= not G20892;
	I29151<= not G20893;
	I29154<= not G20894;
	I29159<= not G20896;
	I29162<= not G20897;
	I29165<= not G20898;
	I29168<= not G20775;
	I29174<= not G20899;
	I29177<= not G20900;
	I29180<= not G20779;
	I29183<= not G21792;
	I29191<= not G20901;
	I29194<= not G20902;
	I29197<= not G20903;
	I29203<= not G20717;
	I29206<= not G20910;
	I29209<= not G20911;
	I29212<= not G20912;
	I29215<= not G20913;
	I29220<= not G20915;
	I29223<= not G20916;
	I29226<= not G20917;
	I29229<= not G20805;
	I29235<= not G20918;
	I29238<= not G20919;
	I29243<= not G20921;
	I29246<= not G20922;
	I29249<= not G20923;
	I29252<= not G20924;
	I29259<= not G20925;
	I29262<= not G20926;
	I29265<= not G20927;
	I29271<= not G20752;
	I29274<= not G20934;
	I29277<= not G20935;
	I29280<= not G20936;
	I29283<= not G20937;
	I29288<= not G20939;
	I29291<= not G20940;
	I29294<= not G20941;
	I29301<= not G20944;
	I29304<= not G20945;
	I29307<= not G20946;
	I29310<= not G20947;
	I29313<= not G20948;
	I29317<= not G20949;
	I29320<= not G20950;
	I29323<= not G20951;
	I29326<= not G20952;
	I29333<= not G20953;
	I29336<= not G20954;
	I29339<= not G20955;
	I29345<= not G20789;
	I29348<= not G20962;
	I29351<= not G20963;
	I29354<= not G20964;
	I29357<= not G20965;
	I29360<= not G21796;
	I29366<= not G20966;
	I29369<= not G20967;
	I29372<= not G20968;
	I29375<= not G20969;
	I29378<= not G20970;
	I29383<= not G20972;
	I29386<= not G20973;
	I29389<= not G20974;
	I29392<= not G20975;
	I29395<= not G20976;
	I29399<= not G20977;
	I29402<= not G20978;
	I29405<= not G20979;
	I29408<= not G20980;
	I29415<= not G20981;
	I29418<= not G20982;
	I29421<= not G20983;
	I29426<= not G20989;
	I29429<= not G20990;
	I29432<= not G20991;
	I29435<= not G20992;
	I29439<= not G20993;
	I29442<= not G20994;
	I29445<= not G20995;
	I29448<= not G20996;
	I29451<= not G20997;
	I29456<= not G20999;
	I29459<= not G21000;
	I29462<= not G21001;
	I29465<= not G21002;
	I29468<= not G21003;
	I29472<= not G21004;
	I29475<= not G21005;
	I29478<= not G21006;
	I29481<= not G21007;
	I29484<= not G21903;
	I29490<= not G21009;
	I29493<= not G21010;
	I29496<= not G21011;
	I29500<= not G21015;
	I29503<= not G21016;
	I29506<= not G21017;
	I29509<= not G21018;
	I29513<= not G21019;
	I29516<= not G21020;
	I29519<= not G21021;
	I29522<= not G21022;
	I29525<= not G21023;
	I29530<= not G21025;
	I29533<= not G21026;
	I29536<= not G21027;
	I29539<= not G21028;
	I29542<= not G21029;
	I29547<= not G21031;
	I29550<= not G21032;
	I29556<= not G21033;
	I29559<= not G21034;
	I29562<= not G21035;
	I29566<= not G21039;
	I29569<= not G21040;
	I29572<= not G21041;
	I29575<= not G21042;
	I29579<= not G21043;
	I29582<= not G21044;
	I29585<= not G21045;
	I29588<= not G21046;
	I29591<= not G21047;
	I29600<= not G21720;
	I29603<= not G21051;
	I29606<= not G21364;
	I29610<= not G21052;
	I29613<= not G21053;
	I29619<= not G21054;
	I29622<= not G21055;
	I29625<= not G21056;
	I29629<= not G21060;
	I29632<= not G21061;
	I29635<= not G21062;
	I29638<= not G21063;
	I29641<= not G20825;
	I29653<= not G21746;
	I29656<= not G21070;
	I29660<= not G21071;
	I29663<= not G21072;
	I29669<= not G21073;
	I29672<= not G21074;
	I29675<= not G21075;
	I29687<= not G21770;
	I29690<= not G21080;
	I29694<= not G21081;
	I29697<= not G21082;
	I29700<= not G20700;
	I29712<= not G21786;
	I29715<= not G21094;
	I29724<= not G21851;
	I29727<= not G20877;
	I29736<= not G20884;
	I29741<= not G21346;
	I29797<= not G21432;
	I29802<= not G21435;
	I29812<= not G21467;
	I29817<= not G21470;
	I29827<= not G21502;
	I29841<= not G21316;
	I29852<= not G21331;
	I29863<= not G21346;
	I29872<= not G21364;
	I29881<= not G21385;
	I29897<= not G23116;
	I29900<= not G23125;
	I29903<= not G23134;
	I29906<= not G21967;
	I29909<= not G23050;
	I29912<= not G23065;
	I29915<= not G23055;
	I29918<= not G23068;
	I29921<= not G23078;
	I29924<= not G23094;
	I29927<= not G23105;
	I29930<= not G22176;
	I29933<= not G22082;
	I29936<= not G22582;
	I29939<= not G22518;
	I29942<= not G22548;
	I29945<= not G22583;
	I29948<= not G22549;
	I29951<= not G22584;
	I29954<= not G22611;
	I29957<= not G22585;
	I29960<= not G22612;
	I29963<= not G22639;
	I29966<= not G22613;
	I29969<= not G22640;
	I29972<= not G22669;
	I29975<= not G22641;
	I29978<= not G22670;
	I29981<= not G22702;
	I29984<= not G22671;
	I29987<= not G22703;
	I29990<= not G22728;
	I29993<= not G22704;
	I29996<= not G22729;
	I29999<= not G22756;
	I30002<= not G22730;
	I30005<= not G22757;
	I30008<= not G22785;
	I30011<= not G22758;
	I30014<= not G22786;
	I30017<= not G22824;
	I30020<= not G22519;
	I30023<= not G22550;
	I30026<= not G22586;
	I30029<= not G22642;
	I30032<= not G22672;
	I30035<= not G22705;
	I30038<= not G22673;
	I30041<= not G22706;
	I30044<= not G22731;
	I30047<= not G22107;
	I30050<= not G22619;
	I30053<= not G22558;
	I30056<= not G22589;
	I30059<= not G22620;
	I30062<= not G22590;
	I30065<= not G22621;
	I30068<= not G22647;
	I30071<= not G22622;
	I30074<= not G22648;
	I30077<= not G22675;
	I30080<= not G22649;
	I30083<= not G22676;
	I30086<= not G22709;
	I30089<= not G22677;
	I30092<= not G22710;
	I30095<= not G22733;
	I30098<= not G22711;
	I30101<= not G22734;
	I30104<= not G22760;
	I30107<= not G22735;
	I30110<= not G22761;
	I30113<= not G22790;
	I30116<= not G22762;
	I30119<= not G22791;
	I30122<= not G22827;
	I30125<= not G22792;
	I30128<= not G22828;
	I30131<= not G22864;
	I30134<= not G22559;
	I30137<= not G22591;
	I30140<= not G22623;
	I30143<= not G22678;
	I30146<= not G22712;
	I30149<= not G22736;
	I30152<= not G22713;
	I30155<= not G22737;
	I30158<= not G22763;
	I30161<= not G22133;
	I30164<= not G22655;
	I30167<= not G22598;
	I30170<= not G22626;
	I30173<= not G22656;
	I30176<= not G22627;
	I30179<= not G22657;
	I30182<= not G22683;
	I30185<= not G22658;
	I30188<= not G22684;
	I30191<= not G22715;
	I30194<= not G22685;
	I30197<= not G22716;
	I30200<= not G22740;
	I30203<= not G22717;
	I30206<= not G22741;
	I30209<= not G22765;
	I30212<= not G22742;
	I30215<= not G22766;
	I30218<= not G22794;
	I30221<= not G22767;
	I30224<= not G22795;
	I30227<= not G22832;
	I30230<= not G22796;
	I30233<= not G22833;
	I30236<= not G22866;
	I30239<= not G22834;
	I30242<= not G22867;
	I30245<= not G22899;
	I30248<= not G22599;
	I30251<= not G22628;
	I30254<= not G22659;
	I30257<= not G22718;
	I30260<= not G22743;
	I30263<= not G22768;
	I30266<= not G22744;
	I30269<= not G22769;
	I30272<= not G22797;
	I30275<= not G22156;
	I30278<= not G22691;
	I30281<= not G22635;
	I30284<= not G22662;
	I30287<= not G22692;
	I30290<= not G22663;
	I30293<= not G22693;
	I30296<= not G22723;
	I30299<= not G22694;
	I30302<= not G22724;
	I30305<= not G22746;
	I30308<= not G22725;
	I30311<= not G22747;
	I30314<= not G22772;
	I30317<= not G22748;
	I30320<= not G22773;
	I30323<= not G22799;
	I30326<= not G22774;
	I30329<= not G22800;
	I30332<= not G22836;
	I30335<= not G22801;
	I30338<= not G22837;
	I30341<= not G22871;
	I30344<= not G22838;
	I30347<= not G22872;
	I30350<= not G22901;
	I30353<= not G22873;
	I30356<= not G22902;
	I30359<= not G22934;
	I30362<= not G22636;
	I30365<= not G22664;
	I30368<= not G22695;
	I30371<= not G22749;
	I30374<= not G22775;
	I30377<= not G22802;
	I30380<= not G22776;
	I30383<= not G22803;
	I30386<= not G22839;
	I30389<= not G22225;
	I30392<= not G22226;
	I30395<= not G22253;
	I30398<= not G22840;
	I30401<= not G22444;
	I30404<= not G22948;
	I30407<= not G22970;
	I30467<= not G23000;
	I30470<= not G23117;
	I30476<= not G22876;
	I30480<= not G23014;
	I30483<= not G23126;
	I30486<= not G23022;
	I30489<= not G22911;
	I30493<= not G23030;
	I30496<= not G23137;
	I30501<= not G23039;
	I30504<= not G22936;
	I30508<= not G23047;
	I30511<= not G21970;
	I30516<= not G23058;
	I30519<= not G22942;
	I30525<= not G23067;
	I30531<= not G23076;
	I30536<= not G23081;
	I30544<= not G23092;
	I30547<= not G23093;
	I30552<= not G23097;
	I30560<= not G23110;
	I30563<= not G23111;
	I30568<= not G23114;
	I30575<= not G23123;
	I30578<= not G23124;
	I30586<= not G23132;
	I30589<= not G23133;
	I30594<= not G22025;
	I30598<= not G22027;
	I30601<= not G22028;
	I30607<= not G22029;
	I30611<= not G22030;
	I30614<= not G22031;
	I30617<= not G22032;
	I30623<= not G22033;
	I30626<= not G22034;
	I30632<= not G22035;
	I30636<= not G22037;
	I30639<= not G22038;
	I30642<= not G22039;
	I30648<= not G22040;
	I30651<= not G22041;
	I30654<= not G22042;
	I30660<= not G22043;
	I30663<= not G22044;
	I30669<= not G22045;
	I30673<= not G22047;
	I30676<= not G22048;
	I30679<= not G22049;
	I30686<= not G23136;
	I30689<= not G22054;
	I30692<= not G22055;
	I30695<= not G22056;
	I30701<= not G22057;
	I30704<= not G22058;
	I30707<= not G22059;
	I30713<= not G22060;
	I30716<= not G22061;
	I30722<= not G22063;
	I30725<= not G22064;
	I30728<= not G22065;
	I30735<= not G22066;
	I30738<= not G22067;
	I30741<= not G22068;
	I30748<= not G21969;
	I30751<= not G22073;
	I30754<= not G22074;
	I30757<= not G22075;
	I30763<= not G22076;
	I30766<= not G22077;
	I30769<= not G22078;
	I30776<= not G22079;
	I30779<= not G22080;
	I30782<= not G22081;
	I30786<= not G22454;
	I30797<= not G22087;
	I30800<= not G22088;
	I30803<= not G22089;
	I30810<= not G22090;
	I30813<= not G22091;
	I30816<= not G22092;
	I30823<= not G21972;
	I30826<= not G22097;
	I30829<= not G22098;
	I30832<= not G22099;
	I30838<= not G22100;
	I30841<= not G22101;
	I30844<= not G22102;
	I30847<= not G22103;
	I30854<= not G22104;
	I30857<= not G22105;
	I30860<= not G22106;
	I30864<= not G22493;
	I30875<= not G22112;
	I30878<= not G22113;
	I30881<= not G22114;
	I30888<= not G22115;
	I30891<= not G22116;
	I30894<= not G22117;
	I30901<= not G21974;
	I30905<= not G22122;
	I30908<= not G22123;
	I30911<= not G22124;
	I30914<= not G22125;
	I30917<= not G22806;
	I30922<= not G22126;
	I30925<= not G22127;
	I30928<= not G22128;
	I30931<= not G22129;
	I30938<= not G22130;
	I30941<= not G22131;
	I30944<= not G22132;
	I30948<= not G22536;
	I30959<= not G22138;
	I30962<= not G22139;
	I30965<= not G22140;
	I30973<= not G22141;
	I30976<= not G22142;
	I30979<= not G22143;
	I30985<= not G22992;
	I30988<= not G22145;
	I30991<= not G22146;
	I30994<= not G22147;
	I30997<= not G22148;
	I31000<= not G22847;
	I31005<= not G22149;
	I31008<= not G22150;
	I31011<= not G22151;
	I31014<= not G22152;
	I31021<= not G22153;
	I31024<= not G22154;
	I31027<= not G22155;
	I31031<= not G22576;
	I31043<= not G22161;
	I31050<= not G22162;
	I31053<= not G22163;
	I31056<= not G22164;
	I31062<= not G23003;
	I31065<= not G22166;
	I31068<= not G22167;
	I31071<= not G22168;
	I31074<= not G22169;
	I31077<= not G22882;
	I31082<= not G22170;
	I31085<= not G22171;
	I31088<= not G22172;
	I31091<= not G22173;
	I31102<= not G22177;
	I31109<= not G22178;
	I31112<= not G22179;
	I31115<= not G22180;
	I31121<= not G23017;
	I31124<= not G22182;
	I31127<= not G22183;
	I31130<= not G22184;
	I31133<= not G22185;
	I31136<= not G22917;
	I31141<= not G22777;
	I31144<= not G22935;
	I31152<= not G22191;
	I31159<= not G22192;
	I31162<= not G22193;
	I31165<= not G22194;
	I31171<= not G23033;
	I31181<= not G22200;
	I31188<= not G21989;
	I31195<= not G22578;
	I31205<= not G22002;
	I31213<= not G22615;
	I31226<= not G22651;
	I31232<= not G22026;
	I31235<= not G22218;
	I31244<= not G22687;
	I31250<= not G22953;
	I31253<= not G22231;
	I31257<= not G22234;
	I31266<= not G22242;
	I31270<= not G22247;
	I31274<= not G22249;
	I31282<= not G22263;
	I31286<= not G22267;
	I31290<= not G22269;
	I31298<= not G22280;
	I31302<= not G22284;
	I31310<= not G22299;
	I31387<= not G22811;
	I31417<= not G22578;
	I31426<= not G22615;
	I31436<= not G22651;
	I31445<= not G22687;
	I31451<= not G23682;
	I31454<= not G23727;
	I31457<= not G23773;
	I31460<= not G23728;
	I31463<= not G23774;
	I31466<= not G23821;
	I31469<= not G23546;
	I31472<= not G23548;
	I31475<= not G23555;
	I31478<= not G23549;
	I31481<= not G23556;
	I31484<= not G23568;
	I31487<= not G23557;
	I31490<= not G23569;
	I31493<= not G23587;
	I31496<= not G23570;
	I31499<= not G23588;
	I31502<= not G23612;
	I31505<= not G23589;
	I31508<= not G23613;
	I31511<= not G23640;
	I31514<= not G23614;
	I31517<= not G23641;
	I31520<= not G23683;
	I31523<= not G23642;
	I31526<= not G23684;
	I31529<= not G23729;
	I31532<= not G23685;
	I31535<= not G23730;
	I31538<= not G23775;
	I31541<= not G23500;
	I31544<= not G23438;
	I31547<= not G23454;
	I31550<= not G23481;
	I31553<= not G23501;
	I31556<= not G23439;
	I31559<= not G24233;
	I31562<= not G23594;
	I31565<= not G24001;
	I31568<= not G24033;
	I31571<= not G24051;
	I31574<= not G23736;
	I31577<= not G23782;
	I31580<= not G23826;
	I31583<= not G23783;
	I31586<= not G23827;
	I31589<= not G23856;
	I31592<= not G23553;
	I31595<= not G23561;
	I31598<= not G23574;
	I31601<= not G23562;
	I31604<= not G23575;
	I31607<= not G23595;
	I31610<= not G23576;
	I31613<= not G23596;
	I31616<= not G23619;
	I31619<= not G23597;
	I31622<= not G23620;
	I31625<= not G23661;
	I31628<= not G23621;
	I31631<= not G23662;
	I31634<= not G23690;
	I31637<= not G23663;
	I31640<= not G23691;
	I31643<= not G23737;
	I31646<= not G23692;
	I31649<= not G23738;
	I31652<= not G23784;
	I31655<= not G23739;
	I31658<= not G23785;
	I31661<= not G23828;
	I31664<= not G23516;
	I31667<= not G23452;
	I31670<= not G23463;
	I31673<= not G23492;
	I31676<= not G23517;
	I31679<= not G23453;
	I31682<= not G24240;
	I31685<= not G23626;
	I31688<= not G24035;
	I31691<= not G24053;
	I31694<= not G24064;
	I31697<= not G23791;
	I31700<= not G23835;
	I31703<= not G23861;
	I31706<= not G23836;
	I31709<= not G23862;
	I31712<= not G23890;
	I31715<= not G23566;
	I31718<= not G23580;
	I31721<= not G23601;
	I31724<= not G23581;
	I31727<= not G23602;
	I31730<= not G23627;
	I31733<= not G23603;
	I31736<= not G23628;
	I31739<= not G23668;
	I31742<= not G23629;
	I31745<= not G23669;
	I31748<= not G23711;
	I31751<= not G23670;
	I31754<= not G23712;
	I31757<= not G23744;
	I31760<= not G23713;
	I31763<= not G23745;
	I31766<= not G23792;
	I31769<= not G23746;
	I31772<= not G23793;
	I31775<= not G23837;
	I31778<= not G23794;
	I31781<= not G23838;
	I31784<= not G23863;
	I31787<= not G23531;
	I31790<= not G23459;
	I31793<= not G23472;
	I31796<= not G23508;
	I31799<= not G23532;
	I31802<= not G23460;
	I31805<= not G24248;
	I31808<= not G23675;
	I31811<= not G24055;
	I31814<= not G24066;
	I31817<= not G24077;
	I31820<= not G23844;
	I31823<= not G23870;
	I31826<= not G23895;
	I31829<= not G23871;
	I31832<= not G23896;
	I31835<= not G23911;
	I31838<= not G23585;
	I31841<= not G23607;
	I31844<= not G23633;
	I31847<= not G23608;
	I31850<= not G23634;
	I31853<= not G23676;
	I31856<= not G23635;
	I31859<= not G23677;
	I31862<= not G23718;
	I31865<= not G23678;
	I31868<= not G23719;
	I31871<= not G23765;
	I31874<= not G23720;
	I31877<= not G23766;
	I31880<= not G23799;
	I31883<= not G23767;
	I31886<= not G23800;
	I31889<= not G23845;
	I31892<= not G23801;
	I31895<= not G23846;
	I31898<= not G23872;
	I31901<= not G23847;
	I31904<= not G23873;
	I31907<= not G23897;
	I31910<= not G23542;
	I31913<= not G23468;
	I31916<= not G23485;
	I31919<= not G23524;
	I31922<= not G23543;
	I31925<= not G23469;
	I31928<= not G24255;
	I31931<= not G23725;
	I31934<= not G24068;
	I31937<= not G24079;
	I31940<= not G24088;
	I31943<= not G24000;
	I31946<= not G23916;
	I31949<= not G23943;
	I32042<= not G23399;
	I32057<= not G23406;
	I32067<= not G24174;
	I32074<= not G23413;
	I32081<= not G24178;
	I32085<= not G24179;
	I32092<= not G23418;
	I32098<= not G24181;
	I32102<= not G24182;
	I32109<= not G24206;
	I32112<= not G24207;
	I32116<= not G24208;
	I32120<= not G24209;
	I32126<= not G24212;
	I32129<= not G24213;
	I32133<= not G24214;
	I32137<= not G24215;
	I32140<= not G24216;
	I32143<= not G24218;
	I32146<= not G24219;
	I32150<= not G24222;
	I32153<= not G24223;
	I32156<= not G24225;
	I32159<= not G24226;
	I32164<= not G24228;
	I32167<= not G24230;
	I32170<= not G24231;
	I32175<= not G24235;
	I32178<= not G24237;
	I32181<= not G24238;
	I32184<= not G23497;
	I32189<= not G24243;
	I32193<= not G23513;
	I32198<= not G24250;
	I32203<= not G23528;
	I32210<= not G23539;
	I32248<= not G23919;
	I32251<= not G23919;
	I32281<= not G23950;
	I32320<= not G23979;
	I32365<= not G24009;
	I32388<= not G23385;
	I32419<= not G24043;
	I32439<= not G23392;
	I32487<= not G23400;
	I32506<= not G23324;
	I32535<= not G23407;
	I32556<= not G23329;
	I32583<= not G23330;
	I32604<= not G23339;
	I32642<= not G23348;
	I32704<= not G23357;
	I32716<= not G23358;
	I32719<= not G23359;
	I32829<= not G24059;
	I32835<= not G24072;
	I32844<= not G23644;
	I32847<= not G24083;
	I32851<= not G23694;
	I32854<= not G24092;
	I32857<= not G23748;
	I32860<= not G23803;
	I32868<= not G25118;
	I32871<= not G24518;
	I32874<= not G24539;
	I32877<= not G24567;
	I32880<= not G24581;
	I32883<= not G24592;
	I32886<= not G24549;
	I32889<= not G24568;
	I32892<= not G24582;
	I32895<= not G24816;
	I32898<= not G24856;
	I32901<= not G25121;
	I32904<= not G24531;
	I32907<= not G24551;
	I32910<= not G24576;
	I32913<= not G24586;
	I32916<= not G24597;
	I32919<= not G24560;
	I32922<= not G24577;
	I32925<= not G24587;
	I32928<= not G24835;
	I32931<= not G24872;
	I32934<= not G25123;
	I32937<= not G24544;
	I32940<= not G24562;
	I32943<= not G24583;
	I32946<= not G24593;
	I32949<= not G24605;
	I32952<= not G24570;
	I32955<= not G24584;
	I32958<= not G24594;
	I32961<= not G24851;
	I32964<= not G24886;
	I32967<= not G25124;
	I32970<= not G24556;
	I32973<= not G24572;
	I32976<= not G24588;
	I32979<= not G24598;
	I32982<= not G24612;
	I32985<= not G24579;
	I32988<= not G24589;
	I32991<= not G24599;
	I32994<= not G24865;
	I32997<= not G24903;
	I33000<= not G24949;
	I33003<= not G24956;
	I33006<= not G24957;
	I33009<= not G24879;
	I33013<= not G25119;
	I33016<= not G25122;
	I33128<= not G24975;
	I33136<= not G24986;
	I33145<= not G24997;
	I33154<= not G25005;
	I33157<= not G25027;
	I33168<= not G25042;
	I33182<= not G25056;
	I33188<= not G24814;
	I33198<= not G25067;
	I33205<= not G24833;
	I33219<= not G24849;
	I33232<= not G24863;
	I33246<= not G24890;
	I33249<= not G24890;
	I33257<= not G24909;
	I33260<= not G24909;
	I33265<= not G24925;
	I33268<= not G24925;
	I33278<= not G25088;
	I33282<= not G25096;
	I33286<= not G24426;
	I33289<= not G25106;
	I33293<= not G25008;
	I33297<= not G24430;
	I33300<= not G25112;
	I33304<= not G25004;
	I33307<= not G25011;
	I33312<= not G25014;
	I33316<= not G24434;
	I33321<= not G24442;
	I33324<= not G25009;
	I33327<= not G25017;
	I33330<= not G25019;
	I33335<= not G25010;
	I33338<= not G25021;
	I33343<= not G25024;
	I33347<= not G24438;
	I33352<= not G24443;
	I33355<= not G25012;
	I33358<= not G25028;
	I33361<= not G25013;
	I33364<= not G25029;
	I33368<= not G24444;
	I33371<= not G25015;
	I33374<= not G25031;
	I33377<= not G25033;
	I33382<= not G25016;
	I33385<= not G25035;
	I33390<= not G25038;
	I33396<= not G24447;
	I33399<= not G25018;
	I33402<= not G24448;
	I33405<= not G25020;
	I33408<= not G25040;
	I33411<= not G24491;
	I33415<= not G24449;
	I33418<= not G25022;
	I33421<= not G25043;
	I33424<= not G25023;
	I33427<= not G25044;
	I33431<= not G24450;
	I33434<= not G25025;
	I33437<= not G25046;
	I33440<= not G25048;
	I33445<= not G25026;
	I33448<= not G25050;
	I33457<= not G24451;
	I33460<= not G24452;
	I33463<= not G25030;
	I33466<= not G25053;
	I33469<= not G24498;
	I33472<= not G24499;
	I33476<= not G24453;
	I33479<= not G25032;
	I33482<= not G24454;
	I33485<= not G25034;
	I33488<= not G25054;
	I33491<= not G24501;
	I33495<= not G24455;
	I33498<= not G25036;
	I33501<= not G25057;
	I33504<= not G25037;
	I33507<= not G25058;
	I33511<= not G24456;
	I33514<= not G25039;
	I33517<= not G25060;
	I33520<= not G25062;
	I33526<= not G24457;
	I33529<= not G25041;
	I33532<= not G24507;
	I33535<= not G24508;
	I33539<= not G24458;
	I33542<= not G24459;
	I33545<= not G25045;
	I33548<= not G25064;
	I33551<= not G24510;
	I33554<= not G24511;
	I33558<= not G24460;
	I33561<= not G25047;
	I33564<= not G24461;
	I33567<= not G25049;
	I33570<= not G25065;
	I33573<= not G24513;
	I33577<= not G24462;
	I33580<= not G25051;
	I33583<= not G25068;
	I33586<= not G25052;
	I33589<= not G25069;
	I33593<= not G24445;
	I33596<= not G24446;
	I33600<= not G24463;
	I33603<= not G24519;
	I33608<= not G24464;
	I33611<= not G25055;
	I33614<= not G24521;
	I33617<= not G24522;
	I33621<= not G24465;
	I33624<= not G24466;
	I33627<= not G25059;
	I33630<= not G25071;
	I33633<= not G24524;
	I33636<= not G24525;
	I33640<= not G24467;
	I33643<= not G25061;
	I33646<= not G24468;
	I33649<= not G25063;
	I33652<= not G25072;
	I33655<= not G24527;
	I33659<= not G24469;
	I33662<= not G24532;
	I33667<= not G24470;
	I33670<= not G25066;
	I33673<= not G24534;
	I33676<= not G24535;
	I33680<= not G24471;
	I33683<= not G24472;
	I33686<= not G25070;
	I33689<= not G25074;
	I33692<= not G24537;
	I33695<= not G24538;
	I33700<= not G24474;
	I33703<= not G24545;
	I33708<= not G24475;
	I33711<= not G25073;
	I33714<= not G24547;
	I33717<= not G24548;
	I33723<= not G24477;
	I33726<= not G24557;
	I33732<= not G24473;
	I33737<= not G24476;
	I33790<= not G25103;
	I33798<= not G25109;
	I33801<= not G25327;
	I33804<= not G25976;
	I33807<= not G25588;
	I33810<= not G25646;
	I33813<= not G25706;
	I33816<= not G25647;
	I33819<= not G25707;
	I33822<= not G25770;
	I33825<= not G25462;
	I33828<= not G25336;
	I33831<= not G25982;
	I33834<= not G25667;
	I33837<= not G25723;
	I33840<= not G25779;
	I33843<= not G25724;
	I33846<= not G25780;
	I33849<= not G25824;
	I33852<= not G25471;
	I33855<= not G25350;
	I33858<= not G25179;
	I33861<= not G25744;
	I33864<= not G25796;
	I33867<= not G25833;
	I33870<= not G25797;
	I33873<= not G25834;
	I33876<= not G25859;
	I33879<= not G25488;
	I33882<= not G25364;
	I33885<= not G25180;
	I33888<= not G25817;
	I33891<= not G25850;
	I33894<= not G25868;
	I33897<= not G25851;
	I33900<= not G25869;
	I33903<= not G25880;
	I33906<= not G25519;
	I33909<= not G25886;
	I33912<= not G25891;
	I33915<= not G25762;
	I33918<= not G25763;
	I33954<= not G25343;
	I33961<= not G25357;
	I33968<= not G25372;
	I33974<= not G25389;
	I33984<= not G25932;
	I33990<= not G25870;
	I33995<= not G25935;
	I33999<= not G25490;
	I34002<= not G25490;
	I34009<= not G25882;
	I34012<= not G25938;
	I34017<= not G25887;
	I34020<= not G25940;
	I34026<= not G25892;
	I34029<= not G25520;
	I34032<= not G25520;
	I34041<= not G25566;
	I34044<= not G25566;
	I34051<= not G25204;
	I34056<= not G25206;
	I34059<= not G25207;
	I34063<= not G25209;
	I34068<= not G25211;
	I34071<= not G25212;
	I34074<= not G25213;
	I34077<= not G25954;
	I34080<= not G25539;
	I34083<= not G25214;
	I34086<= not G25215;
	I34091<= not G25217;
	I34096<= not G25218;
	I34099<= not G25219;
	I34102<= not G25220;
	I34105<= not G25221;
	I34108<= not G25222;
	I34111<= not G25223;
	I34114<= not G25958;
	I34118<= not G25605;
	I34121<= not G25224;
	I34124<= not G25225;
	I34128<= not G25227;
	I34132<= not G25228;
	I34135<= not G25229;
	I34140<= not G25230;
	I34143<= not G25231;
	I34146<= not G25232;
	I34150<= not G25233;
	I34153<= not G25234;
	I34156<= not G25235;
	I34159<= not G25964;
	I34162<= not G25684;
	I34165<= not G25236;
	I34168<= not G25237;
	I34172<= not G25239;
	I34180<= not G25240;
	I34183<= not G25241;
	I34189<= not G25242;
	I34192<= not G25243;
	I34195<= not G25244;
	I34198<= not G25245;
	I34201<= not G25246;
	I34204<= not G25247;
	I34207<= not G25969;
	I34210<= not G25761;
	I34220<= not G25248;
	I34230<= not G25249;
	I34233<= not G25250;
	I34238<= not G25251;
	I34241<= not G25252;
	I34244<= not G25253;
	I34254<= not G25185;
	I34266<= not G25255;
	I34274<= not G25256;
	I34277<= not G25257;
	I34296<= not G25189;
	I34306<= not G25259;
	I34313<= not G25265;
	I34316<= not G25191;
	I34321<= not G25928;
	I34327<= not G25260;
	I34343<= not G25194;
	I34353<= not G25927;
	I34358<= not G25262;
	I34363<= not G25930;
	I34369<= not G25263;
	I34385<= not G25197;
	I34388<= not G25200;
	I34392<= not G25266;
	I34395<= not G25929;
	I34400<= not G25267;
	I34405<= not G25933;
	I34411<= not G25268;
	I34421<= not G25203;
	I34425<= not G25270;
	I34428<= not G25931;
	I34433<= not G25271;
	I34438<= not G25936;
	I34444<= not G25272;
	I34449<= not G25205;
	I34453<= not G25279;
	I34456<= not G25934;
	I34461<= not G25280;
	I34464<= not G25199;
	I34469<= not G25210;
	I34473<= not G25288;
	I34476<= not G25201;
	I34479<= not G25202;
	I34505<= not G25450;
	I34535<= not G25451;
	I34579<= not G25452;
	I34641<= not G26086;
	I34644<= not G26159;
	I34647<= not G26164;
	I34650<= not G26172;
	I34653<= not G26165;
	I34656<= not G26173;
	I34659<= not G26190;
	I34662<= not G26174;
	I34665<= not G26191;
	I34668<= not G26210;
	I34671<= not G26192;
	I34674<= not G26211;
	I34677<= not G26232;
	I34680<= not G26294;
	I34683<= not G26364;
	I34686<= not G26398;
	I34689<= not G26433;
	I34692<= not G26102;
	I34695<= not G26167;
	I34698<= not G26181;
	I34701<= not G26193;
	I34704<= not G26182;
	I34707<= not G26194;
	I34710<= not G26214;
	I34713<= not G26195;
	I34716<= not G26215;
	I34719<= not G26238;
	I34722<= not G26216;
	I34725<= not G26239;
	I34728<= not G26264;
	I34731<= not G26341;
	I34734<= not G26407;
	I34737<= not G26439;
	I34740<= not G26465;
	I34743<= not G26118;
	I34746<= not G26187;
	I34749<= not G26205;
	I34752<= not G26220;
	I34755<= not G26206;
	I34758<= not G26221;
	I34761<= not G26245;
	I34764<= not G26222;
	I34767<= not G26246;
	I34770<= not G26276;
	I34773<= not G26247;
	I34776<= not G26277;
	I34779<= not G26308;
	I34782<= not G26385;
	I34785<= not G26448;
	I34788<= not G26471;
	I34791<= not G26489;
	I34794<= not G26125;
	I34797<= not G26208;
	I34800<= not G26229;
	I34803<= not G26248;
	I34806<= not G26230;
	I34809<= not G26249;
	I34812<= not G26280;
	I34815<= not G26250;
	I34818<= not G26281;
	I34821<= not G26314;
	I34824<= not G26282;
	I34827<= not G26315;
	I34830<= not G26349;
	I34833<= not G26428;
	I34836<= not G26480;
	I34839<= not G26495;
	I34842<= not G26505;
	I34845<= not G26496;
	I34848<= not G26506;
	I34851<= not G26354;
	I34854<= not G26507;
	I34857<= not G26355;
	I34860<= not G26548;
	I34863<= not G26576;
	I34866<= not G26618;
	I34872<= not G26217;
	I34879<= not G26240;
	I34901<= not G26295;
	I34909<= not G26265;
	I34916<= not G26240;
	I34921<= not G26217;
	I34946<= not G26534;
	I34957<= not G26541;
	I34961<= not G26545;
	I34964<= not G26547;
	I34967<= not G26553;
	I34971<= not G26557;
	I34974<= not G26168;
	I34977<= not G26559;
	I34980<= not G26458;
	I34983<= not G26569;
	I34986<= not G26160;
	I34990<= not G26573;
	I34993<= not G26575;
	I34997<= not G26482;
	I35000<= not G26336;
	I35003<= not G26592;
	I35007<= not G26596;
	I35011<= not G26304;
	I35014<= not G26498;
	I35017<= not G26616;
	I35028<= not G26513;
	I35031<= not G26529;
	I35049<= not G26530;
	I35053<= not G26655;
	I35064<= not G26531;
	I35067<= not G26659;
	I35072<= not G26661;
	I35076<= not G26532;
	I35079<= not G26664;
	I35083<= not G26665;
	I35087<= not G26667;
	I35092<= not G26669;
	I35095<= not G26670;
	I35099<= not G26672;
	I35106<= not G26675;
	I35109<= not G26676;
	I35116<= not G26025;
	I35136<= not G26660;
	I35141<= not G26666;
	I35146<= not G26671;
	I35153<= not G26677;
	I35172<= not G26272;
	I35254<= not G26048;
	I35283<= not G26031;
	I35297<= not G26199;
	I35301<= not G26037;
	I35313<= not G26534;
	I35319<= not G26183;
	I35334<= not G26106;
	I35341<= not G26120;
	I35347<= not G26265;
	I35351<= not G26272;
	I35355<= not G26130;
	I35360<= not G26295;
	I35364<= not G26304;
	I35369<= not G26144;
	I35373<= not G26189;
	I35376<= not G26336;
	I35383<= not G26160;
	I35389<= not G26168;
	I35394<= not G26183;
	I35399<= not G26199;
	I35404<= not G26864;
	I35407<= not G27145;
	I35410<= not G26872;
	I35413<= not G26876;
	I35416<= not G26884;
	I35419<= not G26828;
	I35422<= not G26830;
	I35425<= not G26832;
	I35428<= not G26953;
	I35431<= not G26868;
	I35434<= not G27150;
	I35437<= not G27183;
	I35440<= not G27186;
	I35443<= not G26757;
	I35446<= not G26762;
	I35449<= not G27154;
	I35452<= not G27161;
	I35455<= not G26881;
	I35458<= not G26886;
	I35461<= not G26895;
	I35464<= not G26831;
	I35467<= not G26834;
	I35470<= not G26840;
	I35473<= not G27156;
	I35476<= not G27163;
	I35479<= not G27171;
	I35482<= not G27176;
	I35485<= not G27180;
	I35488<= not G26819;
	I35491<= not G26956;
	I35494<= not G26875;
	I35497<= not G27158;
	I35500<= not G26890;
	I35503<= not G26896;
	I35506<= not G26909;
	I35509<= not G26836;
	I35512<= not G26843;
	I35515<= not G26850;
	I35518<= not G26959;
	I35521<= not G26883;
	I35524<= not G27166;
	I35527<= not G26900;
	I35530<= not G26910;
	I35533<= not G26921;
	I35536<= not G26844;
	I35539<= not G26852;
	I35542<= not G26858;
	I35545<= not G26964;
	I35548<= not G27116;
	I35551<= not G27075;
	I35554<= not G27102;
	I35667<= not G27120;
	I35673<= not G27123;
	I35678<= not G27129;
	I35681<= not G26869;
	I35686<= not G27131;
	I35689<= not G26878;
	I35695<= not G26887;
	I35698<= not G26897;
	I35708<= not G26974;
	I35711<= not G26974;
	I35723<= not G27168;
	I35727<= not G26902;
	I35731<= not G26892;
	I35737<= not G26915;
	I35741<= not G27118;
	I35744<= not G26906;
	I35750<= not G26928;
	I35756<= not G27117;
	I35759<= not G27121;
	I35762<= not G26918;
	I35768<= not G26941;
	I35772<= not G26772;
	I35777<= not G27119;
	I35780<= not G27124;
	I35783<= not G26931;
	I35791<= not G26779;
	I35796<= not G27122;
	I35799<= not G27130;
	I35803<= not G26803;
	I35809<= not G26785;
	I35814<= not G27125;
	I35817<= not G26922;
	I35821<= not G26804;
	I35824<= not G26805;
	I35829<= not G26806;
	I35834<= not G26792;
	I35837<= not G26911;
	I35841<= not G26807;
	I35844<= not G26808;
	I35849<= not G26776;
	I35852<= not G26935;
	I35856<= not G26809;
	I35859<= not G26810;
	I35863<= not G26811;
	I35868<= not G26812;
	I35872<= not G26925;
	I35876<= not G26813;
	I35879<= not G26814;
	I35883<= not G26781;
	I35886<= not G26944;
	I35890<= not G26815;
	I35893<= not G26816;
	I35897<= not G26817;
	I35900<= not G26786;
	I35915<= not G26818;
	I35919<= not G26938;
	I35923<= not G26820;
	I35926<= not G26821;
	I35930<= not G26789;
	I35933<= not G26950;
	I35937<= not G26822;
	I35940<= not G26823;
	I35953<= not G26824;
	I35957<= not G26947;
	I35961<= not G26825;
	I35964<= not G26826;
	I35968<= not G26795;
	I35983<= not G26827;
	I36008<= not G26798;
	I36032<= not G27113;
	I36042<= not G26960;
	I36046<= not G26957;
	I36052<= not G26954;
	I36060<= not G27353;
	I36063<= not G27463;
	I36066<= not G27479;
	I36069<= not G27493;
	I36072<= not G27480;
	I36075<= not G27494;
	I36078<= not G27508;
	I36081<= not G27497;
	I36084<= not G27357;
	I36087<= not G27483;
	I36090<= not G27502;
	I36093<= not G27514;
	I36096<= not G27503;
	I36099<= not G27515;
	I36102<= not G27533;
	I36105<= not G27517;
	I36108<= not G27360;
	I36111<= not G27505;
	I36114<= not G27522;
	I36117<= not G27539;
	I36120<= not G27523;
	I36123<= not G27540;
	I36126<= not G27553;
	I36129<= not G27542;
	I36132<= not G27366;
	I36135<= not G27525;
	I36138<= not G27547;
	I36141<= not G27559;
	I36144<= not G27548;
	I36147<= not G27560;
	I36150<= not G27569;
	I36153<= not G27562;
	I36156<= not G27586;
	I36159<= not G27526;
	I36162<= not G27385;
	I36213<= not G27571;
	I36217<= not G27580;
	I36221<= not G27662;
	I36224<= not G27589;
	I36227<= not G27594;
	I36230<= not G27583;
	I36234<= not G27667;
	I36237<= not G27662;
	I36240<= not G27603;
	I36243<= not G27587;
	I36246<= not G27674;
	I36250<= not G27612;
	I36253<= not G27674;
	I36264<= not G27621;
	I36267<= not G27395;
	I36280<= not G27390;
	I36283<= not G27408;
	I36296<= not G27626;
	I36307<= not G27400;
	I36311<= not G27426;
	I36321<= not G27627;
	I36327<= not G27413;
	I36330<= not G27447;
	I36337<= not G27628;
	I36341<= not G27431;
	I36347<= not G27630;
	I36354<= not G27662;
	I36358<= not G27672;
	I36362<= not G27667;
	I36367<= not G27678;
	I36371<= not G27674;
	I36379<= not G27682;
	I36382<= not G27563;
	I36390<= not G27243;
	I36393<= not G27572;
	I36397<= not G27574;
	I36404<= not G27450;
	I36407<= not G27581;
	I36411<= not G27582;
	I36417<= not G27462;
	I36420<= not G27253;
	I36423<= not G27466;
	I36426<= not G27584;
	I36432<= not G27585;
	I36438<= not G27255;
	I36441<= not G27256;
	I36444<= not G27482;
	I36447<= not G27257;
	I36450<= not G27485;
	I36454<= not G27588;
	I36459<= not G27258;
	I36462<= not G27259;
	I36465<= not G27260;
	I36468<= not G27261;
	I36473<= not G27262;
	I36476<= not G27263;
	I36479<= not G27504;
	I36483<= not G27264;
	I36486<= not G27507;
	I36490<= not G27265;
	I36493<= not G27266;
	I36496<= not G27267;
	I36499<= not G27268;
	I36502<= not G27269;
	I36507<= not G27270;
	I36510<= not G27271;
	I36513<= not G27272;
	I36516<= not G27273;
	I36521<= not G27274;
	I36524<= not G27275;
	I36527<= not G27524;
	I36530<= not G27276;
	I36533<= not G27277;
	I36536<= not G27278;
	I36539<= not G27279;
	I36542<= not G27280;
	I36545<= not G27281;
	I36551<= not G27282;
	I36554<= not G27283;
	I36557<= not G27284;
	I36560<= not G27285;
	I36563<= not G27286;
	I36568<= not G27287;
	I36571<= not G27288;
	I36574<= not G27289;
	I36577<= not G27290;
	I36582<= not G27291;
	I36585<= not G27292;
	I36588<= not G27293;
	I36598<= not G27294;
	I36601<= not G27295;
	I36604<= not G27296;
	I36609<= not G27297;
	I36612<= not G27298;
	I36615<= not G27299;
	I36618<= not G27300;
	I36621<= not G27301;
	I36627<= not G27302;
	I36630<= not G27303;
	I36633<= not G27304;
	I36636<= not G27305;
	I36639<= not G27306;
	I36644<= not G27307;
	I36647<= not G27308;
	I36650<= not G27309;
	I36653<= not G27310;
	I36656<= not G27311;
	I36659<= not G27312;
	I36663<= not G27313;
	I36673<= not G27314;
	I36676<= not G27315;
	I36679<= not G27316;
	I36684<= not G27317;
	I36687<= not G27318;
	I36690<= not G27319;
	I36693<= not G27320;
	I36696<= not G27321;
	I36702<= not G27322;
	I36705<= not G27323;
	I36708<= not G27324;
	I36711<= not G27325;
	I36714<= not G27326;
	I36718<= not G27327;
	I36721<= not G27328;
	I36724<= not G27329;
	I36728<= not G27330;
	I36738<= not G27331;
	I36741<= not G27332;
	I36744<= not G27333;
	I36749<= not G27334;
	I36752<= not G27335;
	I36755<= not G27336;
	I36758<= not G27337;
	I36761<= not G27338;
	I36766<= not G27339;
	I36769<= not G27340;
	I36772<= not G27341;
	I36776<= not G27342;
	I36786<= not G27343;
	I36789<= not G27344;
	I36792<= not G27345;
	I36797<= not G27346;
	I36800<= not G27347;
	I36803<= not G27348;
	I36808<= not G27354;
	I36848<= not G27383;
	I36860<= not G27386;
	I36864<= not G27384;
	I36867<= not G27786;
	I36870<= not G27955;
	I36873<= not G27971;
	I36876<= not G27986;
	I36879<= not G27972;
	I36882<= not G27987;
	I36885<= not G28003;
	I36888<= not G27988;
	I36891<= not G28004;
	I36894<= not G28022;
	I36897<= not G28005;
	I36900<= not G28023;
	I36903<= not G28045;
	I36906<= not G27989;
	I36909<= not G28006;
	I36912<= not G28024;
	I36915<= not G28007;
	I36918<= not G28025;
	I36921<= not G28047;
	I36924<= not G28026;
	I36927<= not G28048;
	I36930<= not G28071;
	I36933<= not G28049;
	I36936<= not G28072;
	I36939<= not G28095;
	I36942<= not G27905;
	I36945<= not G27793;
	I36948<= not G27976;
	I36951<= not G27992;
	I36954<= not G28010;
	I36957<= not G27993;
	I36960<= not G28011;
	I36963<= not G28030;
	I36966<= not G28012;
	I36969<= not G28031;
	I36972<= not G28052;
	I36975<= not G28032;
	I36978<= not G28053;
	I36981<= not G28074;
	I36984<= not G28013;
	I36987<= not G28033;
	I36990<= not G28054;
	I36993<= not G28034;
	I36996<= not G28055;
	I36999<= not G28076;
	I37002<= not G28056;
	I37005<= not G28077;
	I37008<= not G28096;
	I37011<= not G28078;
	I37014<= not G28097;
	I37017<= not G28113;
	I37020<= not G27910;
	I37023<= not G27799;
	I37026<= not G27998;
	I37029<= not G28016;
	I37032<= not G28037;
	I37035<= not G28017;
	I37038<= not G28038;
	I37041<= not G28060;
	I37044<= not G28039;
	I37047<= not G28061;
	I37050<= not G28081;
	I37053<= not G28062;
	I37056<= not G28082;
	I37059<= not G28099;
	I37062<= not G28040;
	I37065<= not G28063;
	I37068<= not G28083;
	I37071<= not G28064;
	I37074<= not G28084;
	I37077<= not G28101;
	I37080<= not G28085;
	I37083<= not G28102;
	I37086<= not G28114;
	I37089<= not G28103;
	I37092<= not G28115;
	I37095<= not G28124;
	I37098<= not G27918;
	I37101<= not G27805;
	I37104<= not G28021;
	I37107<= not G28043;
	I37110<= not G28067;
	I37113<= not G28044;
	I37116<= not G28068;
	I37119<= not G28089;
	I37122<= not G28069;
	I37125<= not G28090;
	I37128<= not G28106;
	I37131<= not G28091;
	I37134<= not G28107;
	I37137<= not G28117;
	I37140<= not G28070;
	I37143<= not G28092;
	I37146<= not G28108;
	I37149<= not G28093;
	I37152<= not G28109;
	I37155<= not G28119;
	I37158<= not G28110;
	I37161<= not G28120;
	I37164<= not G28125;
	I37167<= not G28121;
	I37170<= not G28126;
	I37173<= not G28132;
	I37176<= not G27927;
	I37179<= not G27784;
	I37182<= not G27791;
	I37185<= not G27797;
	I37188<= not G27785;
	I37191<= not G27792;
	I37194<= not G27800;
	I37197<= not G27903;
	I37200<= not G27907;
	I37203<= not G27912;
	I37228<= not G28194;
	I37232<= not G28200;
	I37238<= not G28179;
	I37252<= not G28200;
	I37260<= not G28179;
	I37266<= not G28200;
	I37269<= not G28145;
	I37273<= not G28179;
	I37277<= not G28146;
	I37280<= not G28179;
	I37284<= not G28147;
	I37291<= not G28148;
	I37319<= not G28149;
	I37330<= not G28194;
	I37334<= not G28194;
	I37379<= not G28199;
	I37386<= not G28194;
	I37394<= not G27718;
	I37400<= not G28200;
	I37410<= not G27722;
	I37415<= not G28179;
	I37426<= not G27724;
	I37459<= not G27759;
	I37467<= not G27760;
	I37471<= not G27761;
	I37474<= not G27762;
	I37481<= not G27763;
	I37484<= not G27764;
	I37488<= not G27765;
	I37494<= not G27766;
	I37497<= not G27767;
	I37502<= not G27768;
	I37508<= not G27769;
	I37514<= not G27771;
	I37566<= not G28370;
	I37569<= not G28498;
	I37572<= not G28524;
	I37575<= not G28527;
	I37578<= not G28432;
	I37581<= not G28374;
	I37584<= not G28526;
	I37587<= not G28552;
	I37590<= not G28555;
	I37593<= not G28443;
	I37596<= not G28377;
	I37599<= not G28553;
	I37602<= not G28579;
	I37605<= not G28583;
	I37608<= not G28455;
	I37611<= not G28382;
	I37614<= not G28580;
	I37617<= not G28607;
	I37620<= not G28611;
	I37623<= not G28467;
	I37626<= not G28393;
	I37629<= not G28369;
	I37632<= not G28372;
	I37635<= not G28390;
	I37638<= not G28395;
	I37641<= not G28375;
	I37644<= not G28341;
	I37647<= not G28343;
	I37650<= not G28347;
	I37653<= not G28359;
	I37656<= not G28365;
	I37659<= not G28437;
	I37662<= not G28447;
	I37665<= not G28458;
	I37702<= not G28512;
	I37712<= not G28512;
	I37716<= not G28540;
	I37725<= not G28540;
	I37729<= not G28567;
	I37736<= not G28567;
	I37740<= not G28595;
	I37746<= not G28595;
	I37752<= not G28512;
	I37757<= not G28512;
	I37760<= not G28540;
	I37765<= not G28512;
	I37768<= not G28540;
	I37771<= not G28567;
	I37775<= not G28540;
	I37778<= not G28567;
	I37781<= not G28595;
	I37784<= not G28567;
	I37787<= not G28595;
	I37790<= not G28595;
	I37793<= not G28638;
	I37796<= not G28634;
	I37800<= not G28635;
	I37804<= not G28636;
	I37808<= not G28637;
	I37842<= not G28501;
	I37846<= not G28501;
	I37851<= not G28668;
	I37854<= not G28529;
	I37858<= not G28501;
	I37863<= not G28529;
	I37868<= not G28321;
	I37871<= not G28556;
	I37875<= not G28501;
	I37880<= not G28529;
	I37885<= not G28556;
	I37891<= not G28325;
	I37894<= not G28584;
	I37897<= not G28501;
	I37901<= not G28529;
	I37906<= not G28556;
	I37912<= not G28584;
	I37917<= not G28328;
	I37920<= not G28501;
	I37924<= not G28529;
	I37928<= not G28556;
	I37934<= not G28584;
	I37939<= not G28501;
	I37942<= not G28501;
	I37946<= not G28529;
	I37950<= not G28556;
	I37956<= not G28584;
	I37961<= not G28501;
	I37965<= not G28529;
	I37968<= not G28529;
	I37973<= not G28556;
	I37978<= not G28584;
	I37982<= not G28501;
	I37986<= not G28529;
	I37991<= not G28556;
	I37994<= not G28556;
	I37999<= not G28584;
	I38003<= not G28529;
	I38007<= not G28556;
	I38011<= not G28584;
	I38014<= not G28584;
	I38018<= not G28342;
	I38024<= not G28556;
	I38028<= not G28584;
	I38032<= not G28344;
	I38035<= not G28345;
	I38038<= not G28346;
	I38042<= not G28584;
	I38046<= not G28348;
	I38049<= not G28349;
	I38053<= not G28350;
	I38056<= not G28351;
	I38059<= not G28352;
	I38064<= not G28353;
	I38068<= not G28354;
	I38071<= not G28355;
	I38074<= not G28356;
	I38077<= not G28357;
	I38080<= not G28358;
	I38085<= not G28360;
	I38088<= not G28361;
	I38091<= not G28362;
	I38094<= not G28363;
	I38097<= not G28364;
	I38101<= not G28366;
	I38104<= not G28367;
	I38107<= not G28368;
	I38111<= not G28371;
	I38119<= not G28420;
	I38122<= not G28421;
	I38125<= not G28425;
	I38128<= not G28419;
	I38136<= not G28833;
	I38139<= not G29061;
	I38142<= not G29073;
	I38145<= not G29081;
	I38148<= not G29074;
	I38151<= not G29082;
	I38154<= not G29089;
	I38157<= not G28882;
	I38160<= not G28835;
	I38163<= not G29075;
	I38166<= not G29084;
	I38169<= not G29091;
	I38172<= not G29085;
	I38175<= not G29092;
	I38178<= not G29098;
	I38181<= not G28899;
	I38184<= not G28837;
	I38187<= not G29086;
	I38190<= not G29093;
	I38193<= not G29099;
	I38196<= not G29094;
	I38199<= not G29100;
	I38202<= not G29104;
	I38205<= not G28924;
	I38208<= not G28839;
	I38211<= not G29095;
	I38214<= not G29101;
	I38217<= not G29105;
	I38220<= not G29102;
	I38223<= not G29106;
	I38226<= not G29108;
	I38229<= not G28950;
	I38232<= not G29117;
	I38235<= not G29118;
	I38238<= not G29119;
	I38241<= not G28832;
	I38245<= not G28920;
	I38250<= not G28941;
	I38258<= not G28963;
	I38272<= not G29013;
	I38275<= not G28987;
	I38278<= not G28963;
	I38282<= not G28941;
	I38321<= not G29113;
	I38330<= not G29120;
	I38339<= not G29120;
	I38342<= not G28886;
	I38345<= not G29109;
	I38348<= not G28874;
	I38352<= not G29110;
	I38355<= not G29039;
	I38360<= not G29111;
	I38363<= not G29016;
	I38369<= not G29112;
	I38386<= not G28734;
	I38391<= not G28730;
	I38396<= not G28727;
	I38401<= not G28725;
	I38405<= not G28723;
	I38408<= not G28721;
	I38412<= not G28720;
	I38421<= not G28740;
	I38428<= not G28732;
	I38434<= not G28735;
	I38437<= not G28736;
	I38440<= not G28738;
	I38447<= not G28744;
	I38450<= not G28745;
	I38453<= not G28746;
	I38456<= not G28747;
	I38459<= not G28749;
	I38462<= not G29120;
	I38466<= not G28754;
	I38471<= not G28758;
	I38474<= not G28759;
	I38477<= not G28760;
	I38480<= not G28761;
	I38483<= not G28990;
	I38486<= not G28763;
	I38491<= not G28767;
	I38496<= not G28771;
	I38499<= not G28772;
	I38502<= not G28773;
	I38505<= not G28774;
	I38510<= not G28778;
	I38515<= not G28782;
	I38518<= not G28783;
	I38524<= not G28788;
	I38536<= not G28920;
	I38539<= not G29113;
	I38548<= not G28903;
	I38591<= not G28987;
	I38594<= not G28990;
	I38599<= not G29013;
	I38602<= not G29016;
	I38606<= not G29039;
	I38609<= not G28874;
	I38613<= not G28886;
	I38617<= not G28903;
	I38620<= not G29246;
	I38623<= not G29293;
	I38626<= not G29297;
	I38629<= not G29304;
	I38632<= not G29298;
	I38635<= not G29305;
	I38638<= not G29311;
	I38641<= not G29249;
	I38644<= not G29299;
	I38647<= not G29306;
	I38650<= not G29314;
	I38653<= not G29307;
	I38656<= not G29315;
	I38659<= not G29322;
	I38662<= not G29253;
	I38665<= not G29412;
	I38668<= not G29168;
	I38671<= not G29171;
	I38674<= not G29177;
	I38677<= not G29400;
	I38680<= not G29404;
	I38683<= not G29308;
	I38686<= not G29316;
	I38689<= not G29325;
	I38692<= not G29317;
	I38695<= not G29326;
	I38698<= not G29331;
	I38701<= not G29401;
	I38704<= not G29405;
	I38707<= not G29407;
	I38710<= not G29408;
	I38713<= not G29410;
	I38716<= not G29230;
	I38719<= not G29258;
	I38722<= not G29319;
	I38725<= not G29327;
	I38728<= not G29334;
	I38731<= not G29328;
	I38734<= not G29335;
	I38737<= not G29339;
	I38740<= not G29288;
	I38743<= not G29267;
	I38746<= not G29270;
	I38749<= not G29273;
	I38752<= not G29276;
	I38755<= not G29278;
	I38758<= not G29279;
	I38761<= not G29281;
	I38764<= not G29237;
	I38767<= not G29244;
	I38770<= not G29309;
	I38801<= not G29358;
	I38804<= not G29353;
	I38807<= not G29356;
	I38817<= not G29354;
	I38827<= not G29355;
	I38838<= not G29357;
	I38848<= not G29167;
	I38851<= not G29169;
	I38854<= not G29170;
	I38857<= not G29172;
	I38860<= not G29173;
	I38863<= not G29178;
	I38866<= not G29179;
	I38869<= not G29181;
	I38872<= not G29182;
	I38875<= not G29184;
	I38878<= not G29185;
	I38881<= not G29187;
	I38885<= not G29192;
	I38898<= not G29194;
	I38905<= not G29197;
	I38909<= not G29198;
	I38916<= not G29201;
	I38920<= not G29204;
	I38924<= not G29205;
	I38931<= not G29209;
	I38936<= not G29212;
	I38940<= not G29213;
	I38947<= not G29218;
	I38951<= not G29221;
	I38958<= not G29226;
	I38975<= not G29348;
	I38999<= not G29496;
	I39002<= not G29506;
	I39005<= not G29507;
	I39008<= not G29509;
	I39011<= not G29530;
	I39014<= not G29535;
	I39017<= not G29542;
	I39020<= not G29499;
	I39023<= not G29508;
	I39026<= not G29510;
	I39029<= not G29512;
	I39032<= not G29537;
	I39035<= not G29544;
	I39038<= not G29551;
	I39041<= not G29501;
	I39044<= not G29511;
	I39047<= not G29513;
	I39050<= not G29515;
	I39053<= not G29546;
	I39056<= not G29554;
	I39059<= not G29561;
	I39062<= not G29504;
	I39065<= not G29514;
	I39068<= not G29516;
	I39071<= not G29517;
	I39074<= not G29556;
	I39077<= not G29563;
	I39080<= not G29568;
	I39083<= not G29519;
	I39086<= not G29497;
	I39089<= not G29495;
	I39121<= not G29579;
	I39124<= not G29606;
	I39127<= not G29608;
	I39130<= not G29580;
	I39133<= not G29609;
	I39136<= not G29611;
	I39139<= not G29612;
	I39142<= not G29581;
	I39145<= not G29613;
	I39148<= not G29616;
	I39151<= not G29617;
	I39154<= not G29582;
	I39157<= not G29618;
	I39160<= not G29620;
	I39164<= not G29621;
	I39168<= not G29623;
	I39234<= not G29689;
	I39237<= not G29690;
	I39240<= not G29691;
	I39243<= not G29694;
	I39246<= not G29692;
	I39249<= not G29693;
	I39252<= not G29695;
	I39255<= not G29698;
	I39258<= not G29696;
	I39261<= not G29697;
	I39264<= not G29699;
	I39267<= not G29702;
	I39270<= not G29700;
	I39273<= not G29701;
	I39276<= not G29704;
	I39279<= not G29708;
	I39398<= not G29664;
	I39401<= not G29662;
	I39404<= not G29661;
	I39407<= not G29660;
	I39411<= not G29659;
	I39414<= not G29658;
	I39418<= not G29668;
	I39423<= not G29666;
	I39454<= not G29940;
	I39457<= not G29943;
	I39460<= not G29932;
	I39463<= not G29933;
	I39466<= not G29934;
	I39469<= not G29935;
	I39472<= not G29937;
	I39475<= not G29938;
	I39550<= not G29848;
	I39573<= not G29936;
	I39577<= not G29939;
	I39585<= not G29941;
	I39622<= not G30052;
	I39625<= not G30076;
	I39628<= not G30078;
	I39631<= not G30084;
	I39635<= not G30055;
	I39638<= not G30056;
	I39641<= not G30057;
	I39647<= not G30058;
	I39674<= not G30072;
	I39761<= not G30072;
	I39764<= not G30060;
	I39767<= not G30061;
	I39770<= not G30063;
	I39773<= not G30064;
	I39776<= not G30066;
	I39779<= not G30053;
	I39782<= not G30054;
	I39785<= not G30124;
	I39788<= not G30125;
	I39791<= not G30126;
	I39794<= not G30130;
	I39797<= not G30307;
	I39800<= not G30309;
	I39803<= not G30308;
	I39806<= not G30310;
	I39809<= not G30311;
	I39812<= not G30312;
	I39815<= not G30313;
	I39818<= not G30215;
	I39821<= not G30267;
	I39825<= not G30268;
	I39828<= not G30269;
	I39832<= not G30270;
	I39835<= not G30271;
	I39840<= not G30272;
	I39843<= not G30273;
	I39848<= not G30274;
	I39853<= not G30275;
	I39856<= not G30276;
	I39859<= not G30277;
	I39863<= not G30278;
	I39866<= not G30279;
	I39870<= not G30280;
	I39873<= not G30281;
	I39878<= not G30282;
	I39881<= not G30283;
	I39886<= not G30284;
	I39889<= not G30285;
	I39892<= not G30286;
	I39895<= not G30287;
	I39899<= not G30288;
	I39902<= not G30289;
	I39906<= not G30290;
	I39909<= not G30291;
	I39913<= not G30292;
	I39916<= not G30293;
	I39919<= not G30294;
	I39922<= not G30295;
	I39926<= not G30296;
	I39930<= not G30297;
	I39933<= not G30298;
	I39936<= not G30299;
	I39939<= not G30300;
	I39942<= not G30301;
	I39945<= not G30302;
	I39948<= not G30303;
	I39951<= not G30304;
	I39976<= not G30245;
	I39982<= not G30305;
	I39985<= not G30246;
	I39991<= not G30247;
	I39997<= not G30248;
	I40002<= not G30249;
	I40008<= not G30250;
	I40016<= not G30251;
	I40021<= not G30252;
	I40027<= not G30253;
	I40032<= not G30254;
	I40039<= not G30255;
	I40044<= not G30256;
	I40051<= not G30257;
	I40054<= not G30258;
	I40059<= not G30259;
	I40066<= not G30260;
	I40071<= not G30261;
	I40075<= not G30262;
	I40078<= not G30263;
	I40083<= not G30264;
	I40086<= not G30265;
	I40091<= not G30266;
	I40098<= not G30491;
	I40101<= not G30326;
	I40104<= not G30342;
	I40107<= not G30343;
	I40110<= not G30357;
	I40113<= not G30368;
	I40116<= not G30408;
	I40119<= not G30435;
	I40122<= not G30443;
	I40125<= not G30466;
	I40128<= not G30479;
	I40131<= not G30493;
	I40134<= not G30480;
	I40137<= not G30494;
	I40140<= not G30328;
	I40143<= not G30329;
	I40146<= not G30344;
	I40149<= not G30358;
	I40152<= not G30359;
	I40155<= not G30369;
	I40158<= not G30376;
	I40161<= not G30439;
	I40164<= not G30446;
	I40167<= not G30456;
	I40170<= not G30483;
	I40173<= not G30497;
	I40176<= not G30331;
	I40179<= not G30498;
	I40182<= not G30332;
	I40185<= not G30346;
	I40188<= not G30347;
	I40191<= not G30360;
	I40194<= not G30370;
	I40197<= not G30371;
	I40200<= not G30377;
	I40203<= not G30380;
	I40206<= not G30450;
	I40209<= not G30459;
	I40212<= not G30471;
	I40215<= not G30501;
	I40218<= not G30335;
	I40221<= not G30349;
	I40224<= not G30336;
	I40227<= not G30350;
	I40230<= not G30362;
	I40233<= not G30363;
	I40236<= not G30373;
	I40239<= not G30378;
	I40242<= not G30379;
	I40245<= not G30381;
	I40248<= not G30382;
	I40251<= not G30463;
	I40254<= not G30474;
	I40257<= not G30488;
	I40260<= not G30339;
	I40263<= not G30353;
	I40266<= not G30365;
	I40269<= not G30354;
	I40272<= not G30366;
	I40275<= not G30375;
	I40288<= not G30455;
	I40291<= not G30468;
	I40294<= not G30470;
	I40297<= not G30482;
	I40300<= not G30485;
	I40303<= not G30487;
	I40307<= not G30500;
	I40310<= not G30503;
	I40313<= not G30505;
	I40317<= not G30338;
	I40320<= not G30341;
	I40326<= not G30356;
	I40420<= not G30578;
	I40423<= not G30579;
	I40426<= not G30581;
	I40429<= not G30580;
	I40432<= not G30582;
	I40435<= not G30585;
	I40438<= not G30583;
	I40441<= not G30586;
	I40444<= not G30591;
	I40447<= not G30587;
	I40450<= not G30592;
	I40453<= not G30600;
	I40456<= not G30668;
	I40459<= not G30669;
	I40462<= not G30670;
	I40465<= not G30671;
	I40468<= not G30672;
	I40471<= not G30673;
	I40475<= not G30674;
	I40478<= not G30675;
	I40481<= not G30676;
	I40484<= not G30677;
	I40487<= not G30678;
	I40490<= not G30679;
	I40495<= not G30680;
	I40498<= not G30681;
	I40501<= not G30682;
	I40504<= not G30683;
	I40507<= not G30684;
	I40510<= not G30686;
	I40515<= not G30687;
	I40518<= not G30688;
	I40521<= not G30689;
	I40524<= not G30690;
	I40527<= not G30691;
	I40531<= not G30692;
	I40534<= not G30693;
	I40537<= not G30694;
	I40542<= not G30695;
	I40555<= not G30699;
	I40565<= not G30700;
	I40568<= not G30701;
	I40578<= not G30702;
	I40581<= not G30703;
	I40584<= not G30704;
	I40594<= not G30705;
	I40597<= not G30706;
	I40600<= not G30707;
	I40611<= not G30708;
	I40614<= not G30709;
	I40618<= not G30566;
	I40634<= not G30571;
	I40637<= not G30570;
	I40640<= not G30569;
	I40643<= not G30568;
	I40647<= not G30567;
	I40651<= not G30574;
	I40654<= not G30573;
	I40658<= not G30572;
	I40661<= not G30635;
	I40664<= not G30636;
	I40667<= not G30637;
	I40670<= not G30638;
	I40673<= not G30639;
	I40676<= not G30640;
	I40679<= not G30641;
	I40682<= not G30642;
	I40685<= not G30643;
	I40688<= not G30644;
	I40691<= not G30645;
	I40694<= not G30646;
	I40697<= not G30647;
	I40700<= not G30648;
	I40703<= not G30649;
	I40706<= not G30650;
	I40709<= not G30651;
	I40712<= not G30652;
	I40715<= not G30653;
	I40718<= not G30654;
	I40721<= not G30655;
	I40724<= not G30656;
	I40727<= not G30657;
	I40730<= not G30658;
	I40733<= not G30659;
	I40736<= not G30660;
	I40739<= not G30661;
	I40742<= not G30662;
	I40745<= not G30663;
	I40748<= not G30664;
	I40751<= not G30665;
	I40754<= not G30666;
	I40757<= not G30667;
	I40760<= not G30722;
	I40763<= not G30729;
	I40766<= not G30737;
	I40769<= not G30803;
	I40772<= not G30804;
	I40775<= not G30807;
	I40778<= not G30805;
	I40781<= not G30808;
	I40784<= not G30813;
	I40787<= not G30809;
	I40790<= not G30814;
	I40793<= not G30821;
	I40796<= not G30829;
	I40799<= not G30723;
	I40802<= not G30730;
	I40805<= not G30767;
	I40808<= not G30769;
	I40811<= not G30772;
	I40814<= not G30731;
	I40817<= not G30738;
	I40820<= not G30745;
	I40823<= not G30806;
	I40826<= not G30810;
	I40829<= not G30815;
	I40832<= not G30811;
	I40835<= not G30816;
	I40838<= not G30822;
	I40841<= not G30817;
	I40844<= not G30823;
	I40847<= not G30830;
	I40850<= not G30724;
	I40853<= not G30732;
	I40856<= not G30739;
	I40859<= not G30770;
	I40862<= not G30773;
	I40865<= not G30776;
	I40868<= not G30740;
	I40871<= not G30746;
	I40874<= not G30751;
	I40877<= not G30812;
	I40880<= not G30818;
	I40883<= not G30824;
	I40886<= not G30819;
	I40889<= not G30825;
	I40892<= not G30831;
	I40895<= not G30826;
	I40898<= not G30832;
	I40901<= not G30725;
	I40904<= not G30733;
	I40907<= not G30741;
	I40910<= not G30747;
	I40913<= not G30774;
	I40916<= not G30777;
	I40919<= not G30781;
	I40922<= not G30748;
	I40925<= not G30752;
	I40928<= not G30756;
	I40931<= not G30820;
	I40934<= not G30827;
	I40937<= not G30833;
	I40940<= not G30828;
	I40943<= not G30834;
	I40946<= not G30726;
	I40949<= not G30835;
	I40952<= not G30727;
	I40955<= not G30734;
	I40958<= not G30742;
	I40961<= not G30749;
	I40964<= not G30753;
	I40967<= not G30778;
	I40970<= not G30782;
	I40973<= not G30784;
	I40976<= not G30799;
	I40979<= not G30800;
	I40982<= not G30802;
	I40985<= not G30792;
	I40988<= not G30793;
	I40991<= not G30794;
	I40994<= not G30795;
	I40997<= not G30797;
	I41024<= not G30765;
	I41035<= not G30796;
	I41038<= not G30798;
	I41041<= not G30801;
	I41044<= not G30928;
	I41047<= not G30937;
	I41050<= not G30938;
	I41053<= not G30939;
	I41090<= not G30965;
	I41093<= not G30964;
	I41096<= not G30963;
	I41099<= not G30962;
	I41102<= not G30969;
	I41105<= not G30968;
	I41108<= not G30967;
	I41111<= not G30966;
	I41114<= not G30976;
	I41117<= not G30977;
	I41120<= not G30978;
	I41123<= not G30979;
	I41126<= not G30972;
	I41129<= not G30973;
	I41132<= not G30974;
	I41135<= not G30975;
	I41138<= not G30971;
	I41141<= not G30988;
	G5630<=G325 and G349;
	G5649<=G331 and G351;
	G5650<=G325 and G364;
	G5658<=G1012 and G1036;
	G5676<=G337 and G353;
	G5677<=G331 and G366;
	G5678<=G325 and G379;
	G5687<=G1018 and G1038;
	G5688<=G1012 and G1051;
	G5696<=G1706 and G1730;
	G5709<=G337 and G368;
	G5710<=G331 and G381;
	G5711<=G325 and G394;
	G5728<=G1024 and G1040;
	G5729<=G1018 and G1053;
	G5730<=G1012 and G1066;
	G5739<=G1712 and G1732;
	G5740<=G1706 and G1745;
	G5748<=G2400 and G2424;
	G5757<=G337 and G383;
	G5758<=G331 and G396;
	G5767<=G1024 and G1055;
	G5768<=G1018 and G1068;
	G5769<=G1012 and G1081;
	G5786<=G1718 and G1734;
	G5787<=G1712 and G1747;
	G5788<=G1706 and G1760;
	G5797<=G2406 and G2426;
	G5798<=G2400 and G2439;
	G5807<=G337 and G324;
	G5816<=G1024 and G1070;
	G5817<=G1018 and G1083;
	G5826<=G1718 and G1749;
	G5827<=G1712 and G1762;
	G5828<=G1706 and G1775;
	G5845<=G2412 and G2428;
	G5846<=G2406 and G2441;
	G5847<=G2400 and G2454;
	G5863<=G1024 and G1011;
	G5872<=G1718 and G1764;
	G5873<=G1712 and G1777;
	G5882<=G2412 and G2443;
	G5883<=G2406 and G2456;
	G5884<=G2400 and G2469;
	G5910<=G1718 and G1705;
	G5919<=G2412 and G2458;
	G5920<=G2406 and G2471;
	G5949<=G2412 and G2399;
	G8327<=G3254 and G219;
	G8328<=G6314 and G225;
	G8329<=G6232 and G231;
	G8339<=G6519 and G903;
	G8340<=G6369 and G909;
	G8350<=G6574 and G1594;
	G8385<=G3254 and G228;
	G8386<=G6314 and G234;
	G8387<=G6232 and G240;
	G8394<=G3410 and G906;
	G8395<=G6519 and G912;
	G8396<=G6369 and G918;
	G8406<=G6783 and G1597;
	G8407<=G6574 and G1603;
	G8417<=G6838 and G2288;
	G8431<=G3254 and G237;
	G8432<=G6314 and G243;
	G8433<=G6232 and G249;
	G8437<=G3410 and G915;
	G8438<=G6519 and G921;
	G8439<=G6369 and G927;
	G8446<=G3566 and G1600;
	G8447<=G6783 and G1606;
	G8448<=G6574 and G1612;
	G8458<=G7085 and G2291;
	G8459<=G6838 and G2297;
	G8463<=G3254 and G246;
	G8464<=G6314 and G252;
	G8465<=G6232 and G258;
	G8466<=G3410 and G924;
	G8467<=G6519 and G930;
	G8468<=G6369 and G936;
	G8472<=G3566 and G1609;
	G8473<=G6783 and G1615;
	G8474<=G6574 and G1621;
	G8481<=G3722 and G2294;
	G8482<=G7085 and G2300;
	G8483<=G6838 and G2306;
	G8484<=G6232 and G186;
	G8485<=G3254 and G255;
	G8486<=G6314 and G261;
	G8487<=G6232 and G267;
	G8488<=G3410 and G933;
	G8489<=G6519 and G939;
	G8490<=G6369 and G945;
	G8491<=G3566 and G1618;
	G8492<=G6783 and G1624;
	G8493<=G6574 and G1630;
	G8497<=G3722 and G2303;
	G8498<=G7085 and G2309;
	G8499<=G6838 and G2315;
	G8500<=G6314 and G189;
	G8501<=G6232 and G195;
	G8502<=G3254 and G264;
	G8503<=G6314 and G270;
	G8504<=G6369 and G873;
	G8505<=G3410 and G942;
	G8506<=G6519 and G948;
	G8507<=G6369 and G954;
	G8508<=G3566 and G1627;
	G8509<=G6783 and G1633;
	G8510<=G6574 and G1639;
	G8511<=G3722 and G2312;
	G8512<=G7085 and G2318;
	G8513<=G6838 and G2324;
	G8515<=G3254 and G192;
	G8516<=G6314 and G198;
	G8517<=G6232 and G204;
	G8518<=G3254 and G273;
	G8519<=G6519 and G876;
	G8520<=G6369 and G882;
	G8521<=G3410 and G951;
	G8522<=G6519 and G957;
	G8523<=G6574 and G1567;
	G8524<=G3566 and G1636;
	G8525<=G6783 and G1642;
	G8526<=G6574 and G1648;
	G8527<=G3722 and G2321;
	G8528<=G7085 and G2327;
	G8529<=G6838 and G2333;
	G8531<=G3254 and G201;
	G8532<=G6314 and G207;
	G8534<=G3410 and G879;
	G8535<=G6519 and G885;
	G8536<=G6369 and G891;
	G8537<=G3410 and G960;
	G8538<=G6783 and G1570;
	G8539<=G6574 and G1576;
	G8540<=G3566 and G1645;
	G8541<=G6783 and G1651;
	G8542<=G6838 and G2261;
	G8543<=G3722 and G2330;
	G8544<=G7085 and G2336;
	G8545<=G6838 and G2342;
	G8546<=G3254 and G210;
	G8548<=G3410 and G888;
	G8549<=G6519 and G894;
	G8551<=G3566 and G1573;
	G8552<=G6783 and G1579;
	G8553<=G6574 and G1585;
	G8554<=G3566 and G1654;
	G8555<=G7085 and G2264;
	G8556<=G6838 and G2270;
	G8557<=G3722 and G2339;
	G8558<=G7085 and G2345;
	G8559<=G3410 and G897;
	G8561<=G3566 and G1582;
	G8562<=G6783 and G1588;
	G8564<=G3722 and G2267;
	G8565<=G7085 and G2273;
	G8566<=G6838 and G2279;
	G8567<=G3722 and G2348;
	G8570<=G3566 and G1591;
	G8572<=G3722 and G2276;
	G8573<=G7085 and G2282;
	G8576<=G3722 and G2285;
	G8601<=G6643 and G7153;
	G8612<=G3338 and G6908;
	G8613<=G6945 and G7349;
	G8621<=G6486 and G6672;
	G8625<=G3494 and G7158;
	G8626<=G7195 and G7479;
	G8631<=G6751 and G6974;
	G8635<=G3650 and G7354;
	G8636<=G7391 and G7535;
	G8650<=G7053 and G7224;
	G8654<=G3806 and G7484;
	G8666<=G7303 and G7420;
	G8676<=G6643 and G7838;
	G8687<=G3338 and G7827;
	G8688<=G6945 and G7858;
	G8703<=G6486 and G7819;
	G8704<=G6643 and G7996;
	G8705<=G3494 and G7842;
	G8706<=G7195 and G7888;
	G8717<=G3338 and G7953;
	G8722<=G6751 and G7830;
	G8723<=G6945 and G8071;
	G8724<=G3650 and G7862;
	G8725<=G7391 and G7912;
	G8751<=G6486 and G7906;
	G8755<=G3494 and G8004;
	G8760<=G7053 and G7845;
	G8761<=G7195 and G8156;
	G8762<=G3806 and G7892;
	G8774<=G6751 and G7958;
	G8778<=G3650 and G8079;
	G8783<=G7303 and G7865;
	G8784<=G7391 and G8242;
	G8797<=G7053 and G8009;
	G8801<=G3806 and G8164;
	G8816<=G7303 and G8084;
	G8841<=G6486 and G490;
	G8842<=G6512 and G5508;
	G8861<=G6643 and G493;
	G8868<=G6751 and G1177;
	G8869<=G6776 and G5552;
	G8892<=G3338 and G496;
	G8899<=G6945 and G1180;
	G8906<=G7053 and G1871;
	G8907<=G7078 and G5598;
	G8932<=G3494 and G1183;
	G8939<=G7195 and G1874;
	G8946<=G7303 and G2565;
	G8947<=G7328 and G5615;
	G8972<=G3650 and G1877;
	G8979<=G7391 and G2568;
	G9004<=G3806 and G2571;
	G9009<=G6486 and G565;
	G9026<=G5438 and G7610;
	G9033<=G6643 and G567;
	G9034<=G6751 and G1251;
	G9047<=G6448 and G7616;
	G9048<=G3338 and G489;
	G9049<=G5473 and G7619;
	G9056<=G6945 and G1253;
	G9057<=G7053 and G1945;
	G9061<=G3306 and G7623;
	G9062<=G5438 and G7626;
	G9063<=G5438 and G7629;
	G9064<=G6713 and G7632;
	G9065<=G3494 and G1176;
	G9066<=G5512 and G7635;
	G9073<=G7195 and G1947;
	G9074<=G7303 and G2639;
	G9075<=G6448 and G7643;
	G9076<=G5438 and G7646;
	G9077<=G6448 and G7649;
	G9078<=G3462 and G7652;
	G9079<=G5473 and G7655;
	G9080<=G5473 and G7658;
	G9081<=G7015 and G7661;
	G9082<=G3650 and G1870;
	G9083<=G5556 and G7664;
	G9090<=G7391 and G2641;
	G9091<=G3306 and G7670;
	G9092<=G6448 and G7673;
	G9093<=G3306 and G7676;
	G9094<=G6713 and G7679;
	G9095<=G5473 and G7682;
	G9096<=G6713 and G7685;
	G9097<=G3618 and G7688;
	G9098<=G5512 and G7691;
	G9099<=G5512 and G7694;
	G9100<=G7265 and G7697;
	G9101<=G3806 and G2564;
	G9102<=G3306 and G7703;
	G9103<=G3462 and G7706;
	G9104<=G6713 and G7709;
	G9105<=G3462 and G7712;
	G9106<=G7015 and G7715;
	G9107<=G5512 and G7718;
	G9108<=G7015 and G7721;
	G9109<=G3774 and G7724;
	G9110<=G5556 and G7727;
	G9111<=G5556 and G7730;
	G9112<=G3462 and G7733;
	G9113<=G3618 and G7736;
	G9114<=G7015 and G7739;
	G9115<=G3618 and G7742;
	G9116<=G7265 and G7745;
	G9117<=G5556 and G7748;
	G9118<=G7265 and G7751;
	G9119<=G5438 and G7754;
	G9120<=G3618 and G7757;
	G9121<=G3774 and G7760;
	G9122<=G7265 and G7763;
	G9123<=G3774 and G7766;
	G9124<=G6448 and G7769;
	G9125<=G5473 and G7776;
	G9126<=G3774 and G7779;
	G9127<=G3306 and G7782;
	G9131<=G6713 and G7785;
	G9132<=G5512 and G7792;
	G9133<=G3462 and G7796;
	G9137<=G7015 and G7799;
	G9138<=G5556 and G7806;
	G9139<=G3618 and G7809;
	G9143<=G7265 and G7812;
	G9145<=G3774 and G7823;
	G9241<=G6232 and G7950;
	G9301<=G6314 and G7990;
	G9302<=G6232 and G7993;
	G9319<=G6369 and G8001;
	G9364<=G3254 and G8053;
	G9365<=G6314 and G8056;
	G9366<=G6232 and G8059;
	G9367<=G6232 and G8062;
	G9382<=G6519 and G8065;
	G9383<=G6369 and G8068;
	G9400<=G6574 and G8076;
	G9438<=G3254 and G8123;
	G9439<=G6314 and G8126;
	G9440<=G6232 and G8129;
	G9441<=G6314 and G8132;
	G9442<=G6232 and G8135;
	G9461<=G3410 and G8138;
	G9462<=G6519 and G8141;
	G9463<=G6369 and G8144;
	G9464<=G6369 and G8147;
	G9479<=G6783 and G8150;
	G9480<=G6574 and G8153;
	G9497<=G6838 and G8161;
	G9518<=G3254 and G8191;
	G9519<=G6314 and G8194;
	G9520<=G6232 and G8197;
	G9521<=G3254 and G8200;
	G9522<=G6314 and G8203;
	G9523<=G6232 and G8206;
	G9534<=G7772 and G6135 and G538;
	G9580<=G3410 and G8209;
	G9581<=G6519 and G8212;
	G9582<=G6369 and G8215;
	G9583<=G6519 and G8218;
	G9584<=G6369 and G8221;
	G9603<=G3566 and G8224;
	G9604<=G6783 and G8227;
	G9605<=G6574 and G8230;
	G9606<=G6574 and G8233;
	G9621<=G7085 and G8236;
	G9622<=G6838 and G8239;
	G9630<=G3254 and G3922;
	G9631<=G6314 and G3925;
	G9632<=G6232 and G3928;
	G9633<=G3254 and G3931;
	G9634<=G6314 and G3934;
	G9635<=G6232 and G3937;
	G9636<=I16735 and I16736;
	G9639<=G5438 and G408;
	G9647<=G6678 and G3942;
	G9648<=G6678 and G3945;
	G9660<=G3410 and G3948;
	G9661<=G6519 and G3951;
	G9662<=G6369 and G3954;
	G9663<=G3410 and G3957;
	G9664<=G6519 and G3960;
	G9665<=G6369 and G3963;
	G9676<=G7788 and G6145 and G1224;
	G9722<=G3566 and G3966;
	G9723<=G6783 and G3969;
	G9724<=G6574 and G3972;
	G9725<=G6783 and G3975;
	G9726<=G6574 and G3978;
	G9745<=G3722 and G3981;
	G9746<=G7085 and G3984;
	G9747<=G6838 and G3987;
	G9748<=G6838 and G3990;
	G9759<=G3254 and G4000;
	G9760<=G6314 and G4003;
	G9761<=G6232 and G4006;
	G9762<=G3254 and G4009;
	G9763<=G6314 and G4012;
	G9764<=G6448 and G411;
	G9765<=G5438 and G417;
	G9766<=G5438 and G4017;
	G9773<=G6912 and G4020;
	G9774<=G6678 and G4023;
	G9775<=G6912 and G4026;
	G9776<=G3410 and G4029;
	G9777<=G6519 and G4032;
	G9778<=G6369 and G4035;
	G9779<=G3410 and G4038;
	G9780<=G6519 and G4041;
	G9781<=G6369 and G4044;
	G9782<=I16826 and I16827;
	G9785<=G5473 and G1095;
	G9793<=G6980 and G4049;
	G9794<=G6980 and G4052;
	G9806<=G3566 and G4055;
	G9807<=G6783 and G4058;
	G9808<=G6574 and G4061;
	G9809<=G3566 and G4064;
	G9810<=G6783 and G4067;
	G9811<=G6574 and G4070;
	G9822<=G7802 and G6166 and G1918;
	G9868<=G3722 and G4073;
	G9869<=G7085 and G4076;
	G9870<=G6838 and G4079;
	G9871<=G7085 and G4082;
	G9872<=G6838 and G4085;
	G9887<=G6232 and G4095;
	G9888<=G3254 and G4098;
	G9889<=G6314 and G4101;
	G9890<=G6232 and G4104;
	G9891<=G3254 and G4107;
	G9892<=G3306 and G414;
	G9893<=G6448 and G420;
	G9894<=G6448 and G4112;
	G9901<=G3366 and G4115;
	G9902<=G6912 and G4118;
	G9903<=G6678 and G4121;
	G9904<=G3366 and G4124;
	G9905<=G3410 and G4127;
	G9906<=G6519 and G4130;
	G9907<=G6369 and G4133;
	G9908<=G3410 and G4136;
	G9909<=G6519 and G4139;
	G9910<=G6713 and G1098;
	G9911<=G5473 and G1104;
	G9912<=G5473 and G4144;
	G9919<=G7162 and G4147;
	G9920<=G6980 and G4150;
	G9921<=G7162 and G4153;
	G9922<=G3566 and G4156;
	G9923<=G6783 and G4159;
	G9924<=G6574 and G4162;
	G9925<=G3566 and G4165;
	G9926<=G6783 and G4168;
	G9927<=G6574 and G4171;
	G9928<=I16930 and I16931;
	G9931<=G5512 and G1789;
	G9939<=G7230 and G4176;
	G9940<=G7230 and G4179;
	G9952<=G3722 and G4182;
	G9953<=G7085 and G4185;
	G9954<=G6838 and G4188;
	G9955<=G3722 and G4191;
	G9956<=G7085 and G4194;
	G9957<=G6838 and G4197;
	G9968<=G7815 and G6193 and G2612;
	G10007<=G6314 and G4205;
	G10008<=G6232 and G4208;
	G10009<=G3254 and G4211;
	G10010<=G6314 and G4214;
	G10011<=G5438 and G4217;
	G10012<=G3306 and G423;
	G10013<=G3306 and G4221;
	G10014<=G5438 and G429;
	G10024<=G3398 and G6912;
	G10035<=G3366 and G4225;
	G10036<=G6912 and G4228;
	G10037<=G6678 and G4231;
	G10041<=G6369 and G4234;
	G10042<=G3410 and G4237;
	G10043<=G6519 and G4240;
	G10044<=G6369 and G4243;
	G10045<=G3410 and G4246;
	G10046<=G3462 and G1101;
	G10047<=G6713 and G1107;
	G10048<=G6713 and G4251;
	G10055<=G3522 and G4254;
	G10056<=G7162 and G4257;
	G10057<=G6980 and G4260;
	G10058<=G3522 and G4263;
	G10059<=G3566 and G4266;
	G10060<=G6783 and G4269;
	G10061<=G6574 and G4272;
	G10062<=G3566 and G4275;
	G10063<=G6783 and G4278;
	G10064<=G7015 and G1792;
	G10065<=G5512 and G1798;
	G10066<=G5512 and G4283;
	G10073<=G7358 and G4286;
	G10074<=G7230 and G4289;
	G10075<=G7358 and G4292;
	G10076<=G3722 and G4295;
	G10077<=G7085 and G4298;
	G10078<=G6838 and G4301;
	G10079<=G3722 and G4304;
	G10080<=G7085 and G4307;
	G10081<=G6838 and G4310;
	G10082<=I17042 and I17043;
	G10085<=G5556 and G2483;
	G10093<=G7426 and G4315;
	G10094<=G7426 and G4318;
	G10101<=G3254 and G4329;
	G10102<=G6314 and G4332;
	G10103<=G3254 and G4335;
	G10104<=G6448 and G4340;
	G10105<=G5438 and G4343;
	G10106<=G6448 and G432;
	G10107<=G5438 and G438;
	G10108<=G6486 and G569;
	G10112<=G3366 and G4348;
	G10113<=G6912 and G4351;
	G10114<=G6678 and G4354;
	G10115<=G6678 and G4357;
	G10116<=G6519 and G4360;
	G10117<=G6369 and G4363;
	G10118<=G3410 and G4366;
	G10119<=G6519 and G4369;
	G10120<=G5473 and G4372;
	G10121<=G3462 and G1110;
	G10122<=G3462 and G4376;
	G10123<=G5473 and G1116;
	G10133<=G3554 and G7162;
	G10144<=G3522 and G4380;
	G10145<=G7162 and G4383;
	G10146<=G6980 and G4386;
	G10150<=G6574 and G4389;
	G10151<=G3566 and G4392;
	G10152<=G6783 and G4395;
	G10153<=G6574 and G4398;
	G10154<=G3566 and G4401;
	G10155<=G3618 and G1795;
	G10156<=G7015 and G1801;
	G10157<=G7015 and G4406;
	G10164<=G3678 and G4409;
	G10165<=G7358 and G4412;
	G10166<=G7230 and G4415;
	G10167<=G3678 and G4418;
	G10168<=G3722 and G4421;
	G10169<=G7085 and G4424;
	G10170<=G6838 and G4427;
	G10171<=G3722 and G4430;
	G10172<=G7085 and G4433;
	G10173<=G7265 and G2486;
	G10174<=G5556 and G2492;
	G10175<=G5556 and G4438;
	G10182<=G7488 and G4441;
	G10183<=G7426 and G4444;
	G10184<=G7488 and G4447;
	G10186<=G3013 and G7466 and G3024 and I17156;
	G10192<=G3254 and G4453;
	G10193<=G3306 and G4465;
	G10194<=G6448 and G4468;
	G10195<=G5438 and G4471;
	G10196<=G3306 and G435;
	G10197<=G6448 and G441;
	G10198<=G6643 and G571;
	G10199<=G6486 and G4476;
	G10200<=G6486 and G587;
	G10201<=G3366 and G4480;
	G10202<=G6912 and G4483;
	G10203<=G6678 and G4486;
	G10204<=G6912 and G4489;
	G10205<=G6678 and G4492;
	G10206<=G3410 and G4498;
	G10207<=G6519 and G4501;
	G10208<=G3410 and G4504;
	G10209<=G6713 and G4509;
	G10210<=G5473 and G4512;
	G10211<=G6713 and G1119;
	G10212<=G5473 and G1125;
	G10213<=G6751 and G1255;
	G10217<=G3522 and G4517;
	G10218<=G7162 and G4520;
	G10219<=G6980 and G4523;
	G10220<=G6980 and G4526;
	G10221<=G6783 and G4529;
	G10222<=G6574 and G4532;
	G10223<=G3566 and G4535;
	G10224<=G6783 and G4538;
	G10225<=G5512 and G4541;
	G10226<=G3618 and G1804;
	G10227<=G3618 and G4545;
	G10228<=G5512 and G1810;
	G10238<=G3710 and G7358;
	G10249<=G3678 and G4549;
	G10250<=G7358 and G4552;
	G10251<=G7230 and G4555;
	G10255<=G6838 and G4558;
	G10256<=G3722 and G4561;
	G10257<=G7085 and G4564;
	G10258<=G6838 and G4567;
	G10259<=G3722 and G4570;
	G10260<=G3774 and G2489;
	G10261<=G7265 and G2495;
	G10262<=G7265 and G4575;
	G10269<=G3834 and G4578;
	G10270<=G7488 and G4581;
	G10271<=G7426 and G4584;
	G10272<=G3834 and G4587;
	G10279<=G3306 and G4592;
	G10280<=G6448 and G4595;
	G10281<=G5438 and G4598;
	G10282<=G3306 and G444;
	G10283<=G3338 and G573;
	G10284<=G6643 and G4603;
	G10285<=G6486 and G4606;
	G10286<=G6643 and G590;
	G10287<=G6486 and G596;
	G10288<=G3366 and G4611;
	G10289<=G6912 and G4614;
	G10290<=G6678 and G4617;
	G10291<=G3366 and G4620;
	G10292<=G6912 and G4623;
	G10293<=G6678 and G4626;
	G10294<=G3410 and G4629;
	G10295<=G3462 and G4641;
	G10296<=G6713 and G4644;
	G10297<=G5473 and G4647;
	G10298<=G3462 and G1122;
	G10299<=G6713 and G1128;
	G10300<=G6945 and G1257;
	G10301<=G6751 and G4652;
	G10302<=G6751 and G1273;
	G10303<=G3522 and G4656;
	G10304<=G7162 and G4659;
	G10305<=G6980 and G4662;
	G10306<=G7162 and G4665;
	G10307<=G6980 and G4668;
	G10308<=G3566 and G4674;
	G10309<=G6783 and G4677;
	G10310<=G3566 and G4680;
	G10311<=G7015 and G4685;
	G10312<=G5512 and G4688;
	G10313<=G7015 and G1813;
	G10314<=G5512 and G1819;
	G10315<=G7053 and G1949;
	G10319<=G3678 and G4693;
	G10320<=G7358 and G4696;
	G10321<=G7230 and G4699;
	G10322<=G7230 and G4702;
	G10323<=G7085 and G4705;
	G10324<=G6838 and G4708;
	G10325<=G3722 and G4711;
	G10326<=G7085 and G4714;
	G10327<=G5556 and G4717;
	G10328<=G3774 and G2498;
	G10329<=G3774 and G4721;
	G10330<=G5556 and G2504;
	G10340<=G3866 and G7488;
	G10351<=G3834 and G4725;
	G10352<=G7488 and G4728;
	G10353<=G7426 and G4731;
	G10360<=G3306 and G4737;
	G10361<=G6448 and G4740;
	G10362<=G3338 and G4743;
	G10363<=G6643 and G4746;
	G10364<=G6486 and G4749;
	G10365<=G3338 and G593;
	G10366<=G6643 and G599;
	G10367<=G3366 and G4754;
	G10368<=G6912 and G4757;
	G10369<=G6678 and G4760;
	G10370<=G3366 and G4763;
	G10371<=G6912 and G4766;
	G10372<=G3462 and G4769;
	G10373<=G6713 and G4772;
	G10374<=G5473 and G4775;
	G10375<=G3462 and G1131;
	G10376<=G3494 and G1259;
	G10377<=G6945 and G4780;
	G10378<=G6751 and G4783;
	G10379<=G6945 and G1276;
	G10380<=G6751 and G1282;
	G10381<=G3522 and G4788;
	G10382<=G7162 and G4791;
	G10383<=G6980 and G4794;
	G10384<=G3522 and G4797;
	G10385<=G7162 and G4800;
	G10386<=G6980 and G4803;
	G10387<=G3566 and G4806;
	G10388<=G3618 and G4818;
	G10389<=G7015 and G4821;
	G10390<=G5512 and G4824;
	G10391<=G3618 and G1816;
	G10392<=G7015 and G1822;
	G10393<=G7195 and G1951;
	G10394<=G7053 and G4829;
	G10395<=G7053 and G1967;
	G10396<=G3678 and G4833;
	G10397<=G7358 and G4836;
	G10398<=G7230 and G4839;
	G10399<=G7358 and G4842;
	G10400<=G7230 and G4845;
	G10401<=G3722 and G4851;
	G10402<=G7085 and G4854;
	G10403<=G3722 and G4857;
	G10404<=G7265 and G4862;
	G10405<=G5556 and G4865;
	G10406<=G7265 and G2507;
	G10407<=G5556 and G2513;
	G10408<=G7303 and G2643;
	G10412<=G3834 and G4870;
	G10413<=G7488 and G4873;
	G10414<=G7426 and G4876;
	G10415<=G7426 and G4879;
	G10422<=G3306 and G4882;
	G10423<=G5438 and G4885;
	G10430<=G3338 and G4888;
	G10431<=G6643 and G4891;
	G10432<=G6486 and G4894;
	G10433<=G3338 and G602;
	G10434<=G6486 and G605;
	G10435<=G3366 and G4899;
	G10436<=G6912 and G4902;
	G10437<=G6678 and G4905;
	G10438<=G3366 and G4908;
	G10439<=G3462 and G4913;
	G10440<=G6713 and G4916;
	G10441<=G3494 and G4919;
	G10442<=G6945 and G4922;
	G10443<=G6751 and G4925;
	G10444<=G3494 and G1279;
	G10445<=G6945 and G1285;
	G10446<=G3522 and G4930;
	G10447<=G7162 and G4933;
	G10448<=G6980 and G4936;
	G10449<=G3522 and G4939;
	G10450<=G7162 and G4942;
	G10451<=G3618 and G4945;
	G10452<=G7015 and G4948;
	G10453<=G5512 and G4951;
	G10454<=G3618 and G1825;
	G10455<=G3650 and G1953;
	G10456<=G7195 and G4956;
	G10457<=G7053 and G4959;
	G10458<=G7195 and G1970;
	G10459<=G7053 and G1976;
	G10460<=G3678 and G4964;
	G10461<=G7358 and G4967;
	G10462<=G7230 and G4970;
	G10463<=G3678 and G4973;
	G10464<=G7358 and G4976;
	G10465<=G7230 and G4979;
	G10466<=G3722 and G4982;
	G10467<=G3774 and G4994;
	G10468<=G7265 and G4997;
	G10469<=G5556 and G5000;
	G10470<=G3774 and G2510;
	G10471<=G7265 and G2516;
	G10472<=G7391 and G2645;
	G10473<=G7303 and G5005;
	G10474<=G7303 and G2661;
	G10475<=G3834 and G5009;
	G10476<=G7488 and G5012;
	G10477<=G7426 and G5015;
	G10478<=G7488 and G5018;
	G10479<=G7426 and G5021;
	G10480<=G7466 and G7342 and I17429;
	G10485<=G6448 and G5024;
	G10492<=G3338 and G5027;
	G10493<=G6643 and G5030;
	G10494<=G6643 and G608;
	G10495<=G6486 and G614;
	G10496<=G3366 and G5035;
	G10497<=G6912 and G5038;
	G10498<=G3462 and G5041;
	G10499<=G5473 and G5044;
	G10506<=G3494 and G5047;
	G10507<=G6945 and G5050;
	G10508<=G6751 and G5053;
	G10509<=G3494 and G1288;
	G10510<=G6751 and G1291;
	G10511<=G3522 and G5058;
	G10512<=G7162 and G5061;
	G10513<=G6980 and G5064;
	G10514<=G3522 and G5067;
	G10515<=G3618 and G5072;
	G10516<=G7015 and G5075;
	G10517<=G3650 and G5078;
	G10518<=G7195 and G5081;
	G10519<=G7053 and G5084;
	G10520<=G3650 and G1973;
	G10521<=G7195 and G1979;
	G10522<=G3678 and G5089;
	G10523<=G7358 and G5092;
	G10524<=G7230 and G5095;
	G10525<=G3678 and G5098;
	G10526<=G7358 and G5101;
	G10527<=G3774 and G5104;
	G10528<=G7265 and G5107;
	G10529<=G5556 and G5110;
	G10530<=G3774 and G2519;
	G10531<=G3806 and G2647;
	G10532<=G7391 and G5115;
	G10533<=G7303 and G5118;
	G10534<=G7391 and G2664;
	G10535<=G7303 and G2670;
	G10536<=G3834 and G5123;
	G10537<=G7488 and G5126;
	G10538<=G7426 and G5129;
	G10539<=G3834 and G5132;
	G10540<=G7488 and G5135;
	G10541<=G7426 and G5138;
	G10548<=G3306 and G5142;
	G10555<=G3338 and G5145;
	G10556<=G3338 and G611;
	G10557<=G6643 and G617;
	G10558<=G3366 and G5150;
	G10559<=G6713 and G5153;
	G10566<=G3494 and G5156;
	G10567<=G6945 and G5159;
	G10568<=G6945 and G1294;
	G10569<=G6751 and G1300;
	G10570<=G3522 and G5164;
	G10571<=G7162 and G5167;
	G10572<=G3618 and G5170;
	G10573<=G5512 and G5173;
	G10580<=G3650 and G5176;
	G10581<=G7195 and G5179;
	G10582<=G7053 and G5182;
	G10583<=G3650 and G1982;
	G10584<=G7053 and G1985;
	G10585<=G3678 and G5187;
	G10586<=G7358 and G5190;
	G10587<=G7230 and G5193;
	G10588<=G3678 and G5196;
	G10589<=G3774 and G5201;
	G10590<=G7265 and G5204;
	G10591<=G3806 and G5207;
	G10592<=G7391 and G5210;
	G10593<=G7303 and G5213;
	G10594<=G3806 and G2667;
	G10595<=G7391 and G2673;
	G10596<=G3834 and G5218;
	G10597<=G7488 and G5221;
	G10598<=G7426 and G5224;
	G10599<=G3834 and G5227;
	G10600<=G7488 and G5230;
	G10604<=G3338 and G620;
	G10605<=G3462 and G5235;
	G10612<=G3494 and G5238;
	G10613<=G3494 and G1297;
	G10614<=G6945 and G1303;
	G10615<=G3522 and G5243;
	G10616<=G7015 and G5246;
	G10623<=G3650 and G5249;
	G10624<=G7195 and G5252;
	G10625<=G7195 and G1988;
	G10626<=G7053 and G1994;
	G10627<=G3678 and G5257;
	G10628<=G7358 and G5260;
	G10629<=G3774 and G5263;
	G10630<=G5556 and G5266;
	G10637<=G3806 and G5269;
	G10638<=G7391 and G5272;
	G10639<=G7303 and G5275;
	G10640<=G3806 and G2676;
	G10641<=G7303 and G2679;
	G10642<=G3834 and G5280;
	G10643<=G7488 and G5283;
	G10644<=G7426 and G5286;
	G10645<=G3834 and G5289;
	G10650<=G6678 and G5293;
	G10651<=G3494 and G1306;
	G10652<=G3618 and G5298;
	G10659<=G3650 and G5301;
	G10660<=G3650 and G1991;
	G10661<=G7195 and G1997;
	G10662<=G3678 and G5306;
	G10663<=G7265 and G5309;
	G10670<=G3806 and G5312;
	G10671<=G7391 and G5315;
	G10672<=G7391 and G2682;
	G10673<=G7303 and G2688;
	G10674<=G3834 and G5320;
	G10675<=G7488 and G5323;
	G10678<=G6912 and G5327;
	G10680<=G6980 and G5330;
	G10681<=G3650 and G2000;
	G10682<=G3774 and G5335;
	G10689<=G3806 and G5338;
	G10690<=G3806 and G2685;
	G10691<=G7391 and G2691;
	G10692<=G3834 and G5343;
	G10693<=G7462 and G7522 and G2924 and G7545;
	G10704<=G3366 and G5352;
	G10707<=G7162 and G5355;
	G10709<=G7230 and G5358;
	G10710<=G3806 and G2694;
	G10711<=G7595 and G7600 and I17599;
	G10724<=G3522 and G5369;
	G10727<=G7358 and G5372;
	G10729<=G7426 and G5375;
	G10745<=G3678 and G5382;
	G10748<=G7488 and G5385;
	G10764<=G3834 and G5391;
	G11347<=G6232 and G213;
	G11420<=G6314 and G216;
	G11421<=G6232 and G222;
	G11431<=G6369 and G900;
	G11607<=G5871 and G8360;
	G11612<=G5881 and G8378;
	G11637<=G5918 and G8427;
	G11771<=G554 and G8622;
	G11788<=G1240 and G8632;
	G11805<=G6173 and G8643;
	G11814<=G1934 and G8651;
	G11816<=G7869 and G8655;
	G11838<=G6205 and G8659;
	G11847<=G2628 and G8667;
	G11851<=G7849 and G8670;
	G11880<=G6294 and G8678;
	G11885<=G7834 and G8684;
	G11922<=G6431 and G8690;
	G11926<=G8169 and G8696;
	G11966<=G8090 and G8708;
	G11967<=G7967 and G8711;
	G12012<=G8015 and G8745;
	G12069<=G7964 and G8763;
	G12070<=G8018 and G8766;
	G12128<=G7916 and G8785;
	G12129<=G7872 and G8788;
	G12186<=G8093 and G8805;
	G12273<=G8172 and G8829;
	G12274<=G7900 and G8832;
	G12307<=G7919 and G8853;
	G12330<=G8246 and G8879;
	G12331<=G7927 and G8882;
	G12353<=G7852 and G8915;
	G12376<=G7974 and G8949;
	G12419<=G8028 and G9006;
	G12429<=G8101 and G9044;
	G12477<=G7822 and G9128;
	G12494<=G7833 and G9134;
	G12514<=G7848 and G9140;
	G12531<=G7868 and G9146;
	G12650<=G6149 and G9290;
	G12876<=I19937 and I19938;
	G12908<=G7899 and G10004;
	G12916<=I19971 and I19972;
	G12938<=G8179 and G10096;
	G12945<=I19996 and I19997;
	G12966<=G7926 and G10189;
	G12974<=I20021 and I20022;
	G12989<=G8254 and G10273;
	G12990<=G8180 and G10276;
	G13000<=G7973 and G10357;
	G13004<=G10186 and G8317;
	G13009<=G3995 and G10416;
	G13010<=G8255 and G10419;
	G13023<=G8027 and G10482;
	G13031<=G7879 and G10542;
	G13032<=G3996 and G10545;
	G13042<=G8100 and G10601;
	G13055<=G7471 and G7570 and I20100;
	G13056<=G4092 and G10646;
	G13082<=I20131 and I20132;
	G13110<=G10693 and G2883 and G7562 and G10711;
	G13247<=G298 and G11032;
	G13266<=G5628 and G11088;
	G13270<=G985 and G11102;
	G13289<=G5647 and G11141;
	G13291<=G5656 and G11154;
	G13295<=G1679 and G11170;
	G13316<=G5675 and G11210;
	G13320<=G5685 and G11225;
	G13322<=G5694 and G11240;
	G13326<=G2373 and G11256;
	G13335<=G5708 and G11278;
	G13340<=G5727 and G11294;
	G13343<=G5737 and G11309;
	G13345<=G5746 and G11324;
	G13355<=G5756 and G11355;
	G13360<=G5766 and G11373;
	G13365<=G5785 and G11389;
	G13368<=G5795 and G11404;
	G13385<=G5815 and G11441;
	G13390<=G5825 and G11459;
	G13395<=G5844 and G11475;
	G13477<=G6016 and G12191;
	G13479<=G6017 and G12196;
	G13480<=G6018 and G12197;
	G13481<=G5864 and G11603;
	G13483<=G6020 and G12209;
	G13484<=G6021 and G12210;
	G13485<=G6022 and G12211;
	G13486<=G6023 and G12212;
	G13487<=G5874 and G11608;
	G13488<=G6025 and G12218;
	G13489<=G6026 and G12219;
	G13490<=G6027 and G12220;
	G13491<=G6028 and G12221;
	G13492<=G2371 and G12222;
	G13493<=G5887 and G11613;
	G13496<=G6032 and G12246;
	G13498<=G6033 and G12251;
	G13499<=G6034 and G12252;
	G13500<=G5911 and G11633;
	G13502<=G6036 and G12264;
	G13503<=G6037 and G12265;
	G13504<=G6038 and G12266;
	G13505<=G6039 and G12267;
	G13506<=G5921 and G11638;
	G13513<=G6043 and G12289;
	G13515<=G6044 and G12294;
	G13516<=G6045 and G12295;
	G13517<=G5950 and G11656;
	G13527<=G6047 and G12325;
	G13609<=G6141 and G12456;
	G13619<=G6162 and G12466;
	G13623<=G5428 and G12472;
	G13625<=G6173 and G12476;
	G13631<=G6189 and G12481;
	G13634<=G12776 and G8617;
	G13636<=G6205 and G12493;
	G13642<=G6221 and G12498;
	G13643<=G5431 and G12502;
	G13645<=G6281 and G12504;
	G13646<=G7772 and G12505;
	G13648<=G6294 and G12513;
	G13654<=G8093 and G11791;
	G13655<=G7540 and G12518;
	G13656<=G12776 and G8640;
	G13671<=G6418 and G12521;
	G13672<=G7788 and G12522;
	G13674<=G6431 and G12530;
	G13675<=G7561 and G12532;
	G13676<=G5434 and G12533;
	G13701<=G6623 and G12536;
	G13702<=G7802 and G12537;
	G13703<=G8018 and G11848;
	G13704<=G7581 and G12542;
	G13705<=G12776 and G8673;
	G13738<=G6887 and G12545;
	G13739<=G7815 and G12546;
	G13740<=G6636 and G12547;
	G13755<=G7347 and G12551;
	G13787<=G7967 and G11923;
	G13788<=G6897 and G12553;
	G13789<=G7140 and G12554;
	G13790<=G7475 and G12558;
	G13796<=G7477 and G12559;
	G13815<=G7139 and G12560;
	G13816<=G7530 and G12596;
	G13818<=G7531 and G12597;
	G13824<=G7533 and G12598;
	G13833<=G7919 and G12009;
	G13834<=G7336 and G12599;
	G13835<=G7461 and G12600;
	G13837<=G7556 and G12642;
	G13839<=G7557 and G12643;
	G13845<=G7559 and G12644;
	G13846<=G7460 and G12645;
	G13847<=G7521 and G12646;
	G13851<=G7579 and G12688;
	G13853<=G7580 and G12689;
	G13854<=G5349 and G12690;
	G13855<=G7541 and G12691;
	G13860<=G7593 and G12742;
	G13862<=G5366 and G12743;
	G13865<=G548 and G12748;
	G13870<=G7582 and G12768;
	G13871<=G7898 and G12775;
	G13878<=G7610 and G12782;
	G13880<=G1234 and G12790;
	G13884<=G7594 and G12807;
	G13892<=G7616 and G12815;
	G13900<=G7619 and G12821;
	G13902<=G1928 and G12829;
	G13904<=G7337 and G12843;
	G13905<=G7925 and G12847;
	G13913<=G7623 and G12850;
	G13914<=G7626 and G12851;
	G13933<=G7632 and G12853;
	G13941<=G7635 and G12859;
	G13943<=G2622 and G12867;
	G13944<=G7141 and G12874;
	G13952<=G7643 and G12881;
	G13953<=G7646 and G12882;
	G13969<=G7652 and G12891;
	G13970<=G7655 and G12892;
	G13989<=G7661 and G12894;
	G13997<=G7664 and G12900;
	G13998<=G7972 and G12907;
	G14006<=G7670 and G12914;
	G14007<=G7673 and G12915;
	G14022<=G7679 and G12921;
	G14023<=G7682 and G12922;
	G14039<=G7688 and G12931;
	G14040<=G7691 and G12932;
	G14059<=G7697 and G12934;
	G14067<=G7703 and G12940;
	G14097<=G7706 and G12943;
	G14098<=G7709 and G12944;
	G14113<=G7715 and G12950;
	G14114<=G7718 and G12951;
	G14130<=G7724 and G12960;
	G14131<=G7727 and G12961;
	G14143<=G8026 and G12965;
	G14182<=G7733 and G12969;
	G14212<=G7736 and G12972;
	G14213<=G7739 and G12973;
	G14228<=G7745 and G12979;
	G14229<=G7748 and G12980;
	G14297<=G7757 and G12993;
	G14327<=G7760 and G12996;
	G14328<=G7763 and G12997;
	G14336<=G8099 and G12998;
	G14419<=G7779 and G13003;
	G14690<=G7841 and G13101;
	G14724<=G7861 and G13117;
	G14752<=G7891 and G13130;
	G14767<=G13245 and G10765;
	G14773<=G7915 and G13141;
	G14884<=G8169 and G12548;
	G14894<=G3940 and G13148;
	G14956<=G11059 and G13151;
	G14957<=G4015 and G13152;
	G14958<=G4016 and G13153;
	G14975<=G4047 and G13154;
	G15020<=G8090 and G12561;
	G15030<=G4110 and G13158;
	G15031<=G4111 and G13159;
	G15046<=G4142 and G13161;
	G15047<=G4143 and G13162;
	G15064<=G4174 and G13163;
	G15093<=G7869 and G12601;
	G15094<=G7872 and G12604;
	G15104<=G4220 and G13167;
	G15105<=G4224 and G13168;
	G15126<=G4249 and G13169;
	G15127<=G4250 and G13170;
	G15142<=G4281 and G13172;
	G15143<=G4282 and G13173;
	G15160<=G4313 and G13174;
	G15171<=G8015 and G12647;
	G15172<=G4346 and G13176;
	G15173<=G4347 and G13177;
	G15178<=G640 and G12651;
	G15196<=G4375 and G13178;
	G15197<=G4379 and G13179;
	G15218<=G4404 and G13180;
	G15219<=G4405 and G13181;
	G15234<=G4436 and G13183;
	G15235<=G4437 and G13184;
	G15243<=G7849 and G12692;
	G15244<=G7852 and G12695;
	G15245<=G4474 and G13185;
	G15246<=G4475 and G13186;
	G15247<=G4479 and G13187;
	G15257<=G4357 and G12702;
	G15258<=G4515 and G13188;
	G15259<=G4516 and G13189;
	G15264<=G1326 and G12705;
	G15282<=G4544 and G13190;
	G15283<=G4548 and G13191;
	G15304<=G4573 and G13192;
	G15305<=G4574 and G13193;
	G15320<=G7964 and G12744;
	G15321<=G4601 and G13195;
	G15324<=G4609 and G13196;
	G15325<=G4610 and G13197;
	G15335<=G4489 and G12749;
	G15336<=G4492 and G12752;
	G15337<=G4650 and G13198;
	G15338<=G4651 and G13199;
	G15339<=G4655 and G13200;
	G15349<=G4526 and G12759;
	G15350<=G4691 and G13201;
	G15351<=G4692 and G13202;
	G15356<=G2020 and G12762;
	G15374<=G4720 and G13203;
	G15375<=G4724 and G13204;
	G15388<=G7834 and G12769;
	G15389<=G8246 and G12772;
	G15391<=G4752 and G13205;
	G15392<=G4753 and G13206;
	G15402<=G4620 and G12783;
	G15403<=G4623 and G12786;
	G15407<=G4778 and G13207;
	G15410<=G4786 and G13208;
	G15411<=G4787 and G13209;
	G15421<=G4665 and G12791;
	G15422<=G4668 and G12794;
	G15423<=G4827 and G13210;
	G15424<=G4828 and G13211;
	G15425<=G4832 and G13212;
	G15435<=G4702 and G12801;
	G15436<=G4868 and G13213;
	G15437<=G4869 and G13214;
	G15442<=G2714 and G12804;
	G15452<=G7916 and G12808;
	G15453<=G6898 and G12811;
	G15459<=G4897 and G13218;
	G15460<=G4898 and G13219;
	G15470<=G4763 and G12816;
	G15475<=G4928 and G13220;
	G15476<=G4929 and G13221;
	G15486<=G4797 and G12822;
	G15487<=G4800 and G12825;
	G15491<=G4954 and G13222;
	G15494<=G4962 and G13223;
	G15495<=G4963 and G13224;
	G15505<=G4842 and G12830;
	G15506<=G4845 and G12833;
	G15507<=G5003 and G13225;
	G15508<=G5004 and G13226;
	G15509<=G5008 and G13227;
	G15519<=G4879 and G12840;
	G15520<=G8172 and G12844;
	G15526<=G5033 and G13232;
	G15527<=G5034 and G13233;
	G15545<=G5056 and G13237;
	G15546<=G5057 and G13238;
	G15556<=G4939 and G12854;
	G15561<=G5087 and G13239;
	G15562<=G5088 and G13240;
	G15572<=G4973 and G12860;
	G15573<=G4976 and G12863;
	G15577<=G5113 and G13241;
	G15580<=G5121 and G13242;
	G15581<=G5122 and G13243;
	G15591<=G5018 and G12868;
	G15592<=G5021 and G12871;
	G15593<=G7897 and G13244;
	G15594<=G5148 and G13249;
	G15595<=G5149 and G13250;
	G15604<=G5162 and G13255;
	G15605<=G5163 and G13256;
	G15623<=G5185 and G13260;
	G15624<=G5186 and G13261;
	G15634<=G5098 and G12895;
	G15639<=G5216 and G13262;
	G15640<=G5217 and G13263;
	G15650<=G5132 and G12901;
	G15651<=G5135 and G12904;
	G15658<=G8177 and G13264;
	G15666<=G5233 and G13268;
	G15670<=G5241 and G13272;
	G15671<=G5242 and G13273;
	G15680<=G5255 and G13278;
	G15681<=G5256 and G13279;
	G15699<=G5278 and G13283;
	G15700<=G5279 and G13284;
	G15710<=G5227 and G12935;
	G15717<=G7924 and G13285;
	G15725<=G5296 and G13293;
	G15729<=G5304 and G13297;
	G15730<=G5305 and G13298;
	G15739<=G5318 and G13303;
	G15740<=G5319 and G13304;
	G15753<=G7542 and G12962;
	G15754<=G7837 and G13308;
	G15755<=G8178 and G13309;
	G15765<=G5333 and G13324;
	G15769<=G5341 and G13328;
	G15770<=G5342 and G13329;
	G15780<=G7471 and G3032 and I22028;
	G15781<=G7971 and G13330;
	G15793<=G5361 and G13347;
	G15801<=G7856 and G13351;
	G15802<=G8253 and G13352;
	G15817<=G8025 and G13373;
	G15828<=G7877 and G13398;
	G15829<=G7857 and G13400;
	G15840<=G8098 and G11620;
	G15852<=G7878 and G11642;
	G15902<=G7607 and G2920 and I22136;
	G15998<=G5469 and G11732;
	G16003<=G12013 and G10826;
	G16004<=G5587 and G11734;
	G16008<=G5504 and G11735;
	G16009<=G12071 and G10843;
	G16010<=G7639 and G11736;
	G16015<=G12013 and G10859;
	G16016<=G5601 and G11740;
	G16017<=G12130 and G10862;
	G16018<=G6149 and G11741;
	G16019<=G5507 and G11742;
	G16028<=G5543 and G11745;
	G16029<=G12071 and G10877;
	G16030<=G7667 and G11746;
	G16031<=G6227 and G11747;
	G16032<=G12187 and G10883;
	G16033<=G5546 and G11748;
	G16045<=G12013 and G10892;
	G16046<=G5618 and G11761;
	G16047<=G12130 and G10895;
	G16048<=G6170 and G11762;
	G16049<=G6638 and G11763;
	G16050<=G5590 and G11764;
	G16051<=G12235 and G10901;
	G16052<=G5591 and G11765;
	G16053<=G297 and G11770;
	G16066<=G12071 and G10912;
	G16067<=G7700 and G11774;
	G16068<=G6310 and G11775;
	G16069<=G5346 and G11776;
	G16070<=G12187 and G10921;
	G16071<=G5604 and G11777;
	G16072<=G12275 and G10924;
	G16073<=G5605 and G11778;
	G16074<=G5646 and G11782;
	G16081<=G3304 and G11783;
	G16089<=G984 and G11787;
	G16100<=G12130 and G10937;
	G16101<=G6197 and G11794;
	G16102<=G6905 and G11795;
	G16103<=G5621 and G11796;
	G16104<=G12235 and G10946;
	G16105<=G5622 and G11797;
	G16106<=G12308 and G10949;
	G16107<=G5666 and G11801;
	G16108<=G5667 and G11802;
	G16109<=G8277 and G11803;
	G16110<=G516 and G11804;
	G16111<=G5551 and G13215;
	G16112<=G5684 and G11808;
	G16119<=G3460 and G11809;
	G16127<=G1678 and G11813;
	G16133<=G6444 and G11817;
	G16134<=G5363 and G11818;
	G16135<=G12187 and G10980;
	G16136<=G5640 and G11819;
	G16137<=G12275 and G10983;
	G16138<=G5641 and G11820;
	G16139<=G5704 and G11824;
	G16140<=G5705 and G11825;
	G16141<=G5706 and G11826;
	G16152<=G517 and G11829;
	G16153<=G5592 and G13229;
	G16158<=G5718 and G11834;
	G16159<=G5719 and G11835;
	G16160<=G8286 and G11836;
	G16161<=G1202 and G11837;
	G16162<=G5597 and G13234;
	G16163<=G5736 and G11841;
	G16170<=G3616 and G11842;
	G16178<=G2372 and G11846;
	G16182<=G7149 and G11852;
	G16183<=G12235 and G11014;
	G16184<=G5663 and G11853;
	G16185<=G12308 and G11017;
	G16186<=G5753 and G11856;
	G16187<=G5754 and G11857;
	G16188<=G5755 and G11858;
	G16197<=G518 and G11862;
	G16198<=G5762 and G11866;
	G16199<=G5763 and G11867;
	G16200<=G5764 and G11868;
	G16211<=G1203 and G11871;
	G16212<=G5609 and G13252;
	G16217<=G5776 and G11876;
	G16218<=G5777 and G11877;
	G16219<=G8295 and G11878;
	G16220<=G1896 and G11879;
	G16221<=G5614 and G13257;
	G16222<=G5794 and G11883;
	G16229<=G3772 and G11884;
	G16237<=G5379 and G11886;
	G16238<=G12275 and G11066;
	G16239<=G5700 and G11887;
	G16240<=G5804 and G11891;
	G16241<=G5805 and G11892;
	G16242<=G5806 and G11893;
	G16250<=G519 and G11895;
	G16251<=G5812 and G11898;
	G16252<=G5813 and G11899;
	G16253<=G5814 and G11900;
	G16262<=G1204 and G11904;
	G16263<=G5821 and G11908;
	G16264<=G5822 and G11909;
	G16265<=G5823 and G11910;
	G16276<=G1897 and G11913;
	G16277<=G5634 and G13275;
	G16282<=G5835 and G11918;
	G16283<=G5836 and G11919;
	G16284<=G8304 and G11920;
	G16285<=G2590 and G11921;
	G16286<=G5639 and G13280;
	G16288<=G12308 and G11129;
	G16289<=G5853 and G11929;
	G16290<=G5854 and G11930;
	G16291<=G5855 and G11931;
	G16292<=G294 and G11932;
	G16298<=G520 and G11936;
	G16299<=G5860 and G11941;
	G16300<=G5861 and G11942;
	G16301<=G5862 and G11943;
	G16309<=G1205 and G11945;
	G16310<=G5868 and G11948;
	G16311<=G5869 and G11949;
	G16312<=G5870 and G11950;
	G16321<=G1898 and G11954;
	G16322<=G5877 and G11958;
	G16323<=G5878 and G11959;
	G16324<=G5879 and G11960;
	G16335<=G2591 and G11963;
	G16336<=G5662 and G13300;
	G16342<=G5894 and G11968;
	G16343<=G5895 and G11969;
	G16344<=G5896 and G11970;
	G16345<=G5897 and G11971;
	G16346<=G295 and G11972;
	G16347<=G5900 and G11982;
	G16348<=G5901 and G11983;
	G16349<=G5902 and G11984;
	G16350<=G981 and G11985;
	G16356<=G1206 and G11989;
	G16357<=G5907 and G11994;
	G16358<=G5908 and G11995;
	G16359<=G5909 and G11996;
	G16367<=G1899 and G11998;
	G16368<=G5915 and G12001;
	G16369<=G5916 and G12002;
	G16370<=G5917 and G12003;
	G16379<=G2592 and G12007;
	G16380<=G5925 and G12020;
	G16381<=G5926 and G12021;
	G16382<=G5927 and G12022;
	G16383<=G5928 and G12023;
	G16384<=G296 and G12024;
	G16385<=G5714 and G13336;
	G16386<=G5933 and G12037;
	G16387<=G5934 and G12038;
	G16388<=G5935 and G12039;
	G16389<=G5936 and G12040;
	G16390<=G982 and G12041;
	G16391<=G5939 and G12051;
	G16392<=G5940 and G12052;
	G16393<=G5941 and G12053;
	G16394<=G1675 and G12054;
	G16400<=G1900 and G12058;
	G16401<=G5946 and G12063;
	G16402<=G5947 and G12064;
	G16403<=G5948 and G12065;
	G16411<=G2593 and G12067;
	G16413<=G5954 and G12075;
	G16414<=G5955 and G12076;
	G16415<=G5956 and G12077;
	G16416<=G5957 and G12078;
	G16417<=G5759 and G13356;
	G16418<=G5959 and G12084;
	G16419<=G5960 and G12085;
	G16420<=G5961 and G12086;
	G16421<=G5962 and G12087;
	G16422<=G983 and G12088;
	G16423<=G5772 and G13361;
	G16424<=G5967 and G12101;
	G16425<=G5968 and G12102;
	G16426<=G5969 and G12103;
	G16427<=G5970 and G12104;
	G16428<=G1676 and G12105;
	G16429<=G5973 and G12115;
	G16430<=G5974 and G12116;
	G16431<=G5975 and G12117;
	G16432<=G2369 and G12118;
	G16438<=G2594 and G12122;
	G16443<=G5980 and G12134;
	G16444<=G5981 and G12135;
	G16445<=G5808 and G13381;
	G16447<=G5983 and G12147;
	G16448<=G5984 and G12148;
	G16449<=G5985 and G12149;
	G16450<=G5986 and G12150;
	G16451<=G5818 and G13386;
	G16452<=G5988 and G12156;
	G16453<=G5989 and G12157;
	G16454<=G5990 and G12158;
	G16455<=G5991 and G12159;
	G16456<=G1677 and G12160;
	G16457<=G5831 and G13391;
	G16458<=G5996 and G12173;
	G16459<=G5997 and G12174;
	G16460<=G5998 and G12175;
	G16461<=G5999 and G12176;
	G16462<=G2370 and G12177;
	G16505<=G14776 and G14797 and G16142 and G16243;
	G16513<=G15065 and G13724 and G13764 and G13797;
	G16527<=G14811 and G14849 and G16201 and G16302;
	G16535<=G15161 and G13774 and G13805 and G13825;
	G16558<=G14863 and G14922 and G16266 and G16360;
	G16590<=G14936 and G15003 and G16325 and G16404;
	G16607<=G15022 and G15096;
	G16625<=G15118 and G15188;
	G16639<=G15210 and G15274;
	G16650<=G15296 and G15366;
	G16850<=G6226 and G14764;
	G16855<=G15722 and G8646;
	G16856<=G6443 and G14794;
	G16859<=G15762 and G8662;
	G16864<=G15790 and G8681;
	G16865<=G6896 and G14881;
	G16879<=G15813 and G8693;
	G16894<=G7156 and G14959;
	G16907<=G7335 and G15017;
	G16908<=G7838 and G15032;
	G16909<=G6908 and G15033;
	G16923<=G7352 and G15048;
	G16938<=G7858 and G15128;
	G16939<=G7158 and G15129;
	G16953<=G7482 and G15144;
	G16964<=G7520 and G15170;
	G16966<=G7529 and G15174;
	G16967<=G7827 and G15175;
	G16968<=G6672 and G15176;
	G16969<=G7888 and G15220;
	G16970<=G7354 and G15221;
	G16984<=G7538 and G15236;
	G16987<=G7555 and G15260;
	G16988<=G7842 and G15261;
	G16989<=G6974 and G15262;
	G16990<=G7912 and G15306;
	G16991<=G7484 and G15307;
	G16993<=G7576 and G15322;
	G16994<=G7819 and G15323;
	G16997<=G7578 and G15352;
	G16998<=G7862 and G15353;
	G16999<=G7224 and G15354;
	G17001<=G3254 and G10694 and G14144;
	G17015<=G7996 and G15390;
	G17017<=G7590 and G15408;
	G17018<=G7830 and G15409;
	G17021<=G7592 and G15438;
	G17022<=G7892 and G15439;
	G17023<=G7420 and G15440;
	G17028<=G7604 and G15458;
	G17031<=G3410 and G10714 and G14259;
	G17045<=G8071 and G15474;
	G17047<=G7605 and G15492;
	G17048<=G7845 and G15493;
	G17055<=G7153 and G15524;
	G17056<=G7953 and G15525;
	G17062<=G7613 and G15544;
	G17065<=G3566 and G10735 and G14381;
	G17079<=G8156 and G15560;
	G17081<=G7614 and G15578;
	G17082<=G7865 and G15579;
	G17084<=G7629 and G13954;
	G17090<=G7349 and G15602;
	G17091<=G8004 and G15603;
	G17097<=G7622 and G15622;
	G17100<=G3722 and G10754 and G14493;
	G17114<=G8242 and G15638;
	G17116<=G7649 and G14008;
	G17117<=G7906 and G15665;
	G17122<=G7658 and G14024;
	G17128<=G7479 and G15678;
	G17129<=G8079 and G15679;
	G17135<=G7638 and G15698;
	G17138<=G7676 and G14068;
	G17143<=G7685 and G14099;
	G17144<=G7958 and G15724;
	G17149<=G7694 and G14115;
	G17155<=G7535 and G15737;
	G17156<=G8164 and G15738;
	G17161<=G7712 and G14183;
	G17166<=G7721 and G14214;
	G17167<=G8009 and G15764;
	G17172<=G7730 and G14230;
	G17176<=G7742 and G14298;
	G17181<=G7751 and G14329;
	G17182<=G8084 and G15792;
	G17193<=G7766 and G14420;
	G17268<=G8024 and G15991;
	G17301<=G8097 and G15994;
	G17339<=G8176 and G15997;
	G17352<=G3942 and G14960;
	G17353<=G3945 and G14963;
	G17381<=G8250 and G16001;
	G17382<=G8252 and G16002;
	G17393<=G3941 and G16005;
	G17395<=G6177 and G15034;
	G17396<=G4020 and G15037;
	G17397<=G4023 and G15040;
	G17398<=G4026 and G15043;
	G17408<=G4049 and G15049;
	G17409<=G4052 and G15052;
	G17428<=G3994 and G16007;
	G17446<=G6284 and G16011;
	G17447<=G4115 and G15106;
	G17448<=G4118 and G15109;
	G17449<=G4121 and G15112;
	G17450<=G4124 and G15115;
	G17460<=G4048 and G16012;
	G17461<=G6209 and G15130;
	G17462<=G4147 and G15133;
	G17463<=G4150 and G15136;
	G17464<=G4153 and G15139;
	G17474<=G4176 and G15145;
	G17475<=G4179 and G15148;
	G17485<=G4089 and G16013;
	G17486<=G4091 and G16014;
	G17506<=G6675 and G16023;
	G17508<=G4225 and G15179;
	G17509<=G4228 and G15182;
	G17510<=G4231 and G15185;
	G17526<=G6421 and G16025;
	G17527<=G4254 and G15198;
	G17528<=G4257 and G15201;
	G17529<=G4260 and G15204;
	G17530<=G4263 and G15207;
	G17540<=G4175 and G16026;
	G17541<=G6298 and G15222;
	G17542<=G4286 and G15225;
	G17543<=G4289 and G15228;
	G17544<=G4292 and G15231;
	G17554<=G4315 and G15237;
	G17555<=G4318 and G15240;
	G17556<=G4201 and G16027;
	G17576<=G4348 and G15248;
	G17577<=G4351 and G15251;
	G17578<=G4354 and G15254;
	G17597<=G6977 and G16039;
	G17598<=G4380 and G15265;
	G17599<=G4383 and G15268;
	G17600<=G4386 and G15271;
	G17616<=G6626 and G16041;
	G17617<=G4409 and G15284;
	G17618<=G4412 and G15287;
	G17619<=G4415 and G15290;
	G17620<=G4418 and G15293;
	G17630<=G4314 and G16042;
	G17631<=G6435 and G15308;
	G17632<=G4441 and G15311;
	G17633<=G4444 and G15314;
	G17634<=G4447 and G15317;
	G17635<=G4322 and G16043;
	G17636<=G4324 and G16044;
	G17652<=G4480 and G15326;
	G17653<=G4483 and G15329;
	G17654<=G4486 and G15332;
	G17673<=G4517 and G15340;
	G17674<=G4520 and G15343;
	G17675<=G4523 and G15346;
	G17694<=G7227 and G16061;
	G17695<=G4549 and G15357;
	G17696<=G4552 and G15360;
	G17697<=G4555 and G15363;
	G17713<=G6890 and G16063;
	G17714<=G4578 and G15376;
	G17715<=G4581 and G15379;
	G17716<=G4584 and G15382;
	G17717<=G4587 and G15385;
	G17718<=G4451 and G16064;
	G17719<=G2993 and G16065;
	G17734<=G4611 and G15393;
	G17735<=G4614 and G15396;
	G17736<=G4617 and G15399;
	G17737<=G4626 and G15404;
	G17752<=G4656 and G15412;
	G17753<=G4659 and G15415;
	G17754<=G4662 and G15418;
	G17773<=G4693 and G15426;
	G17774<=G4696 and G15429;
	G17775<=G4699 and G15432;
	G17794<=G7423 and G16097;
	G17795<=G4725 and G15443;
	G17796<=G4728 and G15446;
	G17797<=G4731 and G15449;
	G17798<=G4591 and G16099;
	G17812<=G4754 and G15461;
	G17813<=G4757 and G15464;
	G17814<=G4760 and G15467;
	G17824<=G4766 and G15471;
	G17835<=G4788 and G15477;
	G17836<=G4791 and G15480;
	G17837<=G4794 and G15483;
	G17838<=G4803 and G15488;
	G17853<=G4833 and G15496;
	G17854<=G4836 and G15499;
	G17855<=G4839 and G15502;
	G17874<=G4870 and G15510;
	G17875<=G4873 and G15513;
	G17876<=G4876 and G15516;
	G17877<=G2998 and G15521;
	G17900<=G4899 and G15528;
	G17901<=G4902 and G15531;
	G17902<=G4905 and G15534;
	G17912<=G4908 and G15537;
	G17924<=G4930 and G15547;
	G17925<=G4933 and G15550;
	G17926<=G4936 and G15553;
	G17936<=G4942 and G15557;
	G17947<=G4964 and G15563;
	G17948<=G4967 and G15566;
	G17949<=G4970 and G15569;
	G17950<=G4979 and G15574;
	G17965<=G5009 and G15582;
	G17966<=G5012 and G15585;
	G17967<=G5015 and G15588;
	G17989<=G5035 and G15596;
	G17990<=G5038 and G15599;
	G18011<=G5058 and G15606;
	G18012<=G5061 and G15609;
	G18013<=G5064 and G15612;
	G18023<=G5067 and G15615;
	G18035<=G5089 and G15625;
	G18036<=G5092 and G15628;
	G18037<=G5095 and G15631;
	G18047<=G5101 and G15635;
	G18058<=G5123 and G15641;
	G18059<=G5126 and G15644;
	G18060<=G5129 and G15647;
	G18061<=G5138 and G15652;
	G18062<=G7462 and G15655;
	G18088<=G5150 and G15667;
	G18106<=G5164 and G15672;
	G18107<=G5167 and G15675;
	G18128<=G5187 and G15682;
	G18129<=G5190 and G15685;
	G18130<=G5193 and G15688;
	G18140<=G5196 and G15691;
	G18152<=G5218 and G15701;
	G18153<=G5221 and G15704;
	G18154<=G5224 and G15707;
	G18164<=G5230 and G15711;
	G18165<=G2883 and G16287;
	G18169<=G7527 and G15714;
	G18204<=G5243 and G15726;
	G18222<=G5257 and G15731;
	G18223<=G5260 and G15734;
	G18244<=G5280 and G15741;
	G18245<=G5283 and G15744;
	G18246<=G5286 and G15747;
	G18256<=G5289 and G15750;
	G18311<=G5306 and G15766;
	G18329<=G5320 and G15771;
	G18330<=G5323 and G15774;
	G18333<=G2888 and G15777;
	G18404<=G5343 and G15794;
	G18547<=G13677 and G13750 and I24619;
	G18597<=G13714 and G13791 and I24689;
	G18629<=G13764 and G13819 and I24738;
	G18638<=G13805 and G13840 and I24758;
	G18645<=G14776 and G14895 and G16142 and G13750;
	G18647<=G14895 and G16142 and G16243;
	G18648<=G14811 and G14976 and G16201 and G13791;
	G18649<=G14776 and G14837 and G13657 and G16189;
	G18650<=G14976 and G16201 and G16302;
	G18651<=G14863 and G15065 and G16266 and G13819;
	G18652<=G14797 and G13657 and G13677 and G16243;
	G18653<=G14811 and G14910 and G13687 and G16254;
	G18654<=G15065 and G16266 and G16360;
	G18655<=G14936 and G15161 and G16325 and G13840;
	G18665<=G14776 and G14837 and G16189 and G13706;
	G18666<=G14849 and G13687 and G13714 and G16302;
	G18667<=G14863 and G14991 and G13724 and G16313;
	G18668<=G15161 and G16325 and G16404;
	G18688<=G14811 and G14910 and G16254 and G13756;
	G18689<=G14922 and G13724 and G13764 and G16360;
	G18690<=G14936 and G15080 and G13774 and G16371;
	G18717<=G14863 and G14991 and G16313 and G13797;
	G18718<=G15003 and G13774 and G13805 and G16404;
	G18753<=G14936 and G15080 and G16371 and G13825;
	G18982<=G13519 and G16154;
	G18990<=G13530 and G16213;
	G18994<=G14895 and G13657 and G13677 and G13706;
	G18997<=G13541 and G16278;
	G19007<=G14976 and G13687 and G13714 and G13756;
	G19010<=G13552 and G16337;
	G19063<=G18679 and G14910 and G13687 and G16254;
	G19079<=G14797 and G18692 and G16142 and G16189;
	G19080<=G18708 and G14991 and G13724 and G16313;
	G19087<=G17215 and G16540;
	G19088<=G18656 and G14797 and G16189 and G13706;
	G19089<=G14849 and G18728 and G16201 and G16254;
	G19090<=G18744 and G15080 and G13774 and G16371;
	G19092<=G14776 and G18670 and G18692 and G16293;
	G19093<=G17218 and G16572;
	G19094<=G18679 and G14849 and G16254 and G13756;
	G19095<=G14922 and G18765 and G16266 and G16313;
	G19097<=G13657 and G16243 and I25280;
	G19099<=G14811 and G18699 and G18728 and G16351;
	G19100<=G17220 and G16596;
	G19101<=G18708 and G14922 and G16313 and G13797;
	G19102<=G15003 and G18796 and G16325 and G16371;
	G19104<=G13687 and G16302 and I25291;
	G19106<=G14863 and G18735 and G18765 and G16395;
	G19107<=G17223 and G16616;
	G19108<=G18744 and G15003 and G16371 and G13825;
	G19109<=G13724 and G16360 and I25300;
	G19111<=G14936 and G18772 and G18796 and G16433;
	G19112<=G14657 and G16633;
	G19116<=G13774 and G16404 and I25311;
	G19117<=G14691 and G16644;
	G19124<=G14725 and G16656;
	G19131<=G14753 and G16673;
	G19142<=G17159 and G16719;
	G19143<=G17174 and G16761;
	G19146<=G17191 and G16788;
	G19148<=G17202 and G16817;
	G19150<=G17189 and G8602;
	G19155<=G17200 and G8614;
	G19161<=G17207 and G8627;
	G19166<=G17212 and G8637;
	G19228<=G16662 and G12125;
	G19236<=G16935 and G8802;
	G19241<=G16867 and G14158 and G14071;
	G19248<=G16662 and G8817;
	G19252<=G18725 and G9527;
	G19254<=G16895 and G14273 and G14186;
	G19260<=G16749 and G3124;
	G19267<=G16924 and G14395 and G14301;
	G19282<=G16954 and G14507 and G14423;
	G19284<=G18063 and G3111;
	G19285<=G16749 and G7642;
	G19289<=G17029 and G8580;
	G19303<=G16867 and G16543 and G14071;
	G19307<=G17063 and G8587;
	G19316<=G18063 and G3110;
	G19317<=G16749 and G3126;
	G19320<=G16867 and G16515 and G14158;
	G19324<=G16895 and G16575 and G14186;
	G19328<=G17098 and G8594;
	G19347<=G16895 and G16546 and G14273;
	G19351<=G16924 and G16599 and G14301;
	G19355<=G17136 and G8605;
	G19356<=G18063 and G3112;
	G19381<=G16924 and G16578 and G14395;
	G19385<=G16954 and G16619 and G14423;
	G19413<=G16954 and G16602 and G14507;
	G19449<=G16884 and G14797 and G14776;
	G19476<=G16913 and G14849 and G14811;
	G19499<=G16943 and G14922 and G14863;
	G19520<=G16974 and G15003 and G14936;
	G19531<=G16884 and G16722 and G14776;
	G19540<=G16884 and G16697 and G14797;
	G19541<=G16913 and G16764 and G14811;
	G19544<=G16913 and G16728 and G14849;
	G19545<=G16943 and G16791 and G14863;
	G19547<=G16943 and G16770 and G14922;
	G19548<=G16974 and G16820 and G14936;
	G19549<=G7950 and G17230;
	G19551<=G16974 and G16797 and G15003;
	G19552<=G16829 and G6048;
	G19553<=G7990 and G17237;
	G19554<=G7993 and G17240;
	G19555<=G8001 and G17243;
	G19557<=G8053 and G17249;
	G19558<=G8056 and G17252;
	G19559<=G8059 and G17255;
	G19560<=G8065 and G17259;
	G19561<=G8068 and G17262;
	G19562<=G8076 and G17265;
	G19564<=G8123 and G17272;
	G19565<=G8126 and G17275;
	G19566<=G8129 and G17278;
	G19567<=G8138 and G17282;
	G19568<=G8141 and G17285;
	G19569<=G8144 and G17288;
	G19570<=G8150 and G17291;
	G19571<=G8153 and G17294;
	G19572<=G8161 and G17297;
	G19574<=G8191 and G17304;
	G19575<=G8194 and G17307;
	G19576<=G8197 and G17310;
	G19584<=G640 and G18756;
	G19585<=G692 and G18757;
	G19586<=G8209 and G17315;
	G19587<=G8212 and G17318;
	G19588<=G8215 and G17321;
	G19589<=G8224 and G17324;
	G19590<=G8227 and G17327;
	G19591<=G8230 and G17330;
	G19592<=G8236 and G17333;
	G19593<=G8239 and G17336;
	G19594<=G16935 and G12555;
	G19597<=G3922 and G17342;
	G19598<=G3925 and G17345;
	G19599<=G3928 and G17348;
	G19600<=G633 and G18783;
	G19601<=G640 and G18784;
	G19602<=G633 and G18785;
	G19603<=G692 and G18786;
	G19604<=G3948 and G17354;
	G19605<=G3951 and G17357;
	G19606<=G3954 and G17360;
	G19614<=G1326 and G18787;
	G19615<=G1378 and G18788;
	G19616<=G3966 and G17363;
	G19617<=G3969 and G17366;
	G19618<=G3972 and G17369;
	G19619<=G3981 and G17372;
	G19620<=G3984 and G17375;
	G19621<=G3987 and G17378;
	G19623<=G4000 and G17384;
	G19624<=G4003 and G17387;
	G19625<=G4006 and G17390;
	G19626<=G640 and G18805;
	G19627<=G633 and G18806;
	G19628<=G653 and G18807;
	G19629<=G692 and G18808;
	G19630<=G4029 and G17399;
	G19631<=G4032 and G17402;
	G19632<=G4035 and G17405;
	G19633<=G1319 and G18809;
	G19634<=G1326 and G18810;
	G19635<=G1319 and G18811;
	G19636<=G1378 and G18812;
	G19637<=G4055 and G17410;
	G19638<=G4058 and G17413;
	G19639<=G4061 and G17416;
	G19647<=G2020 and G18813;
	G19648<=G2072 and G18814;
	G19649<=G4073 and G17419;
	G19650<=G4076 and G17422;
	G19651<=G4079 and G17425;
	G19653<=G4095 and G17430;
	G19654<=G4098 and G17433;
	G19655<=G4101 and G17436;
	G19656<=G4104 and G17439;
	G19660<=G633 and G18822;
	G19661<=G653 and G18823;
	G19662<=G646 and G18824;
	G19663<=G4127 and G17451;
	G19664<=G4130 and G17454;
	G19665<=G4133 and G17457;
	G19666<=G1326 and G18825;
	G19667<=G1319 and G18826;
	G19668<=G1339 and G18827;
	G19669<=G1378 and G18828;
	G19670<=G4156 and G17465;
	G19671<=G4159 and G17468;
	G19672<=G4162 and G17471;
	G19673<=G2013 and G18829;
	G19674<=G2020 and G18830;
	G19675<=G2013 and G18831;
	G19676<=G2072 and G18832;
	G19677<=G4182 and G17476;
	G19678<=G4185 and G17479;
	G19679<=G4188 and G17482;
	G19687<=G2714 and G18833;
	G19688<=G2766 and G18834;
	G19691<=G16841 and G10865;
	G19692<=G4205 and G17487;
	G19693<=G4208 and G17490;
	G19694<=G4211 and G17493;
	G19695<=G4214 and G17496;
	G19697<=G653 and G18838;
	G19698<=G646 and G18839;
	G19699<=G660 and G18840;
	G19700<=G17815 and G16024;
	G19701<=G4234 and G17511;
	G19702<=G4237 and G17514;
	G19703<=G4240 and G17517;
	G19704<=G4243 and G17520;
	G19708<=G1319 and G18841;
	G19709<=G1339 and G18842;
	G19710<=G1332 and G18843;
	G19711<=G4266 and G17531;
	G19712<=G4269 and G17534;
	G19713<=G4272 and G17537;
	G19714<=G2020 and G18844;
	G19715<=G2013 and G18845;
	G19716<=G2033 and G18846;
	G19717<=G2072 and G18847;
	G19718<=G4295 and G17545;
	G19719<=G4298 and G17548;
	G19720<=G4301 and G17551;
	G19721<=G2707 and G18848;
	G19722<=G2714 and G18849;
	G19723<=G2707 and G18850;
	G19724<=G2766 and G18851;
	G19726<=G16847 and G6131;
	G19727<=G4329 and G17557;
	G19728<=G4332 and G17560;
	G19729<=G4335 and G17563;
	G19730<=G653 and G17573;
	G19731<=G646 and G18853;
	G19732<=G660 and G18854;
	G19733<=G672 and G18855;
	G19734<=G17815 and G16034;
	G19735<=G17903 and G16035;
	G19736<=G4360 and G17579;
	G19737<=G4363 and G17582;
	G19738<=G4366 and G17585;
	G19739<=G4369 and G17588;
	G19741<=G1339 and G18856;
	G19742<=G1332 and G18857;
	G19743<=G1346 and G18858;
	G19744<=G17927 and G16040;
	G19745<=G4389 and G17601;
	G19746<=G4392 and G17604;
	G19747<=G4395 and G17607;
	G19748<=G4398 and G17610;
	G19752<=G2013 and G18859;
	G19753<=G2033 and G18860;
	G19754<=G2026 and G18861;
	G19755<=G4421 and G17621;
	G19756<=G4424 and G17624;
	G19757<=G4427 and G17627;
	G19758<=G2714 and G18862;
	G19759<=G2707 and G18863;
	G19760<=G2727 and G18864;
	G19761<=G2766 and G18865;
	G19764<=G4453 and G17637;
	G19765<=G660 and G18870;
	G19766<=G672 and G18871;
	G19767<=G666 and G18872;
	G19768<=G17815 and G16054;
	G19769<=G17903 and G16055;
	G19770<=G4498 and G17655;
	G19771<=G4501 and G17658;
	G19772<=G4504 and G17661;
	G19773<=G1339 and G17670;
	G19774<=G1332 and G18874;
	G19775<=G1346 and G18875;
	G19776<=G1358 and G18876;
	G19777<=G17927 and G16056;
	G19778<=G18014 and G16057;
	G19779<=G4529 and G17676;
	G19780<=G4532 and G17679;
	G19781<=G4535 and G17682;
	G19782<=G4538 and G17685;
	G19784<=G2033 and G18877;
	G19785<=G2026 and G18878;
	G19786<=G2040 and G18879;
	G19787<=G18038 and G16062;
	G19788<=G4558 and G17698;
	G19789<=G4561 and G17701;
	G19790<=G4564 and G17704;
	G19791<=G4567 and G17707;
	G19795<=G2707 and G18880;
	G19796<=G2727 and G18881;
	G19797<=G2720 and G18882;
	G19799<=G17640 and G18074 and I26240;
	G19802<=G672 and G18891;
	G19803<=G666 and G18892;
	G19804<=G679 and G18893;
	G19805<=G17903 and G16088;
	G19806<=G4629 and G17738;
	G19807<=G1346 and G18896;
	G19808<=G1358 and G18897;
	G19809<=G1352 and G18898;
	G19810<=G17927 and G16090;
	G19811<=G18014 and G16091;
	G19812<=G4674 and G17755;
	G19813<=G4677 and G17758;
	G19814<=G4680 and G17761;
	G19815<=G2033 and G17770;
	G19816<=G2026 and G18900;
	G19817<=G2040 and G18901;
	G19818<=G2052 and G18902;
	G19819<=G18038 and G16092;
	G19820<=G18131 and G16093;
	G19821<=G4705 and G17776;
	G19822<=G4708 and G17779;
	G19823<=G4711 and G17782;
	G19824<=G4714 and G17785;
	G19826<=G2727 and G18903;
	G19827<=G2720 and G18904;
	G19828<=G2734 and G18905;
	G19829<=G18155 and G16098;
	G19836<=G7143 and G18908;
	G19837<=G6901 and G17799;
	G19839<=G666 and G18909;
	G19840<=G679 and G18910;
	G19841<=G686 and G18911;
	G19842<=G14525 and G13922 and I26282;
	G19843<=G17741 and G18190 and I26285;
	G19846<=G1358 and G18914;
	G19847<=G1352 and G18915;
	G19848<=G1365 and G18916;
	G19849<=G18014 and G16126;
	G19850<=G4806 and G17839;
	G19851<=G2040 and G18919;
	G19852<=G2052 and G18920;
	G19853<=G2046 and G18921;
	G19854<=G18038 and G16128;
	G19855<=G18131 and G16129;
	G19856<=G4851 and G17856;
	G19857<=G4854 and G17859;
	G19858<=G4857 and G17862;
	G19859<=G2727 and G17871;
	G19860<=G2720 and G18923;
	G19861<=G2734 and G18924;
	G19862<=G2746 and G18925;
	G19863<=G18155 and G16130;
	G19864<=G18247 and G16131;
	G19868<=G16498 and G16867 and G19001;
	G19869<=G679 and G18926;
	G19870<=G686 and G18927;
	G19871<=G14086 and G18275 and I26311;
	G19872<=G1352 and G18928;
	G19873<=G1365 and G18929;
	G19874<=G1372 and G18930;
	G19875<=G14580 and G13978 and I26317;
	G19876<=G17842 and G18297 and I26320;
	G19879<=G2052 and G18933;
	G19880<=G2046 and G18934;
	G19881<=G2059 and G18935;
	G19882<=G18131 and G16177;
	G19883<=G4982 and G17951;
	G19884<=G2734 and G18938;
	G19885<=G2746 and G18939;
	G19886<=G2740 and G18940;
	G19887<=G18155 and G16179;
	G19888<=G18247 and G16180;
	G19889<=G2912 and G18943;
	G19895<=G686 and G18945;
	G19899<=G16520 and G16895 and G16507;
	G19900<=G1365 and G18946;
	G19901<=G1372 and G18947;
	G19902<=G14201 and G18368 and I26348;
	G19903<=G2046 and G18948;
	G19904<=G2059 and G18949;
	G19905<=G2066 and G18950;
	G19906<=G14614 and G14048 and I26354;
	G19907<=G17954 and G18390 and I26357;
	G19910<=G2746 and G18953;
	G19911<=G2740 and G18954;
	G19912<=G2753 and G18955;
	G19913<=G18247 and G16236;
	G19914<=G3018 and G18958;
	G19920<=G1372 and G18961;
	G19924<=G16551 and G16924 and G16529;
	G19925<=G2059 and G18962;
	G19926<=G2066 and G18963;
	G19927<=G14316 and G18463 and I26377;
	G19928<=G2740 and G18964;
	G19929<=G2753 and G18965;
	G19930<=G2760 and G18966;
	G19931<=G14637 and G14139 and I26383;
	G19932<=G2917 and G18166;
	G19935<=G2066 and G18972;
	G19939<=G16583 and G16954 and G16560;
	G19940<=G2753 and G18973;
	G19941<=G2760 and G18974;
	G19942<=G14438 and G18536 and I26396;
	G19943<=G7562 and G18976;
	G19944<=G3028 and G18258;
	G19949<=G5293 and G18278;
	G19952<=G2760 and G18987;
	G19953<=G7566 and G18334;
	G19970<=G18354 and G18276 and I26416;
	G19971<=G5327 and G18355;
	G19976<=G5330 and G18371;
	G19982<=G17992 and G17913 and I26432;
	G19983<=G5352 and G18432;
	G20000<=G18449 and G18369 and I26440;
	G20001<=G5355 and G18450;
	G20006<=G5358 and G18466;
	G20011<=G18063 and G3113;
	G20012<=G16804 and G3135;
	G20013<=G17720 and G12848;
	G20014<=G7615 and G16749;
	G20020<=G18109 and G18024 and I26464;
	G20021<=G5369 and G18505;
	G20038<=G18522 and G18464 and I26472;
	G20039<=G5372 and G18523;
	G20044<=G5375 and G18539;
	G20048<=G16749 and G3127;
	G20049<=G17878 and G3155;
	G20050<=G18070 and G3161;
	G20051<=G18063 and G3114;
	G20052<=G16804 and G3134;
	G20053<=G17720 and G12875;
	G20062<=G18225 and G18141 and I26500;
	G20063<=G5382 and G18569;
	G20080<=G18586 and G18537 and I26508;
	G20081<=G5385 and G18587;
	G20084<=G17969 and G3158;
	G20085<=G18170 and G3164;
	G20086<=G18337 and G3170;
	G20087<=G16749 and G7574;
	G20088<=G16836 and G3147;
	G20089<=G17969 and G9160;
	G20090<=G18063 and G3120;
	G20091<=G16804 and G3136;
	G20092<=G16749 and G7603;
	G20093<=G13657 and G13677 and G13750 and I26525;
	G20094<=G13677 and G13706 and I26528;
	G20103<=G18332 and G18257 and I26541;
	G20104<=G5391 and G18619;
	G20106<=G18261 and G3167;
	G20107<=G18415 and G3173;
	G20108<=G18543 and G3179;
	G20109<=G17878 and G9504;
	G20110<=G18070 and G9286;
	G20111<=G18261 and G9884;
	G20112<=G16749 and G3132;
	G20113<=G16836 and G3142;
	G20114<=G17969 and G9755;
	G20115<=G16804 and G3139;
	G20116<=G16142 and G13677 and G13706 and I26558;
	G20117<=G16189 and G13706 and I26561;
	G20118<=G13687 and G13714 and G13791 and I26564;
	G20119<=G13714 and G13756 and I26567;
	G20131<=G18486 and G3176;
	G20132<=G18593 and G3182;
	G20133<=G18170 and G9505;
	G20134<=G18337 and G9506;
	G20135<=G18486 and G9885;
	G20136<=G17878 and G9423;
	G20137<=G18070 and G9226;
	G20138<=G18261 and G9756;
	G20139<=G16836 and G3151;
	G20144<=G16679 and G16884 and G16665;
	G20145<=G14776 and G18670 and G16142 and G16189;
	G20146<=G16201 and G13714 and G13756 and I26590;
	G20147<=G16254 and G13756 and I26593;
	G20148<=G13724 and G13764 and G13819 and I26596;
	G20149<=G13764 and G13797 and I26599;
	G20156<=G16809 and G3185;
	G20157<=G18415 and G9287;
	G20158<=G18543 and G9886;
	G20159<=G16809 and G9288;
	G20160<=G18170 and G9424;
	G20161<=G18337 and G9426;
	G20162<=G18486 and G9757;
	G20177<=G13677 and G13750 and I26615;
	G20182<=G16705 and G16913 and G16686;
	G20183<=G14811 and G18699 and G16201 and G16254;
	G20184<=G16266 and G13764 and G13797 and I26621;
	G20185<=G16313 and G13797 and I26624;
	G20186<=G13774 and G13805 and G13840 and I26627;
	G20187<=G13805 and G13825 and I26630;
	G20188<=G18593 and G9425;
	G20189<=G16825 and G9289;
	G20190<=G18415 and G9227;
	G20191<=G18543 and G9758;
	G20192<=G16809 and G9228;
	G20197<=G13677 and G13706 and I26639;
	G20211<=G13714 and G13791 and I26645;
	G20216<=G16736 and G16943 and G16712;
	G20217<=G14863 and G18735 and G16266 and G16313;
	G20218<=G16325 and G13805 and G13825 and I26651;
	G20219<=G16371 and G13825 and I26654;
	G20220<=G18593 and G9355;
	G20221<=G16825 and G10099;
	G20222<=G18656 and G18720 and G13657 and G16293;
	G20227<=G13714 and G13756 and I26661;
	G20241<=G13764 and G13819 and I26667;
	G20246<=G16778 and G16974 and G16743;
	G20247<=G14936 and G18772 and G16325 and G16371;
	G20248<=G18656 and G14837 and G16293;
	G20249<=G18679 and G18758 and G13687 and G16351;
	G20254<=G13764 and G13797 and I26676;
	G20268<=G13805 and G13840 and I26682;
	G20270<=G14797 and G18692 and G13657 and G16243;
	G20271<=G18679 and G14910 and G16351;
	G20272<=G18708 and G18789 and G13724 and G16395;
	G20277<=G13805 and G13825 and I26690;
	G20280<=G13677 and G16243 and I26695;
	G20282<=G14849 and G18728 and G13687 and G16302;
	G20283<=G18708 and G14991 and G16395;
	G20284<=G18744 and G18815 and G13774 and G16433;
	G20285<=G16846 and G8103;
	G20291<=G13714 and G16302 and I26708;
	G20293<=G14922 and G18765 and G13724 and G16360;
	G20294<=G18744 and G15080 and G16433;
	G20307<=G13764 and G16360 and I26726;
	G20309<=G15003 and G18796 and G13774 and G16404;
	G20326<=G13805 and G16404 and I26745;
	G20460<=G17351 and G13644;
	G20472<=G17314 and G13669;
	G20480<=G17313 and G11827;
	G20486<=G17281 and G11859;
	G20492<=G17258 and G11894;
	G20499<=G17648 and G11933;
	G20502<=G17566 and G11973;
	G20503<=G17507 and G13817;
	G20506<=G17499 and G12025;
	G20512<=G17445 and G13836;
	G20525<=G17394 and G13849;
	G20538<=G18656 and G14837 and G13657 and G16189;
	G20640<=G4809 and G19064;
	G20647<=G5888 and G19075;
	G20665<=G4985 and G19081;
	G20809<=G5712 and G19113;
	G20826<=G5770 and G19118;
	G20836<=G5829 and G19125;
	G20840<=G5885 and G19132;
	G21049<=G20016 and G14079 and G14165;
	G21067<=G20193 and G12030;
	G21068<=G20058 and G14194 and G14280;
	G21077<=G20223 and G12094;
	G21078<=G20099 and G14309 and G14402;
	G21085<=G19484 and G14158 and G19001;
	G21086<=G20193 and G12142;
	G21091<=G20250 and G12166;
	G21092<=G20124 and G14431 and G14514;
	G21097<=G19505 and G14273 and G16507;
	G21098<=G20223 and G12204;
	G21103<=G20273 and G12228;
	G21107<=G19444 and G17893 and G14079;
	G21111<=G19524 and G14395 and G16529;
	G21112<=G20250 and G12259;
	G21121<=G20054 and G14244;
	G21122<=G20140 and G12279;
	G21123<=G19970 and G19982;
	G21124<=G19471 and G18004 and G14194;
	G21128<=G19534 and G14507 and G16560;
	G21129<=G20273 and G12302;
	G21136<=G19271 and G19261 and I27695;
	G21137<=G5750 and G19272;
	G21138<=G19484 and G14347;
	G21140<=G20095 and G14366;
	G21141<=G20178 and G12315;
	G21142<=G20000 and G20020;
	G21143<=G19494 and G18121 and G14309;
	G21152<=G19357 and G19334 and I27711;
	G21153<=G20054 and G16543 and G16501;
	G21154<=G20193 and G12333;
	G21155<=G20140 and G12336;
	G21156<=G19290 and G19276 and I27717;
	G21157<=G5809 and G19291;
	G21158<=G19505 and G14459;
	G21160<=G20120 and G14478;
	G21161<=G20212 and G12343;
	G21162<=G20038 and G20062;
	G21163<=G19515 and G18237 and G14431;
	G21172<=G19389 and G19368 and I27733;
	G21173<=G20095 and G16575 and G16523;
	G21174<=G20223 and G12363;
	G21175<=G20178 and G12366;
	G21176<=G19308 and G19295 and I27739;
	G21177<=G5865 and G19309;
	G21178<=G19524 and G14546;
	G21180<=G20150 and G14565;
	G21181<=G20242 and G12373;
	G21182<=G20080 and G20103;
	G21188<=G20140 and G12379;
	G21192<=G19419 and G19400 and I27755;
	G21193<=G20120 and G16599 and G16554;
	G21194<=G20250 and G12382;
	G21195<=G20212 and G12385;
	G21196<=G19329 and G19313 and I27761;
	G21197<=G5912 and G19330;
	G21198<=G19534 and G14601;
	G21203<=G20178 and G12409;
	G21207<=G19456 and G19430 and I27772;
	G21208<=G20150 and G16619 and G16586;
	G21209<=G20273 and G12412;
	G21210<=G20242 and G12415;
	G21218<=G20212 and G12421;
	G21226<=G20242 and G12426;
	G21229<=G19578 and G14797 and G16665;
	G21234<=G19608 and G14849 and G16686;
	G21243<=G19641 and G14922 and G16712;
	G21245<=G20299 and G14837;
	G21251<=G19681 and G15003 and G16743;
	G21252<=G19578 and G14895;
	G21254<=G20318 and G14910;
	G21259<=G20299 and G16722 and G16682;
	G21260<=G19608 and G14976;
	G21262<=G20337 and G14991;
	G21267<=G20318 and G16764 and G16708;
	G21268<=G19641 and G15065;
	G21270<=G20357 and G15080;
	G21276<=G20337 and G16791 and G16739;
	G21277<=G19681 and G15161;
	G21283<=G20357 and G16820 and G16781;
	G21284<=G9356 and G20269;
	G21290<=G9356 and G20278;
	G21291<=G9293 and G20279;
	G21292<=G9453 and G20281;
	G21298<=G9356 and G20286;
	G21299<=G9293 and G20287;
	G21300<=G9232 and G20288;
	G21301<=G9453 and G20289;
	G21302<=G9374 and G20290;
	G21303<=G9595 and G20292;
	G21304<=G9293 and G20296;
	G21305<=G9232 and G20297;
	G21306<=G9187 and G20298;
	G21307<=G9453 and G20302;
	G21308<=G9374 and G20303;
	G21309<=G9310 and G20304;
	G21310<=G9595 and G20305;
	G21311<=G9471 and G20306;
	G21312<=G9737 and G20308;
	G21313<=G9232 and G20311;
	G21314<=G9187 and G20312;
	G21315<=G9161 and G20313;
	G21319<=G9374 and G20315;
	G21320<=G9310 and G20316;
	G21321<=G9248 and G20317;
	G21322<=G9595 and G20321;
	G21323<=G9471 and G20322;
	G21324<=G9391 and G20323;
	G21325<=G9737 and G20324;
	G21326<=G9613 and G20325;
	G21328<=G9187 and G20327;
	G21329<=G9161 and G20328;
	G21330<=G9150 and G20329;
	G21334<=G9310 and G20330;
	G21335<=G9248 and G20331;
	G21336<=G9203 and G20332;
	G21337<=G9471 and G20334;
	G21338<=G9391 and G20335;
	G21339<=G9326 and G20336;
	G21340<=G9737 and G20340;
	G21341<=G9613 and G20341;
	G21342<=G9488 and G20342;
	G21343<=G9161 and G20344;
	G21344<=G9150 and G20345;
	G21345<=G15096 and G20346;
	G21349<=G9248 and G20347;
	G21350<=G9203 and G20348;
	G21351<=G9174 and G20349;
	G21352<=G9391 and G20350;
	G21353<=G9326 and G20351;
	G21354<=G9264 and G20352;
	G21355<=G9613 and G20354;
	G21356<=G9488 and G20355;
	G21357<=G9407 and G20356;
	G21360<=G9507 and G20361;
	G21361<=G9150 and G20362;
	G21362<=G15096 and G20363;
	G21363<=G15022 and G20364;
	G21367<=G9203 and G20366;
	G21368<=G9174 and G20367;
	G21369<=G15188 and G20368;
	G21370<=G9326 and G20369;
	G21371<=G9264 and G20370;
	G21372<=G9216 and G20371;
	G21373<=G9488 and G20372;
	G21374<=G9407 and G20373;
	G21375<=G9342 and G20374;
	G21378<=G9507 and G20378;
	G21379<=G9427 and G20379;
	G21380<=G15096 and G20380;
	G21381<=G15022 and G20381;
	G21388<=G6201 and G19657;
	G21389<=G9649 and G20384;
	G21390<=G9174 and G20385;
	G21391<=G15188 and G20386;
	G21392<=G15118 and G20387;
	G21393<=G9264 and G20389;
	G21394<=G9216 and G20390;
	G21395<=G15274 and G20391;
	G21396<=G9407 and G20392;
	G21397<=G9342 and G20393;
	G21398<=G9277 and G20394;
	G21401<=G9507 and G20397;
	G21402<=G9427 and G20398;
	G21403<=G15022 and G20399;
	G21410<=G6363 and G20402;
	G21411<=G9649 and G20403;
	G21412<=G9569 and G20404;
	G21413<=G15188 and G20405;
	G21414<=G15118 and G20406;
	G21418<=G6290 and G19705;
	G21419<=G9795 and G20409;
	G21420<=G9216 and G20410;
	G21421<=G15274 and G20411;
	G21422<=G15210 and G20412;
	G21423<=G9342 and G20414;
	G21424<=G9277 and G20415;
	G21425<=G15366 and G20416;
	G21428<=G9427 and G20420;
	G21438<=G9649 and G20422;
	G21439<=G9569 and G20423;
	G21440<=G15118 and G20424;
	G21444<=G6568 and G20427;
	G21445<=G9795 and G20428;
	G21446<=G9711 and G20429;
	G21447<=G15274 and G20430;
	G21448<=G15210 and G20431;
	G21452<=G6427 and G19749;
	G21453<=G9941 and G20434;
	G21454<=G9277 and G20435;
	G21455<=G15366 and G20436;
	G21456<=G15296 and G20437;
	G21476<=G9569 and G20442;
	G21480<=G9795 and G20444;
	G21481<=G9711 and G20445;
	G21482<=G15210 and G20446;
	G21486<=G6832 and G20449;
	G21487<=G9941 and G20450;
	G21488<=G9857 and G20451;
	G21489<=G15366 and G20452;
	G21490<=G15296 and G20453;
	G21494<=G6632 and G19792;
	G21497<=G3006 and G20456;
	G21517<=G9711 and G20461;
	G21521<=G9941 and G20463;
	G21522<=G9857 and G20464;
	G21523<=G15296 and G20465;
	G21527<=G7134 and G20468;
	G21533<=G17724 and G18179 and G19799 and I28068;
	G21553<=G9857 and G20476;
	G21564<=G13886 and G14153 and G19799 and I28096;
	G21569<=G17825 and G18286 and G19843 and I28103;
	G21589<=G3002 and G19890;
	G21593<=G16498 and G19484 and G14071;
	G21597<=G13927 and G14268 and G19843 and I28126;
	G21602<=G17937 and G18379 and G19876 and I28133;
	G21610<=G7522 and G20490;
	G21611<=G7471 and G19915;
	G21622<=G16520 and G19505 and G14186;
	G21626<=G13983 and G14390 and G19876 and I28155;
	G21631<=G18048 and G18474 and G19907 and I28162;
	G21635<=G7549 and G20496;
	G21639<=G3398 and G20500;
	G21650<=G16551 and G19524 and G14301;
	G21654<=G14053 and G14502 and G19907 and I28181;
	G21658<=G2896 and G20501;
	G21666<=G3398 and G20504;
	G21670<=G3554 and G20505;
	G21681<=G16583 and G19534 and G14423;
	G21687<=G3398 and G20516;
	G21695<=G3554 and G20517;
	G21699<=G3710 and G20518;
	G21707<=G2892 and G19978;
	G21723<=G3554 and G20534;
	G21731<=G3710 and G20535;
	G21735<=G3866 and G20536;
	G21749<=G3710 and G20553;
	G21757<=G3866 and G20554;
	G21758<=G7607 and G20045;
	G21773<=G3866 and G19078;
	G21805<=G16679 and G19578 and G14776;
	G21812<=G16705 and G19608 and G14811;
	G21818<=G16736 and G19641 and G14863;
	G21822<=G16778 and G19681 and G14936;
	G21891<=G19302 and G11749;
	G21892<=G19288 and G13011;
	G21899<=G19323 and G11749;
	G21900<=G19306 and G13011;
	G21906<=G5715 and G20513;
	G21911<=G19350 and G11749;
	G21912<=G19327 and G13011;
	G21913<=G4456 and G20519;
	G21920<=G5773 and G20531;
	G21925<=G19384 and G11749;
	G21926<=G19354 and G13011;
	G21931<=G4632 and G20539;
	G21938<=G5832 and G20550;
	G21990<=G291 and G21187;
	G22004<=G978 and G21202;
	G22015<=G1672 and G21217;
	G22020<=G2366 and G21225;
	G22036<=G21104 and G21095 and G21084 and I28582;
	G22046<=G21117 and G21105 and G21096 and I28594;
	G22062<=G21135 and G21118 and G21106 and I28609;
	G22187<=G21564 and G20986;
	G22196<=G21597 and G21012;
	G22201<=G21271 and G16881;
	G22202<=G21626 and G21036;
	G22206<=G21895 and G11976;
	G22207<=G21278 and G16910;
	G22208<=G21654 and G21057;
	G22211<=G21661 and G12027;
	G22214<=G21907 and G12045;
	G22215<=G21285 and G16940;
	G22220<=G21690 and G12091;
	G22223<=G21921 and G12109;
	G22224<=G21293 and G16971;
	G22228<=G21716 and G12136;
	G22229<=G21661 and G12139;
	G22235<=G21726 and G12163;
	G22238<=G21939 and G12181;
	G22244<=G21742 and G12198;
	G22245<=G21690 and G12201;
	G22250<=G21752 and G12225;
	G22254<=G21716 and G12239;
	G22255<=G21661 and G12242;
	G22264<=G21766 and G12253;
	G22265<=G21726 and G12256;
	G22270<=G92 and G21529;
	G22272<=G21742 and G12282;
	G22273<=G21690 and G12285;
	G22281<=G21782 and G12296;
	G22282<=G21752 and G12299;
	G22285<=G21716 and G12312;
	G22289<=G780 and G21565;
	G22291<=G21766 and G12318;
	G22292<=G21726 and G12321;
	G22305<=G21742 and G12340;
	G22309<=G1466 and G21598;
	G22311<=G21782 and G12346;
	G22312<=G21752 and G12349;
	G22333<=G21766 and G12370;
	G22337<=G2160 and G21627;
	G22340<=G88 and G21184;
	G22358<=G21782 and G12389;
	G22363<=G776 and G21199;
	G22383<=G1462 and G21214;
	G22398<=G2156 and G21222;
	G22483<=G646 and G21861;
	G22515<=G13873 and G21382;
	G22516<=G20885 and G17442;
	G22517<=G21895 and G12608;
	G22526<=G1332 and G21867;
	G22546<=G13886 and G21404;
	G22555<=G13895 and G21415;
	G22556<=G20904 and G17523;
	G22557<=G21907 and G12654;
	G22566<=G2026 and G21872;
	G22577<=G13907 and G21429;
	G22581<=G21895 and G12699;
	G22587<=G13927 and G21441;
	G22595<=G13936 and G21449;
	G22596<=G20928 and G17613;
	G22597<=G21921 and G12708;
	G22606<=G2720 and G21876;
	G22607<=G13946 and G21458;
	G22610<=G660 and G21473;
	G22614<=G13963 and G21477;
	G22618<=G21907 and G12756;
	G22624<=G13983 and G21483;
	G22632<=G13992 and G21491;
	G22633<=G20956 and G17710;
	G22634<=G21939 and G12765;
	G22637<=G20841 and G10927;
	G22638<=G14001 and G21498;
	G22643<=G14016 and G21505;
	G22646<=G1346 and G21514;
	G22650<=G14033 and G21518;
	G22654<=G21921 and G12798;
	G22660<=G14053 and G21524;
	G22665<=G20920 and G6153;
	G22666<=G21825 and G20014;
	G22667<=G14062 and G21530;
	G22674<=G14092 and G21537;
	G22679<=G14107 and G21541;
	G22682<=G2040 and G21550;
	G22686<=G14124 and G21554;
	G22690<=G21939 and G12837;
	G22699<=G7338 and G21883;
	G22700<=G7146 and G21558;
	G22701<=G18174 and G21561;
	G22707<=G14177 and G21566;
	G22714<=G14207 and G21573;
	G22719<=G14222 and G21577;
	G22722<=G2734 and G21586;
	G22726<=G3036 and G21886;
	G22727<=G14238 and G21590;
	G22732<=G18281 and G21594;
	G22738<=G14292 and G21599;
	G22745<=G14322 and G21606;
	G22754<=G14342 and G21612;
	G22759<=G14360 and G21619;
	G22764<=G18374 and G21623;
	G22770<=G14414 and G21628;
	G22788<=G14454 and G21640;
	G22793<=G14472 and G21647;
	G22798<=G18469 and G21651;
	G22804<=G2920 and G21655;
	G22830<=G14541 and G21671;
	G22835<=G14559 and G21678;
	G22841<=G7583 and G21902;
	G22842<=G3032 and G21682;
	G22869<=G14596 and G21700;
	G22874<=G7587 and G21708;
	G22906<=G2924 and G21927;
	G22984<=G16840 and G21400;
	G23104<=G20842 and G15859;
	G23106<=G5857 and G21050;
	G23118<=G20850 and G15890;
	G23119<=G5904 and G21069;
	G23127<=G20858 and G15923;
	G23128<=G5943 and G21079;
	G23138<=G20866 and G15952;
	G23139<=G5977 and G21093;
	G23409<=G21533 and G22408;
	G23414<=G21569 and G22421;
	G23419<=G22755 and G19577;
	G23423<=G21602 and G22443;
	G23428<=G22789 and G19607;
	G23432<=G21631 and G22476;
	G23434<=G22831 and G19640;
	G23440<=G22870 and G19680;
	G23451<=G18552 and G22547;
	G23458<=G18602 and G22588;
	G23462<=G17988 and G22609;
	G23467<=G18634 and G22625;
	G23471<=G18105 and G22645;
	G23476<=G18643 and G22661;
	G23483<=G22945 and G8847;
	G23484<=G18221 and G22681;
	G23494<=G18328 and G22721;
	G23496<=G5802 and G22300;
	G23510<=G5890 and G22753;
	G23512<=G5858 and G22328;
	G23525<=G5929 and G22787;
	G23527<=G5905 and G22353;
	G23536<=G5963 and G22829;
	G23538<=G5944 and G22376;
	G23544<=G5992 and G22868;
	G23547<=G8062 and G22405;
	G23550<=G8132 and G22409;
	G23551<=G8135 and G22412;
	G23552<=G6136 and G22415;
	G23554<=G8147 and G22418;
	G23558<=G8200 and G22422;
	G23559<=G8203 and G22425;
	G23560<=G8206 and G22428;
	G23563<=G8218 and G22431;
	G23564<=G8221 and G22434;
	G23565<=G6146 and G22437;
	G23567<=G8233 and G22440;
	G23571<=G3931 and G22445;
	G23572<=G3934 and G22448;
	G23573<=G3937 and G22451;
	G23577<=G3957 and G22455;
	G23578<=G3960 and G22458;
	G23579<=G3963 and G22461;
	G23582<=G3975 and G22464;
	G23583<=G3978 and G22467;
	G23584<=G6167 and G22470;
	G23586<=G3990 and G22473;
	G23590<=G4009 and G22477;
	G23591<=G4012 and G22480;
	G23592<=G17640 and G22986;
	G23593<=G22845 and G20365;
	G23598<=G4038 and G22484;
	G23599<=G4041 and G22487;
	G23600<=G4044 and G22490;
	G23604<=G4064 and G22494;
	G23605<=G4067 and G22497;
	G23606<=G4070 and G22500;
	G23609<=G4082 and G22503;
	G23610<=G4085 and G22506;
	G23611<=G6194 and G22509;
	G23615<=G4107 and G22512;
	G23616<=G17724 and G22988;
	G23617<=G22810 and G20382;
	G23618<=G22608 and G20383;
	G23622<=G4136 and G22520;
	G23623<=G4139 and G22523;
	G23624<=G17741 and G22989;
	G23625<=G22880 and G20388;
	G23630<=G4165 and G22527;
	G23631<=G4168 and G22530;
	G23632<=G4171 and G22533;
	G23636<=G4191 and G22537;
	G23637<=G4194 and G22540;
	G23638<=G4197 and G22543;
	G23639<=G21825 and G22805;
	G23643<=G17802 and G22991;
	G23659<=G22784 and G17500;
	G23664<=G4246 and G22552;
	G23665<=G17825 and G22995;
	G23666<=G22851 and G20407;
	G23667<=G22644 and G20408;
	G23671<=G4275 and G22560;
	G23672<=G4278 and G22563;
	G23673<=G17842 and G22996;
	G23674<=G22915 and G20413;
	G23679<=G4304 and G22567;
	G23680<=G4307 and G22570;
	G23681<=G4310 and G22573;
	G23686<=G17882 and G22998;
	G23687<=G22668 and G17570;
	G23689<=G6513 and G23001;
	G23693<=G17914 and G23002;
	G23709<=G22826 and G17591;
	G23714<=G4401 and G22592;
	G23715<=G17937 and G23006;
	G23716<=G22886 and G20432;
	G23717<=G22680 and G20433;
	G23721<=G4430 and G22600;
	G23722<=G4433 and G22603;
	G23723<=G17954 and G23007;
	G23724<=G22940 and G20438;
	G23726<=G21825 and G22843;
	G23734<=G17974 and G23008;
	G23735<=G22949 and G9450;
	G23740<=G17993 and G23012;
	G23741<=G22708 and G17667;
	G23743<=G6777 and G23015;
	G23747<=G18025 and G23016;
	G23763<=G22865 and G17688;
	G23768<=G4570 and G22629;
	G23769<=G18048 and G23020;
	G23770<=G22921 and G20454;
	G23771<=G22720 and G20455;
	G23772<=G21825 and G22875;
	G23776<=G18074 and G23021;
	G23777<=G22949 and G9528;
	G23778<=G22954 and G9531;
	G23789<=G18091 and G23024;
	G23790<=G22958 and G9592;
	G23795<=G18110 and G23028;
	G23796<=G22739 and G17767;
	G23798<=G7079 and G23031;
	G23802<=G18142 and G23032;
	G23818<=G22900 and G17788;
	G23820<=G3013 and G23036;
	G23822<=G14148 and G23037;
	G23824<=G22949 and G9641;
	G23825<=G22954 and G9644;
	G23829<=G18190 and G23038;
	G23830<=G22958 and G9670;
	G23831<=G22962 and G9673;
	G23842<=G18207 and G23041;
	G23843<=G22966 and G9734;
	G23848<=G18226 and G23045;
	G23849<=G22771 and G17868;
	G23851<=G7329 and G23048;
	G23852<=G19179 and G22696;
	G23854<=G18265 and G23049;
	G23855<=G22954 and G9767;
	G23857<=G14263 and G23056;
	G23859<=G22958 and G9787;
	G23860<=G22962 and G9790;
	G23864<=G18297 and G23057;
	G23865<=G22966 and G9816;
	G23866<=G22971 and G9819;
	G23877<=G18314 and G23060;
	G23878<=G22975 and G9880;
	G23886<=G18341 and G23064;
	G23888<=G18358 and G23069;
	G23889<=G22962 and G9913;
	G23891<=G14385 and G23074;
	G23893<=G22966 and G9933;
	G23894<=G22971 and G9936;
	G23898<=G18390 and G23075;
	G23899<=G22975 and G9962;
	G23900<=G22980 and G9965;
	G23904<=G3010 and G22750;
	G23907<=G18436 and G23079;
	G23909<=G18453 and G23082;
	G23910<=G22971 and G10067;
	G23912<=G14497 and G23087;
	G23914<=G22975 and G10087;
	G23915<=G22980 and G10090;
	G23917<=G7545 and G23088;
	G23939<=G18509 and G23095;
	G23941<=G18526 and G23098;
	G23942<=G22980 and G10176;
	G23944<=G7570 and G23103;
	G23971<=G18573 and G23112;
	G23972<=G2903 and G23115;
	G24029<=G2900 and G22903;
	G24211<=G22014 and G10969;
	G24217<=G22825 and G10999;
	G24221<=G22979 and G11042;
	G24224<=G22219 and G11045;
	G24229<=G22232 and G11105;
	G24236<=G22243 and G11157;
	G24241<=G22259 and G11228;
	G24246<=G21982 and G11291;
	G24247<=G22551 and G11297;
	G24253<=G21995 and G11370;
	G24256<=G22003 and G11438;
	G24427<=G17086 and G24134 and G13626;
	G24429<=G24115 and G13614;
	G24431<=G17124 and G24153 and G13637;
	G24432<=G14642 and G15904 and G24115;
	G24433<=G24134 and G13626;
	G24435<=G17151 and G24168 and G13649;
	G24436<=G14669 and G15933 and G24134;
	G24437<=G24153 and G13637;
	G24439<=G14703 and G15962 and G24153;
	G24440<=G24168 and G13649;
	G24441<=G14737 and G15981 and G24168;
	G24478<=G23545 and G21119 and G21227;
	G24529<=G19933 and G17896 and G23403;
	G24540<=G18548 and G23089 and G23403;
	G24541<=G23420 and G17896 and G23052;
	G24542<=G19950 and G18007 and G23410;
	G24550<=G18548 and G23420 and G19948;
	G24552<=G18598 and G23107 and G23410;
	G24553<=G23429 and G18007 and G23071;
	G24554<=G19977 and G18124 and G23415;
	G24559<=G79 and G23448;
	G24561<=G18598 and G23429 and G19975;
	G24563<=G18630 and G23120 and G23415;
	G24564<=G23435 and G18124 and G23084;
	G24565<=G20007 and G18240 and G23424;
	G24569<=G767 and G23455;
	G24571<=G18630 and G23435 and G20005;
	G24573<=G18639 and G23129 and G23424;
	G24574<=G23441 and G18240 and G23100;
	G24578<=G1453 and G23464;
	G24580<=G18639 and G23441 and G20043;
	G24585<=G2147 and G23473;
	G24590<=G23486 and G23478;
	G24591<=G83 and G23853;
	G24595<=G23502 and G23489;
	G24596<=G771 and G23887;
	G24603<=G23518 and G23505;
	G24604<=G1457 and G23908;
	G24610<=G23533 and G23521;
	G24611<=G2151 and G23940;
	G24644<=G17203 and G24115;
	G24664<=G17208 and G24134;
	G24676<=G13568 and G24115;
	G24683<=G17214 and G24153;
	G24695<=G13576 and G24134;
	G24700<=G17217 and G24168;
	G24712<=G13585 and G24153;
	G24723<=G13605 and G24168;
	G24745<=G15454 and G24096;
	G24746<=G15454 and G24098;
	G24747<=G9427 and G24099;
	G24748<=G672 and G24101;
	G24749<=G15540 and G24102;
	G24750<=G15454 and G24104;
	G24751<=G9427 and G24105;
	G24752<=G9507 and G24106;
	G24754<=G15540 and G24107;
	G24755<=G9569 and G24108;
	G24757<=G1358 and G24110;
	G24758<=G15618 and G24111;
	G24759<=G21825 and G23885;
	G24760<=G9427 and G24112;
	G24761<=G9507 and G24113;
	G24762<=G12876 and G24114;
	G24767<=G15540 and G24121;
	G24768<=G9569 and G24122;
	G24769<=G9649 and G24123;
	G24772<=G15618 and G24124;
	G24773<=G9711 and G24125;
	G24774<=G2052 and G24127;
	G24775<=G15694 and G24128;
	G24776<=G9507 and G24129;
	G24777<=G12876 and G24130;
	G24779<=G9569 and G24131;
	G24780<=G9649 and G24132;
	G24781<=G12916 and G24133;
	G24788<=G15618 and G24140;
	G24789<=G9711 and G24141;
	G24790<=G9795 and G24142;
	G24792<=G15694 and G24143;
	G24793<=G9857 and G24144;
	G24794<=G2746 and G24146;
	G24795<=G12017 and G24232;
	G24796<=G12876 and G24147;
	G24798<=G9649 and G24148;
	G24799<=G12916 and G24149;
	G24802<=G9711 and G24150;
	G24803<=G9795 and G24151;
	G24804<=G12945 and G24152;
	G24809<=G15694 and G24159;
	G24810<=G9857 and G24160;
	G24811<=G9941 and G24161;
	G24813<=G21825 and G23905;
	G24818<=G12916 and G24162;
	G24821<=G9795 and G24163;
	G24822<=G12945 and G24164;
	G24824<=G9857 and G24165;
	G24825<=G9941 and G24166;
	G24826<=G12974 and G24167;
	G24831<=G24100 and G20401;
	G24838<=G12945 and G24175;
	G24840<=G9941 and G24176;
	G24841<=G12974 and G24177;
	G24843<=G21825 and G23918;
	G24846<=G24109 and G20426;
	G24853<=G12974 and G24180;
	G24855<=G18174 and G23731;
	G24858<=G24047 and G18873;
	G24861<=G24126 and G20448;
	G24867<=G666 and G23779;
	G24869<=G24047 and G18894;
	G24870<=G18281 and G23786;
	G24874<=G24060 and G18899;
	G24876<=G24145 and G20467;
	G24878<=G19830 and G24210;
	G24881<=G24047 and G18912;
	G24882<=G1352 and G23832;
	G24884<=G24060 and G18917;
	G24885<=G18374 and G23839;
	G24888<=G24073 and G18922;
	G24898<=G24060 and G18931;
	G24899<=G2046 and G23867;
	G24901<=G24073 and G18936;
	G24902<=G18469 and G23874;
	G24905<=G24084 and G18941;
	G24906<=G18886 and G23879;
	G24907<=G7466 and G24220;
	G24908<=G7342 and G23882;
	G24921<=G24073 and G18951;
	G24922<=G2740 and G23901;
	G24924<=G24084 and G18956;
	G24938<=G24084 and G18967;
	G24964<=G7595 and G24251;
	G24974<=G7600 and G24030;
	G25086<=G23444 and G10880;
	G25102<=G23444 and G10915;
	G25117<=G23444 and G10974;
	G25128<=G17051 and G24115 and G13614;
	G25178<=G24623 and G20634;
	G25181<=G24636 and G20673;
	G25182<=G24681 and G20676;
	G25184<=G24694 and G20735;
	G25187<=G24633 and G16608;
	G25188<=G24652 and G20763;
	G25192<=G24711 and G20790;
	G25193<=G24653 and G16626;
	G25196<=G24672 and G16640;
	G25198<=G24691 and G16651;
	G25269<=G24648 and G8700;
	G25277<=G24648 and G8714;
	G25278<=G24668 and G8719;
	G25281<=G5606 and G24815;
	G25282<=G24648 and G8748;
	G25286<=G24668 and G8752;
	G25287<=G24687 and G8757;
	G25289<=G5631 and G24834;
	G25290<=G24668 and G8771;
	G25294<=G24687 and G8775;
	G25295<=G24704 and G8780;
	G25299<=G5659 and G24850;
	G25300<=G24687 and G8794;
	G25304<=G24704 and G8798;
	G25309<=G5697 and G24864;
	G25310<=G24704 and G8813;
	G25318<=G24682 and G19358 and G19335;
	G25321<=G25075 and G9669;
	G25328<=G24644 and G17892;
	G25334<=G24644 and G17984;
	G25337<=G24664 and G18003;
	G25342<=G5851 and G24600;
	G25346<=G24644 and G18084;
	G25348<=G24664 and G18101;
	G25351<=G24683 and G18120;
	G25356<=G5898 and G24607;
	G25360<=G24664 and G18200;
	G25362<=G24683 and G18217;
	G25365<=G24700 and G18236;
	G25371<=G5937 and G24619;
	G25375<=G24683 and G18307;
	G25377<=G24700 and G18324;
	G25388<=G5971 and G24630;
	G25392<=G24700 and G18400;
	G25453<=G6142 and G24763;
	G25457<=G6163 and G24784;
	G25461<=G6190 and G24805;
	G25466<=G6222 and G24827;
	G25470<=G24479 and G20400;
	G25475<=G14148 and G25087;
	G25482<=G24480 and G17567;
	G25483<=G24481 and G20421;
	G25487<=G24485 and G20425;
	G25505<=G6707 and G25094;
	G25506<=G14263 and G25095;
	G25513<=G24487 and G17664;
	G25514<=G24488 and G20443;
	G25518<=G24489 and G20447;
	G25552<=G7009 and G25104;
	G25553<=G14385 and G25105;
	G25560<=G24494 and G17764;
	G25561<=G24495 and G20462;
	G25565<=G24496 and G20466;
	G25618<=G7259 and G25110;
	G25619<=G14497 and G25111;
	G25626<=G24504 and G17865;
	G25627<=G24505 and G20477;
	G25628<=G21008 and G25115;
	G25629<=G3024 and G25116;
	G25697<=G7455 and G25120;
	G25881<=G2908 and G25126;
	G25951<=G24800 and G13670;
	G25953<=G24783 and G13699;
	G25957<=G24782 and G11869;
	G25961<=G24770 and G11901;
	G25963<=G24756 and G11944;
	G25968<=G24871 and G11986;
	G25972<=G24859 and G12042;
	G25973<=G24847 and G13838;
	G25975<=G24606 and G21917;
	G25977<=G24845 and G12089;
	G25978<=G24836 and G13850;
	G25980<=G24663 and G21928;
	G25981<=G24819 and G13858;
	G26023<=G25422 and G24912;
	G26024<=G25301 and G21102;
	G26026<=G25431 and G24929;
	G26027<=G25418 and G22271;
	G26028<=G25438 and G24941;
	G26029<=G25445 and G24952;
	G26030<=G25429 and G22304;
	G26032<=G25379 and G19415;
	G26033<=G25395 and G19452;
	G26034<=G25405 and G19479;
	G26035<=G25523 and G19483;
	G26036<=G25413 and G19502;
	G26038<=G25589 and G19504;
	G26039<=G25668 and G19523;
	G26040<=G25745 and G19533;
	G26051<=G70 and G25296;
	G26052<=G25941 and G21087;
	G26053<=G758 and G25306;
	G26054<=G25944 and G21099;
	G26060<=G25943 and G21108;
	G26061<=G1444 and G25315;
	G26062<=G25947 and G21113;
	G26067<=G25946 and G21125;
	G26068<=G2138 and G25324;
	G26069<=G25949 and G21130;
	G26074<=G25948 and G21144;
	G26075<=G74 and G25698;
	G26080<=G25950 and G21164;
	G26082<=G762 and G25771;
	G26085<=G1448 and G25825;
	G26091<=G2142 and G25860;
	G26157<=G21825 and G25630;
	G26158<=G679 and G25937;
	G26163<=G1365 and G25939;
	G26166<=G686 and G25454;
	G26171<=G2059 and G25942;
	G26186<=G1372 and G25458;
	G26188<=G2753 and G25945;
	G26207<=G2066 and G25463;
	G26212<=G4217 and G25467;
	G26213<=G25895 and G9306;
	G26231<=G2760 and G25472;
	G26233<=G4340 and G25476;
	G26234<=G4343 and G25479;
	G26235<=G25895 and G9368;
	G26236<=G25899 and G9371;
	G26243<=G4372 and G25484;
	G26244<=G25903 and G9387;
	G26257<=G4465 and G25493;
	G26258<=G4468 and G25496;
	G26259<=G4471 and G25499;
	G26260<=G25254 and G17649;
	G26261<=G25895 and G9443;
	G26262<=G25899 and G9446;
	G26263<=G4476 and G25502;
	G26268<=G4509 and G25507;
	G26269<=G4512 and G25510;
	G26270<=G25903 and G9465;
	G26271<=G25907 and G9468;
	G26278<=G4541 and G25515;
	G26279<=G25911 and G9484;
	G26288<=G4592 and G25524;
	G26289<=G4595 and G25527;
	G26290<=G4598 and G25530;
	G26291<=G25899 and G9524;
	G26292<=G4603 and G25533;
	G26293<=G4606 and G25536;
	G26298<=G4641 and G25540;
	G26299<=G4644 and G25543;
	G26300<=G4647 and G25546;
	G26301<=G25258 and G17749;
	G26302<=G25903 and G9585;
	G26303<=G25907 and G9588;
	G26307<=G4652 and G25549;
	G26309<=G4685 and G25554;
	G26310<=G4688 and G25557;
	G26311<=G25911 and G9607;
	G26312<=G25915 and G9610;
	G26316<=G4717 and G25562;
	G26317<=G25919 and G9626;
	G26318<=G4737 and G25573;
	G26319<=G4740 and G25576;
	G26324<=G4743 and G25579;
	G26325<=G4746 and G25582;
	G26326<=G4749 and G25585;
	G26332<=G4769 and G25590;
	G26333<=G4772 and G25593;
	G26334<=G4775 and G25596;
	G26335<=G25907 and G9666;
	G26339<=G4780 and G25599;
	G26340<=G4783 and G25602;
	G26342<=G4818 and G25606;
	G26343<=G4821 and G25609;
	G26344<=G4824 and G25612;
	G26345<=G25261 and G17850;
	G26346<=G25911 and G9727;
	G26347<=G25915 and G9730;
	G26348<=G4829 and G25615;
	G26350<=G4862 and G25620;
	G26351<=G4865 and G25623;
	G26352<=G25919 and G9749;
	G26353<=G25923 and G9752;
	G26357<=G4882 and G25634;
	G26361<=G4888 and G25637;
	G26362<=G4891 and G25640;
	G26363<=G4894 and G25643;
	G26365<=G4913 and G25652;
	G26366<=G4916 and G25655;
	G26371<=G4919 and G25658;
	G26372<=G4922 and G25661;
	G26373<=G4925 and G25664;
	G26379<=G4945 and G25669;
	G26380<=G4948 and G25672;
	G26381<=G4951 and G25675;
	G26382<=G25915 and G9812;
	G26383<=G4956 and G25678;
	G26384<=G4959 and G25681;
	G26386<=G4994 and G25685;
	G26387<=G4997 and G25688;
	G26388<=G5000 and G25691;
	G26389<=G25264 and G17962;
	G26390<=G25919 and G9873;
	G26391<=G25923 and G9876;
	G26392<=G5005 and G25694;
	G26396<=G5027 and G25700;
	G26397<=G5030 and G25703;
	G26400<=G5041 and G25711;
	G26404<=G5047 and G25714;
	G26405<=G5050 and G25717;
	G26406<=G5053 and G25720;
	G26408<=G5072 and G25729;
	G26409<=G5075 and G25732;
	G26414<=G5078 and G25735;
	G26415<=G5081 and G25738;
	G26416<=G5084 and G25741;
	G26422<=G5104 and G25746;
	G26423<=G5107 and G25749;
	G26424<=G5110 and G25752;
	G26425<=G25923 and G9958;
	G26426<=G5115 and G25755;
	G26427<=G5118 and G25758;
	G26432<=G5145 and G25767;
	G26437<=G5156 and G25773;
	G26438<=G5159 and G25776;
	G26441<=G5170 and G25784;
	G26445<=G5176 and G25787;
	G26446<=G5179 and G25790;
	G26447<=G5182 and G25793;
	G26449<=G5201 and G25802;
	G26450<=G5204 and G25805;
	G26455<=G5207 and G25808;
	G26456<=G5210 and G25811;
	G26457<=G5213 and G25814;
	G26464<=G5238 and G25821;
	G26469<=G5249 and G25827;
	G26470<=G5252 and G25830;
	G26473<=G5263 and G25838;
	G26477<=G5269 and G25841;
	G26478<=G5272 and G25844;
	G26479<=G5275 and G25847;
	G26488<=G5301 and G25856;
	G26493<=G5312 and G25862;
	G26494<=G5315 and G25865;
	G26504<=G5338 and G25877;
	G26663<=G25274 and G21066;
	G26668<=G25283 and G21076;
	G26673<=G12431 and G25318;
	G26674<=G25291 and G21090;
	G26754<=G14657 and G26508;
	G26755<=G26083 and G22239;
	G26756<=G26113 and G22240;
	G26758<=G16614 and G26521 and G13637;
	G26759<=G26356 and G19251;
	G26760<=G26137 and G22256;
	G26761<=G26154 and G22257;
	G26763<=G14691 and G26516;
	G26764<=G16632 and G26525 and G13649;
	G26765<=G26399 and G19265;
	G26766<=G14725 and G26521;
	G26767<=G26087 and G22287;
	G26768<=G26440 and G19280;
	G26769<=G14753 and G26525;
	G26770<=G26059 and G19287;
	G26771<=G24912 and G26508 and G13614;
	G26773<=G26145 and G22303;
	G26774<=G26472 and G19299;
	G26775<=G26099 and G22318;
	G26777<=G26066 and G19305;
	G26778<=G24929 and G26516 and G13626;
	G26780<=G26119 and G16622;
	G26783<=G26073 and G19326;
	G26784<=G24941 and G26521 and G13637;
	G26787<=G26129 and G16636;
	G26790<=G26079 and G19353;
	G26791<=G24952 and G26525 and G13649;
	G26794<=G26143 and G16647;
	G26797<=G26148 and G16659;
	G26829<=G5623 and G26209;
	G26833<=G5651 and G26237;
	G26842<=G5689 and G26275;
	G26845<=G5664 and G26056;
	G26851<=G5741 and G26313;
	G26853<=G5716 and G26063;
	G26860<=G5774 and G26070;
	G26866<=G5833 and G26076;
	G26955<=G6157 and G26533;
	G26958<=G6184 and G26538;
	G26961<=G13907 and G26175;
	G26962<=G6180 and G26178;
	G26963<=G6216 and G26539;
	G26965<=G23320 and G26540;
	G26966<=G13963 and G26196;
	G26967<=G6212 and G26202;
	G26968<=G6305 and G26542;
	G26969<=G23320 and G26543;
	G26970<=G21976 and G26544;
	G26971<=G23325 and G26546;
	G26972<=G14033 and G26223;
	G26973<=G6301 and G26226;
	G26977<=G23320 and G26550;
	G26978<=G21976 and G26551;
	G26979<=G23331 and G26552;
	G26980<=G23360 and G26554;
	G26981<=G23325 and G26555;
	G26982<=G21983 and G26556;
	G26984<=G23335 and G26558;
	G26985<=G14124 and G26251;
	G26986<=G6438 and G26254;
	G26993<=G21976 and G26561;
	G26994<=G23331 and G26562;
	G26995<=G21991 and G26563;
	G26996<=G23360 and G26564;
	G26997<=G22050 and G26565;
	G26998<=G23325 and G26566;
	G26999<=G21983 and G26567;
	G27000<=G23340 and G26568;
	G27001<=G23364 and G26570;
	G27002<=G23335 and G26571;
	G27003<=G21996 and G26572;
	G27004<=G23344 and G26574;
	G27005<=G23331 and G26578;
	G27006<=G21991 and G26579;
	G27007<=G23360 and G26580;
	G27008<=G22050 and G26581;
	G27009<=G23368 and G26582;
	G27016<=G21983 and G26584;
	G27017<=G23340 and G26585;
	G27018<=G22005 and G26586;
	G27019<=G23364 and G26587;
	G27020<=G22069 and G26588;
	G27021<=G23335 and G26589;
	G27022<=G21996 and G26590;
	G27023<=G23349 and G26591;
	G27024<=G23372 and G26593;
	G27025<=G23344 and G26594;
	G27026<=G22009 and G26595;
	G27027<=G21991 and G26598;
	G27028<=G22050 and G26599;
	G27029<=G23368 and G26600;
	G27030<=G22083 and G26601;
	G27031<=G23340 and G26602;
	G27032<=G22005 and G26603;
	G27033<=G23364 and G26604;
	G27034<=G22069 and G26605;
	G27035<=G23377 and G26606;
	G27042<=G21996 and G26608;
	G27043<=G23349 and G26609;
	G27044<=G22016 and G26610;
	G27045<=G23372 and G26611;
	G27046<=G22093 and G26612;
	G27047<=G23344 and G26613;
	G27048<=G22009 and G26614;
	G27049<=G23353 and G26615;
	G27050<=G23381 and G26617;
	G27052<=G4885 and G26358;
	G27053<=G23368 and G26619;
	G27054<=G22083 and G26620;
	G27055<=G22005 and G26621;
	G27056<=G22069 and G26622;
	G27057<=G23377 and G26623;
	G27058<=G22108 and G26624;
	G27059<=G23349 and G26625;
	G27060<=G22016 and G26626;
	G27061<=G23372 and G26627;
	G27062<=G22093 and G26628;
	G27063<=G23388 and G26629;
	G27070<=G22009 and G26631;
	G27071<=G23353 and G26632;
	G27072<=G22021 and G26633;
	G27073<=G23381 and G26634;
	G27074<=G22118 and G26635;
	G27076<=G5024 and G26393;
	G27077<=G22083 and G26636;
	G27079<=G5044 and G26401;
	G27080<=G23377 and G26637;
	G27081<=G22108 and G26638;
	G27082<=G22016 and G26639;
	G27083<=G22093 and G26640;
	G27084<=G23388 and G26641;
	G27085<=G22134 and G26642;
	G27086<=G23353 and G26643;
	G27087<=G22021 and G26644;
	G27088<=G23381 and G26645;
	G27089<=G22118 and G26646;
	G27090<=G23395 and G26647;
	G27091<=G5142 and G26429;
	G27092<=G5153 and G26434;
	G27093<=G22108 and G26648;
	G27095<=G5173 and G26442;
	G27096<=G23388 and G26649;
	G27097<=G22134 and G26650;
	G27098<=G22021 and G26651;
	G27099<=G22118 and G26652;
	G27100<=G23395 and G26653;
	G27101<=G22157 and G26654;
	G27103<=G5235 and G26461;
	G27104<=G5246 and G26466;
	G27105<=G22134 and G26656;
	G27107<=G5266 and G26474;
	G27108<=G23395 and G26657;
	G27109<=G22157 and G26658;
	G27110<=G5298 and G26485;
	G27111<=G5309 and G26490;
	G27112<=G22157 and G26662;
	G27115<=G5335 and G26501;
	G27178<=G26110 and G22213;
	G27181<=G16570 and G26508 and G13614;
	G27182<=G26151 and G22217;
	G27185<=G26126 and G22230;
	G27187<=G16594 and G26516 and G13626;
	G27240<=G26905 and G22241;
	G27241<=G10730 and G26934;
	G27242<=G26793 and G8357;
	G27244<=G26914 and G22258;
	G27245<=G26877 and G22286;
	G27246<=G26988 and G16676;
	G27247<=G27011 and G16702;
	G27248<=G27037 and G16733;
	G27249<=G27065 and G16775;
	G27355<=G61 and G26837;
	G27356<=G65 and G26987;
	G27358<=G749 and G26846;
	G27359<=G753 and G27010;
	G27364<=G1435 and G26855;
	G27365<=G1439 and G27036;
	G27370<=G27126 and G8874;
	G27371<=G2129 and G26861;
	G27372<=G2133 and G27064;
	G27394<=G17802 and G27134;
	G27396<=G692 and G27135;
	G27407<=G17914 and G27136;
	G27409<=G1378 and G27137;
	G27425<=G18025 and G27138;
	G27427<=G2072 and G27139;
	G27446<=G18142 and G27141;
	G27448<=G2766 and G27142;
	G27495<=G23945 and G27146;
	G27509<=G23945 and G27148;
	G27516<=G23974 and G27151;
	G27530<=G23945 and G27153;
	G27534<=G23974 and G27155;
	G27541<=G24004 and G27159;
	G27552<=G23974 and G27162;
	G27554<=G24004 and G27164;
	G27561<=G24038 and G27167;
	G27568<=G24004 and G27172;
	G27570<=G24038 and G27173;
	G27578<=G24038 and G27177;
	G27656<=G26796 and G11004;
	G27657<=G27114 and G11051;
	G27659<=G27132 and G11114;
	G27660<=G26835 and G11117;
	G27661<=G26841 and G11173;
	G27666<=G26849 and G11243;
	G27671<=G26885 and G22212;
	G27673<=G26854 and G11312;
	G27679<=G26782 and G11386;
	G27680<=G26983 and G11392;
	G27681<=G26788 and G11456;
	G27719<=G27496 and G20649;
	G27720<=G27481 and G20652;
	G27721<=G27579 and G20655;
	G27723<=G27464 and G20679;
	G27725<=G27532 and G20704;
	G27726<=G27531 and G20732;
	G27727<=G27414 and G19301;
	G27728<=G27564 and G20766;
	G27729<=G27435 and G19322;
	G27730<=G27454 and G19349;
	G27731<=G27470 and G19383;
	G27732<=G27492 and G16758;
	G27733<=G27513 and G16785;
	G27734<=G27538 and G16814;
	G27737<=G27558 and G16832;
	G27770<=G5642 and G27449;
	G27772<=G5680 and G27465;
	G27773<=G5732 and G27484;
	G27774<=G5702 and G27361;
	G27775<=G5790 and G27506;
	G27779<=G5760 and G27367;
	G27783<=G5819 and G27373;
	G27790<=G5875 and G27376;
	G27904<=G13873 and G27387;
	G27908<=G13886 and G27391;
	G27909<=G13895 and G27397;
	G27913<=G4017 and G27401;
	G27914<=G13927 and G27404;
	G27915<=G13936 and G27410;
	G27922<=G4112 and G27416;
	G27923<=G4144 and G27419;
	G27924<=G13983 and G27422;
	G27926<=G13992 and G27428;
	G27931<=G4221 and G27432;
	G27935<=G4251 and G27437;
	G27936<=G4283 and G27440;
	G27938<=G14053 and G27443;
	G27945<=G4376 and G27451;
	G27949<=G4406 and G27456;
	G27951<=G4438 and G27459;
	G27963<=G4545 and G27467;
	G27968<=G4575 and G27472;
	G27970<=G14238 and G27475;
	G27984<=G4721 and G27486;
	G27985<=G14342 and G27489;
	G27991<=G14360 and G27498;
	G28008<=G27590 and G9770;
	G28009<=G14454 and G27510;
	G28015<=G14472 and G27518;
	G28027<=G27590 and G9895;
	G28028<=G27595 and G9898;
	G28035<=G27599 and G9916;
	G28036<=G14541 and G27535;
	G28042<=G14559 and G27543;
	G28050<=G27590 and G10018;
	G28051<=G27595 and G10021;
	G28057<=G27599 and G10049;
	G28058<=G27604 and G10052;
	G28065<=G27608 and G10070;
	G28066<=G14596 and G27555;
	G28073<=G27595 and G10109;
	G28079<=G27599 and G10127;
	G28080<=G27604 and G10130;
	G28086<=G27608 and G10158;
	G28087<=G27613 and G10161;
	G28094<=G27617 and G10179;
	G28098<=G27604 and G10214;
	G28104<=G27608 and G10232;
	G28105<=G27613 and G10235;
	G28111<=G27617 and G10263;
	G28112<=G27622 and G10266;
	G28116<=G27613 and G10316;
	G28122<=G27617 and G10334;
	G28123<=G27622 and G10337;
	G28127<=G27622 and G10409;
	G28171<=G27349 and G10898;
	G28176<=G27349 and G10940;
	G28188<=G27349 and G11008;
	G28193<=G27573 and G21914;
	G28319<=G27855 and G22246;
	G28320<=G27854 and G20637;
	G28322<=G27937 and G13868;
	G28323<=G8580 and G27838;
	G28324<=G27810 and G20659;
	G28326<=G27865 and G22274;
	G28327<=G27900 and G22275;
	G28329<=G27823 and G20708;
	G28330<=G27864 and G20711;
	G28331<=G27802 and G22307;
	G28332<=G27883 and G22331;
	G28333<=G27882 and G20772;
	G28334<=G27842 and G20793;
	G28335<=G27814 and G22343;
	G28336<=G27896 and G20810;
	G28337<=G28002 and G19448;
	G28338<=G28029 and G19475;
	G28339<=G28059 and G19498;
	G28340<=G28088 and G19519;
	G28373<=G56 and G27969;
	G28376<=G744 and G27990;
	G28378<=G52 and G27776;
	G28379<=G27868 and G19390 and G19369;
	G28380<=G1430 and G28014;
	G28381<=G28157 and G9815;
	G28383<=G740 and G27780;
	G28385<=G2124 and G28041;
	G28387<=G1426 and G27787;
	G28389<=G2120 and G27794;
	G28396<=G7754 and G27806;
	G28398<=G7769 and G27817;
	G28399<=G7776 and G27820;
	G28401<=G7782 and G27831;
	G28402<=G7785 and G27839;
	G28404<=G7792 and G27843;
	G28405<=G7796 and G27847;
	G28407<=G7799 and G27858;
	G28408<=G7806 and G27861;
	G28411<=G7809 and G27872;
	G28412<=G7812 and G27879;
	G28416<=G7823 and G27889;
	G28422<=G17640 and G28150;
	G28423<=G17724 and G28152;
	G28424<=G17741 and G28153;
	G28426<=G28128 and G9170;
	G28427<=G26092 and G28154;
	G28428<=G17825 and G28155;
	G28429<=G17842 and G28156;
	G28430<=G28128 and G9196;
	G28431<=G26092 and G28158;
	G28433<=G28133 and G9212;
	G28434<=G26114 and G28159;
	G28435<=G17937 and G28160;
	G28436<=G17954 and G28161;
	G28438<=G17882 and G27919;
	G28439<=G28128 and G9242;
	G28440<=G26092 and G28162;
	G28441<=G28133 and G9257;
	G28442<=G26114 and G28163;
	G28444<=G28137 and G9273;
	G28445<=G26121 and G28164;
	G28446<=G18048 and G28165;
	G28448<=G17974 and G27928;
	G28450<=G17993 and G27932;
	G28451<=G28133 and G9320;
	G28452<=G26114 and G28166;
	G28453<=G28137 and G9335;
	G28454<=G26121 and G28167;
	G28456<=G28141 and G9351;
	G28457<=G26131 and G28168;
	G28459<=G18074 and G27939;
	G28460<=G18091 and G27942;
	G28462<=G18110 and G27946;
	G28463<=G28137 and G9401;
	G28464<=G26121 and G28169;
	G28465<=G28141 and G9416;
	G28466<=G26131 and G28170;
	G28468<=G18265 and G28172;
	G28469<=G18179 and G27952;
	G28471<=G18190 and G27956;
	G28472<=G18207 and G27959;
	G28474<=G18226 and G27965;
	G28475<=G28141 and G9498;
	G28476<=G26131 and G28173;
	G28477<=G18341 and G28174;
	G28478<=G18358 and G28175;
	G28479<=G18286 and G27973;
	G28480<=G18297 and G27977;
	G28481<=G18314 and G27981;
	G28484<=G18436 and G28177;
	G28485<=G18453 and G28178;
	G28486<=G18379 and G27994;
	G28487<=G18390 and G27999;
	G28492<=G18509 and G28186;
	G28493<=G18526 and G28187;
	G28494<=G18474 and G28018;
	G28497<=G18573 and G28190;
	G28657<=G27925 and G13700;
	G28659<=G27917 and G13736;
	G28660<=G27916 and G11911;
	G28662<=G27911 and G11951;
	G28663<=G27906 and G11997;
	G28664<=G27997 and G12055;
	G28665<=G27827 and G22222;
	G28666<=G27980 and G12106;
	G28667<=G27964 and G13852;
	G28669<=G27897 and G22233;
	G28670<=G27798 and G21935;
	G28671<=G27962 and G12161;
	G28672<=G27950 and G13859;
	G28707<=G12436 and G28379;
	G28708<=G28392 and G22260;
	G28709<=G28400 and G22261;
	G28710<=G28403 and G22262;
	G28711<=G10749 and G28415;
	G28712<=G28406 and G22276;
	G28713<=G28410 and G22290;
	G28714<=G28394 and G22306;
	G28715<=G28414 and G22332;
	G28716<=G28449 and G19319;
	G28717<=G28461 and G19346;
	G28718<=G28473 and G19380;
	G28719<=G28482 and G19412;
	G28722<=G28523 and G16694;
	G28724<=G28551 and G16725;
	G28726<=G28578 and G16767;
	G28729<=G28606 and G16794;
	G28834<=G5751 and G28483;
	G28836<=G5810 and G28491;
	G28838<=G5866 and G28496;
	G28840<=G5913 and G28500;
	G28841<=G27834 and G28554;
	G28843<=G27834 and G28581;
	G28844<=G27850 and G28582;
	G28846<=G27834 and G28608;
	G28847<=G27850 and G28609;
	G28848<=G27875 and G28610;
	G28849<=G27850 and G28616;
	G28850<=G27875 and G28617;
	G28851<=G27892 and G28618;
	G28852<=G27875 and G28623;
	G28853<=G27892 and G28624;
	G28854<=G27892 and G28629;
	G28880<=G13946 and G28639;
	G28881<=G28612 and G9199;
	G28892<=G14001 and G28640;
	G28893<=G28612 and G9245;
	G28897<=G14016 and G28641;
	G28898<=G28619 and G9260;
	G28909<=G14062 and G28642;
	G28910<=G28612 and G9303;
	G28914<=G14092 and G28643;
	G28915<=G28619 and G9323;
	G28919<=G14107 and G28644;
	G28923<=G28625 and G9338;
	G28931<=G14153 and G28645;
	G28935<=G14177 and G28646;
	G28936<=G28619 and G9384;
	G28940<=G14207 and G28647;
	G28944<=G28625 and G9404;
	G28948<=G14222 and G28648;
	G28949<=G28630 and G9419;
	G28958<=G14268 and G28649;
	G28962<=G14292 and G28650;
	G28966<=G28625 and G9481;
	G28970<=G14322 and G28651;
	G28971<=G28630 and G9501;
	G28986<=G14390 and G28652;
	G28996<=G14414 and G28653;
	G28997<=G28630 and G9623;
	G29022<=G14502 and G28655;
	G29130<=G28397 and G22221;
	G29174<=G29031 and G20684;
	G29175<=G29009 and G20687;
	G29176<=G29097 and G20690;
	G29180<=G28982 and G20714;
	G29183<=G29064 and G20739;
	G29186<=G29063 and G20769;
	G29188<=G29083 and G20796;
	G29196<=G15022 and G28741;
	G29200<=G15096 and G28751;
	G29203<=G15118 and G28755;
	G29208<=G15188 and G28764;
	G29211<=G15210 and G28768;
	G29217<=G15274 and G28775;
	G29220<=G15296 and G28779;
	G29225<=G15366 and G28785;
	G29229<=G9293 and G28791;
	G29232<=G9356 and G28796;
	G29233<=G9374 and G28799;
	G29234<=G9427 and G28804;
	G29235<=G9453 and G28807;
	G29236<=G9471 and G28810;
	G29238<=G9569 and G28814;
	G29239<=G9595 and G28817;
	G29240<=G9613 and G28820;
	G29241<=G9711 and G28823;
	G29242<=G9737 and G28826;
	G29243<=G9857 and G28829;
	G29248<=G28855 and G8836;
	G29251<=G28855 and G8856;
	G29252<=G28859 and G8863;
	G29255<=G28855 and G8885;
	G29256<=G28859 and G8894;
	G29257<=G28863 and G8901;
	G29259<=G28859 and G8925;
	G29260<=G28863 and G8934;
	G29261<=G28867 and G8941;
	G29262<=G28863 and G8965;
	G29263<=G28867 and G8974;
	G29264<=G28867 and G8997;
	G29284<=G29001 and G28871;
	G29289<=G29030 and G28883;
	G29294<=G29053 and G28900;
	G29300<=G29072 and G28925;
	G29302<=G29026 and G28928;
	G29310<=G28978 and G28951;
	G29312<=G29049 and G28955;
	G29320<=G29088 and G28972;
	G29321<=G29008 and G28979;
	G29323<=G29068 and G28983;
	G29329<=G29096 and G29002;
	G29330<=G29038 and G29010;
	G29332<=G29080 and G29019;
	G29336<=G29045 and G29023;
	G29337<=G29103 and G29032;
	G29338<=G29060 and G29042;
	G29341<=G29062 and G29046;
	G29342<=G29107 and G29054;
	G29344<=G29076 and G29065;
	G29346<=G29087 and G29077;
	G29411<=G29090 and G21932;
	G29464<=G29190 and G8375;
	G29465<=G29191 and G8424;
	G29466<=G8587 and G29265;
	G29467<=G29340 and G19467;
	G29468<=G29343 and G19490;
	G29469<=G29345 and G19511;
	G29470<=G29347 and G19530;
	G29471<=G21461 and G29266;
	G29472<=G21461 and G29268;
	G29473<=G21508 and G29269;
	G29474<=G21508 and G29271;
	G29475<=G21544 and G29272;
	G29476<=G21544 and G29274;
	G29477<=G21580 and G29275;
	G29478<=G21580 and G29277;
	G29479<=G21461 and G29280;
	G29480<=G21461 and G29282;
	G29481<=G21508 and G29283;
	G29482<=G21461 and G29285;
	G29483<=G21508 and G29286;
	G29484<=G21544 and G29287;
	G29485<=G21508 and G29290;
	G29486<=G21544 and G29291;
	G29487<=G21580 and G29292;
	G29488<=G21544 and G29295;
	G29489<=G21580 and G29296;
	G29490<=G21580 and G29301;
	G29502<=G29350 and G8912;
	G29518<=G28728 and G29360;
	G29520<=G28731 and G29361;
	G29521<=G28733 and G29362;
	G29522<=G27735 and G29363;
	G29523<=G28737 and G29364;
	G29524<=G28739 and G29365;
	G29525<=G29195 and G29366;
	G29526<=G27741 and G29367;
	G29527<=G28748 and G29368;
	G29528<=G28750 and G29369;
	G29529<=G29199 and G29370;
	G29531<=G29202 and G29371;
	G29532<=G27746 and G29372;
	G29533<=G28762 and G29373;
	G29534<=G29206 and G29374;
	G29536<=G29207 and G29375;
	G29538<=G29210 and G29376;
	G29539<=G27754 and G29377;
	G29540<=G26041 and G29378;
	G29541<=G29214 and G29379;
	G29543<=G29215 and G29380;
	G29545<=G29216 and G29381;
	G29547<=G29219 and G29382;
	G29548<=G28784 and G29383;
	G29549<=G26043 and G29384;
	G29550<=G29222 and G29385;
	G29553<=G29223 and G29386;
	G29555<=G29224 and G29387;
	G29557<=G28789 and G29388;
	G29558<=G28790 and G29389;
	G29559<=G26045 and G29390;
	G29560<=G29227 and G29391;
	G29562<=G29228 and G29392;
	G29564<=G28794 and G29393;
	G29565<=G28795 and G29394;
	G29566<=G26047 and G29395;
	G29567<=G29231 and G29396;
	G29572<=G28802 and G29397;
	G29573<=G28803 and G29398;
	G29575<=G28813 and G29402;
	G29607<=G29193 and G11056;
	G29610<=G29349 and G11123;
	G29614<=G29359 and G11182;
	G29615<=G29245 and G11185;
	G29619<=G29247 and G11259;
	G29622<=G29250 and G11327;
	G29624<=G29254 and G11407;
	G29625<=G29189 and G11472;
	G29626<=G29318 and G11478;
	G29790<=G29491 and G10918;
	G29792<=G29491 and G10977;
	G29793<=G29491 and G11063;
	G29810<=G29748 and G22248;
	G29811<=G29703 and G20644;
	G29812<=G29762 and G12223;
	G29813<=G29760 and G13869;
	G29814<=G29728 and G22266;
	G29815<=G29727 and G20662;
	G29816<=G29759 and G13883;
	G29817<=G29709 and G20694;
	G29818<=G29732 and G22293;
	G29819<=G29751 and G22294;
	G29820<=G29717 and G20743;
	G29821<=G29731 and G20746;
	G29822<=G29705 and G22335;
	G29827<=G29741 and G22356;
	G29828<=G29740 and G20802;
	G29833<=G29725 and G20813;
	G29834<=G29713 and G22366;
	G29839<=G29747 and G20827;
	G29909<=G29735 and G19420 and G19401;
	G29910<=G29779 and G9961;
	G29942<=G29771 and G28877;
	G29944<=G29782 and G28889;
	G29945<=G29773 and G28894;
	G29946<=G29778 and G28906;
	G29947<=G29785 and G28911;
	G29948<=G29775 and G28916;
	G29949<=G29781 and G28932;
	G29950<=G29788 and G28937;
	G29951<=G29777 and G28945;
	G29952<=G29784 and G28959;
	G29953<=G29791 and G28967;
	G29954<=G29770 and G28975;
	G29955<=G29787 and G28993;
	G29956<=G29780 and G28998;
	G29957<=G29772 and G29005;
	G29958<=G29783 and G29027;
	G29959<=G29774 and G29035;
	G29960<=G29786 and G29050;
	G29961<=G29776 and G29057;
	G29962<=G29789 and G29069;
	G29963<=G29758 and G13737;
	G29964<=G29757 and G13786;
	G29965<=G29756 and G11961;
	G29966<=G29755 and G12004;
	G29967<=G29754 and G12066;
	G29968<=G29765 and G12119;
	G29969<=G29721 and G22237;
	G29970<=G29764 and G12178;
	G29971<=G29763 and G13861;
	G29980<=G29881 and G8324;
	G29981<=G29869 and G8330;
	G29982<=G29893 and G8336;
	G29983<=G29885 and G8344;
	G29984<=G29873 and G8351;
	G29985<=G29897 and G8363;
	G29986<=G29877 and G8366;
	G29987<=G29889 and G8369;
	G29988<=G29881 and G8382;
	G29989<=G29893 and G8391;
	G29990<=G29885 and G8397;
	G29991<=G29901 and G8403;
	G29992<=G12441 and G29909;
	G29993<=G29897 and G8411;
	G29994<=G29889 and G8418;
	G29995<=G29893 and G8434;
	G29996<=G29901 and G8443;
	G29997<=G29918 and G22277;
	G29998<=G29922 and G22278;
	G29999<=G29924 and G22279;
	G30000<=G10767 and G29930;
	G30001<=G29897 and G8449;
	G30002<=G29905 and G8455;
	G30003<=G29901 and G8469;
	G30004<=G29926 and G22295;
	G30005<=G29905 and G8478;
	G30006<=G29928 and G22310;
	G30007<=G29905 and G8494;
	G30008<=G29919 and G22334;
	G30009<=G29929 and G22357;
	G30077<=G29823 and G10963;
	G30079<=G29823 and G10988;
	G30080<=G29829 and G10996;
	G30081<=G29823 and G11022;
	G30082<=G29829 and G11036;
	G30083<=G29835 and G11048;
	G30085<=G29829 and G11092;
	G30086<=G29835 and G11108;
	G30087<=G29840 and G11120;
	G30088<=G29844 and G11138;
	G30089<=G29835 and G11160;
	G30090<=G29840 and G11176;
	G30091<=G29844 and G11202;
	G30092<=G29849 and G11205;
	G30093<=G29853 and G11222;
	G30094<=G29840 and G11246;
	G30095<=G29857 and G11265;
	G30096<=G29844 and G11268;
	G30097<=G29849 and G11271;
	G30098<=G29853 and G11284;
	G30099<=G29861 and G11287;
	G30100<=G29865 and G11306;
	G30101<=G29857 and G11341;
	G30102<=G29849 and G11348;
	G30103<=G29869 and G11358;
	G30104<=G29853 and G11361;
	G30105<=G29861 and G11364;
	G30106<=G29865 and G11379;
	G30107<=G29873 and G11382;
	G30108<=G29877 and G11401;
	G30109<=G29857 and G11411;
	G30110<=G29881 and G11417;
	G30111<=G29869 and G11425;
	G30112<=G29861 and G11432;
	G30113<=G29885 and G11444;
	G30114<=G29865 and G11447;
	G30115<=G29873 and G11450;
	G30116<=G29921 and G22236;
	G30117<=G29877 and G11465;
	G30118<=G29889 and G11468;
	G30123<=G30070 and G20641;
	G30127<=G30065 and G20719;
	G30128<=G30062 and G20722;
	G30129<=G30071 and G20725;
	G30131<=G30059 and G20749;
	G30132<=G30068 and G20776;
	G30133<=G30067 and G20799;
	G30138<=G30069 and G20816;
	G30216<=G30036 and G8921;
	G30217<=G30036 and G8955;
	G30218<=G30040 and G8961;
	G30219<=G30036 and G8980;
	G30220<=G30040 and G8987;
	G30221<=G30044 and G8993;
	G30222<=G30040 and G9010;
	G30223<=G30044 and G9016;
	G30224<=G30048 and G9022;
	G30225<=G30044 and G9035;
	G30226<=G30048 and G9041;
	G30227<=G30048 and G9058;
	G30327<=G30187 and G8321;
	G30330<=G30195 and G8333;
	G30333<=G30191 and G8341;
	G30334<=G30203 and G8347;
	G30337<=G30199 and G8354;
	G30340<=G30207 and G8372;
	G30345<=G30195 and G8388;
	G30348<=G30203 and G8400;
	G30351<=G30199 and G8408;
	G30352<=G30211 and G8414;
	G30355<=G30207 and G8421;
	G30361<=G30203 and G8440;
	G30364<=G30211 and G8452;
	G30367<=G30207 and G8460;
	G30372<=G8594 and G30228;
	G30374<=G30211 and G8475;
	G30387<=G30229 and G8888;
	G30388<=G30229 and G8918;
	G30389<=G30233 and G8928;
	G30390<=G30229 and G8952;
	G30391<=G30233 and G8958;
	G30392<=G30237 and G8968;
	G30393<=G30233 and G8984;
	G30394<=G30237 and G8990;
	G30395<=G30241 and G9000;
	G30396<=G30237 and G9013;
	G30397<=G30241 and G9019;
	G30398<=G30241 and G9038;
	G30407<=G30134 and G10991;
	G30409<=G30134 and G11025;
	G30410<=G30139 and G11028;
	G30411<=G30143 and G11039;
	G30436<=G30134 and G11079;
	G30437<=G30139 and G11082;
	G30438<=G30147 and G11085;
	G30440<=G30143 and G11095;
	G30441<=G30151 and G11098;
	G30442<=G30155 and G11111;
	G30444<=G30139 and G11132;
	G30445<=G30147 and G11135;
	G30447<=G30143 and G11145;
	G30448<=G30151 and G11148;
	G30449<=G30159 and G11151;
	G30451<=G30155 and G11163;
	G30452<=G30163 and G11166;
	G30453<=G30167 and G11179;
	G30454<=G30147 and G11199;
	G30457<=G30151 and G11216;
	G30458<=G30159 and G11219;
	G30460<=G30155 and G11231;
	G30461<=G30163 and G11234;
	G30462<=G30171 and G11237;
	G30464<=G30167 and G11249;
	G30465<=G30175 and G11252;
	G30467<=G30179 and G11274;
	G30469<=G30159 and G11281;
	G30472<=G30163 and G11300;
	G30473<=G30171 and G11303;
	G30475<=G30167 and G11315;
	G30476<=G30175 and G11318;
	G30477<=G30183 and G11321;
	G30478<=G30187 and G11344;
	G30481<=G30179 and G11351;
	G30484<=G30191 and G11367;
	G30486<=G30171 and G11376;
	G30489<=G30175 and G11395;
	G30490<=G30183 and G11398;
	G30492<=G30187 and G11414;
	G30495<=G30179 and G11422;
	G30496<=G30195 and G11428;
	G30499<=G30191 and G11435;
	G30502<=G30199 and G11453;
	G30504<=G30183 and G11462;
	G30696<=G30383 and G10943;
	G30697<=G30383 and G11011;
	G30698<=G30383 and G11126;
	G30728<=G30605 and G22252;
	G30735<=G30629 and G22268;
	G30736<=G30584 and G20669;
	G30743<=G30610 and G22283;
	G30744<=G30609 and G20697;
	G30750<=G30593 and G20729;
	G30754<=G30614 and G22313;
	G30755<=G30632 and G22314;
	G30757<=G30601 and G20780;
	G30758<=G30613 and G20783;
	G30759<=G30588 and G22360;
	G30760<=G30622 and G22379;
	G30761<=G30621 and G20822;
	G30762<=G30608 and G20830;
	G30763<=G30597 and G22386;
	G30764<=G30628 and G20837;
	G30766<=G30617 and G19457 and G19431;
	G30916<=G30785 and G22251;
	G30917<=G12446 and G30766;
	G30918<=G30780 and G22296;
	G30919<=G30786 and G22297;
	G30920<=G30787 and G22298;
	G30921<=G10773 and G30791;
	G30922<=G30788 and G22315;
	G30923<=G30789 and G22338;
	G30924<=G30783 and G22359;
	G30925<=G30790 and G22380;
	G30944<=G30935 and G20666;
	G30945<=G30931 and G20754;
	G30946<=G30930 and G20757;
	G30947<=G30936 and G20760;
	G30948<=G30929 and G20786;
	G30949<=G30933 and G20806;
	G30950<=G30932 and G20819;
	G30951<=G30934 and G20833;
	G30953<=G8605 and G30952;
	I16735<=G5856 and G4338 and G4339 and G5141;
	I16736<=G5713 and G5958 and G4735 and G4736;
	I16826<=G5903 and G4507 and G4508 and G5234;
	I16827<=G5771 and G5987 and G4911 and G4912;
	I16930<=G5942 and G4683 and G4684 and G5297;
	I16931<=G5830 and G6024 and G5070 and G5071;
	I17042<=G5976 and G4860 and G4861 and G5334;
	I17043<=G5886 and G6040 and G5199 and G5200;
	I17156<=G6898 and G2998 and G6901 and G3002;
	I17429<=G6901 and G7338 and G7146;
	I17599<=G7566 and G7583 and G7587;
	I19937<=G9507 and G9427 and G9356 and G9293;
	I19938<=G9232 and G9187 and G9161 and G9150;
	I19971<=G9649 and G9569 and G9453 and G9374;
	I19972<=G9310 and G9248 and G9203 and G9174;
	I19996<=G9795 and G9711 and G9595 and G9471;
	I19997<=G9391 and G9326 and G9264 and G9216;
	I20021<=G9941 and G9857 and G9737 and G9613;
	I20022<=G9488 and G9407 and G9342 and G9277;
	I20100<=G10186 and G3018 and G3028;
	I20131<=G8313 and G7542 and G2888 and G7566;
	I20132<=G2892 and G2903 and G7595 and G2908;
	I22028<=G13004 and G3018 and G7549;
	I22136<=G13082 and G2912 and G7522;
	I24619<=G14776 and G14837 and G16142;
	I24689<=G14811 and G14910 and G16201;
	I24738<=G14863 and G14991 and G16266;
	I24758<=G14936 and G15080 and G16325;
	I25280<=G18656 and G18670 and G18720;
	I25291<=G18679 and G18699 and G18758;
	I25300<=G18708 and G18735 and G18789;
	I25311<=G18744 and G18772 and G18815;
	I26240<=G18174 and G18341 and G17974;
	I26282<=G18188 and G18089 and G17991;
	I26285<=G18281 and G18436 and G18091;
	I26311<=G18353 and G13958 and G14011;
	I26317<=G18295 and G18205 and G18108;
	I26320<=G18374 and G18509 and G18207;
	I26348<=G18448 and G14028 and G14102;
	I26354<=G18388 and G18312 and G18224;
	I26357<=G18469 and G18573 and G18314;
	I26377<=G18521 and G14119 and G14217;
	I26383<=G18483 and G18405 and G18331;
	I26396<=G18585 and G14234 and G14332;
	I26416<=G18553 and G18491 and G18431;
	I26432<=G18277 and G18189 and G18090;
	I26440<=G18603 and G18555 and G18504;
	I26464<=G18370 and G18296 and G18206;
	I26472<=G18635 and G18605 and G18568;
	I26500<=G18465 and G18389 and G18313;
	I26508<=G18644 and G18637 and G18618;
	I26525<=G18656 and G18670 and G18692;
	I26528<=G18656 and G14837 and G13657;
	I26541<=G18538 and G18484 and G18406;
	I26558<=G14776 and G18670 and G18720;
	I26561<=G14776 and G18720 and G13657;
	I26564<=G18679 and G18699 and G18728;
	I26567<=G18679 and G14910 and G13687;
	I26590<=G14811 and G18699 and G18758;
	I26593<=G14811 and G18758 and G13687;
	I26596<=G18708 and G18735 and G18765;
	I26599<=G18708 and G14991 and G13724;
	I26615<=G14797 and G18692 and G13657;
	I26621<=G14863 and G18735 and G18789;
	I26624<=G14863 and G18789 and G13724;
	I26627<=G18744 and G18772 and G18796;
	I26630<=G18744 and G15080 and G13774;
	I26639<=G18656 and G18670 and G16142;
	I26645<=G14849 and G18728 and G13687;
	I26651<=G14936 and G18772 and G18815;
	I26654<=G14936 and G18815 and G13774;
	I26661<=G18679 and G18699 and G16201;
	I26667<=G14922 and G18765 and G13724;
	I26676<=G18708 and G18735 and G16266;
	I26682<=G15003 and G18796 and G13774;
	I26690<=G18744 and G18772 and G16325;
	I26695<=G18670 and G18692 and G16142;
	I26708<=G18699 and G18728 and G16201;
	I26726<=G18735 and G18765 and G16266;
	I26745<=G18772 and G18796 and G16325;
	I27695<=G19318 and G19300 and G19286;
	I27711<=G19262 and G19414 and G19386;
	I27717<=G19345 and G19321 and G19304;
	I27733<=G19277 and G19451 and G19416;
	I27739<=G19379 and G19348 and G19325;
	I27755<=G19296 and G19478 and G19453;
	I27761<=G19411 and G19382 and G19352;
	I27772<=G19314 and G19501 and G19480;
	I28068<=G17802 and G18265 and G17882;
	I28096<=G13907 and G14238 and G13946;
	I28103<=G17914 and G18358 and G17993;
	I28126<=G13963 and G14360 and G14016;
	I28133<=G18025 and G18453 and G18110;
	I28155<=G14033 and G14472 and G14107;
	I28162<=G18142 and G18526 and G18226;
	I28181<=G14124 and G14559 and G14222;
	I28582<=G19141 and G21133 and G21116;
	I28594<=G21167 and G21147 and G21134;
	I28609<=G21183 and G21168 and G21148;
	G7855<= not (I15168 and I15169);
	G7875<= not (I15184 and I15185);
	G7876<= not (I15191 and I15192);
	G7895<= not (I15205 and I15206);
	G7896<= not (I15212 and I15213);
	G7922<= not (I15238 and I15239);
	G7923<= not (I15245 and I15246);
	G7970<= not (I15277 and I15278);
	G8381<= not (G8182 and G8120 and G8044 and G7989);
	G8533<= not (G3398 and G3366);
	G8547<= not (G3398 and G3366);
	G8550<= not (G3554 and G3522);
	G8560<= not (G3554 and G3522);
	G8563<= not (G3710 and G3678);
	G8571<= not (G3710 and G3678);
	G8574<= not (G3866 and G3834);
	G8577<= not (G3866 and G3834);
	G9883<= not (I16880 and I16881);
	G10003<= not (I16966 and I16967);
	G10038<= not (G7772 and G3366);
	G10095<= not (I17060 and I17061);
	G10147<= not (G7788 and G3522);
	G10185<= not (I17150 and I17151);
	G10252<= not (G7802 and G3678);
	G10354<= not (G7815 and G3834);
	G10649<= not (G3398 and G6912);
	G10676<= not (G3398 and G6678);
	G10677<= not (G3398 and G6912);
	G10679<= not (G3554 and G7162);
	G10703<= not (G3398 and G6678);
	G10705<= not (G3554 and G6980);
	G10706<= not (G3554 and G7162);
	G10708<= not (G3710 and G7358);
	G10723<= not (G3554 and G6980);
	G10725<= not (G3710 and G7230);
	G10726<= not (G3710 and G7358);
	G10728<= not (G3866 and G7488);
	G10744<= not (G3710 and G7230);
	G10746<= not (G3866 and G7426);
	G10747<= not (G3866 and G7488);
	G10763<= not (G3866 and G7426);
	G11188<= not (I18107 and I18108);
	G11189<= not (I18114 and I18115);
	G11262<= not (I18191 and I18192);
	G11263<= not (I18198 and I18199);
	G11264<= not (I18205 and I18206);
	G11330<= not (I18281 and I18282);
	G11331<= not (I18288 and I18289);
	G11410<= not (I18369 and I18370);
	G11617<= not (G8313 and G2883);
	G11621<= not (I18800 and I18801);
	G11661<= not (G9534 and G3366);
	G11662<= not (G9534 and G3366);
	G11672<= not (G9534 and G3366);
	G11673<= not (G9676 and G3522);
	G11674<= not (G9676 and G3522);
	G11683<= not (G9534 and G3366);
	G11684<= not (G9676 and G3522);
	G11685<= not (G9822 and G3678);
	G11686<= not (G9822 and G3678);
	G11691<= not (G9534 and G3366);
	G11692<= not (G9676 and G3522);
	G11693<= not (G9822 and G3678);
	G11694<= not (G9968 and G3834);
	G11695<= not (G9968 and G3834);
	G11696<= not (G9534 and G3366);
	G11698<= not (G9676 and G3522);
	G11699<= not (G9822 and G3678);
	G11700<= not (G9968 and G3834);
	G11701<= not (G9534 and G3366);
	G11702<= not (G9676 and G3522);
	G11704<= not (G9822 and G3678);
	G11705<= not (G9968 and G3834);
	G11707<= not (G9534 and G3366);
	G11708<= not (G9534 and G3366);
	G11709<= not (G9676 and G3522);
	G11710<= not (G9822 and G3678);
	G11712<= not (G9968 and G3834);
	G11713<= not (G10481 and G9144);
	G11716<= not (G9534 and G3366);
	G11717<= not (G9676 and G3522);
	G11718<= not (G9676 and G3522);
	G11719<= not (G9822 and G3678);
	G11720<= not (G9968 and G3834);
	G11721<= not (G9534 and G3366);
	G11722<= not (G9676 and G3522);
	G11723<= not (G9822 and G3678);
	G11724<= not (G9822 and G3678);
	G11725<= not (G9968 and G3834);
	G11726<= not (G9676 and G3522);
	G11727<= not (G9822 and G3678);
	G11728<= not (G9968 and G3834);
	G11729<= not (G9968 and G3834);
	G11730<= not (G9822 and G3678);
	G11731<= not (G9968 and G3834);
	G11733<= not (G9968 and G3834);
	G12433<= not (G2879 and G10778);
	G12486<= not (G8278 and G6448);
	G12503<= not (G8278 and G5438);
	G12506<= not (G8287 and G6713);
	G12520<= not (G8287 and G5473);
	G12523<= not (G8296 and G7015);
	G12535<= not (G8296 and G5512);
	G12538<= not (G8305 and G7265);
	G12544<= not (G8305 and G5556);
	G12988<= not (I20032 and I20033);
	G12999<= not (I20049 and I20050);
	G13020<= not (G9534 and G6912);
	G13021<= not (G9534 and G6912);
	G13026<= not (G9534 and G6678);
	G13027<= not (G9534 and G6912);
	G13028<= not (G9534 and G6678);
	G13029<= not (G9676 and G7162);
	G13030<= not (G9676 and G7162);
	G13034<= not (G9534 and G6678);
	G13035<= not (G9534 and G6912);
	G13037<= not (G9676 and G6980);
	G13038<= not (G9676 and G7162);
	G13039<= not (G9676 and G6980);
	G13040<= not (G9822 and G7358);
	G13041<= not (G9822 and G7358);
	G13044<= not (G9534 and G6678);
	G13045<= not (G9534 and G6912);
	G13047<= not (G9676 and G6980);
	G13048<= not (G9676 and G7162);
	G13050<= not (G9822 and G7230);
	G13051<= not (G9822 and G7358);
	G13052<= not (G9822 and G7230);
	G13053<= not (G9968 and G7488);
	G13054<= not (G9968 and G7488);
	G13058<= not (G9534 and G6678);
	G13059<= not (G9534 and G6912);
	G13061<= not (G9676 and G6980);
	G13062<= not (G9676 and G7162);
	G13064<= not (G9822 and G7230);
	G13065<= not (G9822 and G7358);
	G13067<= not (G9968 and G7426);
	G13068<= not (G9968 and G7488);
	G13069<= not (G9968 and G7426);
	G13071<= not (G9534 and G6678);
	G13072<= not (G9534 and G6912);
	G13074<= not (G9676 and G6980);
	G13075<= not (G9676 and G7162);
	G13077<= not (G9822 and G7230);
	G13078<= not (G9822 and G7358);
	G13080<= not (G9968 and G7426);
	G13081<= not (G9968 and G7488);
	G13087<= not (G9534 and G6678);
	G13088<= not (G9534 and G6912);
	G13089<= not (G9534 and G6912);
	G13090<= not (G9676 and G6980);
	G13091<= not (G9676 and G7162);
	G13093<= not (G9822 and G7230);
	G13094<= not (G9822 and G7358);
	G13096<= not (G9968 and G7426);
	G13097<= not (G9968 and G7488);
	G13098<= not (G9534 and G6678);
	G13099<= not (G9534 and G6912);
	G13100<= not (G9534 and G6678);
	G13102<= not (G9676 and G6980);
	G13103<= not (G9676 and G7162);
	G13104<= not (G9676 and G7162);
	G13105<= not (G9822 and G7230);
	G13106<= not (G9822 and G7358);
	G13108<= not (G9968 and G7426);
	G13109<= not (G9968 and G7488);
	G13112<= not (G9534 and G6678);
	G13113<= not (G9534 and G6912);
	G13114<= not (G9676 and G6980);
	G13115<= not (G9676 and G7162);
	G13116<= not (G9676 and G6980);
	G13118<= not (G9822 and G7230);
	G13119<= not (G9822 and G7358);
	G13120<= not (G9822 and G7358);
	G13121<= not (G9968 and G7426);
	G13122<= not (G9968 and G7488);
	G13123<= not (G9534 and G6678);
	G13125<= not (G9676 and G6980);
	G13126<= not (G9676 and G7162);
	G13127<= not (G9822 and G7230);
	G13128<= not (G9822 and G7358);
	G13129<= not (G9822 and G7230);
	G13131<= not (G9968 and G7426);
	G13132<= not (G9968 and G7488);
	G13133<= not (G9968 and G7488);
	G13134<= not (G9676 and G6980);
	G13136<= not (G9822 and G7230);
	G13137<= not (G9822 and G7358);
	G13138<= not (G9968 and G7426);
	G13139<= not (G9968 and G7488);
	G13140<= not (G9968 and G7426);
	G13142<= not (G9822 and G7230);
	G13144<= not (G9968 and G7426);
	G13145<= not (G9968 and G7488);
	G13146<= not (G9968 and G7426);
	G13147<= not (G8278 and G3306);
	G13150<= not (G8287 and G3462);
	G13156<= not (G8296 and G3618);
	G13165<= not (G8305 and G3774);
	G13245<= not (G10779 and G7901);
	G13305<= not (G8317 and G2993);
	G13348<= not (I20430 and I20431);
	G13370<= not (I20466 and I20467);
	G13399<= not (I20505 and I20506);
	G13476<= not (G12565 and G3254);
	G13478<= not (G12611 and G3410);
	G13482<= not (G12657 and G3566);
	G13494<= not (G12565 and G3254);
	G13495<= not (G12611 and G3410);
	G13497<= not (G12657 and G3566);
	G13501<= not (G12711 and G3722);
	G13507<= not (I20744 and I20745);
	G13510<= not (G12565 and G3254);
	G13511<= not (G12611 and G3410);
	G13512<= not (G12657 and G3566);
	G13514<= not (G12711 and G3722);
	G13518<= not (G12565 and G3254);
	G13524<= not (G12611 and G3410);
	G13525<= not (G12657 and G3566);
	G13526<= not (G12711 and G3722);
	G13528<= not (G12565 and G3254);
	G13529<= not (G12611 and G3410);
	G13535<= not (G12657 and G3566);
	G13536<= not (G12711 and G3722);
	G13537<= not (G12565 and G3254);
	G13538<= not (G12565 and G3254);
	G13539<= not (G12611 and G3410);
	G13540<= not (G12657 and G3566);
	G13546<= not (G12711 and G3722);
	G13547<= not (G12565 and G3254);
	G13548<= not (G12611 and G3410);
	G13549<= not (G12611 and G3410);
	G13550<= not (G12657 and G3566);
	G13551<= not (G12711 and G3722);
	G13557<= not (G12611 and G3410);
	G13558<= not (G12657 and G3566);
	G13559<= not (G12657 and G3566);
	G13560<= not (G12711 and G3722);
	G13561<= not (G12657 and G3566);
	G13562<= not (G12711 and G3722);
	G13563<= not (G12711 and G3722);
	G13564<= not (G12711 and G3722);
	G13599<= not (G12886 and G3366);
	G13611<= not (G12926 and G3522);
	G13621<= not (G12955 and G3678);
	G13633<= not (G12984 and G3834);
	G13893<= not (G8580 and G12463);
	G13915<= not (G8822 and G12473 and G12463);
	G13934<= not (G8587 and G12478);
	G13957<= not (G10730 and G12473);
	G13971<= not (G8846 and G12490 and G12478);
	G13990<= not (G8594 and G12495);
	G14027<= not (G10749 and G12490);
	G14041<= not (G8873 and G12510 and G12495);
	G14060<= not (G8605 and G12515);
	G14118<= not (G10767 and G12510);
	G14132<= not (G8911 and G12527 and G12515);
	G14233<= not (G10773 and G12527);
	G15454<= not (G9232 and G9150 and G12780);
	G15540<= not (G9310 and G9174 and G12819);
	G15618<= not (G9391 and G9216 and G12857);
	G15660<= not (G13401 and G12354);
	G15664<= not (G12565 and G6314);
	G15694<= not (G9488 and G9277 and G12898);
	G15718<= not (G13286 and G12354);
	G15719<= not (G13401 and G12392);
	G15720<= not (G12565 and G6232);
	G15721<= not (G12565 and G6314);
	G15723<= not (G12611 and G6519);
	G15756<= not (G13313 and G12354);
	G15757<= not (G11622 and G12392);
	G15758<= not (G12565 and G6232);
	G15759<= not (G12565 and G6314);
	G15760<= not (G12611 and G6369);
	G15761<= not (G12611 and G6519);
	G15763<= not (G12657 and G6783);
	G15782<= not (G13332 and G12354);
	G15783<= not (G11643 and G12392);
	G15784<= not (G12565 and G6232);
	G15785<= not (G12565 and G6314);
	G15786<= not (G12611 and G6369);
	G15787<= not (G12611 and G6519);
	G15788<= not (G12657 and G6574);
	G15789<= not (G12657 and G6783);
	G15791<= not (G12711 and G7085);
	G15803<= not (G13375 and G12354);
	G15804<= not (G11660 and G12392);
	G15805<= not (G12565 and G6232);
	G15806<= not (G12565 and G6314);
	G15807<= not (G12611 and G6369);
	G15808<= not (G12611 and G6519);
	G15809<= not (G12657 and G6574);
	G15810<= not (G12657 and G6783);
	G15811<= not (G12711 and G6838);
	G15812<= not (G12711 and G7085);
	G15814<= not (I22063 and I22064);
	G15818<= not (G13024 and G12354);
	G15819<= not (G13286 and G12392);
	G15820<= not (G12565 and G6232);
	G15821<= not (G12565 and G6314);
	G15822<= not (G12611 and G6369);
	G15823<= not (G12611 and G6519);
	G15824<= not (G12657 and G6574);
	G15825<= not (G12657 and G6783);
	G15826<= not (G12711 and G6838);
	G15827<= not (G12711 and G7085);
	G15830<= not (G13310 and G12392);
	G15831<= not (G13313 and G12392);
	G15832<= not (G12565 and G6232);
	G15833<= not (G12565 and G6314);
	G15834<= not (G12611 and G6369);
	G15835<= not (G12611 and G6519);
	G15836<= not (G12657 and G6574);
	G15837<= not (G12657 and G6783);
	G15838<= not (G12711 and G6838);
	G15839<= not (G12711 and G7085);
	G15841<= not (G13331 and G12392);
	G15842<= not (G13332 and G12392);
	G15843<= not (G12565 and G6314);
	G15844<= not (G12565 and G6232);
	G15845<= not (G12565 and G6314);
	G15846<= not (G12611 and G6369);
	G15847<= not (G12611 and G6519);
	G15848<= not (G12657 and G6574);
	G15849<= not (G12657 and G6783);
	G15850<= not (G12711 and G6838);
	G15851<= not (G12711 and G7085);
	G15853<= not (G13310 and G12354);
	G15854<= not (G13353 and G12392);
	G15855<= not (G13354 and G12392);
	G15856<= not (G12565 and G6232);
	G15857<= not (G12565 and G6314);
	G15858<= not (G12565 and G6232);
	G15866<= not (G12611 and G6519);
	G15867<= not (G12611 and G6369);
	G15868<= not (G12611 and G6519);
	G15869<= not (G12657 and G6574);
	G15870<= not (G12657 and G6783);
	G15871<= not (G12711 and G6838);
	G15872<= not (G12711 and G7085);
	G15877<= not (G13374 and G12392);
	G15878<= not (G13375 and G12392);
	G15879<= not (G12565 and G6232);
	G15887<= not (G12611 and G6369);
	G15888<= not (G12611 and G6519);
	G15889<= not (G12611 and G6369);
	G15897<= not (G12657 and G6783);
	G15898<= not (G12657 and G6574);
	G15899<= not (G12657 and G6783);
	G15900<= not (G12711 and G6838);
	G15901<= not (G12711 and G7085);
	G15903<= not (G13404 and G12392);
	G15912<= not (G12611 and G6369);
	G15920<= not (G12657 and G6574);
	G15921<= not (G12657 and G6783);
	G15922<= not (G12657 and G6574);
	G15930<= not (G12711 and G7085);
	G15931<= not (G12711 and G6838);
	G15932<= not (G12711 and G7085);
	G15941<= not (G12657 and G6574);
	G15949<= not (G12711 and G6838);
	G15950<= not (G12711 and G7085);
	G15951<= not (G12711 and G6838);
	G15970<= not (G12711 and G6838);
	G15990<= not (G12886 and G6912);
	G15992<= not (G12886 and G6678);
	G15993<= not (G12926 and G7162);
	G15995<= not (G12926 and G6980);
	G15996<= not (G12955 and G7358);
	G15999<= not (G12955 and G7230);
	G16000<= not (G12984 and G7488);
	G16006<= not (G12984 and G7426);
	G16085<= not (G12883 and G633);
	G16123<= not (G12923 and G1319);
	G16132<= not (I22283 and I22284);
	G16174<= not (G12952 and G2013);
	G16181<= not (I22317 and I22318);
	G16233<= not (G12981 and G2707);
	G16341<= not (G12377 and G12407);
	G16412<= not (G12565 and G3254);
	G16439<= not (G13082 and G2912);
	G16442<= not (G12565 and G3254);
	G16446<= not (G12611 and G3410);
	G16463<= not (G13004 and G3018);
	G16536<= not (G15873 and G2896);
	G16566<= not (I22631 and I22632);
	G16662<= not (I22706 and I22707);
	G16935<= not (I22885 and I22886);
	G16965<= not (I22901 and I22902);
	G16985<= not (I22918 and I22919);
	G16986<= not (I22925 and I22926);
	G16992<= not (I22937 and I22938);
	G16995<= not (I22946 and I22947);
	G16996<= not (I22953 and I22954);
	G17000<= not (I22963 and I22964);
	G17016<= not (I22973 and I22974);
	G17019<= not (I22982 and I22983);
	G17020<= not (I22989 and I22990);
	G17024<= not (I22999 and I23000);
	G17030<= not (I23009 and I23010);
	G17046<= not (I23019 and I23020);
	G17049<= not (I23028 and I23029);
	G17050<= not (I23035 and I23036);
	G17058<= not (I23046 and I23047);
	G17064<= not (I23056 and I23057);
	G17080<= not (I23066 and I23067);
	G17083<= not (I23075 and I23076);
	G17085<= not (I23083 and I23084);
	G17093<= not (I23094 and I23095);
	G17099<= not (I23104 and I23105);
	G17115<= not (I23114 and I23115);
	G17118<= not (G13915 and G13893);
	G17121<= not (I23124 and I23125);
	G17123<= not (I23132 and I23133);
	G17131<= not (I23143 and I23144);
	G17137<= not (I23153 and I23154);
	G17139<= not (G13957 and G13915);
	G17142<= not (I23162 and I23163);
	G17145<= not (G13971 and G13934);
	G17148<= not (I23172 and I23173);
	G17150<= not (I23180 and I23181);
	G17158<= not (I23191 and I23192);
	G17159<= not (G14642 and G14657);
	G17160<= not (I23199 and I23200);
	G17162<= not (G14027 and G13971);
	G17165<= not (I23208 and I23209);
	G17168<= not (G14041 and G13990);
	G17171<= not (I23218 and I23219);
	G17173<= not (I23226 and I23227);
	G17174<= not (G14669 and G14691);
	G17175<= not (I23234 and I23235);
	G17177<= not (G14118 and G14041);
	G17180<= not (I23243 and I23244);
	G17183<= not (G14132 and G14060);
	G17190<= not (I23257 and I23258);
	G17191<= not (G14703 and G14725);
	G17192<= not (I23265 and I23266);
	G17194<= not (G14233 and G14132);
	G17201<= not (I23278 and I23279);
	G17202<= not (G14737 and G14753);
	G17729<= not (I23807 and I23808);
	G17807<= not (I23879 and I23880);
	G17830<= not (I23894 and I23895);
	G17887<= not (I23942 and I23943);
	G17913<= not (I23959 and I23960);
	G17919<= not (I23967 and I23968);
	G17942<= not (I23982 and I23983);
	G17968<= not (I24006 and I24007);
	G17979<= not (I24016 and I24017);
	G17985<= not (G14641 and G9636);
	G17992<= not (I24029 and I24030);
	G17998<= not (I24037 and I24038);
	G18024<= not (I24054 and I24055);
	G18030<= not (I24062 and I24063);
	G18053<= not (I24077 and I24078);
	G18079<= not (I24092 and I24093);
	G18090<= not (I24103 and I24104);
	G18096<= not (I24111 and I24112);
	G18102<= not (G14668 and G9782);
	G18109<= not (I24124 and I24125);
	G18115<= not (I24132 and I24133);
	G18141<= not (I24149 and I24150);
	G18147<= not (I24157 and I24158);
	G18183<= not (I24179 and I24180);
	G18189<= not (I24187 and I24188);
	G18195<= not (I24195 and I24196);
	G18206<= not (I24206 and I24207);
	G18212<= not (I24214 and I24215);
	G18218<= not (G14702 and G9928);
	G18225<= not (I24227 and I24228);
	G18231<= not (I24235 and I24236);
	G18257<= not (I24252 and I24253);
	G18270<= not (I24264 and I24265);
	G18276<= not (I24272 and I24273);
	G18277<= not (I24279 and I24280);
	G18290<= not (I24291 and I24292);
	G18296<= not (I24299 and I24300);
	G18302<= not (I24307 and I24308);
	G18313<= not (I24318 and I24319);
	G18319<= not (I24326 and I24327);
	G18325<= not (G14736 and G10082);
	G18332<= not (I24339 and I24340);
	G18346<= not (I24352 and I24353);
	G18354<= not (I24362 and I24363);
	G18363<= not (I24373 and I24374);
	G18369<= not (I24381 and I24382);
	G18370<= not (I24388 and I24389);
	G18383<= not (I24400 and I24401);
	G18389<= not (I24408 and I24409);
	G18395<= not (I24416 and I24417);
	G18406<= not (I24427 and I24428);
	G18419<= not (I24437 and I24438);
	G18424<= not (I24444 and I24445);
	G18431<= not (I24453 and I24454);
	G18441<= not (I24465 and I24466);
	G18449<= not (I24475 and I24476);
	G18458<= not (I24486 and I24487);
	G18464<= not (I24494 and I24495);
	G18465<= not (I24501 and I24502);
	G18478<= not (I24513 and I24514);
	G18484<= not (I24521 and I24522);
	G18491<= not (I24531 and I24532);
	G18492<= not (I24538 and I24539);
	G18497<= not (I24545 and I24546);
	G18504<= not (I24554 and I24555);
	G18514<= not (I24566 and I24567);
	G18522<= not (I24576 and I24577);
	G18531<= not (I24587 and I24588);
	G18537<= not (I24595 and I24596);
	G18538<= not (I24602 and I24603);
	G18542<= not (I24612 and I24613);
	G18553<= not (I24625 and I24626);
	G18555<= not (I24633 and I24634);
	G18556<= not (I24640 and I24641);
	G18561<= not (I24647 and I24648);
	G18568<= not (I24656 and I24657);
	G18578<= not (I24668 and I24669);
	G18586<= not (I24678 and I24679);
	G18603<= not (I24695 and I24696);
	G18605<= not (I24703 and I24704);
	G18606<= not (I24710 and I24711);
	G18611<= not (I24717 and I24718);
	G18618<= not (I24726 and I24727);
	G18635<= not (I24744 and I24745);
	G18637<= not (I24752 and I24753);
	G18644<= not (I24764 and I24765);
	G18977<= not (G15797 and G3006);
	G18980<= not (I25031 and I25032);
	G19067<= not (G16554 and G16578);
	G19084<= not (G16586 and G16602);
	G19103<= not (G18590 and G2924);
	G19121<= not (G16682 and G16697);
	G19128<= not (G16708 and G16728);
	G19135<= not (G16739 and G16770);
	G19138<= not (G16781 and G16797);
	G19141<= not (G3088 and G16825);
	G19152<= not (G5378 and G18884);
	G19261<= not (I25533 and I25534);
	G19262<= not (I25540 and I25541);
	G19271<= not (I25561 and I25562);
	G19276<= not (I25572 and I25573);
	G19277<= not (I25579 and I25580);
	G19286<= not (I25596 and I25597);
	G19288<= not (G14685 and G8580 and G17057);
	G19290<= not (I25606 and I25607);
	G19295<= not (I25617 and I25618);
	G19296<= not (I25624 and I25625);
	G19300<= not (I25634 and I25635);
	G19304<= not (I25644 and I25645);
	G19306<= not (G14719 and G8587 and G17092);
	G19308<= not (I25654 and I25655);
	G19313<= not (I25665 and I25666);
	G19314<= not (I25672 and I25673);
	G19318<= not (I25682 and I25683);
	G19321<= not (I25691 and I25692);
	G19325<= not (I25701 and I25702);
	G19327<= not (G14747 and G8594 and G17130);
	G19329<= not (I25711 and I25712);
	G19334<= not (I25722 and I25723);
	G19345<= not (I25732 and I25733);
	G19348<= not (I25741 and I25742);
	G19352<= not (I25751 and I25752);
	G19354<= not (G14768 and G8605 and G17157);
	G19357<= not (I25762 and I25763);
	G19368<= not (I25772 and I25773);
	G19379<= not (I25782 and I25783);
	G19382<= not (I25791 and I25792);
	G19386<= not (I25801 and I25802);
	G19389<= not (I25810 and I25811);
	G19400<= not (I25820 and I25821);
	G19411<= not (I25830 and I25831);
	G19414<= not (I25839 and I25840);
	G19416<= not (I25847 and I25848);
	G19419<= not (I25856 and I25857);
	G19430<= not (I25866 and I25867);
	G19451<= not (I25881 and I25882);
	G19453<= not (I25889 and I25890);
	G19456<= not (I25898 and I25899);
	G19478<= not (I25914 and I25915);
	G19480<= not (I25922 and I25923);
	G19501<= not (I25939 and I25940);
	G19865<= not (G16607 and G9636);
	G19896<= not (G16625 and G9782);
	G19921<= not (G16639 and G9928);
	G19936<= not (G16650 and G10082);
	G19954<= not (G17186 and G92);
	G19984<= not (G17197 and G780);
	G20022<= not (G17204 and G1466);
	G20064<= not (G17209 and G2160);
	G20473<= not (G18085 and G646);
	G20481<= not (G18201 and G1332);
	G20487<= not (G18308 and G2026);
	G20493<= not (G18401 and G2720);
	G20497<= not (G5410 and G18886);
	G20522<= not (G16501 and G16515);
	G20537<= not (G18626 and G3036);
	G20542<= not (G16523 and G16546);
	G20633<= not (G20164 and G3254);
	G20648<= not (G20164 and G3254);
	G20658<= not (G20198 and G3410);
	G20672<= not (G20164 and G3254);
	G20683<= not (G20198 and G3410);
	G20693<= not (G20228 and G3566);
	G20700<= not (G20153 and G2903);
	G20703<= not (G20164 and G3254);
	G20707<= not (G20198 and G3410);
	G20718<= not (G20228 and G3566);
	G20728<= not (G20255 and G3722);
	G20738<= not (G20198 and G3410);
	G20742<= not (G20228 and G3566);
	G20753<= not (G20255 and G3722);
	G20775<= not (G20228 and G3566);
	G20779<= not (G20255 and G3722);
	G20805<= not (G20255 and G3722);
	G20825<= not (G19219 and G15959);
	G21659<= not (G20164 and G6314);
	G21660<= not (I28190 and I28191);
	G21685<= not (G20164 and G6232);
	G21686<= not (G20164 and G6314);
	G21688<= not (G20198 and G6519);
	G21689<= not (I28218 and I28219);
	G21714<= not (G20164 and G6232);
	G21715<= not (G20164 and G6314);
	G21720<= not (G14256 and G15177 and G19871 and G19842);
	G21721<= not (G20198 and G6369);
	G21722<= not (G20198 and G6519);
	G21724<= not (G20228 and G6783);
	G21725<= not (I28248 and I28249);
	G21736<= not (G20164 and G6232);
	G21737<= not (G20164 and G6314);
	G21740<= not (G20198 and G6369);
	G21741<= not (G20198 and G6519);
	G21746<= not (G14378 and G15263 and G19902 and G19875);
	G21747<= not (G20228 and G6574);
	G21748<= not (G20228 and G6783);
	G21750<= not (G20255 and G7085);
	G21751<= not (I28272 and I28273);
	G21759<= not (G20164 and G6232);
	G21760<= not (G20198 and G6369);
	G21761<= not (G20198 and G6519);
	G21764<= not (G20228 and G6574);
	G21765<= not (G20228 and G6783);
	G21770<= not (G14490 and G15355 and G19927 and G19906);
	G21771<= not (G20255 and G6838);
	G21772<= not (G20255 and G7085);
	G21775<= not (G20198 and G6369);
	G21776<= not (G20228 and G6574);
	G21777<= not (G20228 and G6783);
	G21780<= not (G20255 and G6838);
	G21781<= not (G20255 and G7085);
	G21786<= not (G14577 and G15441 and G19942 and G19931);
	G21790<= not (G20228 and G6574);
	G21791<= not (G20255 and G6838);
	G21792<= not (G20255 and G7085);
	G21804<= not (G20255 and G6838);
	G21848<= not (G17807 and G19181 and G19186);
	G21850<= not (G17979 and G19187 and G19191);
	G21855<= not (G17919 and G19188 and G19193);
	G21857<= not (G18079 and G19192 and G19200);
	G21858<= not (G18096 and G19194 and G19202);
	G21859<= not (G18030 and G19195 and G19204);
	G21860<= not (G18270 and G19201 and G19209);
	G21862<= not (G18195 and G19203 and G19211);
	G21863<= not (G18212 and G19205 and G19213);
	G21864<= not (G18147 and G19206 and G19215);
	G21865<= not (G18424 and G19210 and G19221);
	G21866<= not (G18363 and G19212 and G19222);
	G21868<= not (G18302 and G19214 and G19224);
	G21869<= not (G18319 and G19216 and G19226);
	G21870<= not (G18497 and G19223 and G19231);
	G21871<= not (G18458 and G19225 and G19232);
	G21873<= not (G18395 and G19227 and G19234);
	G21874<= not (G18561 and G19233 and G19244);
	G21875<= not (G18531 and G19235 and G19245);
	G21877<= not (G18611 and G19246 and G19257);
	G21879<= not (G18419 and G19250 and G19263);
	G21881<= not (G18492 and G19264 and G19278);
	G21885<= not (G18556 and G19279 and G19297);
	G21888<= not (G18606 and G19298 and G19315);
	G21903<= not (G20008 and G3013);
	G21976<= not (G19242 and G21120 and G19275);
	G21983<= not (G19255 and G21139 and G19294);
	G21989<= not (G21048 and G18623);
	G21991<= not (G21501 and G21536);
	G21996<= not (G19268 and G21159 and G19312);
	G22002<= not (G21065 and G21711);
	G22005<= not (G21540 and G21572);
	G22009<= not (G19283 and G21179 and G19333);
	G22016<= not (G21576 and G21605);
	G22021<= not (G21609 and G21634);
	G22050<= not (G19450 and G21244 and G19503);
	G22069<= not (G19477 and G21253 and G19522);
	G22083<= not (G21774 and G21787);
	G22093<= not (G19500 and G21261 and G19532);
	G22108<= not (G21789 and G21801);
	G22118<= not (G19521 and G21269 and G19542);
	G22134<= not (G21803 and G21809);
	G22157<= not (G21811 and G21816);
	G22188<= not (I28727 and I28728);
	G22197<= not (I28742 and I28743);
	G22203<= not (I28754 and I28755);
	G22209<= not (I28766 and I28767);
	G22317<= not (G21152 and G21241 and G21136);
	G22339<= not (G14442 and G21149 and G10694);
	G22342<= not (G21172 and G21249 and G21156);
	G22362<= not (G14529 and G21169 and G10714);
	G22365<= not (G21192 and G21258 and G21176);
	G22381<= not (G21211 and G14442 and G10694);
	G22382<= not (G14584 and G21189 and G10735);
	G22385<= not (G21207 and G21266 and G21196);
	G22396<= not (G21219 and G14529 and G10714);
	G22397<= not (G14618 and G21204 and G10754);
	G22399<= not (G21230 and G14584 and G10735);
	G22400<= not (G21235 and G14618 and G10754);
	G22608<= not (G20842 and G20885);
	G22644<= not (G20850 and G20904);
	G22668<= not (G16075 and G21271);
	G22680<= not (G20858 and G20928);
	G22708<= not (G16113 and G21278);
	G22720<= not (G20866 and G20956);
	G22739<= not (G16164 and G21285);
	G22771<= not (G16223 and G21293);
	G22809<= not (G21850 and G21848 and G21879);
	G22844<= not (G21865 and G21860 and G21857);
	G22845<= not (G19441 and G20885);
	G22846<= not (G8278 and G21660);
	G22850<= not (G21858 and G21855 and G21881);
	G22876<= not (G21238 and G83);
	G22879<= not (G21870 and G21866 and G21862);
	G22880<= not (G19468 and G20904);
	G22881<= not (G8287 and G21689);
	G22885<= not (G21863 and G21859 and G21885);
	G22911<= not (G21246 and G771);
	G22914<= not (G21874 and G21871 and G21868);
	G22915<= not (G19491 and G20928);
	G22916<= not (G8296 and G21725);
	G22920<= not (G21869 and G21864 and G21888);
	G22936<= not (G21255 and G1457);
	G22939<= not (G21877 and G21875 and G21873);
	G22940<= not (G19512 and G20956);
	G22941<= not (G8305 and G21751);
	G22942<= not (G21263 and G2151);
	G22992<= not (G21636 and G672);
	G23003<= not (G21667 and G1358);
	G23017<= not (G21696 and G2052);
	G23033<= not (G21732 and G2746);
	G23320<= not (G23066 and G23051);
	G23325<= not (G23080 and G23070);
	G23331<= not (G22999 and G22174);
	G23335<= not (G23096 and G23083);
	G23340<= not (G23013 and G22189);
	G23344<= not (G23113 and G23099);
	G23349<= not (G23029 and G22198);
	G23353<= not (G23046 and G22204);
	G23360<= not (G21980 and G21975);
	G23364<= not (G21987 and G21981);
	G23368<= not (G23135 and G22288);
	G23372<= not (G22000 and G21988);
	G23376<= not (G18435 and G22812);
	G23377<= not (G21968 and G22308);
	G23381<= not (G22013 and G22001);
	G23387<= not (G18508 and G22852);
	G23388<= not (G21971 and G22336);
	G23394<= not (G18572 and G22887);
	G23395<= not (G21973 and G22361);
	G23402<= not (G18622 and G22922);
	G23478<= not (G22809 and G14442 and G10694);
	G23486<= not (G22844 and G14442 and G10694);
	G23489<= not (G22850 and G14529 and G10714);
	G23495<= not (G10694 and G14442 and G22316);
	G23502<= not (G22879 and G14529 and G10714);
	G23505<= not (G22885 and G14584 and G10735);
	G23511<= not (G10714 and G14529 and G22341);
	G23518<= not (G22914 and G14584 and G10735);
	G23521<= not (G22920 and G14618 and G10754);
	G23526<= not (G10735 and G14584 and G22364);
	G23533<= not (G22939 and G14618 and G10754);
	G23537<= not (G10754 and G14618 and G22384);
	G23660<= not (I30791 and I30792);
	G23710<= not (I30869 and I30870);
	G23764<= not (I30953 and I30954);
	G23819<= not (I31036 and I31037);
	G23906<= not (G22812 and G13958);
	G23936<= not (G22812 and G13922);
	G23937<= not (G22812 and G13918);
	G23938<= not (G22852 and G14028);
	G23953<= not (G22812 and G14525);
	G23968<= not (G22852 and G13978);
	G23969<= not (G22852 and G13974);
	G23970<= not (G22887 and G14119);
	G23973<= not (G22812 and G14450);
	G23982<= not (G22852 and G14580);
	G23997<= not (G22887 and G14048);
	G23998<= not (G22887 and G14044);
	G23999<= not (G22922 and G14234);
	G24002<= not (G22812 and G14355);
	G24003<= not (G22852 and G14537);
	G24012<= not (G22887 and G14614);
	G24027<= not (G22922 and G14139);
	G24028<= not (G22922 and G14135);
	G24034<= not (G22812 and G14252);
	G24036<= not (G22852 and G14467);
	G24037<= not (G22887 and G14592);
	G24046<= not (G22922 and G14637);
	G24052<= not (G22812 and G14171);
	G24054<= not (G22852 and G14374);
	G24056<= not (G22887 and G14554);
	G24057<= not (G22922 and G14626);
	G24058<= not (G22812 and G14086);
	G24065<= not (G22852 and G14286);
	G24067<= not (G22887 and G14486);
	G24069<= not (G22922 and G14609);
	G24070<= not (G22812 and G14011);
	G24071<= not (G22852 and G14201);
	G24078<= not (G22887 and G14408);
	G24080<= not (G22922 and G14573);
	G24081<= not (G22852 and G14102);
	G24082<= not (G22887 and G14316);
	G24089<= not (G22922 and G14520);
	G24090<= not (G22887 and G14217);
	G24091<= not (G22922 and G14438);
	G24093<= not (G22922 and G14332);
	G24100<= not (G20885 and G22175);
	G24109<= not (G20904 and G22190);
	G24126<= not (G20928 and G22199);
	G24145<= not (G20956 and G22205);
	G24442<= not (G23644 and G3306);
	G24443<= not (G23644 and G3306);
	G24444<= not (G23694 and G3462);
	G24447<= not (G23644 and G3306);
	G24448<= not (G23923 and G3338);
	G24449<= not (G23694 and G3462);
	G24450<= not (G23748 and G3618);
	G24451<= not (G23644 and G3306);
	G24452<= not (G23923 and G3338);
	G24453<= not (G23694 and G3462);
	G24454<= not (G23955 and G3494);
	G24455<= not (G23748 and G3618);
	G24456<= not (G23803 and G3774);
	G24457<= not (G23923 and G3338);
	G24458<= not (G23694 and G3462);
	G24459<= not (G23955 and G3494);
	G24460<= not (G23748 and G3618);
	G24461<= not (G23984 and G3650);
	G24462<= not (G23803 and G3774);
	G24463<= not (G23923 and G3338);
	G24464<= not (G23955 and G3494);
	G24465<= not (G23748 and G3618);
	G24466<= not (G23984 and G3650);
	G24467<= not (G23803 and G3774);
	G24468<= not (G24014 and G3806);
	G24469<= not (G23955 and G3494);
	G24470<= not (G23984 and G3650);
	G24471<= not (G23803 and G3774);
	G24472<= not (G24014 and G3806);
	G24474<= not (G23984 and G3650);
	G24475<= not (G24014 and G3806);
	G24477<= not (G24014 and G3806);
	G24616<= not (G499 and G23376);
	G24627<= not (G1186 and G23387);
	G24641<= not (G1880 and G23394);
	G24660<= not (G2574 and G23402);
	G24753<= not (I32266 and I32267);
	G24766<= not (I32285 and I32286);
	G24771<= not (I32296 and I32297);
	G24778<= not (I32309 and I32310);
	G24787<= not (I32324 and I32325);
	G24791<= not (I32334 and I32335);
	G24797<= not (I32346 and I32347);
	G24801<= not (I32356 and I32357);
	G24808<= not (I32369 and I32370);
	G24812<= not (I32379 and I32380);
	G24814<= not (G24239 and G24244);
	G24817<= not (I32392 and I32393);
	G24820<= not (I32401 and I32402);
	G24823<= not (I32410 and I32411);
	G24830<= not (I32423 and I32424);
	G24832<= not (I32431 and I32432);
	G24833<= not (G24245 and G24252);
	G24837<= not (I32444 and I32445);
	G24839<= not (I32452 and I32453);
	G24842<= not (I32461 and I32462);
	G24844<= not (I32469 and I32470);
	G24848<= not (I32479 and I32480);
	G24849<= not (G24254 and G24257);
	G24852<= not (I32491 and I32492);
	G24854<= not (I32499 and I32500);
	G24857<= not (I32510 and I32511);
	G24860<= not (I32519 and I32520);
	G24862<= not (I32527 and I32528);
	G24863<= not (G24258 and G23319);
	G24866<= not (I32539 and I32540);
	G24868<= not (I32547 and I32548);
	G24873<= not (I32560 and I32561);
	G24875<= not (I32568 and I32569);
	G24877<= not (I32576 and I32577);
	G24880<= not (I32587 and I32588);
	G24883<= not (I32596 and I32597);
	G24887<= not (I32608 and I32609);
	G24889<= not (I32616 and I32617);
	G24897<= not (I32625 and I32626);
	G24900<= not (I32634 and I32635);
	G24904<= not (I32646 and I32647);
	G24920<= not (I32660 and I32661);
	G24923<= not (I32669 and I32670);
	G24928<= not (I32678 and I32679);
	G24937<= not (I32687 and I32688);
	G24940<= not (I32696 and I32697);
	G24951<= not (I32709 and I32710);
	G24963<= not (I32725 and I32726);
	G24975<= not (G23497 and G74);
	G24986<= not (G23513 and G762);
	G24997<= not (G23528 and G1448);
	G25004<= not (G23644 and G6448);
	G25005<= not (G23539 and G2142);
	G25008<= not (G23644 and G5438);
	G25009<= not (G23644 and G6448);
	G25010<= not (G23694 and G6713);
	G25011<= not (G23644 and G5438);
	G25012<= not (G23644 and G6448);
	G25013<= not (G23923 and G6643);
	G25014<= not (G23694 and G5473);
	G25015<= not (G23694 and G6713);
	G25016<= not (G23748 and G7015);
	G25017<= not (G23644 and G5438);
	G25018<= not (G23644 and G6448);
	G25019<= not (G23923 and G6486);
	G25020<= not (G23923 and G6643);
	G25021<= not (G23694 and G5473);
	G25022<= not (G23694 and G6713);
	G25023<= not (G23955 and G6945);
	G25024<= not (G23748 and G5512);
	G25025<= not (G23748 and G7015);
	G25026<= not (G23803 and G7265);
	G25028<= not (G23644 and G5438);
	G25029<= not (G23923 and G6486);
	G25030<= not (G23923 and G6643);
	G25031<= not (G23694 and G5473);
	G25032<= not (G23694 and G6713);
	G25033<= not (G23955 and G6751);
	G25034<= not (G23955 and G6945);
	G25035<= not (G23748 and G5512);
	G25036<= not (G23748 and G7015);
	G25037<= not (G23984 and G7195);
	G25038<= not (G23803 and G5556);
	G25039<= not (G23803 and G7265);
	G25040<= not (G23923 and G6486);
	G25041<= not (G23923 and G6643);
	G25043<= not (G23694 and G5473);
	G25044<= not (G23955 and G6751);
	G25045<= not (G23955 and G6945);
	G25046<= not (G23748 and G5512);
	G25047<= not (G23748 and G7015);
	G25048<= not (G23984 and G7053);
	G25049<= not (G23984 and G7195);
	G25050<= not (G23803 and G5556);
	G25051<= not (G23803 and G7265);
	G25052<= not (G24014 and G7391);
	G25053<= not (G23923 and G6486);
	G25054<= not (G23955 and G6751);
	G25055<= not (G23955 and G6945);
	G25057<= not (G23748 and G5512);
	G25058<= not (G23984 and G7053);
	G25059<= not (G23984 and G7195);
	G25060<= not (G23803 and G5556);
	G25061<= not (G23803 and G7265);
	G25062<= not (G24014 and G7303);
	G25063<= not (G24014 and G7391);
	G25064<= not (G23955 and G6751);
	G25065<= not (G23984 and G7053);
	G25066<= not (G23984 and G7195);
	G25068<= not (G23803 and G5556);
	G25069<= not (G24014 and G7303);
	G25070<= not (G24014 and G7391);
	G25071<= not (G23984 and G7053);
	G25072<= not (G24014 and G7303);
	G25073<= not (G24014 and G7391);
	G25074<= not (G24014 and G7303);
	G25088<= not (G23950 and G679);
	G25096<= not (G23979 and G1365);
	G25106<= not (G24009 and G2059);
	G25112<= not (G24043 and G2753);
	G25200<= not (G24965 and G3306);
	G25203<= not (G24978 and G3462);
	G25205<= not (G24989 and G3618);
	G25210<= not (G25000 and G3774);
	G25312<= not (G21211 and G14442 and G10694 and G24590);
	G25320<= not (G21219 and G14529 and G10714 and G24595);
	G25331<= not (G21230 and G14584 and G10735 and G24603);
	G25340<= not (G21235 and G14618 and G10754 and G24610);
	G25927<= not (G24965 and G6448);
	G25928<= not (G24965 and G5438);
	G25929<= not (G24978 and G6713);
	G25930<= not (G24978 and G5473);
	G25931<= not (G24989 and G7015);
	G25933<= not (G24989 and G5512);
	G25934<= not (G25000 and G7265);
	G25936<= not (G25000 and G5556);
	G25954<= not (G22806 and G24517);
	G25958<= not (G22847 and G24530);
	G25964<= not (G22882 and G24543);
	G25969<= not (G22917 and G24555);
	G26059<= not (G25422 and G25379 and G25274);
	G26066<= not (G25431 and G25395 and G25283);
	G26073<= not (G25438 and G25405 and G25291);
	G26079<= not (G25445 and G25413 and G25301);
	G26106<= not (G23644 and G25354);
	G26119<= not (G8278 and G14657 and G25422 and G25379);
	G26120<= not (G23694 and G25369);
	G26129<= not (G8287 and G14691 and G25431 and G25395);
	G26130<= not (G23748 and G25386);
	G26143<= not (G8296 and G14725 and G25438 and G25405);
	G26144<= not (G23803 and G25402);
	G26148<= not (G8305 and G14753 and G25445 and G25413);
	G26356<= not (G16539 and G25183);
	G26399<= not (G16571 and G25186);
	G26440<= not (G16595 and G25190);
	G26458<= not (G25343 and G65);
	G26472<= not (G16615 and G25195);
	G26482<= not (G25357 and G753);
	G26498<= not (G25372 and G1439);
	G26513<= not (G25389 and G2133);
	G26772<= not (G26320 and G3306);
	G26779<= not (G26367 and G3462);
	G26785<= not (G26410 and G3618);
	G26792<= not (G26451 and G3774);
	G26859<= not (I35021 and I35022);
	G26865<= not (I35035 and I35036);
	G26867<= not (I35043 and I35044);
	G26874<= not (I35058 and I35059);
	G26892<= not (G25699 and G26283 and G25569 and G25631);
	G26902<= not (G25631 and G26283 and G25569);
	G26906<= not (G25772 and G26327 and G25648 and G25708);
	G26911<= not (G25569 and G26283);
	G26915<= not (G25708 and G26327 and G25648);
	G26918<= not (G25826 and G26374 and G25725 and G25781);
	G26925<= not (G25648 and G26327);
	G26928<= not (G25781 and G26374 and G25725);
	G26931<= not (G25861 and G26417 and G25798 and G25835);
	G26934<= not (I35124 and I35125);
	G26938<= not (G25725 and G26374);
	G26941<= not (G25835 and G26417 and G25798);
	G26947<= not (G25798 and G26417);
	G27117<= not (G26320 and G6448);
	G27118<= not (G26320 and G5438);
	G27119<= not (G26367 and G6713);
	G27121<= not (G26367 and G5473);
	G27122<= not (G26410 and G7015);
	G27124<= not (G26410 and G5512);
	G27125<= not (G26451 and G7265);
	G27130<= not (G26451 and G5556);
	G27379<= not (I35702 and I35703);
	G27382<= not (I35715 and I35716);
	G27390<= not (G26989 and G6448);
	G27395<= not (G26989 and G5438);
	G27400<= not (G27012 and G6713);
	G27408<= not (G27012 and G5473);
	G27413<= not (G27038 and G7015);
	G27426<= not (G27038 and G5512);
	G27431<= not (G27066 and G7265);
	G27447<= not (G27066 and G5556);
	G27528<= not (I35905 and I35906);
	G27550<= not (I35945 and I35946);
	G27566<= not (I35975 and I35976);
	G27571<= not (G26869 and G56);
	G27576<= not (I35993 and I35994);
	G27580<= not (G26878 and G744);
	G27583<= not (G26887 and G1430);
	G27587<= not (G26897 and G2124);
	G27626<= not (G26989 and G3306);
	G27627<= not (G27012 and G3462);
	G27628<= not (G27038 and G3618);
	G27630<= not (G27066 and G3774);
	G27738<= not (G25367 and G27415);
	G27743<= not (G25384 and G27436);
	G27751<= not (G25400 and G27455);
	G27756<= not (G25410 and G27471);
	G27801<= not (I36257 and I36258);
	G27809<= not (I36271 and I36272);
	G27830<= not (I36290 and I36291);
	G27838<= not (I36301 and I36302);
	G27846<= not (I36315 and I36316);
	G28046<= not (I36592 and I36593);
	G28075<= not (I36667 and I36668);
	G28100<= not (I36732 and I36733);
	G28118<= not (I36780 and I36781);
	G28384<= not (I37296 and I37297);
	G28386<= not (I37304 and I37305);
	G28388<= not (I37312 and I37313);
	G28391<= not (I37323 and I37324);
	G28415<= not (I37357 and I37358);
	G28842<= not (I37814 and I37815);
	G28845<= not (I37823 and I37824);
	G28978<= not (G9150 and G28512);
	G29001<= not (G9161 and G28512);
	G29008<= not (G9174 and G28540);
	G29026<= not (G9187 and G28512);
	G29030<= not (G9203 and G28540);
	G29038<= not (G9216 and G28567);
	G29045<= not (G9232 and G28512);
	G29049<= not (G9248 and G28540);
	G29053<= not (G9264 and G28567);
	G29060<= not (G9277 and G28595);
	G29062<= not (G9310 and G28540);
	G29068<= not (G9326 and G28567);
	G29072<= not (G9342 and G28595);
	G29076<= not (G9391 and G28567);
	G29080<= not (G9407 and G28595);
	G29087<= not (G9488 and G28595);
	G29088<= not (G9507 and G28512);
	G29096<= not (G9649 and G28540);
	G29103<= not (G9795 and G28567);
	G29107<= not (G9941 and G28595);
	G29265<= not (I38379 and I38380);
	G29498<= not (I38811 and I38812);
	G29500<= not (I38821 and I38822);
	G29503<= not (I38832 and I38833);
	G29505<= not (I38842 and I38843);
	G29911<= not (I39324 and I39325);
	G29913<= not (I39332 and I39333);
	G29915<= not (I39340 and I39341);
	G29917<= not (I39348 and I39349);
	G29923<= not (I39360 and I39361);
	G29925<= not (I39368 and I39369);
	G29927<= not (I39376 and I39377);
	G29930<= not (I39385 and I39386);
	G29931<= not (I39392 and I39393);
	G30034<= not (I39533 and I39534);
	G30035<= not (I39540 and I39541);
	G30228<= not (I39690 and I39691);
	G30768<= not (I40559 and I40560);
	G30771<= not (I40572 and I40573);
	G30775<= not (I40588 and I40589);
	G30779<= not (I40604 and I40605);
	G30791<= not (I40628 and I40629);
	G30926<= not (I41011 and I41012);
	G30927<= not (I41018 and I41019);
	G30952<= not (I41065 and I41066);
	I15167<= not (G2981 and G2874);
	I15168<= not (G2981 and I15167);
	I15169<= not (G2874 and I15167);
	I15183<= not (G2975 and G2978);
	I15184<= not (G2975 and I15183);
	I15185<= not (G2978 and I15183);
	I15190<= not (G2956 and G2959);
	I15191<= not (G2956 and I15190);
	I15192<= not (G2959 and I15190);
	I15204<= not (G2969 and G2972);
	I15205<= not (G2969 and I15204);
	I15206<= not (G2972 and I15204);
	I15211<= not (G2947 and G2953);
	I15212<= not (G2947 and I15211);
	I15213<= not (G2953 and I15211);
	I15237<= not (G2963 and G2966);
	I15238<= not (G2963 and I15237);
	I15239<= not (G2966 and I15237);
	I15244<= not (G2941 and G2944);
	I15245<= not (G2941 and I15244);
	I15246<= not (G2944 and I15244);
	I15276<= not (G2935 and G2938);
	I15277<= not (G2935 and I15276);
	I15278<= not (G2938 and I15276);
	I16879<= not (G4203 and G3998);
	I16880<= not (G4203 and I16879);
	I16881<= not (G3998 and I16879);
	I16965<= not (G4734 and G4452);
	I16966<= not (G4734 and I16965);
	I16967<= not (G4452 and I16965);
	I17059<= not (G6637 and G6309);
	I17060<= not (G6637 and I17059);
	I17061<= not (G6309 and I17059);
	I17149<= not (G7465 and G7142);
	I17150<= not (G7465 and I17149);
	I17151<= not (G7142 and I17149);
	I18106<= not (G7875 and G7855);
	I18107<= not (G7875 and I18106);
	I18108<= not (G7855 and I18106);
	I18113<= not (G3997 and G8181);
	I18114<= not (G3997 and I18113);
	I18115<= not (G8181 and I18113);
	I18190<= not (G7922 and G7895);
	I18191<= not (G7922 and I18190);
	I18192<= not (G7895 and I18190);
	I18197<= not (G7896 and G7876);
	I18198<= not (G7896 and I18197);
	I18199<= not (G7876 and I18197);
	I18204<= not (G7975 and G4202);
	I18205<= not (G7975 and I18204);
	I18206<= not (G4202 and I18204);
	I18280<= not (G7970 and G7923);
	I18281<= not (G7970 and I18280);
	I18282<= not (G7923 and I18280);
	I18287<= not (G8256 and G8102);
	I18288<= not (G8256 and I18287);
	I18289<= not (G8102 and I18287);
	I18368<= not (G4325 and G4093);
	I18369<= not (G4325 and I18368);
	I18370<= not (G4093 and I18368);
	I18799<= not (G11410 and G11331);
	I18800<= not (G11410 and I18799);
	I18801<= not (G11331 and I18799);
	I20031<= not (G10003 and G9883);
	I20032<= not (G10003 and I20031);
	I20033<= not (G9883 and I20031);
	I20048<= not (G10185 and G10095);
	I20049<= not (G10185 and I20048);
	I20050<= not (G10095 and I20048);
	I20429<= not (G11262 and G11188);
	I20430<= not (G11262 and I20429);
	I20431<= not (G11188 and I20429);
	I20465<= not (G11330 and G11263);
	I20466<= not (G11330 and I20465);
	I20467<= not (G11263 and I20465);
	I20504<= not (G11264 and G11189);
	I20505<= not (G11264 and I20504);
	I20506<= not (G11189 and I20504);
	I20743<= not (G11621 and G13399);
	I20744<= not (G11621 and I20743);
	I20745<= not (G13399 and I20743);
	I22062<= not (G12999 and G12988);
	I22063<= not (G12999 and I22062);
	I22064<= not (G12988 and I22062);
	I22282<= not (G2962 and G13348);
	I22283<= not (G2962 and I22282);
	I22284<= not (G13348 and I22282);
	I22316<= not (G2934 and G13370);
	I22317<= not (G2934 and I22316);
	I22318<= not (G13370 and I22316);
	I22630<= not (G13507 and G15978);
	I22631<= not (G13507 and I22630);
	I22632<= not (G15978 and I22630);
	I22705<= not (G13348 and G15661);
	I22706<= not (G13348 and I22705);
	I22707<= not (G15661 and I22705);
	I22884<= not (G13370 and G15661);
	I22885<= not (G13370 and I22884);
	I22886<= not (G15661 and I22884);
	I22900<= not (G15022 and G14000);
	I22901<= not (G15022 and I22900);
	I22902<= not (G14000 and I22900);
	I22917<= not (G15096 and G13945);
	I22918<= not (G15096 and I22917);
	I22919<= not (G13945 and I22917);
	I22924<= not (G15118 and G14091);
	I22925<= not (G15118 and I22924);
	I22926<= not (G14091 and I22924);
	I22936<= not (G9150 and G13906);
	I22937<= not (G9150 and I22936);
	I22938<= not (G13906 and I22936);
	I22945<= not (G15188 and G14015);
	I22946<= not (G15188 and I22945);
	I22947<= not (G14015 and I22945);
	I22952<= not (G15210 and G14206);
	I22953<= not (G15210 and I22952);
	I22954<= not (G14206 and I22952);
	I22962<= not (G9161 and G13885);
	I22963<= not (G9161 and I22962);
	I22964<= not (G13885 and I22962);
	I22972<= not (G9174 and G13962);
	I22973<= not (G9174 and I22972);
	I22974<= not (G13962 and I22972);
	I22981<= not (G15274 and G14106);
	I22982<= not (G15274 and I22981);
	I22983<= not (G14106 and I22981);
	I22988<= not (G15296 and G14321);
	I22989<= not (G15296 and I22988);
	I22990<= not (G14321 and I22988);
	I22998<= not (G9187 and G13872);
	I22999<= not (G9187 and I22998);
	I23000<= not (G13872 and I22998);
	I23008<= not (G9203 and G13926);
	I23009<= not (G9203 and I23008);
	I23010<= not (G13926 and I23008);
	I23018<= not (G9216 and G14032);
	I23019<= not (G9216 and I23018);
	I23020<= not (G14032 and I23018);
	I23027<= not (G15366 and G14221);
	I23028<= not (G15366 and I23027);
	I23029<= not (G14221 and I23027);
	I23034<= not (G9232 and G13864);
	I23035<= not (G9232 and I23034);
	I23036<= not (G13864 and I23034);
	I23045<= not (G9248 and G13894);
	I23046<= not (G9248 and I23045);
	I23047<= not (G13894 and I23045);
	I23055<= not (G9264 and G13982);
	I23056<= not (G9264 and I23055);
	I23057<= not (G13982 and I23055);
	I23065<= not (G9277 and G14123);
	I23066<= not (G9277 and I23065);
	I23067<= not (G14123 and I23065);
	I23074<= not (G9293 and G13856);
	I23075<= not (G9293 and I23074);
	I23076<= not (G13856 and I23074);
	I23082<= not (G9310 and G13879);
	I23083<= not (G9310 and I23082);
	I23084<= not (G13879 and I23082);
	I23093<= not (G9326 and G13935);
	I23094<= not (G9326 and I23093);
	I23095<= not (G13935 and I23093);
	I23103<= not (G9342 and G14052);
	I23104<= not (G9342 and I23103);
	I23105<= not (G14052 and I23103);
	I23113<= not (G9356 and G13848);
	I23114<= not (G9356 and I23113);
	I23115<= not (G13848 and I23113);
	I23123<= not (G9374 and G13866);
	I23124<= not (G9374 and I23123);
	I23125<= not (G13866 and I23123);
	I23131<= not (G9391 and G13901);
	I23132<= not (G9391 and I23131);
	I23133<= not (G13901 and I23131);
	I23142<= not (G9407 and G13991);
	I23143<= not (G9407 and I23142);
	I23144<= not (G13991 and I23142);
	I23152<= not (G9427 and G14061);
	I23153<= not (G9427 and I23152);
	I23154<= not (G14061 and I23152);
	I23161<= not (G9453 and G13857);
	I23162<= not (G9453 and I23161);
	I23163<= not (G13857 and I23161);
	I23171<= not (G9471 and G13881);
	I23172<= not (G9471 and I23171);
	I23173<= not (G13881 and I23171);
	I23179<= not (G9488 and G13942);
	I23180<= not (G9488 and I23179);
	I23181<= not (G13942 and I23179);
	I23190<= not (G9507 and G13999);
	I23191<= not (G9507 and I23190);
	I23192<= not (G13999 and I23190);
	I23198<= not (G9569 and G14176);
	I23199<= not (G9569 and I23198);
	I23200<= not (G14176 and I23198);
	I23207<= not (G9595 and G13867);
	I23208<= not (G9595 and I23207);
	I23209<= not (G13867 and I23207);
	I23217<= not (G9613 and G13903);
	I23218<= not (G9613 and I23217);
	I23219<= not (G13903 and I23217);
	I23225<= not (G9649 and G14090);
	I23226<= not (G9649 and I23225);
	I23227<= not (G14090 and I23225);
	I23233<= not (G9711 and G14291);
	I23234<= not (G9711 and I23233);
	I23235<= not (G14291 and I23233);
	I23242<= not (G9737 and G13882);
	I23243<= not (G9737 and I23242);
	I23244<= not (G13882 and I23242);
	I23256<= not (G9795 and G14205);
	I23257<= not (G9795 and I23256);
	I23258<= not (G14205 and I23256);
	I23264<= not (G9857 and G14413);
	I23265<= not (G9857 and I23264);
	I23266<= not (G14413 and I23264);
	I23277<= not (G9941 and G14320);
	I23278<= not (G9941 and I23277);
	I23279<= not (G14320 and I23277);
	I23806<= not (G14062 and G9150);
	I23807<= not (G14062 and I23806);
	I23808<= not (G9150 and I23806);
	I23878<= not (G14001 and G9187);
	I23879<= not (G14001 and I23878);
	I23880<= not (G9187 and I23878);
	I23893<= not (G14177 and G9174);
	I23894<= not (G14177 and I23893);
	I23895<= not (G9174 and I23893);
	I23941<= not (G13946 and G9293);
	I23942<= not (G13946 and I23941);
	I23943<= not (G9293 and I23941);
	I23958<= not (G6513 and G14171);
	I23959<= not (G6513 and I23958);
	I23960<= not (G14171 and I23958);
	I23966<= not (G14092 and G9248);
	I23967<= not (G14092 and I23966);
	I23968<= not (G9248 and I23966);
	I23981<= not (G14292 and G9216);
	I23982<= not (G14292 and I23981);
	I23983<= not (G9216 and I23981);
	I24005<= not (G7548 and G15814);
	I24006<= not (G7548 and I24005);
	I24007<= not (G15814 and I24005);
	I24015<= not (G13907 and G9427);
	I24016<= not (G13907 and I24015);
	I24017<= not (G9427 and I24015);
	I24028<= not (G6201 and G14086);
	I24029<= not (G6201 and I24028);
	I24030<= not (G14086 and I24028);
	I24036<= not (G14016 and G9374);
	I24037<= not (G14016 and I24036);
	I24038<= not (G9374 and I24036);
	I24053<= not (G6777 and G14286);
	I24054<= not (G6777 and I24053);
	I24055<= not (G14286 and I24053);
	I24061<= not (G14207 and G9326);
	I24062<= not (G14207 and I24061);
	I24063<= not (G9326 and I24061);
	I24076<= not (G14414 and G9277);
	I24077<= not (G14414 and I24076);
	I24078<= not (G9277 and I24076);
	I24091<= not (G13886 and G15096);
	I24092<= not (G13886 and I24091);
	I24093<= not (G15096 and I24091);
	I24102<= not (G6363 and G14011);
	I24103<= not (G6363 and I24102);
	I24104<= not (G14011 and I24102);
	I24110<= not (G13963 and G9569);
	I24111<= not (G13963 and I24110);
	I24112<= not (G9569 and I24110);
	I24123<= not (G6290 and G14201);
	I24124<= not (G6290 and I24123);
	I24125<= not (G14201 and I24123);
	I24131<= not (G14107 and G9471);
	I24132<= not (G14107 and I24131);
	I24133<= not (G9471 and I24131);
	I24148<= not (G7079 and G14408);
	I24149<= not (G7079 and I24148);
	I24150<= not (G14408 and I24148);
	I24156<= not (G14322 and G9407);
	I24157<= not (G14322 and I24156);
	I24158<= not (G9407 and I24156);
	I24178<= not (G13873 and G9161);
	I24179<= not (G13873 and I24178);
	I24180<= not (G9161 and I24178);
	I24186<= not (G6177 and G13958);
	I24187<= not (G6177 and I24186);
	I24188<= not (G13958 and I24186);
	I24194<= not (G13927 and G15188);
	I24195<= not (G13927 and I24194);
	I24196<= not (G15188 and I24194);
	I24205<= not (G6568 and G14102);
	I24206<= not (G6568 and I24205);
	I24207<= not (G14102 and I24205);
	I24213<= not (G14033 and G9711);
	I24214<= not (G14033 and I24213);
	I24215<= not (G9711 and I24213);
	I24226<= not (G6427 and G14316);
	I24227<= not (G6427 and I24226);
	I24228<= not (G14316 and I24226);
	I24234<= not (G14222 and G9613);
	I24235<= not (G14222 and I24234);
	I24236<= not (G9613 and I24234);
	I24251<= not (G7329 and G14520);
	I24252<= not (G7329 and I24251);
	I24253<= not (G14520 and I24251);
	I24263<= not (G14342 and G9232);
	I24264<= not (G14342 and I24263);
	I24265<= not (G9232 and I24263);
	I24271<= not (G6180 and G13922);
	I24272<= not (G6180 and I24271);
	I24273<= not (G13922 and I24271);
	I24278<= not (G6284 and G13918);
	I24279<= not (G6284 and I24278);
	I24280<= not (G13918 and I24278);
	I24290<= not (G13895 and G9203);
	I24291<= not (G13895 and I24290);
	I24292<= not (G9203 and I24290);
	I24298<= not (G6209 and G14028);
	I24299<= not (G6209 and I24298);
	I24300<= not (G14028 and I24298);
	I24306<= not (G13983 and G15274);
	I24307<= not (G13983 and I24306);
	I24308<= not (G15274 and I24306);
	I24317<= not (G6832 and G14217);
	I24318<= not (G6832 and I24317);
	I24319<= not (G14217 and I24317);
	I24325<= not (G14124 and G9857);
	I24326<= not (G14124 and I24325);
	I24327<= not (G9857 and I24325);
	I24338<= not (G6632 and G14438);
	I24339<= not (G6632 and I24338);
	I24340<= not (G14438 and I24338);
	I24351<= not (G14238 and G9356);
	I24352<= not (G14238 and I24351);
	I24353<= not (G9356 and I24351);
	I24361<= not (G6157 and G14525);
	I24362<= not (G6157 and I24361);
	I24363<= not (G14525 and I24361);
	I24372<= not (G14454 and G9310);
	I24373<= not (G14454 and I24372);
	I24374<= not (G9310 and I24372);
	I24380<= not (G6212 and G13978);
	I24381<= not (G6212 and I24380);
	I24382<= not (G13978 and I24380);
	I24387<= not (G6421 and G13974);
	I24388<= not (G6421 and I24387);
	I24389<= not (G13974 and I24387);
	I24399<= not (G13936 and G9264);
	I24400<= not (G13936 and I24399);
	I24401<= not (G9264 and I24399);
	I24407<= not (G6298 and G14119);
	I24408<= not (G6298 and I24407);
	I24409<= not (G14119 and I24407);
	I24415<= not (G14053 and G15366);
	I24416<= not (G14053 and I24415);
	I24417<= not (G15366 and I24415);
	I24426<= not (G7134 and G14332);
	I24427<= not (G7134 and I24426);
	I24428<= not (G14332 and I24426);
	I24436<= not (G14153 and G15022);
	I24437<= not (G14153 and I24436);
	I24438<= not (G15022 and I24436);
	I24443<= not (G14148 and G9507);
	I24444<= not (G14148 and I24443);
	I24445<= not (G9507 and I24443);
	I24452<= not (G6142 and G14450);
	I24453<= not (G6142 and I24452);
	I24454<= not (G14450 and I24452);
	I24464<= not (G14360 and G9453);
	I24465<= not (G14360 and I24464);
	I24466<= not (G9453 and I24464);
	I24474<= not (G6184 and G14580);
	I24475<= not (G6184 and I24474);
	I24476<= not (G14580 and I24474);
	I24485<= not (G14541 and G9391);
	I24486<= not (G14541 and I24485);
	I24487<= not (G9391 and I24485);
	I24493<= not (G6301 and G14048);
	I24494<= not (G6301 and I24493);
	I24495<= not (G14048 and I24493);
	I24500<= not (G6626 and G14044);
	I24501<= not (G6626 and I24500);
	I24502<= not (G14044 and I24500);
	I24512<= not (G13992 and G9342);
	I24513<= not (G13992 and I24512);
	I24514<= not (G9342 and I24512);
	I24520<= not (G6435 and G14234);
	I24521<= not (G6435 and I24520);
	I24522<= not (G14234 and I24520);
	I24530<= not (G6707 and G14355);
	I24531<= not (G6707 and I24530);
	I24532<= not (G14355 and I24530);
	I24537<= not (G14268 and G15118);
	I24538<= not (G14268 and I24537);
	I24539<= not (G15118 and I24537);
	I24544<= not (G14263 and G9649);
	I24545<= not (G14263 and I24544);
	I24546<= not (G9649 and I24544);
	I24553<= not (G6163 and G14537);
	I24554<= not (G6163 and I24553);
	I24555<= not (G14537 and I24553);
	I24565<= not (G14472 and G9595);
	I24566<= not (G14472 and I24565);
	I24567<= not (G9595 and I24565);
	I24575<= not (G6216 and G14614);
	I24576<= not (G6216 and I24575);
	I24577<= not (G14614 and I24575);
	I24586<= not (G14596 and G9488);
	I24587<= not (G14596 and I24586);
	I24588<= not (G9488 and I24586);
	I24594<= not (G6438 and G14139);
	I24595<= not (G6438 and I24594);
	I24596<= not (G14139 and I24594);
	I24601<= not (G6890 and G14135);
	I24602<= not (G6890 and I24601);
	I24603<= not (G14135 and I24601);
	I24611<= not (G15814 and G15978);
	I24612<= not (G15814 and I24611);
	I24613<= not (G15978 and I24611);
	I24624<= not (G6136 and G14252);
	I24625<= not (G6136 and I24624);
	I24626<= not (G14252 and I24624);
	I24632<= not (G7009 and G14467);
	I24633<= not (G7009 and I24632);
	I24634<= not (G14467 and I24632);
	I24639<= not (G14390 and G15210);
	I24640<= not (G14390 and I24639);
	I24641<= not (G15210 and I24639);
	I24646<= not (G14385 and G9795);
	I24647<= not (G14385 and I24646);
	I24648<= not (G9795 and I24646);
	I24655<= not (G6190 and G14592);
	I24656<= not (G6190 and I24655);
	I24657<= not (G14592 and I24655);
	I24667<= not (G14559 and G9737);
	I24668<= not (G14559 and I24667);
	I24669<= not (G9737 and I24667);
	I24677<= not (G6305 and G14637);
	I24678<= not (G6305 and I24677);
	I24679<= not (G14637 and I24677);
	I24694<= not (G6146 and G14374);
	I24695<= not (G6146 and I24694);
	I24696<= not (G14374 and I24694);
	I24702<= not (G7259 and G14554);
	I24703<= not (G7259 and I24702);
	I24704<= not (G14554 and I24702);
	I24709<= not (G14502 and G15296);
	I24710<= not (G14502 and I24709);
	I24711<= not (G15296 and I24709);
	I24716<= not (G14497 and G9941);
	I24717<= not (G14497 and I24716);
	I24718<= not (G9941 and I24716);
	I24725<= not (G6222 and G14626);
	I24726<= not (G6222 and I24725);
	I24727<= not (G14626 and I24725);
	I24743<= not (G6167 and G14486);
	I24744<= not (G6167 and I24743);
	I24745<= not (G14486 and I24743);
	I24751<= not (G7455 and G14609);
	I24752<= not (G7455 and I24751);
	I24753<= not (G14609 and I24751);
	I24763<= not (G6194 and G14573);
	I24764<= not (G6194 and I24763);
	I24765<= not (G14573 and I24763);
	I25030<= not (G8029 and G13507);
	I25031<= not (G8029 and I25030);
	I25032<= not (G13507 and I25030);
	I25532<= not (G52 and G18179);
	I25533<= not (G52 and I25532);
	I25534<= not (G18179 and I25532);
	I25539<= not (G92 and G18174);
	I25540<= not (G92 and I25539);
	I25541<= not (G18174 and I25539);
	I25560<= not (G56 and G17724);
	I25561<= not (G56 and I25560);
	I25562<= not (G17724 and I25560);
	I25571<= not (G740 and G18286);
	I25572<= not (G740 and I25571);
	I25573<= not (G18286 and I25571);
	I25578<= not (G780 and G18281);
	I25579<= not (G780 and I25578);
	I25580<= not (G18281 and I25578);
	I25595<= not (G61 and G18074);
	I25596<= not (G61 and I25595);
	I25597<= not (G18074 and I25595);
	I25605<= not (G744 and G17825);
	I25606<= not (G744 and I25605);
	I25607<= not (G17825 and I25605);
	I25616<= not (G1426 and G18379);
	I25617<= not (G1426 and I25616);
	I25618<= not (G18379 and I25616);
	I25623<= not (G1466 and G18374);
	I25624<= not (G1466 and I25623);
	I25625<= not (G18374 and I25623);
	I25633<= not (G65 and G17640);
	I25634<= not (G65 and I25633);
	I25635<= not (G17640 and I25633);
	I25643<= not (G749 and G18190);
	I25644<= not (G749 and I25643);
	I25645<= not (G18190 and I25643);
	I25653<= not (G1430 and G17937);
	I25654<= not (G1430 and I25653);
	I25655<= not (G17937 and I25653);
	I25664<= not (G2120 and G18474);
	I25665<= not (G2120 and I25664);
	I25666<= not (G18474 and I25664);
	I25671<= not (G2160 and G18469);
	I25672<= not (G2160 and I25671);
	I25673<= not (G18469 and I25671);
	I25681<= not (G70 and G17974);
	I25682<= not (G70 and I25681);
	I25683<= not (G17974 and I25681);
	I25690<= not (G753 and G17741);
	I25691<= not (G753 and I25690);
	I25692<= not (G17741 and I25690);
	I25700<= not (G1435 and G18297);
	I25701<= not (G1435 and I25700);
	I25702<= not (G18297 and I25700);
	I25710<= not (G2124 and G18048);
	I25711<= not (G2124 and I25710);
	I25712<= not (G18048 and I25710);
	I25721<= not (G74 and G18341);
	I25722<= not (G74 and I25721);
	I25723<= not (G18341 and I25721);
	I25731<= not (G758 and G18091);
	I25732<= not (G758 and I25731);
	I25733<= not (G18091 and I25731);
	I25740<= not (G1439 and G17842);
	I25741<= not (G1439 and I25740);
	I25742<= not (G17842 and I25740);
	I25750<= not (G2129 and G18390);
	I25751<= not (G2129 and I25750);
	I25752<= not (G18390 and I25750);
	I25761<= not (G79 and G17882);
	I25762<= not (G79 and I25761);
	I25763<= not (G17882 and I25761);
	I25771<= not (G762 and G18436);
	I25772<= not (G762 and I25771);
	I25773<= not (G18436 and I25771);
	I25781<= not (G1444 and G18207);
	I25782<= not (G1444 and I25781);
	I25783<= not (G18207 and I25781);
	I25790<= not (G2133 and G17954);
	I25791<= not (G2133 and I25790);
	I25792<= not (G17954 and I25790);
	I25800<= not (G83 and G18265);
	I25801<= not (G83 and I25800);
	I25802<= not (G18265 and I25800);
	I25809<= not (G767 and G17993);
	I25810<= not (G767 and I25809);
	I25811<= not (G17993 and I25809);
	I25819<= not (G1448 and G18509);
	I25820<= not (G1448 and I25819);
	I25821<= not (G18509 and I25819);
	I25829<= not (G2138 and G18314);
	I25830<= not (G2138 and I25829);
	I25831<= not (G18314 and I25829);
	I25838<= not (G88 and G17802);
	I25839<= not (G88 and I25838);
	I25840<= not (G17802 and I25838);
	I25846<= not (G771 and G18358);
	I25847<= not (G771 and I25846);
	I25848<= not (G18358 and I25846);
	I25855<= not (G1453 and G18110);
	I25856<= not (G1453 and I25855);
	I25857<= not (G18110 and I25855);
	I25865<= not (G2142 and G18573);
	I25866<= not (G2142 and I25865);
	I25867<= not (G18573 and I25865);
	I25880<= not (G776 and G17914);
	I25881<= not (G776 and I25880);
	I25882<= not (G17914 and I25880);
	I25888<= not (G1457 and G18453);
	I25889<= not (G1457 and I25888);
	I25890<= not (G18453 and I25888);
	I25897<= not (G2147 and G18226);
	I25898<= not (G2147 and I25897);
	I25899<= not (G18226 and I25897);
	I25913<= not (G1462 and G18025);
	I25914<= not (G1462 and I25913);
	I25915<= not (G18025 and I25913);
	I25921<= not (G2151 and G18526);
	I25922<= not (G2151 and I25921);
	I25923<= not (G18526 and I25921);
	I25938<= not (G2156 and G18142);
	I25939<= not (G2156 and I25938);
	I25940<= not (G18142 and I25938);
	I28189<= not (G14079 and G19444);
	I28190<= not (G14079 and I28189);
	I28191<= not (G19444 and I28189);
	I28217<= not (G14194 and G19471);
	I28218<= not (G14194 and I28217);
	I28219<= not (G19471 and I28217);
	I28247<= not (G14309 and G19494);
	I28248<= not (G14309 and I28247);
	I28249<= not (G19494 and I28247);
	I28271<= not (G14431 and G19515);
	I28272<= not (G14431 and I28271);
	I28273<= not (G19515 and I28271);
	I28726<= not (G21887 and G13519);
	I28727<= not (G21887 and I28726);
	I28728<= not (G13519 and I28726);
	I28741<= not (G21890 and G13530);
	I28742<= not (G21890 and I28741);
	I28743<= not (G13530 and I28741);
	I28753<= not (G21893 and G13541);
	I28754<= not (G21893 and I28753);
	I28755<= not (G13541 and I28753);
	I28765<= not (G21901 and G13552);
	I28766<= not (G21901 and I28765);
	I28767<= not (G13552 and I28765);
	I30790<= not (G22846 and G14079);
	I30791<= not (G22846 and I30790);
	I30792<= not (G14079 and I30790);
	I30868<= not (G22881 and G14194);
	I30869<= not (G22881 and I30868);
	I30870<= not (G14194 and I30868);
	I30952<= not (G22916 and G14309);
	I30953<= not (G22916 and I30952);
	I30954<= not (G14309 and I30952);
	I31035<= not (G22941 and G14431);
	I31036<= not (G22941 and I31035);
	I31037<= not (G14431 and I31035);
	I32265<= not (G17903 and G23936);
	I32266<= not (G17903 and I32265);
	I32267<= not (G23936 and I32265);
	I32284<= not (G17815 and G23953);
	I32285<= not (G17815 and I32284);
	I32286<= not (G23953 and I32284);
	I32295<= not (G18014 and G23968);
	I32296<= not (G18014 and I32295);
	I32297<= not (G23968 and I32295);
	I32308<= not (G17903 and G23973);
	I32309<= not (G17903 and I32308);
	I32310<= not (G23973 and I32308);
	I32323<= not (G17927 and G23982);
	I32324<= not (G17927 and I32323);
	I32325<= not (G23982 and I32323);
	I32333<= not (G18131 and G23997);
	I32334<= not (G18131 and I32333);
	I32335<= not (G23997 and I32333);
	I32345<= not (G17815 and G24002);
	I32346<= not (G17815 and I32345);
	I32347<= not (G24002 and I32345);
	I32355<= not (G18014 and G24003);
	I32356<= not (G18014 and I32355);
	I32357<= not (G24003 and I32355);
	I32368<= not (G18038 and G24012);
	I32369<= not (G18038 and I32368);
	I32370<= not (G24012 and I32368);
	I32378<= not (G18247 and G24027);
	I32379<= not (G18247 and I32378);
	I32380<= not (G24027 and I32378);
	I32391<= not (G17903 and G24034);
	I32392<= not (G17903 and I32391);
	I32393<= not (G24034 and I32391);
	I32400<= not (G17927 and G24036);
	I32401<= not (G17927 and I32400);
	I32402<= not (G24036 and I32400);
	I32409<= not (G18131 and G24037);
	I32410<= not (G18131 and I32409);
	I32411<= not (G24037 and I32409);
	I32422<= not (G18155 and G24046);
	I32423<= not (G18155 and I32422);
	I32424<= not (G24046 and I32422);
	I32430<= not (G17815 and G24052);
	I32431<= not (G17815 and I32430);
	I32432<= not (G24052 and I32430);
	I32443<= not (G18014 and G24054);
	I32444<= not (G18014 and I32443);
	I32445<= not (G24054 and I32443);
	I32451<= not (G18038 and G24056);
	I32452<= not (G18038 and I32451);
	I32453<= not (G24056 and I32451);
	I32460<= not (G18247 and G24057);
	I32461<= not (G18247 and I32460);
	I32462<= not (G24057 and I32460);
	I32468<= not (G17903 and G24058);
	I32469<= not (G17903 and I32468);
	I32470<= not (G24058 and I32468);
	I32478<= not (G17927 and G24065);
	I32479<= not (G17927 and I32478);
	I32480<= not (G24065 and I32478);
	I32490<= not (G18131 and G24067);
	I32491<= not (G18131 and I32490);
	I32492<= not (G24067 and I32490);
	I32498<= not (G18155 and G24069);
	I32499<= not (G18155 and I32498);
	I32500<= not (G24069 and I32498);
	I32509<= not (G17815 and G24070);
	I32510<= not (G17815 and I32509);
	I32511<= not (G24070 and I32509);
	I32518<= not (G18014 and G24071);
	I32519<= not (G18014 and I32518);
	I32520<= not (G24071 and I32518);
	I32526<= not (G18038 and G24078);
	I32527<= not (G18038 and I32526);
	I32528<= not (G24078 and I32526);
	I32538<= not (G18247 and G24080);
	I32539<= not (G18247 and I32538);
	I32540<= not (G24080 and I32538);
	I32546<= not (G17903 and G23906);
	I32547<= not (G17903 and I32546);
	I32548<= not (G23906 and I32546);
	I32559<= not (G17927 and G24081);
	I32560<= not (G17927 and I32559);
	I32561<= not (G24081 and I32559);
	I32567<= not (G18131 and G24082);
	I32568<= not (G18131 and I32567);
	I32569<= not (G24082 and I32567);
	I32575<= not (G18155 and G24089);
	I32576<= not (G18155 and I32575);
	I32577<= not (G24089 and I32575);
	I32586<= not (G17815 and G23937);
	I32587<= not (G17815 and I32586);
	I32588<= not (G23937 and I32586);
	I32595<= not (G18014 and G23938);
	I32596<= not (G18014 and I32595);
	I32597<= not (G23938 and I32595);
	I32607<= not (G18038 and G24090);
	I32608<= not (G18038 and I32607);
	I32609<= not (G24090 and I32607);
	I32615<= not (G18247 and G24091);
	I32616<= not (G18247 and I32615);
	I32617<= not (G24091 and I32615);
	I32624<= not (G17927 and G23969);
	I32625<= not (G17927 and I32624);
	I32626<= not (G23969 and I32624);
	I32633<= not (G18131 and G23970);
	I32634<= not (G18131 and I32633);
	I32635<= not (G23970 and I32633);
	I32645<= not (G18155 and G24093);
	I32646<= not (G18155 and I32645);
	I32647<= not (G24093 and I32645);
	I32659<= not (G18038 and G23998);
	I32660<= not (G18038 and I32659);
	I32661<= not (G23998 and I32659);
	I32668<= not (G18247 and G23999);
	I32669<= not (G18247 and I32668);
	I32670<= not (G23999 and I32668);
	I32677<= not (G23823 and G14165);
	I32678<= not (G23823 and I32677);
	I32679<= not (G14165 and I32677);
	I32686<= not (G18155 and G24028);
	I32687<= not (G18155 and I32686);
	I32688<= not (G24028 and I32686);
	I32695<= not (G23858 and G14280);
	I32696<= not (G23858 and I32695);
	I32697<= not (G14280 and I32695);
	I32708<= not (G23892 and G14402);
	I32709<= not (G23892 and I32708);
	I32710<= not (G14402 and I32708);
	I32724<= not (G23913 and G14514);
	I32725<= not (G23913 and I32724);
	I32726<= not (G14514 and I32724);
	I35020<= not (G26110 and G26099);
	I35021<= not (G26110 and I35020);
	I35022<= not (G26099 and I35020);
	I35034<= not (G26087 and G26154);
	I35035<= not (G26087 and I35034);
	I35036<= not (G26154 and I35034);
	I35042<= not (G26151 and G26145);
	I35043<= not (G26151 and I35042);
	I35044<= not (G26145 and I35042);
	I35057<= not (G26137 and G26126);
	I35058<= not (G26137 and I35057);
	I35059<= not (G26126 and I35057);
	I35123<= not (G26107 and G26096);
	I35124<= not (G26107 and I35123);
	I35125<= not (G26096 and I35123);
	I35701<= not (G26867 and G26874);
	I35702<= not (G26867 and I35701);
	I35703<= not (G26874 and I35701);
	I35714<= not (G26859 and G26865);
	I35715<= not (G26859 and I35714);
	I35716<= not (G26865 and I35714);
	I35904<= not (G27051 and G14831);
	I35905<= not (G27051 and I35904);
	I35906<= not (G14831 and I35904);
	I35944<= not (G27078 and G14904);
	I35945<= not (G27078 and I35944);
	I35946<= not (G14904 and I35944);
	I35974<= not (G27094 and G14985);
	I35975<= not (G27094 and I35974);
	I35976<= not (G14985 and I35974);
	I35992<= not (G27106 and G15074);
	I35993<= not (G27106 and I35992);
	I35994<= not (G15074 and I35992);
	I36256<= not (G27527 and G15859);
	I36257<= not (G27527 and I36256);
	I36258<= not (G15859 and I36256);
	I36270<= not (G27549 and G15890);
	I36271<= not (G27549 and I36270);
	I36272<= not (G15890 and I36270);
	I36289<= not (G27565 and G15923);
	I36290<= not (G27565 and I36289);
	I36291<= not (G15923 and I36289);
	I36300<= not (G27382 and G27379);
	I36301<= not (G27382 and I36300);
	I36302<= not (G27379 and I36300);
	I36314<= not (G27575 and G15952);
	I36315<= not (G27575 and I36314);
	I36316<= not (G15952 and I36314);
	I36591<= not (G27529 and G14885);
	I36592<= not (G27529 and I36591);
	I36593<= not (G14885 and I36591);
	I36666<= not (G27551 and G14966);
	I36667<= not (G27551 and I36666);
	I36668<= not (G14966 and I36666);
	I36731<= not (G27567 and G15055);
	I36732<= not (G27567 and I36731);
	I36733<= not (G15055 and I36731);
	I36779<= not (G27577 and G15151);
	I36780<= not (G27577 and I36779);
	I36781<= not (G15151 and I36779);
	I37295<= not (G27827 and G27814);
	I37296<= not (G27827 and I37295);
	I37297<= not (G27814 and I37295);
	I37303<= not (G27802 and G27900);
	I37304<= not (G27802 and I37303);
	I37305<= not (G27900 and I37303);
	I37311<= not (G27897 and G27883);
	I37312<= not (G27897 and I37311);
	I37313<= not (G27883 and I37311);
	I37322<= not (G27865 and G27855);
	I37323<= not (G27865 and I37322);
	I37324<= not (G27855 and I37322);
	I37356<= not (G27824 and G27811);
	I37357<= not (G27824 and I37356);
	I37358<= not (G27811 and I37356);
	I37813<= not (G28388 and G28391);
	I37814<= not (G28388 and I37813);
	I37815<= not (G28391 and I37813);
	I37822<= not (G28384 and G28386);
	I37823<= not (G28384 and I37822);
	I37824<= not (G28386 and I37822);
	I38378<= not (G28845 and G28842);
	I38379<= not (G28845 and I38378);
	I38380<= not (G28842 and I38378);
	I38810<= not (G29303 and G15904);
	I38811<= not (G29303 and I38810);
	I38812<= not (G15904 and I38810);
	I38820<= not (G29313 and G15933);
	I38821<= not (G29313 and I38820);
	I38822<= not (G15933 and I38820);
	I38831<= not (G29324 and G15962);
	I38832<= not (G29324 and I38831);
	I38833<= not (G15962 and I38831);
	I38841<= not (G29333 and G15981);
	I38842<= not (G29333 and I38841);
	I38843<= not (G15981 and I38841);
	I39323<= not (G29721 and G29713);
	I39324<= not (G29721 and I39323);
	I39325<= not (G29713 and I39323);
	I39331<= not (G29705 and G29751);
	I39332<= not (G29705 and I39331);
	I39333<= not (G29751 and I39331);
	I39339<= not (G29748 and G29741);
	I39340<= not (G29748 and I39339);
	I39341<= not (G29741 and I39339);
	I39347<= not (G29732 and G29728);
	I39348<= not (G29732 and I39347);
	I39349<= not (G29728 and I39347);
	I39359<= not (G29766 and G15880);
	I39360<= not (G29766 and I39359);
	I39361<= not (G15880 and I39359);
	I39367<= not (G29767 and G15913);
	I39368<= not (G29767 and I39367);
	I39369<= not (G15913 and I39367);
	I39375<= not (G29768 and G15942);
	I39376<= not (G29768 and I39375);
	I39377<= not (G15942 and I39375);
	I39384<= not (G29718 and G29710);
	I39385<= not (G29718 and I39384);
	I39386<= not (G29710 and I39384);
	I39391<= not (G29769 and G15971);
	I39392<= not (G29769 and I39391);
	I39393<= not (G15971 and I39391);
	I39532<= not (G29915 and G29917);
	I39533<= not (G29915 and I39532);
	I39534<= not (G29917 and I39532);
	I39539<= not (G29911 and G29913);
	I39540<= not (G29911 and I39539);
	I39541<= not (G29913 and I39539);
	I39689<= not (G30035 and G30034);
	I39690<= not (G30035 and I39689);
	I39691<= not (G30034 and I39689);
	I40558<= not (G30605 and G30597);
	I40559<= not (G30605 and I40558);
	I40560<= not (G30597 and I40558);
	I40571<= not (G30588 and G30632);
	I40572<= not (G30588 and I40571);
	I40573<= not (G30632 and I40571);
	I40587<= not (G30629 and G30622);
	I40588<= not (G30629 and I40587);
	I40589<= not (G30622 and I40587);
	I40603<= not (G30614 and G30610);
	I40604<= not (G30614 and I40603);
	I40605<= not (G30610 and I40603);
	I40627<= not (G30602 and G30594);
	I40628<= not (G30602 and I40627);
	I40629<= not (G30594 and I40627);
	I41010<= not (G30775 and G30779);
	I41011<= not (G30775 and I41010);
	I41012<= not (G30779 and I41010);
	I41017<= not (G30768 and G30771);
	I41018<= not (G30768 and I41017);
	I41019<= not (G30771 and I41017);
	I41064<= not (G30927 and G30926);
	I41065<= not (G30927 and I41064);
	I41066<= not (G30926 and I41064);
	G9144<=G2986 or G5389;
	G10778<=G2929 or G8022;
	G12377<=G7553 or G11059;
	G12407<=G7573 or G10779;
	G12886<=G9534 or G3398;
	G12926<=G9676 or G3554;
	G12955<=G9822 or G3710;
	G12984<=G9968 or G3866;
	G16539<=G15880 or G14657;
	G16571<=G15913 or G14691;
	G16595<=G15942 or G14725;
	G16615<=G15971 or G14753;
	G17973<=G11623 or G15659;
	G19181<=G17729 or G17979;
	G19186<=G18419 or G17887;
	G19187<=G18419 or G17729;
	G19188<=G17830 or G18096;
	G19191<=G17807 or G17887;
	G19192<=G18183 or G18270;
	G19193<=G18492 or G17998;
	G19194<=G18492 or G17830;
	G19195<=G17942 or G18212;
	G19200<=G18346 or G18424;
	G19201<=G18183 or G18424;
	G19202<=G17919 or G17998;
	G19203<=G18290 or G18363;
	G19204<=G18556 or G18115;
	G19205<=G18556 or G17942;
	G19206<=G18053 or G18319;
	G19209<=G18079 or G18346;
	G19210<=G18079 or G18183;
	G19211<=G18441 or G18497;
	G19212<=G18290 or G18497;
	G19213<=G18030 or G18115;
	G19214<=G18383 or G18458;
	G19215<=G18606 or G18231;
	G19216<=G18606 or G18053;
	G19221<=G18270 or G18346;
	G19222<=G18195 or G18441;
	G19223<=G18195 or G18290;
	G19224<=G18514 or G18561;
	G19225<=G18383 or G18561;
	G19226<=G18147 or G18231;
	G19227<=G18478 or G18531;
	G19230<=G16985 or G16965 or I25477;
	G19231<=G18363 or G18441;
	G19232<=G18302 or G18514;
	G19233<=G18302 or G18383;
	G19234<=G18578 or G18611;
	G19235<=G18478 or G18611;
	G19240<=G17083 or G17050 or I25495;
	G19242<=G14244 or G16501;
	G19243<=G16995 or G16986 or I25500;
	G19244<=G18458 or G18514;
	G19245<=G18395 or G18578;
	G19246<=G18395 or G18478;
	G19250<=G17729 or G17807;
	G19253<=G17121 or G17085 or I25516;
	G19255<=G14366 or G16523;
	G19256<=G17019 or G16996 or I25521;
	G19257<=G18531 or G18578;
	G19263<=G17887 or G17979;
	G19264<=G17830 or G17919;
	G19266<=G17148 or G17123 or I25549;
	G19268<=G14478 or G16554;
	G19269<=G17049 or G17020 or I25554;
	G19275<=G16867 or G16515 or G19001;
	G19278<=G17998 or G18096;
	G19279<=G17942 or G18030;
	G19281<=G17171 or G17150 or I25588;
	G19283<=G14565 or G16586;
	G19294<=G16895 or G16546 or G16507;
	G19297<=G18115 or G18212;
	G19298<=G18053 or G18147;
	G19312<=G16924 or G16578 or G16529;
	G19315<=G18231 or G18319;
	G19333<=G16954 or G16602 or G16560;
	G19450<=G14837 or G16682;
	G19477<=G14910 or G16708;
	G19500<=G14991 or G16739;
	G19503<=G16884 or G16697 or G16665;
	G19521<=G15080 or G16781;
	G19522<=G16913 or G16728 or G16686;
	G19532<=G16943 or G16770 or G16712;
	G19542<=G16974 or G16797 or G16743;
	G19981<=G17729 or G18419 or I26429;
	G20015<=G18183 or G18079 or I26455;
	G20019<=G17830 or G18492 or I26461;
	G20057<=G18290 or G18195 or I26491;
	G20061<=G17942 or G18556 or I26497;
	G20098<=G18383 or G18302 or I26532;
	G20102<=G18053 or G18606 or I26538;
	G20123<=G18478 or G18395 or I26571;
	G21120<=G19484 or G16515 or G14071;
	G21139<=G19505 or G16546 or G14186;
	G21159<=G19524 or G16578 or G14301;
	G21179<=G19534 or G16602 or G14423;
	G21244<=G19578 or G16697 or G14776;
	G21253<=G19608 or G16728 or G14811;
	G21261<=G19641 or G16770 or G14863;
	G21269<=G19681 or G16797 or G14936;
	G21501<=G20522 or G16867 or G14071;
	G21536<=G20522 or G19484 or G19001;
	G21540<=G20542 or G16895 or G14186;
	G21572<=G20542 or G19505 or G16507;
	G21576<=G19067 or G16924 or G14301;
	G21605<=G19067 or G19524 or G16529;
	G21609<=G19084 or G16954 or G14423;
	G21634<=G19084 or G19534 or G16560;
	G21774<=G19121 or G16884 or G14776;
	G21787<=G19121 or G19578 or G16665;
	G21788<=G20117 or G20094 or I28305;
	G21789<=G19128 or G16913 or G14811;
	G21799<=G16505 or G20538 or G18994 or I28318;
	G21800<=G18665 or G20270 or G20248 or G18647;
	G21801<=G19128 or G19608 or G16686;
	G21802<=G20147 or G20119 or I28323;
	G21803<=G19135 or G16943 or G14863;
	G21806<=G20116 or G20093 or G18547 or G19097;
	G21807<=G16527 or G19063 or G19007 or I28330;
	G21808<=G18688 or G20282 or G20271 or G18650;
	G21809<=G19135 or G19641 or G16712;
	G21810<=G20185 or G20149 or I28335;
	G21811<=G19138 or G16974 or G14936;
	G21813<=G20146 or G20118 or G18597 or G19104;
	G21814<=G16558 or G19080 or G16513 or I28341;
	G21815<=G18717 or G20293 or G20283 or G18654;
	G21816<=G19138 or G19681 or G16743;
	G21817<=G20219 or G20187 or I28346;
	G21819<=G20184 or G20148 or G18629 or G19109;
	G21820<=G16590 or G19090 or G16535 or I28351;
	G21821<=G18753 or G20309 or G20294 or G18668;
	G21823<=G20218 or G20186 or G18638 or G19116;
	G21844<=G20222 or G18645 or I28365;
	G21846<=G20249 or G18648 or I28369;
	G21849<=G20272 or G18651 or I28374;
	G21856<=G20284 or G18655 or I28380;
	G22175<=G16075 or G20842;
	G22190<=G16113 or G20850;
	G22199<=G16164 or G20858;
	G22205<=G16223 or G20866;
	G22811<=G562 or G559 or G12451 or G21851;
	G23052<=G21800 or G21788 or G21844;
	G23071<=G21808 or G21802 or G21846;
	G23084<=G21815 or G21810 or G21849;
	G23089<=G21806 or G21799;
	G23100<=G21821 or G21817 or G21856;
	G23107<=G21813 or G21807;
	G23120<=G21819 or G21814;
	G23129<=G21823 or G21820;
	G23319<=G14493 or G22385;
	G23688<=G23106 or G21906;
	G23742<=G23119 or G21920;
	G23797<=G23128 or G21938;
	G23850<=G23139 or G20647;
	G23919<=G22666 or G23140;
	G24239<=G19387 or G22401;
	G24244<=G14144 or G22317;
	G24245<=G19417 or G22402;
	G24252<=G14259 or G22342;
	G24254<=G19454 or G22403;
	G24257<=G14381 or G22365;
	G24258<=G19481 or G22404;
	G24633<=G24094 or G20842;
	G24653<=G24095 or G20850;
	G24672<=G24097 or G20858;
	G24691<=G24103 or G20866;
	G24890<=G23639 or G23144;
	G24909<=G23726 or G23142;
	G24925<=G23772 or G23141;
	G24965<=G23922 or G23945;
	G24978<=G23954 or G23974;
	G24989<=G23983 or G24004;
	G25000<=G24013 or G24038;
	G25183<=G24958 or G24893;
	G25186<=G24969 or G24916;
	G25190<=G24982 or G24933;
	G25195<=G24993 or G24945;
	G25489<=G24795 or G16466;
	G25490<=G24759 or G23146;
	G25520<=G24813 or G23145;
	G25566<=G24843 or G23143;
	G26320<=G25852 or G25870;
	G26367<=G25873 or G25882;
	G26410<=G25885 or G25887;
	G26451<=G25890 or G25892;
	G26974<=G26157 or G23147;
	G27113<=G1248 or G1245 or G26534;
	G28501<=G27738 or G25764;
	G28512<=G26481 or G27738;
	G28529<=G27743 or G25818;
	G28540<=G26497 or G27743;
	G28556<=G27751 or G25853;
	G28567<=G26512 or G27751;
	G28584<=G27756 or G25874;
	G28595<=G26520 or G27756;
	G29348<=G1942 or G1939 or G29113;
	G30305<=G2636 or G2633 or G30072;
	I25477<=G17024 or G17000 or G16992;
	I25495<=G17158 or G17137 or G17115;
	I25500<=G17058 or G17030 or G17016;
	I25516<=G17173 or G17160 or G17142;
	I25521<=G17093 or G17064 or G17046;
	I25549<=G17190 or G17175 or G17165;
	I25554<=G17131 or G17099 or G17080;
	I25588<=G17201 or G17192 or G17180;
	I26429<=G17979 or G17887 or G17807;
	I26455<=G18424 or G18346 or G18270;
	I26461<=G18096 or G17998 or G17919;
	I26491<=G18497 or G18441 or G18363;
	I26497<=G18212 or G18115 or G18030;
	I26532<=G18561 or G18514 or G18458;
	I26538<=G18319 or G18231 or G18147;
	I26571<=G18611 or G18578 or G18531;
	I28305<=G20197 or G20177 or G20145;
	I28318<=G19092 or G19088 or G19079;
	I28323<=G20227 or G20211 or G20183;
	I28330<=G19099 or G19094 or G19089;
	I28335<=G20254 or G20241 or G20217;
	I28341<=G19106 or G19101 or G19095;
	I28346<=G20277 or G20268 or G20247;
	I28351<=G19111 or G19108 or G19102;
	I28365<=G20280 or G18652 or G18649;
	I28369<=G20291 or G18666 or G18653;
	I28374<=G20307 or G18689 or G18667;
	I28380<=G20326 or G18718 or G18690;
	G7528<= not (G3151 or G3142 or G3147);
	G7575<= not (G2984 or G2985);
	G7795<= not (G2992 or G2991);
	G8430<= not (G3198 or G8120 or G3194 or G3191);
	G10784<= not (G5630 or G5649 or G5676);
	G10789<= not (G5650 or G5677 or G5709);
	G10793<= not (G5658 or G5687 or G5728);
	G10797<= not (G5678 or G5710 or G5757);
	G10801<= not (G5688 or G5729 or G5767);
	G10805<= not (G5696 or G5739 or G5786);
	G10810<= not (G5711 or G5758 or G5807);
	G10814<= not (G5730 or G5768 or G5816);
	G10818<= not (G5740 or G5787 or G5826);
	G10822<= not (G5748 or G5797 or G5845);
	G10831<= not (G5769 or G5817 or G5863);
	G10835<= not (G5788 or G5827 or G5872);
	G10839<= not (G5798 or G5846 or G5882);
	G10851<= not (G5828 or G5873 or G5910);
	G10855<= not (G5847 or G5883 or G5919);
	G10872<= not (G5884 or G5920 or G5949);
	G11600<= not (G9049 or G9064 or G9078);
	G11622<= not (G8183 or G11332 or G7928 or G11069);
	G11624<= not (G9062 or G9075 or G9091);
	G11627<= not (G9063 or G9077 or G9093);
	G11630<= not (G9066 or G9081 or G9097);
	G11643<= not (G11481 or G8045 or G7928 or G11069);
	G11644<= not (G9076 or G9092 or G9102);
	G11647<= not (G9079 or G9094 or G9103);
	G11650<= not (G9080 or G9096 or G9105);
	G11653<= not (G9083 or G9100 or G9109);
	G11660<= not (G8183 or G8045 or G7928 or G11069);
	G11663<= not (G9095 or G9104 or G9112);
	G11666<= not (G9098 or G9106 or G9113);
	G11669<= not (G9099 or G9108 or G9115);
	G11675<= not (G9107 or G9114 or G9120);
	G11678<= not (G9110 or G9116 or G9121);
	G11681<= not (G9111 or G9118 or G9123);
	G11687<= not (G9117 or G9122 or G9126);
	G11690<= not (G9119 or G9124 or G9127);
	G11697<= not (G9125 or G9131 or G9133);
	G11703<= not (G9132 or G9137 or G9139);
	G11711<= not (G9138 or G9143 or G9145);
	G11744<= not (G9241 or G9301 or G9364);
	G11759<= not (G9302 or G9365 or G9438);
	G11760<= not (G9319 or G9382 or G9461);
	G11767<= not (G9366 or G9439 or G9518);
	G11768<= not (G9367 or G9441 or G9521);
	G11772<= not (G9383 or G9462 or G9580);
	G11773<= not (G9400 or G9479 or G9603);
	G11780<= not (G9440 or G9519 or G9630);
	G11781<= not (G9442 or G9522 or G9633);
	G11784<= not (G9463 or G9581 or G9660);
	G11785<= not (G9464 or G9583 or G9663);
	G11789<= not (G9480 or G9604 or G9722);
	G11790<= not (G9497 or G9621 or G9745);
	G11799<= not (G9520 or G9631 or G9759);
	G11800<= not (G9523 or G9634 or G9762);
	G11806<= not (G9582 or G9661 or G9776);
	G11807<= not (G9584 or G9664 or G9779);
	G11810<= not (G9605 or G9723 or G9806);
	G11811<= not (G9606 or G9725 or G9809);
	G11815<= not (G9622 or G9746 or G9868);
	G11822<= not (G9632 or G9760 or G9888);
	G11823<= not (G9635 or G9763 or G9891);
	G11828<= not (G9639 or G9764 or G9892);
	G11830<= not (G9647 or G9773 or G9901);
	G11831<= not (G9648 or G9775 or G9904);
	G11832<= not (G9662 or G9777 or G9905);
	G11833<= not (G9665 or G9780 or G9908);
	G11839<= not (G9724 or G9807 or G9922);
	G11840<= not (G9726 or G9810 or G9925);
	G11843<= not (G9747 or G9869 or G9952);
	G11844<= not (G9748 or G9871 or G9955);
	G11855<= not (G9761 or G9889 or G10009);
	G11860<= not (G9765 or G9893 or G10012);
	G11861<= not (G9766 or G9894 or G10013);
	G11863<= not (G9774 or G9902 or G10035);
	G11864<= not (G9778 or G9906 or G10042);
	G11865<= not (G9781 or G9909 or G10045);
	G11870<= not (G9785 or G9910 or G10046);
	G11872<= not (G9793 or G9919 or G10055);
	G11873<= not (G9794 or G9921 or G10058);
	G11874<= not (G9808 or G9923 or G10059);
	G11875<= not (G9811 or G9926 or G10062);
	G11881<= not (G9870 or G9953 or G10076);
	G11882<= not (G9872 or G9956 or G10079);
	G11889<= not (G9887 or G10007 or G10101);
	G11890<= not (G9890 or G10010 or G10103);
	G11896<= not (G9903 or G10036 or G10112);
	G11897<= not (G9907 or G10043 or G10118);
	G11902<= not (G9911 or G10047 or G10121);
	G11903<= not (G9912 or G10048 or G10122);
	G11905<= not (G9920 or G10056 or G10144);
	G11906<= not (G9924 or G10060 or G10151);
	G11907<= not (G9927 or G10063 or G10154);
	G11912<= not (G9931 or G10064 or G10155);
	G11914<= not (G9939 or G10073 or G10164);
	G11915<= not (G9940 or G10075 or G10167);
	G11916<= not (G9954 or G10077 or G10168);
	G11917<= not (G9957 or G10080 or G10171);
	G11928<= not (G10008 or G10102 or G10192);
	G11934<= not (G10011 or G10104 or G10193);
	G11935<= not (G10014 or G10106 or G10196);
	G11938<= not (G10037 or G10113 or G10201);
	G11939<= not (G10041 or G10116 or G10206);
	G11940<= not (G10044 or G10119 or G10208);
	G11946<= not (G10057 or G10145 or G10217);
	G11947<= not (G10061 or G10152 or G10223);
	G11952<= not (G10065 or G10156 or G10226);
	G11953<= not (G10066 or G10157 or G10227);
	G11955<= not (G10074 or G10165 or G10249);
	G11956<= not (G10078 or G10169 or G10256);
	G11957<= not (G10081 or G10172 or G10259);
	G11962<= not (G10085 or G10173 or G10260);
	G11964<= not (G10093 or G10182 or G10269);
	G11965<= not (G10094 or G10184 or G10272);
	G11974<= not (G10105 or G10194 or G10279);
	G11975<= not (G10107 or G10197 or G10282);
	G11979<= not (G10114 or G10202 or G10288);
	G11980<= not (G10115 or G10204 or G10291);
	G11981<= not (G10117 or G10207 or G10294);
	G11987<= not (G10120 or G10209 or G10295);
	G11988<= not (G10123 or G10211 or G10298);
	G11991<= not (G10146 or G10218 or G10303);
	G11992<= not (G10150 or G10221 or G10308);
	G11993<= not (G10153 or G10224 or G10310);
	G11999<= not (G10166 or G10250 or G10319);
	G12000<= not (G10170 or G10257 or G10325);
	G12005<= not (G10174 or G10261 or G10328);
	G12006<= not (G10175 or G10262 or G10329);
	G12008<= not (G10183 or G10270 or G10351);
	G12026<= not (G10195 or G10280 or G10360);
	G12033<= not (G10199 or G10284 or G10362);
	G12034<= not (G10200 or G10286 or G10365);
	G12035<= not (G10203 or G10289 or G10367);
	G12036<= not (G10205 or G10292 or G10370);
	G12043<= not (G10210 or G10296 or G10372);
	G12044<= not (G10212 or G10299 or G10375);
	G12048<= not (G10219 or G10304 or G10381);
	G12049<= not (G10220 or G10306 or G10384);
	G12050<= not (G10222 or G10309 or G10387);
	G12056<= not (G10225 or G10311 or G10388);
	G12057<= not (G10228 or G10313 or G10391);
	G12060<= not (G10251 or G10320 or G10396);
	G12061<= not (G10255 or G10323 or G10401);
	G12062<= not (G10258 or G10326 or G10403);
	G12068<= not (G10271 or G10352 or G10412);
	G12079<= not (G10281 or G10361 or G10422);
	G12080<= not (G10285 or G10363 or G10430);
	G12081<= not (G10287 or G10366 or G10433);
	G12082<= not (G10290 or G10368 or G10435);
	G12083<= not (G10293 or G10371 or G10438);
	G12090<= not (G10297 or G10373 or G10439);
	G12097<= not (G10301 or G10377 or G10441);
	G12098<= not (G10302 or G10379 or G10444);
	G12099<= not (G10305 or G10382 or G10446);
	G12100<= not (G10307 or G10385 or G10449);
	G12107<= not (G10312 or G10389 or G10451);
	G12108<= not (G10314 or G10392 or G10454);
	G12112<= not (G10321 or G10397 or G10460);
	G12113<= not (G10322 or G10399 or G10463);
	G12114<= not (G10324 or G10402 or G10466);
	G12120<= not (G10327 or G10404 or G10467);
	G12121<= not (G10330 or G10406 or G10470);
	G12124<= not (G10353 or G10413 or G10475);
	G12145<= not (G10364 or G10431 or G10492);
	G12146<= not (G10369 or G10436 or G10496);
	G12151<= not (G10374 or G10440 or G10498);
	G12152<= not (G10378 or G10442 or G10506);
	G12153<= not (G10380 or G10445 or G10509);
	G12154<= not (G10383 or G10447 or G10511);
	G12155<= not (G10386 or G10450 or G10514);
	G12162<= not (G10390 or G10452 or G10515);
	G12169<= not (G10394 or G10456 or G10517);
	G12170<= not (G10395 or G10458 or G10520);
	G12171<= not (G10398 or G10461 or G10522);
	G12172<= not (G10400 or G10464 or G10525);
	G12179<= not (G10405 or G10468 or G10527);
	G12180<= not (G10407 or G10471 or G10530);
	G12184<= not (G10414 or G10476 or G10536);
	G12185<= not (G10415 or G10478 or G10539);
	G12192<= not (G10423 or G10485 or G10548);
	G12193<= not (G10432 or G10493 or G10555);
	G12194<= not (G10434 or G10494 or G10556);
	G12195<= not (G10437 or G10497 or G10558);
	G12207<= not (G10443 or G10507 or G10566);
	G12208<= not (G10448 or G10512 or G10570);
	G12213<= not (G10453 or G10516 or G10572);
	G12214<= not (G10457 or G10518 or G10580);
	G12215<= not (G10459 or G10521 or G10583);
	G12216<= not (G10462 or G10523 or G10585);
	G12217<= not (G10465 or G10526 or G10588);
	G12224<= not (G10469 or G10528 or G10589);
	G12231<= not (G10473 or G10532 or G10591);
	G12232<= not (G10474 or G10534 or G10594);
	G12233<= not (G10477 or G10537 or G10596);
	G12234<= not (G10479 or G10540 or G10599);
	G12245<= not (G10495 or G10557 or G10604);
	G12247<= not (G10499 or G10559 or G10605);
	G12248<= not (G10508 or G10567 or G10612);
	G12249<= not (G10510 or G10568 or G10613);
	G12250<= not (G10513 or G10571 or G10615);
	G12262<= not (G10519 or G10581 or G10623);
	G12263<= not (G10524 or G10586 or G10627);
	G12268<= not (G10529 or G10590 or G10629);
	G12269<= not (G10533 or G10592 or G10637);
	G12270<= not (G10535 or G10595 or G10640);
	G12271<= not (G10538 or G10597 or G10642);
	G12272<= not (G10541 or G10600 or G10645);
	G12288<= not (G10569 or G10614 or G10651);
	G12290<= not (G10573 or G10616 or G10652);
	G12291<= not (G10582 or G10624 or G10659);
	G12292<= not (G10584 or G10625 or G10660);
	G12293<= not (G10587 or G10628 or G10662);
	G12305<= not (G10593 or G10638 or G10670);
	G12306<= not (G10598 or G10643 or G10674);
	G12324<= not (G10626 or G10661 or G10681);
	G12326<= not (G10630 or G10663 or G10682);
	G12327<= not (G10639 or G10671 or G10689);
	G12328<= not (G10641 or G10672 or G10690);
	G12329<= not (G10644 or G10675 or G10692);
	G12339<= not (G10650 or G10678 or G10704);
	G12352<= not (G10673 or G10691 or G10710);
	G12369<= not (G10680 or G10707 or G10724);
	G12388<= not (G10709 or G10727 or G10745);
	G12418<= not (G10729 or G10748 or G10764);
	G12431<= not (G8580 or G10730);
	G12436<= not (G8587 or G10749);
	G12441<= not (G8594 or G10767);
	G12446<= not (G8605 or G10773);
	G12451<= not (G499 or G8983);
	G12457<= not (G9009 or G9033 or G9048);
	G12467<= not (G9034 or G9056 or G9065);
	G12482<= not (G9057 or G9073 or G9082);
	G12487<= not (G10108 or G10198 or G10283);
	G12499<= not (G9074 or G9090 or G9101);
	G12507<= not (G10213 or G10300 or G10376);
	G12524<= not (G10315 or G10393 or G10455);
	G12539<= not (G10408 or G10472 or G10531);
	G12698<= not (G11347 or G11420 or G8327);
	G12747<= not (G11421 or G8328 or G8385);
	G12755<= not (G11431 or G8339 or G8394);
	G12780<= not (G9187 or G9161);
	G12781<= not (G8329 or G8386 or G8431);
	G12789<= not (G8340 or G8395 or G8437);
	G12797<= not (G8350 or G8406 or G8446);
	G12814<= not (G8387 or G8432 or G8463);
	G12819<= not (G9248 or G9203);
	G12820<= not (G8396 or G8438 or G8466);
	G12828<= not (G8407 or G8447 or G8472);
	G12836<= not (G8417 or G8458 or G8481);
	G12849<= not (G8433 or G8464 or G8485);
	G12852<= not (G8439 or G8467 or G8488);
	G12857<= not (G9326 or G9264);
	G12858<= not (G8448 or G8473 or G8491);
	G12866<= not (G8459 or G8482 or G8497);
	G12880<= not (G8465 or G8486 or G8502);
	G12883<= not (G10038 or G6284);
	G12890<= not (G8468 or G8489 or G8505);
	G12893<= not (G8474 or G8492 or G8508);
	G12898<= not (G9407 or G9342);
	G12899<= not (G8483 or G8498 or G8511);
	G12912<= not (G8484 or G8500 or G8515);
	G12913<= not (G8487 or G8503 or G8518);
	G12920<= not (G8490 or G8506 or G8521);
	G12923<= not (G10147 or G6421);
	G12930<= not (G8493 or G8509 or G8524);
	G12933<= not (G8499 or G8512 or G8527);
	G12939<= not (G8501 or G8516 or G8531);
	G12941<= not (G8504 or G8519 or G8534);
	G12942<= not (G8507 or G8522 or G8537);
	G12949<= not (G8510 or G8525 or G8540);
	G12952<= not (G10252 or G6626);
	G12959<= not (G8513 or G8528 or G8543);
	G12967<= not (G8517 or G8532 or G8546);
	G12968<= not (G8520 or G8535 or G8548);
	G12970<= not (G8523 or G8538 or G8551);
	G12971<= not (G8526 or G8541 or G8554);
	G12978<= not (G8529 or G8544 or G8557);
	G12981<= not (G10354 or G6890);
	G12991<= not (G8536 or G8549 or G8559);
	G12992<= not (G8539 or G8552 or G8561);
	G12994<= not (G8542 or G8555 or G8564);
	G12995<= not (G8545 or G8558 or G8567);
	G13001<= not (G8553 or G8562 or G8570);
	G13002<= not (G8556 or G8565 or G8572);
	G13022<= not (G8566 or G8573 or G8576);
	G13024<= not (G11481 or G8045 or G7928 or G7880);
	G13111<= not (G8601 or G8612 or G8621);
	G13124<= not (G8613 or G8625 or G8631);
	G13135<= not (G8626 or G8635 or G8650);
	G13143<= not (G8636 or G8654 or G8666);
	G13149<= not (G8676 or G8687 or G8703);
	G13155<= not (G8688 or G8705 or G8722);
	G13160<= not (G8704 or G8717 or G8751);
	G13164<= not (G8706 or G8724 or G8760);
	G13171<= not (G8723 or G8755 or G8774);
	G13175<= not (G8725 or G8762 or G8783);
	G13182<= not (G8761 or G8778 or G8797);
	G13194<= not (G8784 or G8801 or G8816);
	G13228<= not (G8841 or G8861 or G8892);
	G13251<= not (G8868 or G8899 or G8932);
	G13274<= not (G8906 or G8939 or G8972);
	G13286<= not (G11481 or G11332 or G11190 or G7880);
	G13299<= not (G8946 or G8979 or G9004);
	G13310<= not (G11481 or G11332 or G11190 or G11069);
	G13313<= not (G8183 or G11332 or G11190 or G7880);
	G13331<= not (G8183 or G11332 or G11190 or G11069);
	G13332<= not (G11481 or G8045 or G11190 or G7880);
	G13353<= not (G11481 or G8045 or G11190 or G11069);
	G13354<= not (G8183 or G8045 or G11190 or G7880);
	G13374<= not (G8183 or G8045 or G11190 or G11069);
	G13375<= not (G11481 or G11332 or G7928 or G7880);
	G13378<= not (G9026 or G9047 or G9061);
	G13401<= not (G11481 or G11332 or G7928 or G11069);
	G13404<= not (G8183 or G11332 or G7928 or G7880);
	G15661<= not (G11737 or G7345);
	G15797<= not (G13305 or G7143);
	G15873<= not (G11617 or G7562);
	G15959<= not (G2814 or G13082);
	G15978<= not (G11737 or G7152);
	G16020<= not (G6200 or G12457 or G10952);
	G16036<= not (G6289 or G12467 or G10952);
	G16058<= not (G6426 or G12482 or G10952);
	G16082<= not (G10952 or G6140 or G12487);
	G16094<= not (G6631 or G12499 or G10952);
	G16120<= not (G10952 or G6161 or G12507);
	G16171<= not (G10952 or G6188 or G12524);
	G16230<= not (G10952 or G6220 or G12539);
	G16498<= not (G14158 or G14347);
	G16520<= not (G14273 or G14459);
	G16551<= not (G14395 or G14546);
	G16567<= not (G15904 or G15880 or G15859);
	G16570<= not (G15904 or G15880 or G14630);
	G16583<= not (G14507 or G14601);
	G16591<= not (G15933 or G15913 or G15890);
	G16594<= not (G15933 or G15913 or G14650);
	G16611<= not (G15962 or G15942 or G15923);
	G16614<= not (G15962 or G15942 or G14677);
	G16629<= not (G15981 or G15971 or G15952);
	G16632<= not (G15981 or G15971 or G14711);
	G16643<= not (G15904 or G14642 or G15859);
	G16654<= not (G14690 or G12477);
	G16655<= not (G15933 or G14669 or G15890);
	G16671<= not (G14724 or G12494);
	G16672<= not (G15962 or G14703 or G15923);
	G16679<= not (G14797 or G14895);
	G16692<= not (G14752 or G12514);
	G16693<= not (G15981 or G14737 or G15952);
	G16705<= not (G14849 or G14976);
	G16718<= not (G14773 or G12531);
	G16736<= not (G14922 or G15065);
	G16778<= not (G15003 or G15161);
	G16802<= not (G13469 or G3897);
	G16803<= not (G15593 or G12908);
	G16823<= not (G5362 or G13469);
	G16824<= not (G15658 or G12938);
	G16829<= not (G14956 or G12564);
	G16835<= not (G15717 or G12966);
	G16841<= not (G15021 or G12607);
	G16844<= not (G15754 or G12989);
	G16845<= not (G15755 or G12990);
	G16847<= not (G15095 or G12650);
	G16851<= not (G15781 or G13000);
	G16853<= not (G15801 or G13009);
	G16854<= not (G15802 or G13010);
	G16857<= not (G15817 or G13023);
	G16860<= not (G15828 or G13031);
	G16861<= not (G15829 or G13032);
	G16866<= not (G15840 or G13042);
	G16880<= not (G15852 or G13056);
	G17012<= not (G14657 or G14642 or G15859);
	G17025<= not (G15904 or G15880 or G15859);
	G17042<= not (G14691 or G14669 or G15890);
	G17051<= not (G14657 or G15880 or G14630);
	G17059<= not (G15933 or G15913 or G15890);
	G17076<= not (G14725 or G14703 or G15923);
	G17086<= not (G14691 or G15913 or G14650);
	G17094<= not (G15962 or G15942 or G15923);
	G17111<= not (G14753 or G14737 or G15952);
	G17124<= not (G14725 or G15942 or G14677);
	G17132<= not (G15981 or G15971 or G15952);
	G17151<= not (G14753 or G15971 or G14711);
	G17186<= not (G7949 or G14144);
	G17197<= not (G8000 or G14259);
	G17204<= not (G8075 or G14381);
	G17209<= not (G8160 or G14493);
	G17213<= not (G4326 or G14442);
	G17215<= not (G15904 or G14642);
	G17216<= not (G4495 or G14529);
	G17218<= not (G15933 or G14669);
	G17219<= not (G4671 or G14584);
	G17220<= not (G15962 or G14703);
	G17221<= not (G4848 or G14618);
	G17222<= not (G15998 or G16003);
	G17223<= not (G15981 or G14737);
	G17224<= not (G16004 or G16009);
	G17225<= not (G16008 or G16015);
	G17226<= not (G16010 or G16017);
	G17228<= not (G16016 or G16029);
	G17229<= not (G16019 or G16032);
	G17234<= not (G16028 or G16045);
	G17235<= not (G16030 or G16047);
	G17236<= not (G16033 or G16051);
	G17246<= not (G16046 or G16066);
	G17247<= not (G16050 or G16070);
	G17248<= not (G16052 or G16072);
	G17269<= not (G16067 or G16100);
	G17270<= not (G16071 or G16104);
	G17271<= not (G16073 or G16106);
	G17302<= not (G16103 or G16135);
	G17303<= not (G16105 or G16137);
	G17340<= not (G16136 or G16183);
	G17341<= not (G16138 or G16185);
	G17383<= not (G16184 or G16238);
	G17429<= not (G16239 or G16288);
	G17507<= not (G16298 or G13318);
	G17896<= not (G14352 or G16020);
	G18007<= not (G14464 or G16036);
	G18085<= not (G16085 or G6363);
	G18124<= not (G14551 or G16058);
	G18201<= not (G16123 or G6568);
	G18240<= not (G14606 or G16094);
	G18308<= not (G16174 or G6832);
	G18352<= not (G16082 or G14249);
	G18401<= not (G16233 or G7134);
	G18430<= not (G16020 or G14352);
	G18447<= not (G16120 or G14371);
	G18503<= not (G16036 or G14464);
	G18520<= not (G16171 or G14483);
	G18548<= not (G14249 or G16082);
	G18567<= not (G16058 or G14551);
	G18584<= not (G16230 or G14570);
	G18590<= not (G16439 or G7522);
	G18598<= not (G14371 or G16120);
	G18617<= not (G16094 or G14606);
	G18623<= not (G15902 or G2814);
	G18626<= not (G16463 or G7549);
	G18630<= not (G14483 or G16171);
	G18639<= not (G14570 or G16230);
	G18669<= not (G13623 or G13634);
	G18678<= not (G13625 or G11771);
	G18707<= not (G13636 or G11788);
	G18719<= not (G13643 or G13656);
	G18726<= not (G13645 or G11805);
	G18743<= not (G13648 or G11814);
	G18754<= not (G13655 or G11816);
	G18755<= not (G13871 or G12274);
	G18763<= not (G13671 or G11838);
	G18780<= not (G13674 or G11847);
	G18781<= not (G13675 or G11851);
	G18782<= not (G13676 or G13705);
	G18794<= not (G13701 or G11880);
	G18803<= not (G13704 or G11885);
	G18804<= not (G13905 or G12331);
	G18820<= not (G13738 or G11922);
	G18821<= not (G13740 or G11926);
	G18835<= not (G13788 or G11966);
	G18836<= not (G13789 or G11967);
	G18837<= not (G13998 or G12376);
	G18852<= not (G13815 or G12012);
	G18866<= not (G13834 or G12069);
	G18867<= not (G13835 or G12070);
	G18868<= not (G14143 or G12419);
	G18883<= not (G13846 or G12128);
	G18885<= not (G13847 or G12129);
	G18906<= not (G13855 or G12186);
	G18907<= not (G14336 or G12429);
	G18942<= not (G13870 or G12273);
	G18957<= not (G13884 or G12307);
	G18968<= not (G13904 or G12330);
	G18975<= not (G13944 or G12353);
	G19144<= not (G17268 or G14884);
	G19149<= not (G17339 or G15020);
	G19153<= not (G17381 or G15093);
	G19154<= not (G17382 or G15094);
	G19157<= not (G17428 or G15171);
	G19160<= not (G17446 or G15178);
	G19162<= not (G17485 or G15243);
	G19163<= not (G17486 or G15244);
	G19165<= not (G17526 or G15264);
	G19167<= not (G17556 or G15320);
	G19171<= not (G17616 or G15356);
	G19172<= not (G17635 or G15388);
	G19173<= not (G17636 or G15389);
	G19177<= not (G17713 or G15442);
	G19178<= not (G17718 or G15452);
	G19179<= not (G17719 or G15453);
	G19184<= not (G17798 or G15520);
	G19219<= not (G18165 or G15753);
	G20008<= not (G18977 or G7338);
	G20054<= not (G19001 or G16867);
	G20095<= not (G16507 or G16895);
	G20120<= not (G16529 or G16924);
	G20150<= not (G16560 or G16954);
	G20153<= not (G16536 or G7583);
	G20299<= not (G16665 or G16884);
	G20310<= not (G16850 or G13654);
	G20314<= not (G13646 or G16855);
	G20318<= not (G16686 or G16913);
	G20333<= not (G13672 or G16859);
	G20337<= not (G16712 or G16943);
	G20343<= not (G16856 or G13703);
	G20353<= not (G13702 or G16864);
	G20357<= not (G16743 or G16974);
	G20375<= not (G13739 or G16879);
	G20376<= not (G16865 or G13787);
	G20417<= not (G16907 or G13833);
	G20682<= not (G19160 or G10024);
	G20717<= not (G19165 or G10133);
	G20752<= not (G19171 or G10238);
	G20789<= not (G19177 or G10340);
	G20841<= not (G14767 or G19552);
	G20874<= not (G17301 or G19594);
	G20875<= not (G19584 or G17352);
	G20876<= not (G19585 or G17353);
	G20877<= not (G3919 or G19830);
	G20878<= not (G19600 or G17395);
	G20879<= not (G19601 or G17396);
	G20880<= not (G19602 or G17397);
	G20881<= not (G19603 or G17398);
	G20882<= not (G19614 or G17408);
	G20883<= not (G19615 or G17409);
	G20884<= not (G5394 or G19830);
	G20891<= not (G19626 or G17447);
	G20892<= not (G19627 or G17448);
	G20893<= not (G19628 or G17449);
	G20894<= not (G19629 or G17450);
	G20895<= not (G19633 or G17461);
	G20896<= not (G19634 or G17462);
	G20897<= not (G19635 or G17463);
	G20898<= not (G19636 or G17464);
	G20899<= not (G19647 or G17474);
	G20900<= not (G19648 or G17475);
	G20901<= not (G19660 or G17508);
	G20902<= not (G19661 or G17509);
	G20903<= not (G19662 or G17510);
	G20910<= not (G19666 or G17527);
	G20911<= not (G19667 or G17528);
	G20912<= not (G19668 or G17529);
	G20913<= not (G19669 or G17530);
	G20914<= not (G19673 or G17541);
	G20915<= not (G19674 or G17542);
	G20916<= not (G19675 or G17543);
	G20917<= not (G19676 or G17544);
	G20918<= not (G19687 or G17554);
	G20919<= not (G19688 or G17555);
	G20920<= not (G19691 or G19726);
	G20921<= not (G19697 or G17576);
	G20922<= not (G19698 or G17577);
	G20923<= not (G19699 or G17578);
	G20924<= not (G19700 or G15257);
	G20925<= not (G19708 or G17598);
	G20926<= not (G19709 or G17599);
	G20927<= not (G19710 or G17600);
	G20934<= not (G19714 or G17617);
	G20935<= not (G19715 or G17618);
	G20936<= not (G19716 or G17619);
	G20937<= not (G19717 or G17620);
	G20938<= not (G19721 or G17631);
	G20939<= not (G19722 or G17632);
	G20940<= not (G19723 or G17633);
	G20941<= not (G19724 or G17634);
	G20944<= not (G19731 or G17652);
	G20945<= not (G19732 or G17653);
	G20946<= not (G19733 or G17654);
	G20947<= not (G19734 or G15335);
	G20948<= not (G19735 or G15336);
	G20949<= not (G19741 or G17673);
	G20950<= not (G19742 or G17674);
	G20951<= not (G19743 or G17675);
	G20952<= not (G19744 or G15349);
	G20953<= not (G19752 or G17695);
	G20954<= not (G19753 or G17696);
	G20955<= not (G19754 or G17697);
	G20962<= not (G19758 or G17714);
	G20963<= not (G19759 or G17715);
	G20964<= not (G19760 or G17716);
	G20965<= not (G19761 or G17717);
	G20966<= not (G19765 or G17734);
	G20967<= not (G19766 or G17735);
	G20968<= not (G19767 or G17736);
	G20969<= not (G19768 or G15402);
	G20970<= not (G19769 or G15403);
	G20972<= not (G19774 or G17752);
	G20973<= not (G19775 or G17753);
	G20974<= not (G19776 or G17754);
	G20975<= not (G19777 or G15421);
	G20976<= not (G19778 or G15422);
	G20977<= not (G19784 or G17773);
	G20978<= not (G19785 or G17774);
	G20979<= not (G19786 or G17775);
	G20980<= not (G19787 or G15435);
	G20981<= not (G19795 or G17795);
	G20982<= not (G19796 or G17796);
	G20983<= not (G19797 or G17797);
	G20989<= not (G19802 or G17812);
	G20990<= not (G19803 or G17813);
	G20991<= not (G19804 or G17814);
	G20992<= not (G19805 or G15470);
	G20993<= not (G19807 or G17835);
	G20994<= not (G19808 or G17836);
	G20995<= not (G19809 or G17837);
	G20996<= not (G19810 or G15486);
	G20997<= not (G19811 or G15487);
	G20999<= not (G19816 or G17853);
	G21000<= not (G19817 or G17854);
	G21001<= not (G19818 or G17855);
	G21002<= not (G19819 or G15505);
	G21003<= not (G19820 or G15506);
	G21004<= not (G19826 or G17874);
	G21005<= not (G19827 or G17875);
	G21006<= not (G19828 or G17876);
	G21007<= not (G19829 or G15519);
	G21008<= not (G19836 or G17877);
	G21009<= not (G19839 or G17900);
	G21010<= not (G19840 or G17901);
	G21011<= not (G19841 or G17902);
	G21015<= not (G19846 or G17924);
	G21016<= not (G19847 or G17925);
	G21017<= not (G19848 or G17926);
	G21018<= not (G19849 or G15556);
	G21019<= not (G19851 or G17947);
	G21020<= not (G19852 or G17948);
	G21021<= not (G19853 or G17949);
	G21022<= not (G19854 or G15572);
	G21023<= not (G19855 or G15573);
	G21025<= not (G19860 or G17965);
	G21026<= not (G19861 or G17966);
	G21027<= not (G19862 or G17967);
	G21028<= not (G19863 or G15591);
	G21029<= not (G19864 or G15592);
	G21031<= not (G19869 or G17989);
	G21032<= not (G19870 or G17990);
	G21033<= not (G19872 or G18011);
	G21034<= not (G19873 or G18012);
	G21035<= not (G19874 or G18013);
	G21039<= not (G19879 or G18035);
	G21040<= not (G19880 or G18036);
	G21041<= not (G19881 or G18037);
	G21042<= not (G19882 or G15634);
	G21043<= not (G19884 or G18058);
	G21044<= not (G19885 or G18059);
	G21045<= not (G19886 or G18060);
	G21046<= not (G19887 or G15650);
	G21047<= not (G19888 or G15651);
	G21048<= not (G19889 or G18062);
	G21051<= not (G19895 or G18088);
	G21052<= not (G19900 or G18106);
	G21053<= not (G19901 or G18107);
	G21054<= not (G19903 or G18128);
	G21055<= not (G19904 or G18129);
	G21056<= not (G19905 or G18130);
	G21060<= not (G19910 or G18152);
	G21061<= not (G19911 or G18153);
	G21062<= not (G19912 or G18154);
	G21063<= not (G19913 or G15710);
	G21065<= not (G19914 or G18169);
	G21070<= not (G19920 or G18204);
	G21071<= not (G19925 or G18222);
	G21072<= not (G19926 or G18223);
	G21073<= not (G19928 or G18244);
	G21074<= not (G19929 or G18245);
	G21075<= not (G19930 or G18246);
	G21080<= not (G19935 or G18311);
	G21081<= not (G19940 or G18329);
	G21082<= not (G19941 or G18330);
	G21083<= not (G19943 or G18333);
	G21084<= not (G20011 or G20048);
	G21094<= not (G19952 or G18404);
	G21095<= not (G20012 or G20049 or G20084);
	G21096<= not (G20013 or G20051 or G20087);
	G21104<= not (G20050 or G20085 or G20106);
	G21105<= not (G20052 or G20088 or G20109);
	G21106<= not (G20053 or G20090 or G20112);
	G21116<= not (G20086 or G20107 or G20131);
	G21117<= not (G20089 or G20110 or G20133);
	G21118<= not (G20091 or G20113 or G20136);
	G21119<= not (G20092 or G20115 or G20139);
	G21133<= not (G20108 or G20132 or G20156);
	G21134<= not (G20111 or G20134 or G20157);
	G21135<= not (G20114 or G20137 or G20160);
	G21147<= not (G20135 or G20158 or G20188);
	G21148<= not (G20138 or G20161 or G20190);
	G21149<= not (G20015 or G19981);
	G21167<= not (G20159 or G20189);
	G21168<= not (G20162 or G20191 or G20220);
	G21169<= not (G20057 or G20019);
	G21183<= not (G20192 or G20221);
	G21189<= not (G20098 or G20061);
	G21204<= not (G20123 or G20102);
	G21211<= not (G19240 or G19230);
	G21219<= not (G19253 or G19243);
	G21227<= not (G18414 or G18485 or G20295);
	G21228<= not (G19388 or G17118);
	G21230<= not (G19266 or G19256);
	G21233<= not (G19418 or G17145);
	G21235<= not (G19281 or G19269);
	G21238<= not (G19954 or G5890);
	G21242<= not (G19455 or G17168);
	G21246<= not (G19984 or G5929);
	G21250<= not (G19482 or G17183);
	G21255<= not (G20022 or G5963);
	G21263<= not (G20064 or G5992);
	G21316<= not (G20460 or G16111);
	G21331<= not (G20472 or G16153);
	G21346<= not (G20480 or G13247);
	G21364<= not (G20486 or G13266);
	G21385<= not (G20492 or G13289);
	G21407<= not (G20499 or G13316);
	G21432<= not (G20502 or G13335);
	G21435<= not (G20503 or G16385);
	G21467<= not (G20506 or G13355);
	G21470<= not (G20512 or G16417);
	G21502<= not (G20525 or G16445);
	G21615<= not (G16567 or G19957);
	G21618<= not (G20016 or G14079 or G14165);
	G21636<= not (G20473 or G6513);
	G21643<= not (G16591 or G19987);
	G21646<= not (G20058 or G14194 or G14280);
	G21665<= not (G20507 or G18352);
	G21667<= not (G20481 or G6777);
	G21674<= not (G16611 or G20025);
	G21677<= not (G20099 or G14309 or G14402);
	G21694<= not (G20526 or G18447);
	G21696<= not (G20487 or G7079);
	G21703<= not (G16629 or G20067);
	G21706<= not (G20124 or G14431 or G14514);
	G21711<= not (G19830 or G15780);
	G21730<= not (G20545 or G18520);
	G21732<= not (G20493 or G7329);
	G21738<= not (G19444 or G17893 or G14079);
	G21739<= not (G20507 or G18430);
	G21756<= not (G19070 or G18584);
	G21762<= not (G19471 or G18004 or G14194);
	G21763<= not (G20526 or G18503);
	G21778<= not (G19494 or G18121 or G14309);
	G21779<= not (G20545 or G18567);
	G21793<= not (G19515 or G18237 or G14431);
	G21794<= not (G19070 or G18617);
	G21796<= not (G19830 or G13004);
	G21842<= not (G13609 or G19150);
	G21843<= not (G13619 or G19155);
	G21845<= not (G13631 or G19161);
	G21847<= not (G13642 or G19166);
	G21851<= not (G19252 or G8842);
	G21878<= not (G16964 or G19228);
	G21880<= not (G13854 or G19236);
	G21882<= not (G13862 or G19248);
	G21884<= not (G19260 or G19284);
	G21887<= not (G13519 or G19289);
	G21889<= not (G19285 or G19316);
	G21890<= not (G13530 or G19307);
	G21893<= not (G13541 or G19328);
	G21894<= not (G19317 or G19356);
	G21901<= not (G13552 or G19355);
	G21968<= not (G21234 or G19476);
	G21969<= not (G20895 or G10133);
	G21970<= not (G17182 or G21226);
	G21971<= not (G21243 or G19499);
	G21972<= not (G20914 or G10238);
	G21973<= not (G21251 or G19520);
	G21974<= not (G20938 or G10340);
	G21975<= not (G21245 or G21259);
	G21980<= not (G21252 or G19531 or G19540);
	G21981<= not (G21254 or G21267);
	G21987<= not (G21260 or G19541 or G19544);
	G21988<= not (G21262 or G21276);
	G22000<= not (G21268 or G19545 or G19547);
	G22001<= not (G21270 or G21283);
	G22013<= not (G21277 or G19548 or G19551);
	G22025<= not (G21284 or G19549);
	G22026<= not (G21083 or G18407);
	G22027<= not (G21290 or G19553);
	G22028<= not (G21291 or G19554);
	G22029<= not (G21292 or G19555);
	G22030<= not (G21298 or G19557);
	G22031<= not (G21299 or G19558);
	G22032<= not (G21300 or G19559);
	G22033<= not (G21301 or G19560);
	G22034<= not (G21302 or G19561);
	G22035<= not (G21303 or G19562);
	G22037<= not (G21304 or G19564);
	G22038<= not (G21305 or G19565);
	G22039<= not (G21306 or G19566);
	G22040<= not (G21307 or G19567);
	G22041<= not (G21308 or G19568);
	G22042<= not (G21309 or G19569);
	G22043<= not (G21310 or G19570);
	G22044<= not (G21311 or G19571);
	G22045<= not (G21312 or G19572);
	G22047<= not (G21313 or G19574);
	G22048<= not (G21314 or G19575);
	G22049<= not (G21315 or G19576);
	G22054<= not (G21319 or G19586);
	G22055<= not (G21320 or G19587);
	G22056<= not (G21321 or G19588);
	G22057<= not (G21322 or G19589);
	G22058<= not (G21323 or G19590);
	G22059<= not (G21324 or G19591);
	G22060<= not (G21325 or G19592);
	G22061<= not (G21326 or G19593);
	G22063<= not (G21328 or G19597);
	G22064<= not (G21329 or G19598);
	G22065<= not (G21330 or G19599);
	G22066<= not (G21334 or G19604);
	G22067<= not (G21335 or G19605);
	G22068<= not (G21336 or G19606);
	G22073<= not (G21337 or G19616);
	G22074<= not (G21338 or G19617);
	G22075<= not (G21339 or G19618);
	G22076<= not (G21340 or G19619);
	G22077<= not (G21341 or G19620);
	G22078<= not (G21342 or G19621);
	G22079<= not (G21343 or G19623);
	G22080<= not (G21344 or G19624);
	G22081<= not (G21345 or G19625);
	G22087<= not (G21349 or G19630);
	G22088<= not (G21350 or G19631);
	G22089<= not (G21351 or G19632);
	G22090<= not (G21352 or G19637);
	G22091<= not (G21353 or G19638);
	G22092<= not (G21354 or G19639);
	G22097<= not (G21355 or G19649);
	G22098<= not (G21356 or G19650);
	G22099<= not (G21357 or G19651);
	G22100<= not (G21360 or G19653);
	G22101<= not (G21361 or G19654);
	G22102<= not (G21362 or G19655);
	G22103<= not (G21363 or G19656);
	G22104<= not (G21367 or G19663);
	G22105<= not (G21368 or G19664);
	G22106<= not (G21369 or G19665);
	G22112<= not (G21370 or G19670);
	G22113<= not (G21371 or G19671);
	G22114<= not (G21372 or G19672);
	G22115<= not (G21373 or G19677);
	G22116<= not (G21374 or G19678);
	G22117<= not (G21375 or G19679);
	G22122<= not (G21378 or G19692);
	G22123<= not (G21379 or G19693);
	G22124<= not (G21380 or G19694);
	G22125<= not (G21381 or G19695);
	G22126<= not (G21389 or G19701);
	G22127<= not (G21390 or G19702);
	G22128<= not (G21391 or G19703);
	G22129<= not (G21392 or G19704);
	G22130<= not (G21393 or G19711);
	G22131<= not (G21394 or G19712);
	G22132<= not (G21395 or G19713);
	G22138<= not (G21396 or G19718);
	G22139<= not (G21397 or G19719);
	G22140<= not (G21398 or G19720);
	G22141<= not (G21401 or G19727);
	G22142<= not (G21402 or G19728);
	G22143<= not (G21403 or G19729);
	G22144<= not (G21410 or G19730);
	G22145<= not (G21411 or G19736);
	G22146<= not (G21412 or G19737);
	G22147<= not (G21413 or G19738);
	G22148<= not (G21414 or G19739);
	G22149<= not (G21419 or G19745);
	G22150<= not (G21420 or G19746);
	G22151<= not (G21421 or G19747);
	G22152<= not (G21422 or G19748);
	G22153<= not (G21423 or G19755);
	G22154<= not (G21424 or G19756);
	G22155<= not (G21425 or G19757);
	G22161<= not (G21428 or G19764);
	G22162<= not (G21438 or G19770);
	G22163<= not (G21439 or G19771);
	G22164<= not (G21440 or G19772);
	G22165<= not (G21444 or G19773);
	G22166<= not (G21445 or G19779);
	G22167<= not (G21446 or G19780);
	G22168<= not (G21447 or G19781);
	G22169<= not (G21448 or G19782);
	G22170<= not (G21453 or G19788);
	G22171<= not (G21454 or G19789);
	G22172<= not (G21455 or G19790);
	G22173<= not (G21456 or G19791);
	G22174<= not (G19868 or G21593);
	G22177<= not (G21476 or G19806);
	G22178<= not (G21480 or G19812);
	G22179<= not (G21481 or G19813);
	G22180<= not (G21482 or G19814);
	G22181<= not (G21486 or G19815);
	G22182<= not (G21487 or G19821);
	G22183<= not (G21488 or G19822);
	G22184<= not (G21489 or G19823);
	G22185<= not (G21490 or G19824);
	G22186<= not (G21497 or G19837);
	G22189<= not (G19899 or G21622);
	G22191<= not (G21517 or G19850);
	G22192<= not (G21521 or G19856);
	G22193<= not (G21522 or G19857);
	G22194<= not (G21523 or G19858);
	G22195<= not (G21527 or G19859);
	G22198<= not (G19924 or G21650);
	G22200<= not (G21553 or G19883);
	G22204<= not (G19939 or G21681);
	G22210<= not (G21610 or G19932);
	G22216<= not (G21635 or G19944);
	G22218<= not (G21639 or G19949);
	G22227<= not (G21658 or G19953);
	G22231<= not (G21666 or G19971);
	G22234<= not (G21670 or G19976);
	G22242<= not (G21687 or G19983);
	G22247<= not (G21695 or G20001);
	G22249<= not (G21699 or G20006);
	G22263<= not (G21723 or G20021);
	G22267<= not (G21731 or G20039);
	G22269<= not (G21735 or G20044);
	G22280<= not (G21749 or G20063);
	G22284<= not (G21757 or G20081);
	G22288<= not (G20144 or G21805);
	G22299<= not (G21773 or G20104);
	G22308<= not (G20182 or G21812);
	G22336<= not (G20216 or G21818);
	G22361<= not (G20246 or G21822);
	G22454<= not (G17012 or G21891);
	G22493<= not (G17042 or G21899);
	G22536<= not (G17076 or G21911);
	G22576<= not (G17111 or G21925);
	G22578<= not (G21892 or G18982);
	G22615<= not (G21900 or G18990);
	G22651<= not (G21912 or G18997);
	G22687<= not (G21926 or G19010);
	G22755<= not (G21271 or G20842);
	G22784<= not (G16075 or G20885);
	G22789<= not (G21278 or G20850);
	G22810<= not (G16075 or G20842 or G21271);
	G22826<= not (G16113 or G20904);
	G22831<= not (G21285 or G20858);
	G22851<= not (G16113 or G20850 or G21278);
	G22865<= not (G16164 or G20928);
	G22870<= not (G21293 or G20866);
	G22886<= not (G16164 or G20858 or G21285);
	G22900<= not (G16223 or G20956);
	G22921<= not (G16223 or G20866 or G21293);
	G22935<= not (G21903 or G7466);
	G22953<= not (G20700 or G7595);
	G22985<= not (G21618 or G21049);
	G22987<= not (G21646 or G21068);
	G22990<= not (G21677 or G21078);
	G22997<= not (G21706 or G21092);
	G22999<= not (G21085 or G19241);
	G23000<= not (G16909 or G21067);
	G23009<= not (G21738 or G21107);
	G23013<= not (G21097 or G19254);
	G23014<= not (G16939 or G21077);
	G23022<= not (G16968 or G21086);
	G23023<= not (G14256 or G14175 or G21123);
	G23025<= not (G21762 or G21124);
	G23029<= not (G21111 or G19267);
	G23030<= not (G16970 or G21091);
	G23039<= not (G16989 or G21098);
	G23040<= not (G14378 or G14290 or G21142);
	G23042<= not (G21778 or G21143);
	G23046<= not (G21128 or G19282);
	G23047<= not (G16991 or G21103);
	G23051<= not (G21121 or G21153);
	G23058<= not (G16999 or G21112);
	G23059<= not (G14490 or G14412 or G21162);
	G23061<= not (G21793 or G21163);
	G23066<= not (G21138 or G19303 or G19320);
	G23067<= not (G17015 or G21122);
	G23070<= not (G21140 or G21173);
	G23076<= not (G17023 or G21129);
	G23077<= not (G14577 or G14524 or G21182);
	G23080<= not (G21158 or G19324 or G19347);
	G23081<= not (G17045 or G21141);
	G23083<= not (G21160 or G21193);
	G23092<= not (G17055 or G21154);
	G23093<= not (G17056 or G21155);
	G23096<= not (G21178 or G19351 or G19381);
	G23097<= not (G17079 or G21161);
	G23099<= not (G21180 or G21208);
	G23110<= not (G17090 or G21174);
	G23111<= not (G17091 or G21175);
	G23113<= not (G21198 or G19385 or G19413);
	G23114<= not (G17114 or G21181);
	G23117<= not (G17117 or G21188);
	G23123<= not (G17128 or G21194);
	G23124<= not (G17129 or G21195);
	G23126<= not (G17144 or G21203);
	G23132<= not (G17155 or G21209);
	G23133<= not (G17156 or G21210);
	G23135<= not (G21229 or G19449);
	G23136<= not (G20878 or G10024);
	G23137<= not (G17167 or G21218);
	G23324<= not (G22144 or G10024);
	G23329<= not (G22165 or G10133);
	G23330<= not (G22186 or G22777);
	G23339<= not (G22181 or G10238);
	G23348<= not (G22195 or G10340);
	G23357<= not (G22210 or G20127);
	G23358<= not (G22227 or G18407);
	G23359<= not (G22216 or G22907);
	G23385<= not (G17393 or G22517);
	G23386<= not (G22483 or G21388);
	G23392<= not (G17460 or G22557);
	G23393<= not (G22526 or G21418);
	G23399<= not (G17506 or G22581);
	G23400<= not (G17540 or G22597);
	G23401<= not (G22566 or G21452);
	G23406<= not (G17597 or G22618);
	G23407<= not (G17630 or G22634);
	G23408<= not (G22606 or G21494);
	G23413<= not (G17694 or G22654);
	G23418<= not (G17794 or G22690);
	G23427<= not (G22699 or G21589);
	G23433<= not (G22726 or G21611);
	G23461<= not (G22841 or G21707);
	G23477<= not (G22906 or G21758);
	G23497<= not (G22876 or G5606);
	G23513<= not (G22911 or G5631);
	G23528<= not (G22936 or G5659);
	G23539<= not (G22942 or G5697);
	G23545<= not (G22984 or G20285);
	G23823<= not (G23009 or G18490 or G4456);
	G23858<= not (G23025 or G18554 or G4632);
	G23892<= not (G23042 or G18604 or G4809);
	G23913<= not (G23061 or G18636 or G4985);
	G23922<= not (G4456 or G22985);
	G23945<= not (G4456 or G13565 or G23009);
	G23950<= not (G22992 or G6707);
	G23954<= not (G4632 or G22987);
	G23974<= not (G4632 or G13573 or G23025);
	G23979<= not (G23003 or G7009);
	G23983<= not (G4809 or G22990);
	G24004<= not (G4809 or G13582 or G23042);
	G24009<= not (G23017 or G7259);
	G24013<= not (G4985 or G22997);
	G24038<= not (G4985 or G13602 or G23061);
	G24043<= not (G23033 or G7455);
	G24059<= not (G21990 or G20809);
	G24072<= not (G22004 or G20826);
	G24083<= not (G22015 or G20836);
	G24092<= not (G22020 or G20840);
	G24174<= not (G16894 or G22206);
	G24178<= not (G16908 or G22211);
	G24179<= not (G16923 or G22214);
	G24181<= not (G16938 or G22220);
	G24182<= not (G16953 or G22223);
	G24206<= not (G16966 or G22228);
	G24207<= not (G16967 or G22229);
	G24208<= not (G16969 or G22235);
	G24209<= not (G16984 or G22238);
	G24212<= not (G16987 or G22244);
	G24213<= not (G16988 or G22245);
	G24214<= not (G16990 or G22250);
	G24215<= not (G16993 or G22254);
	G24216<= not (G16994 or G22255);
	G24218<= not (G16997 or G22264);
	G24219<= not (G16998 or G22265);
	G24222<= not (G17017 or G22272);
	G24223<= not (G17018 or G22273);
	G24225<= not (G17021 or G22281);
	G24226<= not (G17022 or G22282);
	G24227<= not (G22270 or G21137);
	G24228<= not (G17028 or G22285);
	G24230<= not (G17047 or G22291);
	G24231<= not (G17048 or G22292);
	G24232<= not (G22637 or G22665);
	G24234<= not (G22289 or G21157);
	G24235<= not (G17062 or G22305);
	G24237<= not (G17081 or G22311);
	G24238<= not (G17082 or G22312);
	G24242<= not (G22309 or G21177);
	G24243<= not (G17097 or G22333);
	G24249<= not (G22337 or G21197);
	G24250<= not (G17135 or G22358);
	G24426<= not (G23386 or G10024);
	G24428<= not (G23544 or G22398);
	G24430<= not (G23393 or G10133);
	G24434<= not (G23401 or G10238);
	G24438<= not (G23408 or G10340);
	G24445<= not (G23427 or G22777);
	G24446<= not (G23433 or G22907);
	G24473<= not (G23461 or G18407);
	G24476<= not (G23477 or G20127);
	G24479<= not (G23593 or G22516);
	G24480<= not (G23617 or G23659);
	G24481<= not (G23618 or G19696);
	G24485<= not (G23625 or G22556);
	G24486<= not (G23643 or G22577);
	G24487<= not (G23666 or G23709);
	G24488<= not (G23667 or G19740);
	G24489<= not (G23674 or G22596);
	G24490<= not (G23686 or G22607);
	G24491<= not (G15247 or G23735);
	G24492<= not (G23689 or G22610);
	G24493<= not (G23693 or G22614);
	G24494<= not (G23716 or G23763);
	G24495<= not (G23717 or G19783);
	G24496<= not (G23724 or G22633);
	G24497<= not (G23734 or G22638);
	G24498<= not (G15324 or G23777);
	G24499<= not (G15325 or G23778);
	G24500<= not (G23740 or G22643);
	G24501<= not (G15339 or G23790);
	G24502<= not (G23743 or G22646);
	G24503<= not (G23747 or G22650);
	G24504<= not (G23770 or G23818);
	G24505<= not (G23771 or G19825);
	G24506<= not (G23776 or G22667);
	G24507<= not (G15391 or G23824);
	G24508<= not (G15392 or G23825);
	G24509<= not (G23789 or G22674);
	G24510<= not (G15410 or G23830);
	G24511<= not (G15411 or G23831);
	G24512<= not (G23795 or G22679);
	G24513<= not (G15425 or G23843);
	G24514<= not (G23798 or G22682);
	G24515<= not (G23802 or G22686);
	G24516<= not (G23820 or G22700);
	G24517<= not (G23822 or G22701);
	G24519<= not (G15459 or G23855);
	G24520<= not (G23829 or G22707);
	G24521<= not (G15475 or G23859);
	G24522<= not (G15476 or G23860);
	G24523<= not (G23842 or G22714);
	G24524<= not (G15494 or G23865);
	G24525<= not (G15495 or G23866);
	G24526<= not (G23848 or G22719);
	G24527<= not (G15509 or G23878);
	G24528<= not (G23851 or G22722);
	G24530<= not (G23857 or G22732);
	G24532<= not (G15545 or G23889);
	G24533<= not (G23864 or G22738);
	G24534<= not (G15561 or G23893);
	G24535<= not (G15562 or G23894);
	G24536<= not (G23877 or G22745);
	G24537<= not (G15580 or G23899);
	G24538<= not (G15581 or G23900);
	G24543<= not (G23891 or G22764);
	G24545<= not (G15623 or G23910);
	G24546<= not (G23898 or G22770);
	G24547<= not (G15639 or G23914);
	G24548<= not (G15640 or G23915);
	G24555<= not (G23912 or G22798);
	G24557<= not (G15699 or G23942);
	G24558<= not (G23917 or G22804);
	G24566<= not (G23944 or G22842);
	G24575<= not (G23972 or G22874);
	G24606<= not (G24183 or G537);
	G24613<= not (G23592 or G22515);
	G24622<= not (G23616 or G22546);
	G24623<= not (G24183 or G529);
	G24624<= not (G23624 or G22555);
	G24636<= not (G24183 or G530);
	G24637<= not (G23665 or G22587);
	G24638<= not (G23673 or G22595);
	G24652<= not (G24183 or G531);
	G24656<= not (G23715 or G22624);
	G24657<= not (G23723 or G22632);
	G24663<= not (G24183 or G532);
	G24675<= not (G23769 or G22660);
	G24681<= not (G24183 or G533);
	G24682<= not (G23688 or G24183);
	G24694<= not (G24183 or G534);
	G24708<= not (G23854 or G22727);
	G24711<= not (G24183 or G536);
	G24717<= not (G23886 or G22754);
	G24720<= not (G23888 or G22759);
	G24728<= not (G23907 or G22788);
	G24731<= not (G23909 or G22793);
	G24736<= not (G23939 or G22830);
	G24739<= not (G23941 or G22835);
	G24742<= not (G23971 or G22869);
	G24756<= not (G16089 or G24211);
	G24770<= not (G16119 or G24217);
	G24782<= not (G16160 or G24221);
	G24783<= not (G16161 or G24224);
	G24800<= not (G16211 or G24229);
	G24819<= not (G16262 or G24236);
	G24836<= not (G16309 or G24241);
	G24845<= not (G16350 or G24246);
	G24847<= not (G16356 or G24247);
	G24859<= not (G16390 or G24253);
	G24871<= not (G16422 or G24256);
	G25027<= not (G24227 or G17001);
	G25042<= not (G24234 or G17031);
	G25056<= not (G24242 or G17065);
	G25067<= not (G24249 or G17100);
	G25075<= not (G13880 or G23483);
	G25076<= not (G23409 or G22187);
	G25077<= not (G23414 or G22196);
	G25078<= not (G23419 or G22201);
	G25081<= not (G23423 or G22202);
	G25082<= not (G23428 or G22207);
	G25085<= not (G23432 or G22208);
	G25091<= not (G23434 or G22215);
	G25099<= not (G23440 or G22224);
	G25125<= not (G23510 or G22340);
	G25127<= not (G23525 or G22363);
	G25129<= not (G23536 or G22383);
	G25185<= not (G24492 or G10024);
	G25189<= not (G24502 or G10133);
	G25191<= not (G24516 or G22777);
	G25194<= not (G24514 or G10238);
	G25197<= not (G24528 or G10340);
	G25199<= not (G24558 or G20127);
	G25201<= not (G24575 or G18407);
	G25202<= not (G24566 or G22907);
	G25204<= not (G24745 or G23547);
	G25206<= not (G24746 or G23550);
	G25207<= not (G24747 or G23551);
	G25208<= not (G24748 or G23552);
	G25209<= not (G24749 or G23554);
	G25211<= not (G24750 or G23558);
	G25212<= not (G24751 or G23559);
	G25213<= not (G24752 or G23560);
	G25214<= not (G24754 or G23563);
	G25215<= not (G24755 or G23564);
	G25216<= not (G24757 or G23565);
	G25217<= not (G24758 or G23567);
	G25218<= not (G24760 or G23571);
	G25219<= not (G24761 or G23572);
	G25220<= not (G24762 or G23573);
	G25221<= not (G24767 or G23577);
	G25222<= not (G24768 or G23578);
	G25223<= not (G24769 or G23579);
	G25224<= not (G24772 or G23582);
	G25225<= not (G24773 or G23583);
	G25226<= not (G24774 or G23584);
	G25227<= not (G24775 or G23586);
	G25228<= not (G24776 or G23590);
	G25229<= not (G24777 or G23591);
	G25230<= not (G24779 or G23598);
	G25231<= not (G24780 or G23599);
	G25232<= not (G24781 or G23600);
	G25233<= not (G24788 or G23604);
	G25234<= not (G24789 or G23605);
	G25235<= not (G24790 or G23606);
	G25236<= not (G24792 or G23609);
	G25237<= not (G24793 or G23610);
	G25238<= not (G24794 or G23611);
	G25239<= not (G24796 or G23615);
	G25240<= not (G24798 or G23622);
	G25241<= not (G24799 or G23623);
	G25242<= not (G24802 or G23630);
	G25243<= not (G24803 or G23631);
	G25244<= not (G24804 or G23632);
	G25245<= not (G24809 or G23636);
	G25246<= not (G24810 or G23637);
	G25247<= not (G24811 or G23638);
	G25248<= not (G24818 or G23664);
	G25249<= not (G24821 or G23671);
	G25250<= not (G24822 or G23672);
	G25251<= not (G24824 or G23679);
	G25252<= not (G24825 or G23680);
	G25253<= not (G24826 or G23681);
	G25254<= not (G24831 or G23687);
	G25255<= not (G24838 or G23714);
	G25256<= not (G24840 or G23721);
	G25257<= not (G24841 or G23722);
	G25258<= not (G24846 or G23741);
	G25259<= not (G24853 or G23768);
	G25260<= not (G24858 or G17737);
	G25261<= not (G24861 or G23796);
	G25262<= not (G24869 or G17824);
	G25263<= not (G24874 or G17838);
	G25264<= not (G24876 or G23849);
	G25265<= not (G24878 or G23852);
	G25266<= not (G24881 or G17912);
	G25267<= not (G24884 or G17936);
	G25268<= not (G24888 or G17950);
	G25270<= not (G24898 or G18023);
	G25271<= not (G24901 or G18047);
	G25272<= not (G24905 or G18061);
	G25273<= not (G24907 or G23904);
	G25279<= not (G24921 or G18140);
	G25280<= not (G24924 or G18164);
	G25288<= not (G24938 or G18256);
	G25311<= not (G24964 or G24029);
	G25343<= not (G24975 or G5623);
	G25357<= not (G24986 or G5651);
	G25372<= not (G24997 or G5689);
	G25389<= not (G25005 or G5741);
	G25418<= not (G24482 or G22319);
	G25426<= not (G24183 or G24616);
	G25429<= not (G24482 or G22319);
	G25450<= not (G16018 or G25086);
	G25451<= not (G16048 or G25102);
	G25452<= not (G16101 or G25117);
	G25523<= not (G20842 or G24429);
	G25539<= not (G25088 or G6157);
	G25569<= not (G24708 or G24490);
	G25589<= not (G20850 or G24433);
	G25605<= not (G25096 or G6184);
	G25631<= not (G24717 or G24497);
	G25648<= not (G24720 or G24500);
	G25668<= not (G20858 or G24437);
	G25684<= not (G25106 or G6216);
	G25699<= not (G24613 or G24506);
	G25708<= not (G24728 or G24509);
	G25725<= not (G24731 or G24512);
	G25745<= not (G20866 or G24440);
	G25761<= not (G25112 or G6305);
	G25764<= not (G25076 or G21615);
	G25772<= not (G24624 or G24520);
	G25781<= not (G24736 or G24523);
	G25798<= not (G24739 or G24526);
	G25818<= not (G25077 or G21643);
	G25826<= not (G24638 or G24533);
	G25835<= not (G24742 or G24536);
	G25852<= not (G4456 or G14831 or G25078);
	G25853<= not (G25081 or G21674);
	G25861<= not (G24657 or G24546);
	G25870<= not (G4456 or G25078 or G18429 or G16075);
	G25873<= not (G4632 or G14904 or G25082);
	G25874<= not (G25085 or G21703);
	G25882<= not (G4632 or G25082 or G18502 or G16113);
	G25885<= not (G4809 or G14985 or G25091);
	G25887<= not (G4809 or G25091 or G18566 or G16164);
	G25890<= not (G4985 or G15074 or G25099);
	G25892<= not (G4985 or G25099 or G18616 or G16223);
	G25932<= not (G25125 or G17001);
	G25935<= not (G25127 or G17031);
	G25938<= not (G25129 or G17065);
	G25940<= not (G24428 or G17100);
	G25941<= not (G24529 or G24540);
	G25943<= not (G24541 or G24550);
	G25944<= not (G24542 or G24552);
	G25946<= not (G24553 or G24561);
	G25947<= not (G24554 or G24563);
	G25948<= not (G24564 or G24571);
	G25949<= not (G24565 or G24573);
	G25950<= not (G24574 or G24580);
	G25962<= not (G24591 or G23496);
	G25967<= not (G24596 or G23512);
	G25974<= not (G24604 or G23527);
	G25979<= not (G24611 or G23538);
	G26025<= not (G25392 or G17193);
	G26031<= not (G25273 or G22777);
	G26037<= not (G25311 or G18407);
	G26041<= not (G25475 or G24855);
	G26042<= not (G25505 or G24867);
	G26043<= not (G25506 or G24870);
	G26044<= not (G25552 or G24882);
	G26045<= not (G25553 or G24885);
	G26046<= not (G25618 or G24899);
	G26047<= not (G25619 or G24902);
	G26048<= not (G25628 or G24906);
	G26049<= not (G25629 or G24908);
	G26050<= not (G25697 or G24922);
	G26055<= not (G25881 or G24974);
	G26081<= not (G25470 or G25482);
	G26083<= not (G25426 or G22319);
	G26084<= not (G25487 or G25513);
	G26087<= not (G6068 or G24183 or G25319);
	G26090<= not (G25518 or G25560);
	G26096<= not (G6068 or G24183 or G25394);
	G26099<= not (G6068 or G24183 or G25313);
	G26103<= not (G25565 or G25626);
	G26107<= not (G6068 or G24183 or G25383);
	G26110<= not (G6068 or G24183 or G25305);
	G26113<= not (G25426 or G22319);
	G26126<= not (G6068 or G24183 or G25368);
	G26137<= not (G6068 or G24183 or G25355);
	G26140<= not (G24183 or G25430);
	G26145<= not (G6068 or G24183 or G25347);
	G26151<= not (G6068 or G24183 or G25335);
	G26154<= not (G6068 or G24183 or G25329);
	G26160<= not (G25951 or G16162);
	G26168<= not (G25953 or G16212);
	G26183<= not (G25957 or G13270);
	G26199<= not (G25961 or G13291);
	G26217<= not (G25963 or G13320);
	G26240<= not (G25968 or G13340);
	G26265<= not (G25972 or G13360);
	G26272<= not (G25973 or G16423);
	G26283<= not (G25954 or G24486);
	G26295<= not (G25977 or G13385);
	G26304<= not (G25978 or G16451);
	G26327<= not (G25958 or G24493);
	G26336<= not (G25981 or G13481);
	G26374<= not (G25964 or G24503);
	G26417<= not (G25969 or G24515);
	G26529<= not (G25962 or G17001);
	G26530<= not (G25967 or G17031);
	G26531<= not (G25974 or G17065);
	G26532<= not (G25979 or G17100);
	G26534<= not (G25321 or G8869);
	G26541<= not (G13755 or G25269);
	G26545<= not (G13790 or G25277);
	G26547<= not (G13796 or G25278);
	G26553<= not (G13816 or G25282);
	G26557<= not (G13818 or G25286);
	G26559<= not (G13824 or G25287);
	G26560<= not (G25281 or G24559);
	G26569<= not (G13837 or G25290);
	G26573<= not (G13839 or G25294);
	G26575<= not (G13845 or G25295);
	G26583<= not (G25289 or G24569);
	G26592<= not (G13851 or G25300);
	G26596<= not (G13853 or G25304);
	G26607<= not (G25299 or G24578);
	G26616<= not (G13860 or G25310);
	G26630<= not (G25309 or G24585);
	G26655<= not (G25328 or G17084);
	G26659<= not (G25334 or G17116);
	G26660<= not (G25208 or G10024);
	G26661<= not (G25337 or G17122);
	G26664<= not (G25346 or G17138);
	G26665<= not (G25348 or G17143);
	G26666<= not (G25216 or G10133);
	G26667<= not (G25351 or G17149);
	G26669<= not (G25360 or G17161);
	G26670<= not (G25362 or G17166);
	G26671<= not (G25226 or G10238);
	G26672<= not (G25365 or G17172);
	G26675<= not (G25375 or G17176);
	G26676<= not (G25377 or G17181);
	G26677<= not (G25238 or G10340);
	G26776<= not (G26042 or G10024);
	G26781<= not (G26044 or G10133);
	G26786<= not (G26049 or G22777);
	G26789<= not (G26046 or G10238);
	G26795<= not (G26050 or G10340);
	G26798<= not (G26055 or G18407);
	G26799<= not (G26158 or G25453);
	G26800<= not (G26163 or G25457);
	G26801<= not (G26171 or G25461);
	G26802<= not (G26188 or G25466);
	G26803<= not (G15105 or G26213);
	G26804<= not (G15172 or G26235);
	G26805<= not (G15173 or G26236);
	G26806<= not (G15197 or G26244);
	G26807<= not (G15245 or G26261);
	G26808<= not (G15246 or G26262);
	G26809<= not (G15258 or G26270);
	G26810<= not (G15259 or G26271);
	G26811<= not (G15283 or G26279);
	G26812<= not (G15321 or G26291);
	G26813<= not (G15337 or G26302);
	G26814<= not (G15338 or G26303);
	G26815<= not (G15350 or G26311);
	G26816<= not (G15351 or G26312);
	G26817<= not (G15375 or G26317);
	G26818<= not (G15407 or G26335);
	G26820<= not (G15423 or G26346);
	G26821<= not (G15424 or G26347);
	G26822<= not (G15436 or G26352);
	G26823<= not (G15437 or G26353);
	G26824<= not (G15491 or G26382);
	G26825<= not (G15507 or G26390);
	G26826<= not (G15508 or G26391);
	G26827<= not (G15577 or G26425);
	G26869<= not (G26458 or G5642);
	G26873<= not (G25483 or G26260);
	G26877<= not (G26140 or G22319);
	G26878<= not (G26482 or G5680);
	G26882<= not (G25514 or G26301);
	G26885<= not (G26140 or G22319);
	G26887<= not (G26498 or G5732);
	G26891<= not (G25561 or G26345);
	G26897<= not (G26513 or G5790);
	G26901<= not (G25627 or G26389);
	G26905<= not (G26096 or G22319);
	G26914<= not (G26107 or G22319);
	G26988<= not (G24893 or G26023);
	G26989<= not (G26663 or G21913);
	G27011<= not (G24916 or G26026);
	G27012<= not (G26668 or G21931);
	G27037<= not (G24933 or G26028);
	G27038<= not (G26674 or G20640);
	G27051<= not (G4456 or G26081);
	G27065<= not (G24945 or G26029);
	G27066<= not (G26024 or G20665);
	G27078<= not (G4632 or G26084);
	G27094<= not (G4809 or G26090);
	G27106<= not (G4985 or G26103);
	G27120<= not (G26560 or G17001);
	G27123<= not (G26583 or G17031);
	G27129<= not (G26607 or G17065);
	G27131<= not (G26630 or G17100);
	G27144<= not (G23451 or G26052);
	G27147<= not (G23458 or G26054);
	G27149<= not (G23462 or G26060);
	G27152<= not (G23467 or G26062);
	G27157<= not (G23471 or G26067);
	G27160<= not (G23476 or G26069);
	G27165<= not (G23484 or G26074);
	G27174<= not (G23494 or G26080);
	G27175<= not (G26075 or G25342);
	G27179<= not (G26082 or G25356);
	G27184<= not (G26085 or G25371);
	G27188<= not (G26091 or G25388);
	G27243<= not (G26802 or G10340);
	G27250<= not (G26955 or G26166);
	G27251<= not (G26958 or G26186);
	G27252<= not (G26963 or G26207);
	G27253<= not (G26965 or G26212);
	G27254<= not (G26968 or G26231);
	G27255<= not (G26969 or G26233);
	G27256<= not (G26970 or G26234);
	G27257<= not (G26971 or G26243);
	G27258<= not (G26977 or G26257);
	G27259<= not (G26978 or G26258);
	G27260<= not (G26979 or G26259);
	G27261<= not (G26980 or G26263);
	G27262<= not (G26981 or G26268);
	G27263<= not (G26982 or G26269);
	G27264<= not (G26984 or G26278);
	G27265<= not (G26993 or G26288);
	G27266<= not (G26994 or G26289);
	G27267<= not (G26995 or G26290);
	G27268<= not (G26996 or G26292);
	G27269<= not (G26997 or G26293);
	G27270<= not (G26998 or G26298);
	G27271<= not (G26999 or G26299);
	G27272<= not (G27000 or G26300);
	G27273<= not (G27001 or G26307);
	G27274<= not (G27002 or G26309);
	G27275<= not (G27003 or G26310);
	G27276<= not (G27004 or G26316);
	G27277<= not (G27005 or G26318);
	G27278<= not (G27006 or G26319);
	G27279<= not (G27007 or G26324);
	G27280<= not (G27008 or G26325);
	G27281<= not (G27009 or G26326);
	G27282<= not (G27016 or G26332);
	G27283<= not (G27017 or G26333);
	G27284<= not (G27018 or G26334);
	G27285<= not (G27019 or G26339);
	G27286<= not (G27020 or G26340);
	G27287<= not (G27021 or G26342);
	G27288<= not (G27022 or G26343);
	G27289<= not (G27023 or G26344);
	G27290<= not (G27024 or G26348);
	G27291<= not (G27025 or G26350);
	G27292<= not (G27026 or G26351);
	G27293<= not (G27027 or G26357);
	G27294<= not (G27028 or G26361);
	G27295<= not (G27029 or G26362);
	G27296<= not (G27030 or G26363);
	G27297<= not (G27031 or G26365);
	G27298<= not (G27032 or G26366);
	G27299<= not (G27033 or G26371);
	G27300<= not (G27034 or G26372);
	G27301<= not (G27035 or G26373);
	G27302<= not (G27042 or G26379);
	G27303<= not (G27043 or G26380);
	G27304<= not (G27044 or G26381);
	G27305<= not (G27045 or G26383);
	G27306<= not (G27046 or G26384);
	G27307<= not (G27047 or G26386);
	G27308<= not (G27048 or G26387);
	G27309<= not (G27049 or G26388);
	G27310<= not (G27050 or G26392);
	G27311<= not (G27053 or G26396);
	G27312<= not (G27054 or G26397);
	G27313<= not (G27055 or G26400);
	G27314<= not (G27056 or G26404);
	G27315<= not (G27057 or G26405);
	G27316<= not (G27058 or G26406);
	G27317<= not (G27059 or G26408);
	G27318<= not (G27060 or G26409);
	G27319<= not (G27061 or G26414);
	G27320<= not (G27062 or G26415);
	G27321<= not (G27063 or G26416);
	G27322<= not (G27070 or G26422);
	G27323<= not (G27071 or G26423);
	G27324<= not (G27072 or G26424);
	G27325<= not (G27073 or G26426);
	G27326<= not (G27074 or G26427);
	G27327<= not (G27077 or G26432);
	G27328<= not (G27080 or G26437);
	G27329<= not (G27081 or G26438);
	G27330<= not (G27082 or G26441);
	G27331<= not (G27083 or G26445);
	G27332<= not (G27084 or G26446);
	G27333<= not (G27085 or G26447);
	G27334<= not (G27086 or G26449);
	G27335<= not (G27087 or G26450);
	G27336<= not (G27088 or G26455);
	G27337<= not (G27089 or G26456);
	G27338<= not (G27090 or G26457);
	G27339<= not (G27093 or G26464);
	G27340<= not (G27096 or G26469);
	G27341<= not (G27097 or G26470);
	G27342<= not (G27098 or G26473);
	G27343<= not (G27099 or G26477);
	G27344<= not (G27100 or G26478);
	G27345<= not (G27101 or G26479);
	G27346<= not (G27105 or G26488);
	G27347<= not (G27108 or G26493);
	G27348<= not (G27109 or G26494);
	G27354<= not (G27112 or G26504);
	G27414<= not (G26770 or G25187);
	G27415<= not (G23104 or G27181 or G25128);
	G27435<= not (G26777 or G25193);
	G27436<= not (G23118 or G27187 or G24427);
	G27450<= not (G26902 or G24613);
	G27454<= not (G26783 or G25196);
	G27455<= not (G23127 or G26758 or G24431);
	G27462<= not (G26892 or G24622);
	G27464<= not (G27178 or G25975);
	G27466<= not (G26915 or G24624);
	G27470<= not (G26790 or G25198);
	G27471<= not (G23138 or G26764 or G24435);
	G27478<= not (G26754 or G24432);
	G27481<= not (G27182 or G25980);
	G27482<= not (G26906 or G24637);
	G27485<= not (G26928 or G24638);
	G27492<= not (G24958 or G24633 or G26771);
	G27496<= not (G27185 or G25178);
	G27501<= not (G26763 or G24436);
	G27504<= not (G26918 or G24656);
	G27507<= not (G26941 or G24657);
	G27513<= not (G24969 or G24653 or G26778);
	G27521<= not (G26766 or G24439);
	G27524<= not (G26931 or G24675);
	G27527<= not (G26759 or G19087);
	G27529<= not (G4456 or G26873);
	G27531<= not (G26760 or G25181);
	G27532<= not (G26761 or G25182);
	G27538<= not (G24982 or G24672 or G26784);
	G27546<= not (G26769 or G24441);
	G27549<= not (G26765 or G19093);
	G27551<= not (G4632 or G26882);
	G27558<= not (G24993 or G24691 or G26791);
	G27563<= not (G26922 or G24708);
	G27564<= not (G26767 or G25184);
	G27565<= not (G26768 or G19100);
	G27567<= not (G4809 or G26891);
	G27572<= not (G26911 or G24717);
	G27573<= not (G26773 or G25188);
	G27574<= not (G26935 or G24720);
	G27575<= not (G26774 or G19107);
	G27577<= not (G4985 or G26901);
	G27579<= not (G26775 or G25192);
	G27581<= not (G26925 or G24728);
	G27582<= not (G26944 or G24731);
	G27584<= not (G26938 or G24736);
	G27585<= not (G26950 or G24739);
	G27588<= not (G26947 or G24742);
	G27594<= not (G27175 or G17001);
	G27603<= not (G27179 or G17031);
	G27612<= not (G27184 or G17065);
	G27621<= not (G27188 or G17100);
	G27629<= not (G26829 or G26051);
	G27631<= not (G26833 or G26053);
	G27655<= not (G26842 or G26061);
	G27658<= not (G26851 or G26068);
	G27672<= not (G26799 or G10024);
	G27678<= not (G26800 or G10133);
	G27682<= not (G26801 or G10238);
	G27718<= not (G27251 or G10133);
	G27722<= not (G27252 or G10238);
	G27724<= not (G27254 or G10340);
	G27735<= not (G27394 or G26961);
	G27736<= not (G27396 or G26962);
	G27741<= not (G27407 or G26966);
	G27742<= not (G27409 or G26967);
	G27746<= not (G27425 or G26972);
	G27747<= not (G27427 or G26973);
	G27754<= not (G27446 or G26985);
	G27755<= not (G27448 or G26986);
	G27759<= not (G27495 or G27052);
	G27760<= not (G27509 or G27076);
	G27761<= not (G27516 or G27079);
	G27762<= not (G27530 or G27091);
	G27763<= not (G27534 or G27092);
	G27764<= not (G27541 or G27095);
	G27765<= not (G27552 or G27103);
	G27766<= not (G27554 or G27104);
	G27767<= not (G27561 or G27107);
	G27768<= not (G27568 or G27110);
	G27769<= not (G27570 or G27111);
	G27771<= not (G27578 or G27115);
	G27798<= not (G27632 or G1223);
	G27802<= not (G6087 or G27632 or G25330);
	G27810<= not (G27632 or G1215);
	G27811<= not (G6087 or G27632 or G25404);
	G27814<= not (G6087 or G27632 or G25322);
	G27823<= not (G27632 or G1216);
	G27824<= not (G6087 or G27632 or G25399);
	G27827<= not (G6087 or G27632 or G25314);
	G27834<= not (G27478 or G14630);
	G27842<= not (G27632 or G1217);
	G27850<= not (G27501 or G14650);
	G27854<= not (G27632 or G1218);
	G27855<= not (G6087 or G27632 or G25385);
	G27864<= not (G27632 or G1219);
	G27865<= not (G6087 or G27632 or G25370);
	G27868<= not (G23742 or G27632);
	G27869<= not (G27632 or G25437);
	G27875<= not (G27521 or G14677);
	G27882<= not (G27632 or G1220);
	G27883<= not (G6087 or G27632 or G25361);
	G27886<= not (G27632 or G24627);
	G27892<= not (G27546 or G14711);
	G27896<= not (G27632 or G1222);
	G27897<= not (G6087 or G27632 or G25349);
	G27900<= not (G6087 or G27632 or G25338);
	G27906<= not (G16127 or G27656);
	G27911<= not (G16170 or G27657);
	G27916<= not (G16219 or G27659);
	G27917<= not (G16220 or G27660);
	G27925<= not (G16276 or G27661);
	G27937<= not (G16321 or G27666);
	G27950<= not (G16367 or G27673);
	G27962<= not (G16394 or G27679);
	G27964<= not (G16400 or G27680);
	G27980<= not (G16428 or G27681);
	G27997<= not (G16456 or G27242);
	G28002<= not (G26032 or G27246);
	G28029<= not (G26033 or G27247);
	G28059<= not (G26034 or G27248);
	G28088<= not (G26036 or G27249);
	G28145<= not (G27629 or G17001);
	G28146<= not (G27631 or G17031);
	G28147<= not (G27655 or G17065);
	G28148<= not (G27658 or G17100);
	G28157<= not (G13902 or G27370);
	G28185<= not (G27356 or G26845);
	G28189<= not (G27359 or G26853);
	G28191<= not (G27365 or G26860);
	G28192<= not (G27372 or G26866);
	G28199<= not (G27250 or G10024);
	G28321<= not (G27742 or G10133);
	G28325<= not (G27747 or G10238);
	G28328<= not (G27755 or G10340);
	G28342<= not (G15460 or G28008);
	G28344<= not (G15526 or G28027);
	G28345<= not (G15527 or G28028);
	G28346<= not (G15546 or G28035);
	G28348<= not (G15594 or G28050);
	G28349<= not (G15595 or G28051);
	G28350<= not (G15604 or G28057);
	G28351<= not (G15605 or G28058);
	G28352<= not (G15624 or G28065);
	G28353<= not (G15666 or G28073);
	G28354<= not (G15670 or G28079);
	G28355<= not (G15671 or G28080);
	G28356<= not (G15680 or G28086);
	G28357<= not (G15681 or G28087);
	G28358<= not (G15700 or G28094);
	G28360<= not (G15725 or G28098);
	G28361<= not (G15729 or G28104);
	G28362<= not (G15730 or G28105);
	G28363<= not (G15739 or G28111);
	G28364<= not (G15740 or G28112);
	G28366<= not (G15765 or G28116);
	G28367<= not (G15769 or G28122);
	G28368<= not (G15770 or G28123);
	G28371<= not (G15793 or G28127);
	G28392<= not (G27886 or G22344);
	G28394<= not (G27869 or G22344);
	G28397<= not (G27869 or G22344);
	G28400<= not (G27886 or G22344);
	G28403<= not (G27811 or G22344);
	G28406<= not (G27824 or G22344);
	G28409<= not (G24676 or G27801);
	G28410<= not (G27748 or G22344);
	G28413<= not (G24695 or G27809);
	G28414<= not (G27748 or G22344);
	G28417<= not (G24712 or G27830);
	G28418<= not (G24723 or G27846);
	G28420<= not (G16031 or G28171);
	G28421<= not (G16068 or G28176);
	G28425<= not (G16133 or G28188);
	G28449<= not (G27727 or G26780);
	G28461<= not (G27729 or G26787);
	G28470<= not (G27671 or G28193);
	G28473<= not (G27730 or G26794);
	G28482<= not (G27731 or G26797);
	G28488<= not (G26755 or G27719);
	G28489<= not (G26756 or G27720);
	G28490<= not (G27240 or G27721);
	G28495<= not (G27244 or G27723);
	G28499<= not (G26027 or G27725);
	G28523<= not (G26035 or G27732);
	G28525<= not (G27245 or G27726);
	G28528<= not (G26030 or G27728);
	G28551<= not (G26038 or G27733);
	G28578<= not (G26039 or G27734);
	G28606<= not (G26040 or G27737);
	G28634<= not (G28185 or G17001);
	G28635<= not (G28189 or G17031);
	G28636<= not (G28191 or G17065);
	G28637<= not (G28192 or G17100);
	G28654<= not (G27770 or G27355);
	G28656<= not (G27772 or G27358);
	G28658<= not (G27773 or G27364);
	G28661<= not (G27775 or G27371);
	G28668<= not (G27736 or G10024);
	G28728<= not (G28422 or G27904);
	G28731<= not (G28423 or G27908);
	G28732<= not (G14894 or G28426);
	G28733<= not (G28424 or G27909);
	G28735<= not (G14957 or G28430);
	G28736<= not (G28427 or G27913);
	G28737<= not (G28428 or G27914);
	G28738<= not (G14975 or G28433);
	G28739<= not (G28429 or G27915);
	G28744<= not (G15030 or G28439);
	G28745<= not (G28431 or G27922);
	G28746<= not (G15046 or G28441);
	G28747<= not (G28434 or G27923);
	G28748<= not (G28435 or G27924);
	G28749<= not (G15064 or G28444);
	G28750<= not (G28436 or G27926);
	G28754<= not (G28440 or G27931);
	G28758<= not (G15126 or G28451);
	G28759<= not (G28442 or G27935);
	G28760<= not (G15142 or G28453);
	G28761<= not (G28445 or G27936);
	G28762<= not (G28446 or G27938);
	G28763<= not (G15160 or G28456);
	G28767<= not (G28452 or G27945);
	G28771<= not (G15218 or G28463);
	G28772<= not (G28454 or G27949);
	G28773<= not (G15234 or G28465);
	G28774<= not (G28457 or G27951);
	G28778<= not (G28464 or G27963);
	G28782<= not (G15304 or G28475);
	G28783<= not (G28466 or G27968);
	G28784<= not (G28468 or G27970);
	G28788<= not (G28476 or G27984);
	G28789<= not (G28477 or G27985);
	G28790<= not (G28478 or G27991);
	G28794<= not (G28484 or G28009);
	G28795<= not (G28485 or G28015);
	G28802<= not (G28492 or G28036);
	G28803<= not (G28493 or G28042);
	G28813<= not (G28497 or G28066);
	G28874<= not (G28657 or G16221);
	G28886<= not (G28659 or G16277);
	G28903<= not (G28660 or G13295);
	G28920<= not (G28662 or G13322);
	G28941<= not (G28663 or G13343);
	G28954<= not (G26673 or G27241 or G28323);
	G28963<= not (G28664 or G13365);
	G28982<= not (G28665 or G28670);
	G28987<= not (G28666 or G13390);
	G28990<= not (G28667 or G16457);
	G29009<= not (G28669 or G28320);
	G29013<= not (G28671 or G11607);
	G29016<= not (G28672 or G13487);
	G29031<= not (G28319 or G28324);
	G29039<= not (G28322 or G13500);
	G29063<= not (G28326 or G28329);
	G29064<= not (G28327 or G28330);
	G29083<= not (G28331 or G28333);
	G29090<= not (G28332 or G28334);
	G29097<= not (G28335 or G28336);
	G29109<= not (G28654 or G17001);
	G29110<= not (G28656 or G17031);
	G29111<= not (G28658 or G17065);
	G29112<= not (G28661 or G17100);
	G29113<= not (G28381 or G8907);
	G29126<= not (G28373 or G27774);
	G29127<= not (G28376 or G27779);
	G29128<= not (G28380 or G27783);
	G29129<= not (G28385 or G27790);
	G29167<= not (G28841 or G28396);
	G29169<= not (G28843 or G28398);
	G29170<= not (G28844 or G28399);
	G29172<= not (G28846 or G28401);
	G29173<= not (G28847 or G28402);
	G29178<= not (G28848 or G28404);
	G29179<= not (G28849 or G28405);
	G29181<= not (G28850 or G28407);
	G29182<= not (G28851 or G28408);
	G29184<= not (G28852 or G28411);
	G29185<= not (G28853 or G28412);
	G29187<= not (G28854 or G28416);
	G29194<= not (G14958 or G28881);
	G29195<= not (G28880 or G28438);
	G29197<= not (G15031 or G28893);
	G29198<= not (G15047 or G28898);
	G29199<= not (G28892 or G28448);
	G29201<= not (G15104 or G28910);
	G29202<= not (G28897 or G28450);
	G29204<= not (G15127 or G28915);
	G29205<= not (G15143 or G28923);
	G29206<= not (G28909 or G28459);
	G29207<= not (G28914 or G28460);
	G29209<= not (G15196 or G28936);
	G29210<= not (G28919 or G28462);
	G29212<= not (G15219 or G28944);
	G29213<= not (G15235 or G28949);
	G29214<= not (G28931 or G28469);
	G29215<= not (G28935 or G28471);
	G29216<= not (G28940 or G28472);
	G29218<= not (G15282 or G28966);
	G29219<= not (G28948 or G28474);
	G29221<= not (G15305 or G28971);
	G29222<= not (G28958 or G28479);
	G29223<= not (G28962 or G28480);
	G29224<= not (G28970 or G28481);
	G29226<= not (G15374 or G28997);
	G29227<= not (G28986 or G28486);
	G29228<= not (G28996 or G28487);
	G29231<= not (G29022 or G28494);
	G29303<= not (G28716 or G19112);
	G29313<= not (G28717 or G19117);
	G29324<= not (G28718 or G19124);
	G29333<= not (G28719 or G19131);
	G29340<= not (G28337 or G28722);
	G29343<= not (G28338 or G28724);
	G29345<= not (G28339 or G28726);
	G29347<= not (G28340 or G28729);
	G29353<= not (G29126 or G17001);
	G29354<= not (G29127 or G17031);
	G29355<= not (G29128 or G17065);
	G29357<= not (G29129 or G17100);
	G29399<= not (G28834 or G28378);
	G29403<= not (G28836 or G28383);
	G29406<= not (G28838 or G28387);
	G29409<= not (G28840 or G28389);
	G29552<= not (G29130 or G29411);
	G29569<= not (G28708 or G29174);
	G29570<= not (G28709 or G29175);
	G29571<= not (G28710 or G29176);
	G29574<= not (G28712 or G29180);
	G29576<= not (G28713 or G29183);
	G29577<= not (G28714 or G29186);
	G29578<= not (G28715 or G29188);
	G29579<= not (G29399 or G17001);
	G29580<= not (G29403 or G17031);
	G29581<= not (G29406 or G17065);
	G29582<= not (G29409 or G17100);
	G29606<= not (G13878 or G29248);
	G29608<= not (G13892 or G29251);
	G29609<= not (G13900 or G29252);
	G29611<= not (G13913 or G29255);
	G29612<= not (G13933 or G29256);
	G29613<= not (G13941 or G29257);
	G29616<= not (G13969 or G29259);
	G29617<= not (G13989 or G29260);
	G29618<= not (G13997 or G29261);
	G29620<= not (G14039 or G29262);
	G29621<= not (G14059 or G29263);
	G29623<= not (G14130 or G29264);
	G29663<= not (G29518 or G29284);
	G29665<= not (G29521 or G29289);
	G29667<= not (G29524 or G29294);
	G29669<= not (G29528 or G29300);
	G29670<= not (G29529 or G29302);
	G29671<= not (G29534 or G29310);
	G29672<= not (G29536 or G29312);
	G29676<= not (G29540 or G29320);
	G29677<= not (G29543 or G29321);
	G29678<= not (G29545 or G29323);
	G29679<= not (G29549 or G29329);
	G29680<= not (G29553 or G29330);
	G29681<= not (G29555 or G29332);
	G29682<= not (G29557 or G29336);
	G29683<= not (G29559 or G29337);
	G29684<= not (G29562 or G29338);
	G29685<= not (G29564 or G29341);
	G29686<= not (G29566 or G29342);
	G29687<= not (G29572 or G29344);
	G29688<= not (G29575 or G29346);
	G29703<= not (G29583 or G1917);
	G29705<= not (G6104 or G29583 or G25339);
	G29709<= not (G29583 or G1909);
	G29710<= not (G6104 or G29583 or G25412);
	G29713<= not (G6104 or G29583 or G25332);
	G29717<= not (G29583 or G1910);
	G29718<= not (G6104 or G29583 or G25409);
	G29721<= not (G6104 or G29583 or G25323);
	G29725<= not (G29583 or G1911);
	G29727<= not (G29583 or G1912);
	G29728<= not (G6104 or G29583 or G25401);
	G29731<= not (G29583 or G1913);
	G29732<= not (G6104 or G29583 or G25387);
	G29735<= not (G23797 or G29583);
	G29736<= not (G29583 or G25444);
	G29740<= not (G29583 or G1914);
	G29741<= not (G6104 or G29583 or G25376);
	G29744<= not (G29583 or G24641);
	G29747<= not (G29583 or G1916);
	G29748<= not (G6104 or G29583 or G25363);
	G29751<= not (G6104 or G29583 or G25352);
	G29754<= not (G16178 or G29607);
	G29755<= not (G16229 or G29610);
	G29756<= not (G16284 or G29614);
	G29757<= not (G16285 or G29615);
	G29758<= not (G16335 or G29619);
	G29759<= not (G16379 or G29622);
	G29760<= not (G16411 or G29624);
	G29761<= not (G28707 or G28711 or G29466);
	G29762<= not (G16432 or G29625);
	G29763<= not (G16438 or G29626);
	G29764<= not (G16462 or G29464);
	G29765<= not (G13492 or G29465);
	G29766<= not (G29467 or G19142);
	G29767<= not (G29468 or G19143);
	G29768<= not (G29469 or G19146);
	G29769<= not (G29470 or G19148);
	G29770<= not (G29471 or G29196);
	G29771<= not (G29472 or G29200);
	G29772<= not (G29473 or G29203);
	G29773<= not (G29474 or G29208);
	G29774<= not (G29475 or G29211);
	G29775<= not (G29476 or G29217);
	G29776<= not (G29477 or G29220);
	G29777<= not (G29478 or G29225);
	G29778<= not (G29479 or G29229);
	G29779<= not (G13943 or G29502);
	G29780<= not (G29480 or G29232);
	G29781<= not (G29481 or G29233);
	G29782<= not (G29482 or G29234);
	G29783<= not (G29483 or G29235);
	G29784<= not (G29484 or G29236);
	G29785<= not (G29485 or G29238);
	G29786<= not (G29486 or G29239);
	G29787<= not (G29487 or G29240);
	G29788<= not (G29488 or G29241);
	G29789<= not (G29489 or G29242);
	G29791<= not (G29490 or G29243);
	G29912<= not (G24676 or G29716);
	G29914<= not (G24695 or G29724);
	G29916<= not (G24712 or G29726);
	G29918<= not (G29744 or G22367);
	G29919<= not (G29736 or G22367);
	G29920<= not (G24723 or G29739);
	G29921<= not (G29736 or G22367);
	G29922<= not (G29744 or G22367);
	G29924<= not (G29710 or G22367);
	G29926<= not (G29718 or G22367);
	G29928<= not (G29673 or G22367);
	G29929<= not (G29673 or G22367);
	G29936<= not (G16049 or G29790);
	G29939<= not (G16102 or G29792);
	G29941<= not (G16182 or G29793);
	G30010<= not (G29520 or G29942);
	G30011<= not (G29522 or G29944);
	G30012<= not (G29523 or G29945);
	G30013<= not (G29525 or G29946);
	G30014<= not (G29526 or G29947);
	G30015<= not (G29527 or G29948);
	G30016<= not (G29531 or G29949);
	G30017<= not (G29532 or G29950);
	G30018<= not (G29533 or G29951);
	G30019<= not (G29538 or G29952);
	G30020<= not (G29539 or G29953);
	G30021<= not (G29541 or G29954);
	G30022<= not (G29547 or G29955);
	G30023<= not (G29548 or G29956);
	G30024<= not (G29550 or G29957);
	G30025<= not (G29558 or G29958);
	G30026<= not (G29560 or G29959);
	G30027<= not (G29565 or G29960);
	G30028<= not (G29567 or G29961);
	G30029<= not (G29573 or G29962);
	G30030<= not (G24676 or G29923);
	G30031<= not (G24695 or G29925);
	G30032<= not (G24712 or G29927);
	G30033<= not (G24723 or G29931);
	G30053<= not (G29963 or G16286);
	G30054<= not (G29964 or G16336);
	G30055<= not (G29965 or G13326);
	G30056<= not (G29966 or G13345);
	G30057<= not (G29967 or G13368);
	G30058<= not (G29968 or G13395);
	G30059<= not (G29969 or G29811);
	G30060<= not (G29970 or G11612);
	G30061<= not (G29971 or G13493);
	G30062<= not (G29810 or G29815);
	G30063<= not (G29812 or G11637);
	G30064<= not (G29813 or G13506);
	G30065<= not (G29814 or G29817);
	G30066<= not (G29816 or G13517);
	G30067<= not (G29818 or G29820);
	G30068<= not (G29819 or G29821);
	G30069<= not (G29822 or G29828);
	G30070<= not (G29827 or G29833);
	G30071<= not (G29834 or G29839);
	G30072<= not (G29910 or G8947);
	G30245<= not (G16074 or G30077);
	G30246<= not (G16107 or G30079);
	G30247<= not (G16112 or G30080);
	G30248<= not (G16139 or G30081);
	G30249<= not (G16158 or G30082);
	G30250<= not (G16163 or G30083);
	G30251<= not (G16198 or G30085);
	G30252<= not (G16217 or G30086);
	G30253<= not (G16222 or G30087);
	G30254<= not (G16242 or G30088);
	G30255<= not (G16263 or G30089);
	G30256<= not (G16282 or G30090);
	G30257<= not (G16290 or G30091);
	G30258<= not (G16291 or G30092);
	G30259<= not (G16301 or G30093);
	G30260<= not (G16322 or G30094);
	G30261<= not (G16342 or G30095);
	G30262<= not (G16343 or G30096);
	G30263<= not (G16344 or G30097);
	G30264<= not (G16348 or G30098);
	G30265<= not (G16349 or G30099);
	G30266<= not (G16359 or G30100);
	G30267<= not (G16380 or G30101);
	G30268<= not (G16382 or G30102);
	G30269<= not (G16386 or G30103);
	G30270<= not (G16387 or G30104);
	G30271<= not (G16388 or G30105);
	G30272<= not (G16392 or G30106);
	G30273<= not (G16393 or G30107);
	G30274<= not (G16403 or G30108);
	G30275<= not (G16413 or G30109);
	G30276<= not (G16415 or G30110);
	G30277<= not (G16418 or G30111);
	G30278<= not (G16420 or G30112);
	G30279<= not (G16424 or G30113);
	G30280<= not (G16425 or G30114);
	G30281<= not (G16426 or G30115);
	G30282<= not (G16430 or G30117);
	G30283<= not (G16431 or G30118);
	G30284<= not (G16444 or G29980);
	G30285<= not (G16447 or G29981);
	G30286<= not (G16449 or G29982);
	G30287<= not (G16452 or G29983);
	G30288<= not (G16454 or G29984);
	G30289<= not (G16458 or G29985);
	G30290<= not (G16459 or G29986);
	G30291<= not (G16460 or G29987);
	G30292<= not (G13477 or G29988);
	G30293<= not (G13480 or G29989);
	G30294<= not (G13483 or G29990);
	G30295<= not (G13485 or G29991);
	G30296<= not (G13488 or G29993);
	G30297<= not (G13490 or G29994);
	G30298<= not (G13496 or G29995);
	G30299<= not (G13499 or G29996);
	G30300<= not (G13502 or G30001);
	G30301<= not (G13504 or G30002);
	G30302<= not (G13513 or G30003);
	G30303<= not (G13516 or G30005);
	G30304<= not (G13527 or G30007);
	G30338<= not (G14297 or G30225);
	G30341<= not (G14328 or G30226);
	G30356<= not (G14419 or G30227);
	G30399<= not (G30116 or G30123);
	G30400<= not (G29997 or G30127);
	G30401<= not (G29998 or G30128);
	G30402<= not (G29999 or G30129);
	G30403<= not (G30004 or G30131);
	G30404<= not (G30006 or G30132);
	G30405<= not (G30008 or G30133);
	G30406<= not (G30009 or G30138);
	G30455<= not (G13953 or G30216);
	G30468<= not (G14007 or G30217);
	G30470<= not (G14023 or G30218);
	G30482<= not (G14067 or G30219);
	G30485<= not (G14098 or G30220);
	G30487<= not (G14114 or G30221);
	G30500<= not (G14182 or G30222);
	G30503<= not (G14213 or G30223);
	G30505<= not (G14229 or G30224);
	G30566<= not (G14327 or G30398);
	G30584<= not (G30412 or G2611);
	G30588<= not (G6119 or G30412 or G25353);
	G30593<= not (G30412 or G2603);
	G30594<= not (G6119 or G30412 or G25419);
	G30597<= not (G6119 or G30412 or G25341);
	G30601<= not (G30412 or G2604);
	G30602<= not (G6119 or G30412 or G25417);
	G30605<= not (G6119 or G30412 or G25333);
	G30608<= not (G30412 or G2605);
	G30609<= not (G30412 or G2606);
	G30610<= not (G6119 or G30412 or G25411);
	G30613<= not (G30412 or G2607);
	G30614<= not (G6119 or G30412 or G25403);
	G30617<= not (G23850 or G30412);
	G30618<= not (G30412 or G25449);
	G30621<= not (G30412 or G2608);
	G30622<= not (G6119 or G30412 or G25393);
	G30625<= not (G30412 or G24660);
	G30628<= not (G30412 or G2610);
	G30629<= not (G6119 or G30412 or G25378);
	G30632<= not (G6119 or G30412 or G25366);
	G30635<= not (G16108 or G30407);
	G30636<= not (G16140 or G30409);
	G30637<= not (G16141 or G30410);
	G30638<= not (G16159 or G30411);
	G30639<= not (G16186 or G30436);
	G30640<= not (G16187 or G30437);
	G30641<= not (G16188 or G30438);
	G30642<= not (G16199 or G30440);
	G30643<= not (G16200 or G30441);
	G30644<= not (G16218 or G30442);
	G30645<= not (G16240 or G30444);
	G30646<= not (G16241 or G30445);
	G30647<= not (G16251 or G30447);
	G30648<= not (G16252 or G30448);
	G30649<= not (G16253 or G30449);
	G30650<= not (G16264 or G30451);
	G30651<= not (G16265 or G30452);
	G30652<= not (G16283 or G30453);
	G30653<= not (G16289 or G30454);
	G30654<= not (G16299 or G30457);
	G30655<= not (G16300 or G30458);
	G30656<= not (G16310 or G30460);
	G30657<= not (G16311 or G30461);
	G30658<= not (G16312 or G30462);
	G30659<= not (G16323 or G30464);
	G30660<= not (G16324 or G30465);
	G30661<= not (G16345 or G30467);
	G30662<= not (G16347 or G30469);
	G30663<= not (G16357 or G30472);
	G30664<= not (G16358 or G30473);
	G30665<= not (G16368 or G30475);
	G30666<= not (G16369 or G30476);
	G30667<= not (G16370 or G30477);
	G30668<= not (G16381 or G30478);
	G30669<= not (G16383 or G30481);
	G30670<= not (G16389 or G30484);
	G30671<= not (G16391 or G30486);
	G30672<= not (G16401 or G30489);
	G30673<= not (G16402 or G30490);
	G30674<= not (G16414 or G30492);
	G30675<= not (G16416 or G30495);
	G30676<= not (G16419 or G30496);
	G30677<= not (G16421 or G30499);
	G30678<= not (G16427 or G30502);
	G30679<= not (G16429 or G30504);
	G30680<= not (G16443 or G30327);
	G30681<= not (G16448 or G30330);
	G30682<= not (G16450 or G30333);
	G30683<= not (G16453 or G30334);
	G30684<= not (G16455 or G30337);
	G30685<= not (G29992 or G30000 or G30372);
	G30686<= not (G16461 or G30340);
	G30687<= not (G13479 or G30345);
	G30688<= not (G13484 or G30348);
	G30689<= not (G13486 or G30351);
	G30690<= not (G13489 or G30352);
	G30691<= not (G13491 or G30355);
	G30692<= not (G13498 or G30361);
	G30693<= not (G13503 or G30364);
	G30694<= not (G13505 or G30367);
	G30695<= not (G13515 or G30374);
	G30699<= not (G13914 or G30387);
	G30700<= not (G13952 or G30388);
	G30701<= not (G13970 or G30389);
	G30702<= not (G14006 or G30390);
	G30703<= not (G14022 or G30391);
	G30704<= not (G14040 or G30392);
	G30705<= not (G14097 or G30393);
	G30706<= not (G14113 or G30394);
	G30707<= not (G14131 or G30395);
	G30708<= not (G14212 or G30396);
	G30709<= not (G14228 or G30397);
	G30780<= not (G30625 or G22387);
	G30783<= not (G30618 or G22387);
	G30785<= not (G30618 or G22387);
	G30786<= not (G30625 or G22387);
	G30787<= not (G30594 or G22387);
	G30788<= not (G30602 or G22387);
	G30789<= not (G30575 or G22387);
	G30790<= not (G30575 or G22387);
	G30796<= not (G16069 or G30696);
	G30798<= not (G16134 or G30697);
	G30801<= not (G16237 or G30698);
	G30929<= not (G30728 or G30736);
	G30930<= not (G30735 or G30744);
	G30931<= not (G30743 or G30750);
	G30932<= not (G30754 or G30757);
	G30933<= not (G30755 or G30758);
	G30934<= not (G30759 or G30761);
	G30935<= not (G30760 or G30762);
	G30936<= not (G30763 or G30764);
	G30954<= not (G30916 or G30944);
	G30955<= not (G30918 or G30945);
	G30956<= not (G30919 or G30946);
	G30957<= not (G30920 or G30947);
	G30958<= not (G30922 or G30948);
	G30959<= not (G30923 or G30949);
	G30960<= not (G30924 or G30950);
	G30961<= not (G30925 or G30951);
	G30970<= not (G30917 or G30921 or G30953);
end RTL;
