-- File created by Bench2VHDL
-- Name: s1494
-- File: bench/s1494.bench
-- Timestamp: 2019-05-21T22:08:28.936857
--
-- Original File
-- =============
--	# s1494
--	# 8 inputs
--	# 19 outputs
--	# 6 D-type flipflops
--	# 89 inverters
--	# 558 gates (354 ANDs + 0 NANDs + 204 ORs + 0 NORs)
--	
--	INPUT(CLR)
--	INPUT(v6)
--	INPUT(v5)
--	INPUT(v4)
--	INPUT(v3)
--	INPUT(v2)
--	INPUT(v1)
--	INPUT(v0)
--	
--	OUTPUT(v13_D_24)
--	OUTPUT(v13_D_23)
--	OUTPUT(v13_D_22)
--	OUTPUT(v13_D_21)
--	OUTPUT(v13_D_20)
--	OUTPUT(v13_D_19)
--	OUTPUT(v13_D_18)
--	OUTPUT(v13_D_17)
--	OUTPUT(v13_D_16)
--	OUTPUT(v13_D_15)
--	OUTPUT(v13_D_14)
--	OUTPUT(v13_D_13)
--	OUTPUT(v13_D_12)
--	OUTPUT(v13_D_11)
--	OUTPUT(v13_D_10)
--	OUTPUT(v13_D_9)
--	OUTPUT(v13_D_8)
--	OUTPUT(v13_D_7)
--	OUTPUT(v13_D_6)
--	
--	v12 = DFF(v13_D_5C)
--	v11 = DFF(v13_D_4C)
--	v10 = DFF(v13_D_3C)
--	v9 = DFF(v13_D_2C)
--	v8 = DFF(v13_D_1C)
--	v7 = DFF(v13_D_0C)
--	
--	v4E = NOT(v4)
--	C70DE = NOT(C70D)
--	C104DE = NOT(C104D)
--	C141DE = NOT(C141D)
--	C191DE = NOT(C191D)
--	C218DE = NOT(C218D)
--	C180DE = NOT(C180D)
--	C90DE = NOT(C90D)
--	v3E = NOT(v3)
--	v1E = NOT(v1)
--	C30DE = NOT(C30D)
--	C194DE = NOT(C194D)
--	C117DE = NOT(C117D)
--	C195DE = NOT(C195D)
--	C208DE = NOT(C208D)
--	C118DE = NOT(C118D)
--	C138DE = NOT(C138D)
--	C220DE = NOT(C220D)
--	C166DE = NOT(C166D)
--	C49DE = NOT(C49D)
--	v5E = NOT(v5)
--	C81DE = NOT(C81D)
--	C131DE = NOT(C131D)
--	v0E = NOT(v0)
--	C144DE = NOT(C144D)
--	C157DE = NOT(C157D)
--	v11E = NOT(v11)
--	v6E = NOT(v6)
--	C129DE = NOT(C129D)
--	v9E = NOT(v9)
--	v2E = NOT(v2)
--	v10E = NOT(v10)
--	v12E = NOT(v12)
--	C165DE = NOT(C165D)
--	C83DE = NOT(C83D)
--	C108DE = NOT(C108D)
--	C124DE = NOT(C124D)
--	v8E = NOT(v8)
--	v7E = NOT(v7)
--	I650 = NOT(Av13_D_24B)
--	v13_D_24 = NOT(I650)
--	I653 = NOT(Av13_D_23B)
--	v13_D_23 = NOT(I653)
--	I656 = NOT(Av13_D_22B)
--	v13_D_22 = NOT(I656)
--	I659 = NOT(Av13_D_21B)
--	v13_D_21 = NOT(I659)
--	I662 = NOT(Av13_D_20B)
--	v13_D_20 = NOT(I662)
--	I665 = NOT(Av13_D_19B)
--	v13_D_19 = NOT(I665)
--	I668 = NOT(Av13_D_18B)
--	v13_D_18 = NOT(I668)
--	I671 = NOT(Av13_D_17B)
--	v13_D_17 = NOT(I671)
--	I674 = NOT(Av13_D_16B)
--	v13_D_16 = NOT(I674)
--	I677 = NOT(Av13_D_15B)
--	v13_D_15 = NOT(I677)
--	I680 = NOT(Av13_D_14B)
--	v13_D_14 = NOT(I680)
--	I683 = NOT(Av13_D_13B)
--	v13_D_13 = NOT(I683)
--	I686 = NOT(Av13_D_12B)
--	v13_D_12 = NOT(I686)
--	I689 = NOT(Av13_D_11B)
--	v13_D_11 = NOT(I689)
--	I692 = NOT(Av13_D_10B)
--	v13_D_10 = NOT(I692)
--	I695 = NOT(Av13_D_9B)
--	v13_D_9 = NOT(I695)
--	I698 = NOT(Av13_D_8B)
--	v13_D_8 = NOT(I698)
--	I701 = NOT(Av13_D_7B)
--	v13_D_7 = NOT(I701)
--	I704 = NOT(Av13_D_6B)
--	v13_D_6 = NOT(I704)
--	I707 = NOT(Av13_D_5B)
--	v13_D_5 = NOT(I707)
--	I710 = NOT(Av13_D_4B)
--	v13_D_4 = NOT(I710)
--	I713 = NOT(Av13_D_3B)
--	v13_D_3 = NOT(I713)
--	I716 = NOT(Av13_D_2B)
--	v13_D_2 = NOT(I716)
--	I719 = NOT(Av13_D_1B)
--	v13_D_1 = NOT(I719)
--	I722 = NOT(Av13_D_0B)
--	v13_D_0 = NOT(I722)
--	
--	v13_D_5C = AND(v13_D_5, CLR)
--	v13_D_4C = AND(v13_D_4, CLR)
--	v13_D_3C = AND(v13_D_3, CLR)
--	v13_D_2C = AND(v13_D_2, CLR)
--	v13_D_1C = AND(v13_D_1, CLR)
--	v13_D_0C = AND(v13_D_0, CLR)
--	I560 = AND(v7E, v12E)
--	I559 = AND(v8, v11)
--	I555 = AND(v0, v8E, v11)
--	I554 = AND(v2E, v8, v9E)
--	I547 = AND(v10, v11E)
--	I546 = AND(v0, v11)
--	I538 = AND(v8, v12E)
--	I537 = AND(v6E, v7E, v8E, v12)
--	I534 = AND(v8E, v10E)
--	I533 = AND(v9, v10)
--	I528 = AND(v9E, v11)
--	I524 = AND(v6, v11E)
--	I520 = AND(v3E, v6E)
--	I518 = AND(v9, v10E)
--	I516 = AND(v1, v12)
--	I514 = AND(v2, v7, v9E, C138DE)
--	I142 = AND(v7E, v9, v11E)
--	I513 = AND(v12E, C166DE, I142)
--	I510 = AND(v9, v10)
--	I508 = AND(v9E, v11E)
--	I506 = AND(v7E, v9, v10E, v12E)
--	I505 = AND(v7, v8, C138DE, C191DE)
--	I503 = AND(v9E, C30DE)
--	I501 = AND(v8E, v11E)
--	I500 = AND(v8, v11, C83DE)
--	I498 = AND(v8, C117DE)
--	II497 = AND(v8E, v9E, C194DE)
--	I495 = AND(v9, v11, C131DE)
--	I494 = AND(v8E, v10, C108DE)
--	I492 = AND(v10, v11E)
--	II491 = AND(v10E, C138DE)
--	I489 = AND(v8E, v11)
--	I486 = AND(v6E, v8E, v12, C129DE)
--	I485 = AND(v6, C141DE, C220DE)
--	I483 = AND(v8E, v9E, v11E, C83DE)
--	I482 = AND(v2, C220DE)
--	I479 = AND(v0, v11)
--	I478 = AND(v10E, C83DE)
--	I476 = AND(v8E, v9, v11E, v12E)
--	I475 = AND(v2E, v8, C138DE)
--	I473 = AND(v0E, C30DE)
--	I471 = AND(v1, v10E, v12)
--	I470 = AND(v8, v12E, C83DE)
--	I468 = AND(v9, C83DE)
--	I466 = AND(v8E, v11E, v12E)
--	I464 = AND(v8E, v10E, v11)
--	I463 = AND(C165DE, C191DE)
--	I461 = AND(v8E, v9, v12)
--	I460 = AND(v2E, v12E, C165DE)
--	I457 = AND(v6, C124DE, C90DE)
--	I456 = AND(v9, C30DE)
--	I453 = AND(v8E, v10E, v12)
--	I452 = AND(v12E, C220DE)
--	I450 = AND(v3, v8, C138DE, C104DE)
--	I449 = AND(C108DE, C83DE)
--	I447 = AND(v8E, v9, v10E, v12E)
--	I446 = AND(v11E, C90DE)
--	I444 = AND(v3E, v9E)
--	I442 = AND(v7E, v8E, v9E)
--	I441 = AND(v11, C220DE)
--	I439 = AND(v6, v12, C124DE)
--	I438 = AND(v0, v10, C144DE)
--	I436 = AND(v8E, v9, C144DE)
--	I435 = AND(v12, C165DE)
--	I433 = AND(v10, C144DE)
--	I432 = AND(v7, C90DE)
--	I430 = AND(v1E, v9, v10E)
--	I429 = AND(v9E, C30DE)
--	I427 = AND(v8E, v9, v10)
--	I425 = AND(v8E, v10E)
--	I423 = AND(v3E, C157DE)
--	I420 = AND(v2E, v7, C131DE)
--	I419 = AND(v5E, v7E, v8E, C30DE)
--	I417 = AND(v5E, v11E, v12E)
--	I415 = AND(v8E, v11E, v12E)
--	I414 = AND(v6, C138DE)
--	I412 = AND(v3, v10E, v12E)
--	I409 = AND(v9, v11E)
--	I406 = AND(v8, v11, C117DE)
--	I405 = AND(v8E, v9E, C194DE)
--	I254 = AND(v1, v6, v7E, v8E)
--	I403 = AND(v9, v12E, C124DE, I254)
--	I402 = AND(v8, v9E, C30DE)
--	I399 = AND(v8, C141D)
--	I398 = AND(v12E, C118DE)
--	I396 = AND(v10E, v12E)
--	I395 = AND(C157D, v9E)
--	I393 = AND(v10E, v12E)
--	I392 = AND(C81D, v11E)
--	I390 = AND(C220D, v10E)
--	I389 = AND(v8, v9, v10)
--	I387 = AND(v8E, v9E, C124DE)
--	I386 = AND(v0, C104D, v8, C30DE)
--	I384 = AND(v10E, C138DE)
--	I383 = AND(C70D, C141DE)
--	I381 = AND(C166D, v11E)
--	I380 = AND(v2, v11)
--	I378 = AND(C218D, v5E, v9, v12E)
--	I377 = AND(v7, v10, C90DE)
--	I375 = AND(C86D, v10E)
--	I374 = AND(v9E, C30DE)
--	I372 = AND(C129D, v12E)
--	I371 = AND(v10E, C90DE)
--	I369 = AND(v9, C124DE)
--	II368 = AND(C30D, C90DE)
--	I366 = AND(v8E, v9, v11E, v12E)
--	I365 = AND(C56D, v8, v11)
--	I363 = AND(v1E, C178D)
--	I362 = AND(v8, C138DE)
--	I360 = AND(v3E, C59D)
--	I359 = AND(v12E, C165DE)
--	I357 = AND(v10, v11E)
--	I356 = AND(C50D, v10E)
--	I354 = AND(C191D, v11)
--	I352 = AND(v8, C124D)
--	I350 = AND(v11, C117D)
--	I349 = AND(C118D, v11E)
--	I347 = AND(C90D, v10E)
--	I346 = AND(v12, C191DE)
--	I344 = AND(C83D, v12E)
--	I342 = AND(C159D, v8E)
--	I341 = AND(v11E, C118DE)
--	I339 = AND(v8E, C144DE)
--	I338 = AND(C108D, C165DE)
--	I336 = AND(C124D, v12)
--	I335 = AND(v12E, C218DE)
--	I333 = AND(v11E, v12E)
--	I332 = AND(C138D, v9E)
--	I329 = AND(v3, v7E, v10)
--	Av13_D_20B = AND(C138DE, C220DE, C104D, I329)
--	II329 = AND(v9, v12, C30D)
--	I328 = AND(v3, v12E, C124DE)
--	I326 = AND(C81DE, C129D)
--	I325 = AND(v10, C90DE)
--	I323 = AND(v10E, C127D)
--	I321 = AND(C33D, v11E, v12E)
--	I320 = AND(v11, C141D)
--	I318 = AND(v11, C118D)
--	I317 = AND(v10, v11E)
--	I315 = AND(C155D, v12E, C129D)
--	I314 = AND(v10, C90DE)
--	I311 = AND(C71D, v9E)
--	I310 = AND(v6E, v9, v12E, C124DE)
--	I308 = AND(C111D, C144DE)
--	I306 = AND(C129DE, C138D)
--	I305 = AND(v9, C49DE)
--	I303 = AND(C172D, v12E)
--	I302 = AND(v11E, C157DE)
--	I300 = AND(v0E, C105D)
--	I299 = AND(v11E, C108DE)
--	I297 = AND(C209D, C208D, v11)
--	I296 = AND(v8E, v9E, C124DE, C83DE)
--	I294 = AND(C211D, v3, v7E, v11E)
--	I368 = AND(v7, v8, v9E)
--	I293 = AND(C138DE, C118DE, I368)
--	I291 = AND(C142D, v11)
--	Av13_D_21B = AND(C213D, v7E, v10E, v12E)
--	I288 = AND(v7E, C203D)
--	I287 = AND(v9, v11)
--	I285 = AND(C222D, v10E)
--	I284 = AND(v11E, C157DE)
--	I282 = AND(C36D, v12)
--	I281 = AND(v3E, C29D)
--	I280 = AND(v1E, C26D)
--	I278 = AND(v10E, C138DE)
--	I276 = AND(C27D, v7E, v9, v12E)
--	I275 = AND(v7, v8, C90DE)
--	I273 = AND(C201D, v8)
--	I272 = AND(v10E, C144DE)
--	I270 = AND(v1E, C55D)
--	I269 = AND(v11E, C108DE, C83DE)
--	I267 = AND(C214D, v7E, v10E)
--	I266 = AND(v7, C49DE, C220DE)
--	Av13_D_16B = AND(C200D, v8, v10)
--	I263 = AND(v7E, v11, C41D)
--	I262 = AND(C42D, v8)
--	I260 = AND(v3E, C78D)
--	I259 = AND(v12E, C129DE, C83DE)
--	I257 = AND(C215D, v9E)
--	I256 = AND(v9, v10, C138DE)
--	II254 = AND(C39D, v8E)
--	I253 = AND(v1E, v10E, C138DE)
--	I251 = AND(v6E, v11E, v12E)
--	I250 = AND(C77D, v3, C138DE)
--	I248 = AND(C45D, v10E)
--	I247 = AND(v10, C144DE)
--	I245 = AND(C185D, v8E)
--	I243 = AND(C131D, v9, C144DE)
--	I242 = AND(C130D, C165DE)
--	I240 = AND(C125D, v9E)
--	I239 = AND(v9, v12, C124DE)
--	I237 = AND(v7, v12E, C221D)
--	I236 = AND(v2E, v8, C219D)
--	I234 = AND(v8, C167D)
--	I233 = AND(C168D, v8E)
--	I232 = AND(C165D, C83DE)
--	I230 = AND(C109D, v10E)
--	I229 = AND(v9, v10, C144DE)
--	I227 = AND(C139D, v8, v10)
--	I226 = AND(v8E, v10E, C144DE)
--	I224 = AND(C163D, v8E, v11)
--	I223 = AND(v7E, C160D, v9E)
--	I222 = AND(C156D, C83DE)
--	I220 = AND(C51D, v12)
--	I219 = AND(C49D, v9)
--	I218 = AND(v12E, C44D, C83DE)
--	I216 = AND(C189D, v9E)
--	I215 = AND(v1, v9, C144DE)
--	I213 = AND(C57D, v10E)
--	I212 = AND(v9E, C49DE)
--	I210 = AND(v9, C120D)
--	I209 = AND(v8, C119D)
--	I208 = AND(C122D, v11E)
--	I206 = AND(v7, C150D)
--	I205 = AND(v8E, C30DE)
--	I203 = AND(C34D, v9)
--	I202 = AND(v9E, C144DE, C83DE, C194DE)
--	I200 = AND(v12E, C124D)
--	I199 = AND(v9E, C63D)
--	I197 = AND(C158D, v7, v11E)
--	I196 = AND(C161D, v11)
--	I194 = AND(v3, v12, C77D)
--	I192 = AND(v8E, v9E, C44D)
--	I191 = AND(v8, v11, C117DE)
--	I189 = AND(v7, v12E)
--	I188 = AND(C175D, v11)
--	I186 = AND(v8, v11, C117DE)
--	I185 = AND(v8E, C195DE)
--	I183 = AND(C183D, v8)
--	I182 = AND(v8E, v10E, C144DE)
--	I180 = AND(C173D, v9E)
--	I179 = AND(v9, v10, C144DE)
--	I177 = AND(C137D, C127D)
--	I176 = AND(v10E, C145D)
--	I175 = AND(v9, C144D)
--	I174 = AND(v8E, C143D)
--	I173 = AND(C146D, v11E)
--	I171 = AND(v8, C193D)
--	I170 = AND(v10, v11E)
--	I169 = AND(C195D, v8E)
--	I167 = AND(v8, v11, C129D)
--	I166 = AND(C205D, v10)
--	I164 = AND(C133D, v8E)
--	I163 = AND(v11E, v12E, C118DE)
--	I161 = AND(C144DE, C191D)
--	I160 = AND(v8, C65D)
--	I158 = AND(C84D, v10E)
--	I157 = AND(C82D, v9E)
--	I156 = AND(C80D, v9)
--	I154 = AND(v2, C40D)
--	I153 = AND(C52D, v8E)
--	I152 = AND(v8, v12E, C129DE)
--	I151 = AND(v9, C138DE)
--	I149 = AND(C112D, v10)
--	I148 = AND(v9, v10E, C144DE)
--	I146 = AND(C223D, v8E, v9E)
--	I145 = AND(C49DE, C166DE, C220DE)
--	Av13_D_23B = AND(C216D, v7E, v8E)
--	II142 = AND(v7E, C169D)
--	I141 = AND(C170D, v8)
--	I140 = AND(v8E, v10E, C144DE)
--	Av13_D_18B = AND(C210D, v7E, v12E)
--	I137 = AND(v8, C46D)
--	I136 = AND(C47D, C144DE)
--	I134 = AND(v7E, v10, C151D)
--	I133 = AND(C152D, v9)
--	I131 = AND(v9, v11E, C157DE)
--	I130 = AND(C60D, C83D)
--	I129 = AND(v8E, C72D)
--	I128 = AND(v8, C69D)
--	I127 = AND(C73D, v10E)
--	I126 = AND(v2, C58D)
--	I124 = AND(C164D, v12E)
--	I123 = AND(v8, C162D)
--	I548 = AND(C199D, v4, v5E)
--	Av13_D_15B = AND(v7E, v12E, I548)
--	I120 = AND(v7E, C123D)
--	I119 = AND(C126D, v8)
--	I117 = AND(v8E, C35D)
--	I116 = AND(C37D, v9)
--	I114 = AND(v9, C97D)
--	I113 = AND(v2E, v12E, C93D)
--	I112 = AND(v11E, v12)
--	I111 = AND(C98D, v10E)
--	I109 = AND(C179D, v2, v8, v11)
--	I108 = AND(C181D, C83DE)
--	I106 = AND(v8E, C114D)
--	I105 = AND(v8, C113D)
--	I104 = AND(v3, C107D, v12)
--	I103 = AND(C115D, v10)
--	I101 = AND(C127D, C128D, v12E)
--	I100 = AND(C134D, v9E)
--	I98 = AND(v8E, v12, C87D)
--	I97 = AND(C88D, v11E)
--	I96 = AND(v8, C85D)
--	I95 = AND(C76D, C81DE)
--	I93 = AND(v7E, C147D)
--	I92 = AND(v7, C140D)
--	I91 = AND(C148D, C131DE)
--	I89 = AND(v7, C48D)
--	I88 = AND(v2E, C43D)
--	I87 = AND(C53D, v7E)
--	I86 = AND(C54D, C165DE)
--	I84 = AND(v7E, C224D)
--	I83 = AND(C225D, v11)
--	I82 = AND(v0E, C217D, C108DE)
--	I80 = AND(v7, v12E, C192D)
--	I79 = AND(v8, C170D)
--	I78 = AND(v7E, C196D)
--	I76 = AND(v7E, C174D)
--	I75 = AND(C129DE, C144DE)
--	I73 = AND(v7, C31D, v8)
--	I72 = AND(C38D, v7E)
--	I71 = AND(v2E, C28D)
--	I69 = AND(v7, C202D)
--	I68 = AND(C206D, v12E)
--	I66 = AND(v8E, v12E, C100D)
--	I65 = AND(v9, C185D)
--	I64 = AND(v11E, C157DE)
--	I63 = AND(v8, C99D)
--	I62 = AND(v6E, C95D)
--	I60 = AND(v7E, C74D)
--	I59 = AND(v7, C67D)
--	I58 = AND(C75D, C129DE)
--	Av13_D_9B = AND(C153D, v12E)
--	I55 = AND(C187D, v12E)
--	I54 = AND(C186D, v9E)
--	I52 = AND(C135D, v7E)
--	I51 = AND(C132D, v7)
--	I49 = AND(v8, C176D)
--	I48 = AND(C177D, v8E)
--	I46 = AND(v7, C110D)
--	I45 = AND(C116D, v7E)
--	I44 = AND(v2E, C106D)
--	I43 = AND(v8, v10, C108DE)
--	I41 = AND(v7, v12E, C96D)
--	I40 = AND(v2, C92D)
--	I39 = AND(C103D, v10E)
--	I38 = AND(C102D, v7E)
--	I36 = AND(v7E, C89D)
--	I35 = AND(C79D, v7, v9, v12E)
--	I34 = AND(C91D, C165DE)
--	I32 = AND(C207D, v2)
--	I642 = AND(v7E, v8E, C124DE)
--	I31 = AND(C108DE, C83DE, I642)
--	I29 = AND(C190D, v10)
--	I28 = AND(v7E, C188D)
--	I27 = AND(C184D, v7)
--	
--	C138D = OR(v11E, v12E)
--	C218D = OR(v7E, v10)
--	C131D = OR(v8E, v10)
--	C220D = OR(v8E, v9E)
--	C155D = OR(v2, v7)
--	C83D = OR(v4E, v5E)
--	C117D = OR(v9E, v2)
--	C178D = OR(I559, I560)
--	C70D = OR(v0, v11E)
--	C157D = OR(v10E, v12E)
--	C151D = OR(I554, I555)
--	C127D = OR(v5E, v4)
--	C142D = OR(v0, v12)
--	C166D = OR(v3E, v6E)
--	C165D = OR(v8E, v11)
--	C30D = OR(v10E, v11E)
--	C159D = OR(I546, I547)
--	C194D = OR(v0, v10E)
--	C193D = OR(v2, v11E)
--	C81D = OR(v2E, v12)
--	C124D = OR(v10, v11)
--	C208D = OR(v5, v4)
--	C191D = OR(v10E, v9)
--	C59D = OR(I537, I538)
--	C108D = OR(v9, v12)
--	C47D = OR(I533, I534)
--	C33D = OR(v6E, v10)
--	C104D = OR(v1, v6E)
--	C144D = OR(v11E, v12)
--	C145D = OR(I528, v12)
--	C90D = OR(v9, v12E)
--	C141D = OR(v10E, v12)
--	C86D = OR(v9, I524)
--	C118D = OR(v2E, v10E)
--	C129D = OR(v9, v10)
--	C50D = OR(I520, v11)
--	C179D = OR(v10, I518)
--	C56D = OR(v9, I516)
--	C200D = OR(I513, I514)
--	C36D = OR(C165DE, v10E)
--	C163D = OR(C129DE, I510)
--	C203D = OR(C70DE, I508)
--	C92D = OR(I505, I506)
--	C201D = OR(I503, v12E)
--	C27D = OR(I500, I501)
--	C209D = OR(II497, I498)
--	C60D = OR(I494, I495)
--	C185D = OR(II491, I492)
--	C137D = OR(C117DE, I489)
--	C45D = OR(C90DE, v11E)
--	C211D = OR(I485, I486)
--	C213D = OR(I482, I483)
--	C79D = OR(C131DE, v11)
--	C172D = OR(I478, I479)
--	C55D = OR(I475, I476)
--	C44D = OR(I473, C124DE)
--	C41D = OR(I470, I471)
--	C93D = OR(C191DE, I468)
--	C29D = OR(C138DE, I466)
--	C96D = OR(I463, I464)
--	C214D = OR(I460, I461)
--	C168D = OR(C159D, v9)
--	C114D = OR(I456, I457)
--	C170D = OR(C124DE, v9E)
--	C78D = OR(I452, I453)
--	C105D = OR(I449, I450)
--	C95D = OR(I446, I447)
--	C98D = OR(C144D, I444)
--	C156D = OR(I441, I442)
--	C215D = OR(I438, I439)
--	C103D = OR(I435, I436)
--	C42D = OR(I432, I433)
--	C100D = OR(I429, I430)
--	C76D = OR(C131DE, I427)
--	C120D = OR(C144D, I425)
--	C39D = OR(I423, v9)
--	C49D = OR(C141D, v11)
--	C217D = OR(I419, I420)
--	C222D = OR(C138DE, I417)
--	C26D = OR(I414, I415)
--	C54D = OR(C90DE, I412)
--	C77D = OR(C104D, v0E)
--	C148D = OR(C90DE, I409)
--	C180D = OR(C194DE, v11E)
--	C128D = OR(I405, I406)
--	C106D = OR(I402, I403)
--	C111D = OR(C83DE, v2)
--	C146D = OR(I398, I399)
--	C158D = OR(I395, I396)
--	C82D = OR(I392, I393)
--	C221D = OR(I389, I390)
--	C107D = OR(I386, I387)
--	C71D = OR(I383, I384)
--	C167D = OR(I380, I381)
--	C219D = OR(I377, I378)
--	C87D = OR(I374, I375)
--	C130D = OR(I371, I372)
--	C31D = OR(II368, I369)
--	C57D = OR(I365, I366)
--	C189D = OR(I362, I363)
--	C75D = OR(I359, I360)
--	C51D = OR(I356, I357)
--	C192D = OR(v8, I354)
--	C150D = OR(C30DE, I352)
--	C119D = OR(I349, v12, I350)
--	C91D = OR(I346, I347)
--	C84D = OR(C138DE, I344)
--	C160D = OR(I341, I342)
--	C109D = OR(I338, I339)
--	C125D = OR(I335, I336)
--	C139D = OR(I332, I333)
--	C69D = OR(I328, II329)
--	C175D = OR(I325, I326)
--	C122D = OR(v12, I323)
--	C34D = OR(I320, I321)
--	C63D = OR(v12E, I317, I318)
--	C161D = OR(I314, I315)
--	C195D = OR(C180DE, v9)
--	C72D = OR(I310, I311)
--	C112D = OR(I308, v9E)
--	C183D = OR(I305, I306)
--	C173D = OR(I302, I303)
--	C115D = OR(I299, I300)
--	C210D = OR(I296, I297)
--	Av13_D_19B = OR(I293, I294)
--	C143D = OR(C49DE, v9, I291)
--	C205D = OR(I287, I288)
--	C223D = OR(I284, I285)
--	C37D = OR(I280, I281, I282)
--	C133D = OR(C49DE, I278)
--	C28D = OR(I275, I276)
--	C202D = OR(I272, I273)
--	C73D = OR(I269, I270)
--	Av13_D_22B = OR(I266, I267)
--	C43D = OR(I262, I263)
--	C88D = OR(I259, I260)
--	C216D = OR(I256, I257)
--	C40D = OR(I253, II254)
--	C80D = OR(I250, I251)
--	C46D = OR(I247, I248)
--	C186D = OR(C49DE, I245)
--	C132D = OR(I242, I243)
--	C126D = OR(I239, I240)
--	C225D = OR(I236, I237)
--	C169D = OR(I232, I233, v12, I234)
--	C110D = OR(I229, I230)
--	C140D = OR(I226, I227)
--	C164D = OR(I222, I223, I224)
--	C52D = OR(I218, I219, I220)
--	C190D = OR(I215, I216)
--	C58D = OR(I212, I213)
--	C123D = OR(C157DE, I208, I209, I210)
--	C152D = OR(I205, I206)
--	C35D = OR(I202, I203)
--	C65D = OR(I199, I200)
--	C162D = OR(I196, I197)
--	C97D = OR(v11E, I194)
--	C199D = OR(I191, I192)
--	C176D = OR(I188, I189)
--	C181D = OR(I185, I186)
--	C184D = OR(I182, I183)
--	C174D = OR(I179, I180)
--	I491 = OR(I173, I174, I175)
--	C147D = OR(I176, I177, I491)
--	I497 = OR(C208DE, C83DE, I169)
--	C196D = OR(I170, v12, I171, I497)
--	C206D = OR(I166, I167)
--	C134D = OR(I163, I164)
--	C67D = OR(I160, I161)
--	C85D = OR(I156, I157, I158)
--	C53D = OR(I151, I152, I153, I154)
--	C113D = OR(I148, I149)
--	C224D = OR(I145, I146)
--	Av13_D_11B = OR(I140, I141, II142)
--	C48D = OR(I136, I137)
--	C153D = OR(I133, I134)
--	I542 = OR(I126, I127, I128)
--	C74D = OR(I129, I130, I131, I542)
--	Av13_D_10B = OR(I123, I124)
--	Av13_D_6B = OR(I119, I120)
--	C38D = OR(I116, I117)
--	C99D = OR(I111, I112, I113, I114)
--	C187D = OR(I108, I109)
--	C116D = OR(I103, I104, I105, I106)
--	C135D = OR(I100, I101)
--	C89D = OR(I95, I96, I97, I98)
--	Av13_D_8B = OR(I91, I92, I93)
--	Av13_D_1B = OR(I86, I87, I88, I89)
--	Av13_D_24B = OR(I82, I83, I84)
--	Av13_D_14B = OR(I78, I79, I80)
--	C177D = OR(I75, I76)
--	Av13_D_0B = OR(I71, I72, I73)
--	C207D = OR(I68, I69)
--	I610 = OR(I62, I63, I64)
--	C102D = OR(I65, I66, I610)
--	Av13_D_2B = OR(I58, I59, I60)
--	C188D = OR(I54, I55)
--	Av13_D_7B = OR(I51, I52)
--	Av13_D_12B = OR(I48, I49)
--	Av13_D_5B = OR(I43, I44, I45, I46)
--	Av13_D_4B = OR(I38, I39, I40, I41)
--	Av13_D_3B = OR(I34, I35, I36)
--	Av13_D_17B = OR(I31, I32)
--	Av13_D_13B = OR(I27, I28, I29)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s1494 is
	port (
		CLK: in std_logic;
		CLR: in std_logic;
		V0: in std_logic;
		V1: in std_logic;
		V2: in std_logic;
		V3: in std_logic;
		V4: in std_logic;
		V5: in std_logic;
		V6: in std_logic;
		V13_D_6: out std_logic;
		V13_D_7: out std_logic;
		V13_D_8: out std_logic;
		V13_D_9: out std_logic;
		V13_D_10: out std_logic;
		V13_D_11: out std_logic;
		V13_D_12: out std_logic;
		V13_D_13: out std_logic;
		V13_D_14: out std_logic;
		V13_D_15: out std_logic;
		V13_D_16: out std_logic;
		V13_D_17: out std_logic;
		V13_D_18: out std_logic;
		V13_D_19: out std_logic;
		V13_D_20: out std_logic;
		V13_D_21: out std_logic;
		V13_D_22: out std_logic;
		V13_D_23: out std_logic;
		V13_D_24: out std_logic
	);
end entity;

architecture RTL of s1494 is
	attribute dont_touch: boolean;

	signal AV13_D_0B: std_logic; attribute dont_touch of AV13_D_0B: signal is true;
	signal AV13_D_1B: std_logic; attribute dont_touch of AV13_D_1B: signal is true;
	signal AV13_D_2B: std_logic; attribute dont_touch of AV13_D_2B: signal is true;
	signal AV13_D_3B: std_logic; attribute dont_touch of AV13_D_3B: signal is true;
	signal AV13_D_4B: std_logic; attribute dont_touch of AV13_D_4B: signal is true;
	signal AV13_D_5B: std_logic; attribute dont_touch of AV13_D_5B: signal is true;
	signal AV13_D_6B: std_logic; attribute dont_touch of AV13_D_6B: signal is true;
	signal AV13_D_7B: std_logic; attribute dont_touch of AV13_D_7B: signal is true;
	signal AV13_D_8B: std_logic; attribute dont_touch of AV13_D_8B: signal is true;
	signal AV13_D_9B: std_logic; attribute dont_touch of AV13_D_9B: signal is true;
	signal AV13_D_10B: std_logic; attribute dont_touch of AV13_D_10B: signal is true;
	signal AV13_D_11B: std_logic; attribute dont_touch of AV13_D_11B: signal is true;
	signal AV13_D_12B: std_logic; attribute dont_touch of AV13_D_12B: signal is true;
	signal AV13_D_13B: std_logic; attribute dont_touch of AV13_D_13B: signal is true;
	signal AV13_D_14B: std_logic; attribute dont_touch of AV13_D_14B: signal is true;
	signal AV13_D_15B: std_logic; attribute dont_touch of AV13_D_15B: signal is true;
	signal AV13_D_16B: std_logic; attribute dont_touch of AV13_D_16B: signal is true;
	signal AV13_D_17B: std_logic; attribute dont_touch of AV13_D_17B: signal is true;
	signal AV13_D_18B: std_logic; attribute dont_touch of AV13_D_18B: signal is true;
	signal AV13_D_19B: std_logic; attribute dont_touch of AV13_D_19B: signal is true;
	signal AV13_D_20B: std_logic; attribute dont_touch of AV13_D_20B: signal is true;
	signal AV13_D_21B: std_logic; attribute dont_touch of AV13_D_21B: signal is true;
	signal AV13_D_22B: std_logic; attribute dont_touch of AV13_D_22B: signal is true;
	signal AV13_D_23B: std_logic; attribute dont_touch of AV13_D_23B: signal is true;
	signal AV13_D_24B: std_logic; attribute dont_touch of AV13_D_24B: signal is true;
	signal C26D: std_logic; attribute dont_touch of C26D: signal is true;
	signal C27D: std_logic; attribute dont_touch of C27D: signal is true;
	signal C28D: std_logic; attribute dont_touch of C28D: signal is true;
	signal C29D: std_logic; attribute dont_touch of C29D: signal is true;
	signal C30D: std_logic; attribute dont_touch of C30D: signal is true;
	signal C30DE: std_logic; attribute dont_touch of C30DE: signal is true;
	signal C31D: std_logic; attribute dont_touch of C31D: signal is true;
	signal C33D: std_logic; attribute dont_touch of C33D: signal is true;
	signal C34D: std_logic; attribute dont_touch of C34D: signal is true;
	signal C35D: std_logic; attribute dont_touch of C35D: signal is true;
	signal C36D: std_logic; attribute dont_touch of C36D: signal is true;
	signal C37D: std_logic; attribute dont_touch of C37D: signal is true;
	signal C38D: std_logic; attribute dont_touch of C38D: signal is true;
	signal C39D: std_logic; attribute dont_touch of C39D: signal is true;
	signal C40D: std_logic; attribute dont_touch of C40D: signal is true;
	signal C41D: std_logic; attribute dont_touch of C41D: signal is true;
	signal C42D: std_logic; attribute dont_touch of C42D: signal is true;
	signal C43D: std_logic; attribute dont_touch of C43D: signal is true;
	signal C44D: std_logic; attribute dont_touch of C44D: signal is true;
	signal C45D: std_logic; attribute dont_touch of C45D: signal is true;
	signal C46D: std_logic; attribute dont_touch of C46D: signal is true;
	signal C47D: std_logic; attribute dont_touch of C47D: signal is true;
	signal C48D: std_logic; attribute dont_touch of C48D: signal is true;
	signal C49D: std_logic; attribute dont_touch of C49D: signal is true;
	signal C49DE: std_logic; attribute dont_touch of C49DE: signal is true;
	signal C50D: std_logic; attribute dont_touch of C50D: signal is true;
	signal C51D: std_logic; attribute dont_touch of C51D: signal is true;
	signal C52D: std_logic; attribute dont_touch of C52D: signal is true;
	signal C53D: std_logic; attribute dont_touch of C53D: signal is true;
	signal C54D: std_logic; attribute dont_touch of C54D: signal is true;
	signal C55D: std_logic; attribute dont_touch of C55D: signal is true;
	signal C56D: std_logic; attribute dont_touch of C56D: signal is true;
	signal C57D: std_logic; attribute dont_touch of C57D: signal is true;
	signal C58D: std_logic; attribute dont_touch of C58D: signal is true;
	signal C59D: std_logic; attribute dont_touch of C59D: signal is true;
	signal C60D: std_logic; attribute dont_touch of C60D: signal is true;
	signal C63D: std_logic; attribute dont_touch of C63D: signal is true;
	signal C65D: std_logic; attribute dont_touch of C65D: signal is true;
	signal C67D: std_logic; attribute dont_touch of C67D: signal is true;
	signal C69D: std_logic; attribute dont_touch of C69D: signal is true;
	signal C70D: std_logic; attribute dont_touch of C70D: signal is true;
	signal C70DE: std_logic; attribute dont_touch of C70DE: signal is true;
	signal C71D: std_logic; attribute dont_touch of C71D: signal is true;
	signal C72D: std_logic; attribute dont_touch of C72D: signal is true;
	signal C73D: std_logic; attribute dont_touch of C73D: signal is true;
	signal C74D: std_logic; attribute dont_touch of C74D: signal is true;
	signal C75D: std_logic; attribute dont_touch of C75D: signal is true;
	signal C76D: std_logic; attribute dont_touch of C76D: signal is true;
	signal C77D: std_logic; attribute dont_touch of C77D: signal is true;
	signal C78D: std_logic; attribute dont_touch of C78D: signal is true;
	signal C79D: std_logic; attribute dont_touch of C79D: signal is true;
	signal C80D: std_logic; attribute dont_touch of C80D: signal is true;
	signal C81D: std_logic; attribute dont_touch of C81D: signal is true;
	signal C81DE: std_logic; attribute dont_touch of C81DE: signal is true;
	signal C82D: std_logic; attribute dont_touch of C82D: signal is true;
	signal C83D: std_logic; attribute dont_touch of C83D: signal is true;
	signal C83DE: std_logic; attribute dont_touch of C83DE: signal is true;
	signal C84D: std_logic; attribute dont_touch of C84D: signal is true;
	signal C85D: std_logic; attribute dont_touch of C85D: signal is true;
	signal C86D: std_logic; attribute dont_touch of C86D: signal is true;
	signal C87D: std_logic; attribute dont_touch of C87D: signal is true;
	signal C88D: std_logic; attribute dont_touch of C88D: signal is true;
	signal C89D: std_logic; attribute dont_touch of C89D: signal is true;
	signal C90D: std_logic; attribute dont_touch of C90D: signal is true;
	signal C90DE: std_logic; attribute dont_touch of C90DE: signal is true;
	signal C91D: std_logic; attribute dont_touch of C91D: signal is true;
	signal C92D: std_logic; attribute dont_touch of C92D: signal is true;
	signal C93D: std_logic; attribute dont_touch of C93D: signal is true;
	signal C95D: std_logic; attribute dont_touch of C95D: signal is true;
	signal C96D: std_logic; attribute dont_touch of C96D: signal is true;
	signal C97D: std_logic; attribute dont_touch of C97D: signal is true;
	signal C98D: std_logic; attribute dont_touch of C98D: signal is true;
	signal C99D: std_logic; attribute dont_touch of C99D: signal is true;
	signal C100D: std_logic; attribute dont_touch of C100D: signal is true;
	signal C102D: std_logic; attribute dont_touch of C102D: signal is true;
	signal C103D: std_logic; attribute dont_touch of C103D: signal is true;
	signal C104D: std_logic; attribute dont_touch of C104D: signal is true;
	signal C104DE: std_logic; attribute dont_touch of C104DE: signal is true;
	signal C105D: std_logic; attribute dont_touch of C105D: signal is true;
	signal C106D: std_logic; attribute dont_touch of C106D: signal is true;
	signal C107D: std_logic; attribute dont_touch of C107D: signal is true;
	signal C108D: std_logic; attribute dont_touch of C108D: signal is true;
	signal C108DE: std_logic; attribute dont_touch of C108DE: signal is true;
	signal C109D: std_logic; attribute dont_touch of C109D: signal is true;
	signal C110D: std_logic; attribute dont_touch of C110D: signal is true;
	signal C111D: std_logic; attribute dont_touch of C111D: signal is true;
	signal C112D: std_logic; attribute dont_touch of C112D: signal is true;
	signal C113D: std_logic; attribute dont_touch of C113D: signal is true;
	signal C114D: std_logic; attribute dont_touch of C114D: signal is true;
	signal C115D: std_logic; attribute dont_touch of C115D: signal is true;
	signal C116D: std_logic; attribute dont_touch of C116D: signal is true;
	signal C117D: std_logic; attribute dont_touch of C117D: signal is true;
	signal C117DE: std_logic; attribute dont_touch of C117DE: signal is true;
	signal C118D: std_logic; attribute dont_touch of C118D: signal is true;
	signal C118DE: std_logic; attribute dont_touch of C118DE: signal is true;
	signal C119D: std_logic; attribute dont_touch of C119D: signal is true;
	signal C120D: std_logic; attribute dont_touch of C120D: signal is true;
	signal C122D: std_logic; attribute dont_touch of C122D: signal is true;
	signal C123D: std_logic; attribute dont_touch of C123D: signal is true;
	signal C124D: std_logic; attribute dont_touch of C124D: signal is true;
	signal C124DE: std_logic; attribute dont_touch of C124DE: signal is true;
	signal C125D: std_logic; attribute dont_touch of C125D: signal is true;
	signal C126D: std_logic; attribute dont_touch of C126D: signal is true;
	signal C127D: std_logic; attribute dont_touch of C127D: signal is true;
	signal C128D: std_logic; attribute dont_touch of C128D: signal is true;
	signal C129D: std_logic; attribute dont_touch of C129D: signal is true;
	signal C129DE: std_logic; attribute dont_touch of C129DE: signal is true;
	signal C130D: std_logic; attribute dont_touch of C130D: signal is true;
	signal C131D: std_logic; attribute dont_touch of C131D: signal is true;
	signal C131DE: std_logic; attribute dont_touch of C131DE: signal is true;
	signal C132D: std_logic; attribute dont_touch of C132D: signal is true;
	signal C133D: std_logic; attribute dont_touch of C133D: signal is true;
	signal C134D: std_logic; attribute dont_touch of C134D: signal is true;
	signal C135D: std_logic; attribute dont_touch of C135D: signal is true;
	signal C137D: std_logic; attribute dont_touch of C137D: signal is true;
	signal C138D: std_logic; attribute dont_touch of C138D: signal is true;
	signal C138DE: std_logic; attribute dont_touch of C138DE: signal is true;
	signal C139D: std_logic; attribute dont_touch of C139D: signal is true;
	signal C140D: std_logic; attribute dont_touch of C140D: signal is true;
	signal C141D: std_logic; attribute dont_touch of C141D: signal is true;
	signal C141DE: std_logic; attribute dont_touch of C141DE: signal is true;
	signal C142D: std_logic; attribute dont_touch of C142D: signal is true;
	signal C143D: std_logic; attribute dont_touch of C143D: signal is true;
	signal C144D: std_logic; attribute dont_touch of C144D: signal is true;
	signal C144DE: std_logic; attribute dont_touch of C144DE: signal is true;
	signal C145D: std_logic; attribute dont_touch of C145D: signal is true;
	signal C146D: std_logic; attribute dont_touch of C146D: signal is true;
	signal C147D: std_logic; attribute dont_touch of C147D: signal is true;
	signal C148D: std_logic; attribute dont_touch of C148D: signal is true;
	signal C150D: std_logic; attribute dont_touch of C150D: signal is true;
	signal C151D: std_logic; attribute dont_touch of C151D: signal is true;
	signal C152D: std_logic; attribute dont_touch of C152D: signal is true;
	signal C153D: std_logic; attribute dont_touch of C153D: signal is true;
	signal C155D: std_logic; attribute dont_touch of C155D: signal is true;
	signal C156D: std_logic; attribute dont_touch of C156D: signal is true;
	signal C157D: std_logic; attribute dont_touch of C157D: signal is true;
	signal C157DE: std_logic; attribute dont_touch of C157DE: signal is true;
	signal C158D: std_logic; attribute dont_touch of C158D: signal is true;
	signal C159D: std_logic; attribute dont_touch of C159D: signal is true;
	signal C160D: std_logic; attribute dont_touch of C160D: signal is true;
	signal C161D: std_logic; attribute dont_touch of C161D: signal is true;
	signal C162D: std_logic; attribute dont_touch of C162D: signal is true;
	signal C163D: std_logic; attribute dont_touch of C163D: signal is true;
	signal C164D: std_logic; attribute dont_touch of C164D: signal is true;
	signal C165D: std_logic; attribute dont_touch of C165D: signal is true;
	signal C165DE: std_logic; attribute dont_touch of C165DE: signal is true;
	signal C166D: std_logic; attribute dont_touch of C166D: signal is true;
	signal C166DE: std_logic; attribute dont_touch of C166DE: signal is true;
	signal C167D: std_logic; attribute dont_touch of C167D: signal is true;
	signal C168D: std_logic; attribute dont_touch of C168D: signal is true;
	signal C169D: std_logic; attribute dont_touch of C169D: signal is true;
	signal C170D: std_logic; attribute dont_touch of C170D: signal is true;
	signal C172D: std_logic; attribute dont_touch of C172D: signal is true;
	signal C173D: std_logic; attribute dont_touch of C173D: signal is true;
	signal C174D: std_logic; attribute dont_touch of C174D: signal is true;
	signal C175D: std_logic; attribute dont_touch of C175D: signal is true;
	signal C176D: std_logic; attribute dont_touch of C176D: signal is true;
	signal C177D: std_logic; attribute dont_touch of C177D: signal is true;
	signal C178D: std_logic; attribute dont_touch of C178D: signal is true;
	signal C179D: std_logic; attribute dont_touch of C179D: signal is true;
	signal C180D: std_logic; attribute dont_touch of C180D: signal is true;
	signal C180DE: std_logic; attribute dont_touch of C180DE: signal is true;
	signal C181D: std_logic; attribute dont_touch of C181D: signal is true;
	signal C183D: std_logic; attribute dont_touch of C183D: signal is true;
	signal C184D: std_logic; attribute dont_touch of C184D: signal is true;
	signal C185D: std_logic; attribute dont_touch of C185D: signal is true;
	signal C186D: std_logic; attribute dont_touch of C186D: signal is true;
	signal C187D: std_logic; attribute dont_touch of C187D: signal is true;
	signal C188D: std_logic; attribute dont_touch of C188D: signal is true;
	signal C189D: std_logic; attribute dont_touch of C189D: signal is true;
	signal C190D: std_logic; attribute dont_touch of C190D: signal is true;
	signal C191D: std_logic; attribute dont_touch of C191D: signal is true;
	signal C191DE: std_logic; attribute dont_touch of C191DE: signal is true;
	signal C192D: std_logic; attribute dont_touch of C192D: signal is true;
	signal C193D: std_logic; attribute dont_touch of C193D: signal is true;
	signal C194D: std_logic; attribute dont_touch of C194D: signal is true;
	signal C194DE: std_logic; attribute dont_touch of C194DE: signal is true;
	signal C195D: std_logic; attribute dont_touch of C195D: signal is true;
	signal C195DE: std_logic; attribute dont_touch of C195DE: signal is true;
	signal C196D: std_logic; attribute dont_touch of C196D: signal is true;
	signal C199D: std_logic; attribute dont_touch of C199D: signal is true;
	signal C200D: std_logic; attribute dont_touch of C200D: signal is true;
	signal C201D: std_logic; attribute dont_touch of C201D: signal is true;
	signal C202D: std_logic; attribute dont_touch of C202D: signal is true;
	signal C203D: std_logic; attribute dont_touch of C203D: signal is true;
	signal C205D: std_logic; attribute dont_touch of C205D: signal is true;
	signal C206D: std_logic; attribute dont_touch of C206D: signal is true;
	signal C207D: std_logic; attribute dont_touch of C207D: signal is true;
	signal C208D: std_logic; attribute dont_touch of C208D: signal is true;
	signal C208DE: std_logic; attribute dont_touch of C208DE: signal is true;
	signal C209D: std_logic; attribute dont_touch of C209D: signal is true;
	signal C210D: std_logic; attribute dont_touch of C210D: signal is true;
	signal C211D: std_logic; attribute dont_touch of C211D: signal is true;
	signal C213D: std_logic; attribute dont_touch of C213D: signal is true;
	signal C214D: std_logic; attribute dont_touch of C214D: signal is true;
	signal C215D: std_logic; attribute dont_touch of C215D: signal is true;
	signal C216D: std_logic; attribute dont_touch of C216D: signal is true;
	signal C217D: std_logic; attribute dont_touch of C217D: signal is true;
	signal C218D: std_logic; attribute dont_touch of C218D: signal is true;
	signal C218DE: std_logic; attribute dont_touch of C218DE: signal is true;
	signal C219D: std_logic; attribute dont_touch of C219D: signal is true;
	signal C220D: std_logic; attribute dont_touch of C220D: signal is true;
	signal C220DE: std_logic; attribute dont_touch of C220DE: signal is true;
	signal C221D: std_logic; attribute dont_touch of C221D: signal is true;
	signal C222D: std_logic; attribute dont_touch of C222D: signal is true;
	signal C223D: std_logic; attribute dont_touch of C223D: signal is true;
	signal C224D: std_logic; attribute dont_touch of C224D: signal is true;
	signal C225D: std_logic; attribute dont_touch of C225D: signal is true;
	signal I27: std_logic; attribute dont_touch of I27: signal is true;
	signal I28: std_logic; attribute dont_touch of I28: signal is true;
	signal I29: std_logic; attribute dont_touch of I29: signal is true;
	signal I31: std_logic; attribute dont_touch of I31: signal is true;
	signal I32: std_logic; attribute dont_touch of I32: signal is true;
	signal I34: std_logic; attribute dont_touch of I34: signal is true;
	signal I35: std_logic; attribute dont_touch of I35: signal is true;
	signal I36: std_logic; attribute dont_touch of I36: signal is true;
	signal I38: std_logic; attribute dont_touch of I38: signal is true;
	signal I39: std_logic; attribute dont_touch of I39: signal is true;
	signal I40: std_logic; attribute dont_touch of I40: signal is true;
	signal I41: std_logic; attribute dont_touch of I41: signal is true;
	signal I43: std_logic; attribute dont_touch of I43: signal is true;
	signal I44: std_logic; attribute dont_touch of I44: signal is true;
	signal I45: std_logic; attribute dont_touch of I45: signal is true;
	signal I46: std_logic; attribute dont_touch of I46: signal is true;
	signal I48: std_logic; attribute dont_touch of I48: signal is true;
	signal I49: std_logic; attribute dont_touch of I49: signal is true;
	signal I51: std_logic; attribute dont_touch of I51: signal is true;
	signal I52: std_logic; attribute dont_touch of I52: signal is true;
	signal I54: std_logic; attribute dont_touch of I54: signal is true;
	signal I55: std_logic; attribute dont_touch of I55: signal is true;
	signal I58: std_logic; attribute dont_touch of I58: signal is true;
	signal I59: std_logic; attribute dont_touch of I59: signal is true;
	signal I60: std_logic; attribute dont_touch of I60: signal is true;
	signal I62: std_logic; attribute dont_touch of I62: signal is true;
	signal I63: std_logic; attribute dont_touch of I63: signal is true;
	signal I64: std_logic; attribute dont_touch of I64: signal is true;
	signal I65: std_logic; attribute dont_touch of I65: signal is true;
	signal I66: std_logic; attribute dont_touch of I66: signal is true;
	signal I68: std_logic; attribute dont_touch of I68: signal is true;
	signal I69: std_logic; attribute dont_touch of I69: signal is true;
	signal I71: std_logic; attribute dont_touch of I71: signal is true;
	signal I72: std_logic; attribute dont_touch of I72: signal is true;
	signal I73: std_logic; attribute dont_touch of I73: signal is true;
	signal I75: std_logic; attribute dont_touch of I75: signal is true;
	signal I76: std_logic; attribute dont_touch of I76: signal is true;
	signal I78: std_logic; attribute dont_touch of I78: signal is true;
	signal I79: std_logic; attribute dont_touch of I79: signal is true;
	signal I80: std_logic; attribute dont_touch of I80: signal is true;
	signal I82: std_logic; attribute dont_touch of I82: signal is true;
	signal I83: std_logic; attribute dont_touch of I83: signal is true;
	signal I84: std_logic; attribute dont_touch of I84: signal is true;
	signal I86: std_logic; attribute dont_touch of I86: signal is true;
	signal I87: std_logic; attribute dont_touch of I87: signal is true;
	signal I88: std_logic; attribute dont_touch of I88: signal is true;
	signal I89: std_logic; attribute dont_touch of I89: signal is true;
	signal I91: std_logic; attribute dont_touch of I91: signal is true;
	signal I92: std_logic; attribute dont_touch of I92: signal is true;
	signal I93: std_logic; attribute dont_touch of I93: signal is true;
	signal I95: std_logic; attribute dont_touch of I95: signal is true;
	signal I96: std_logic; attribute dont_touch of I96: signal is true;
	signal I97: std_logic; attribute dont_touch of I97: signal is true;
	signal I98: std_logic; attribute dont_touch of I98: signal is true;
	signal I100: std_logic; attribute dont_touch of I100: signal is true;
	signal I101: std_logic; attribute dont_touch of I101: signal is true;
	signal I103: std_logic; attribute dont_touch of I103: signal is true;
	signal I104: std_logic; attribute dont_touch of I104: signal is true;
	signal I105: std_logic; attribute dont_touch of I105: signal is true;
	signal I106: std_logic; attribute dont_touch of I106: signal is true;
	signal I108: std_logic; attribute dont_touch of I108: signal is true;
	signal I109: std_logic; attribute dont_touch of I109: signal is true;
	signal I111: std_logic; attribute dont_touch of I111: signal is true;
	signal I112: std_logic; attribute dont_touch of I112: signal is true;
	signal I113: std_logic; attribute dont_touch of I113: signal is true;
	signal I114: std_logic; attribute dont_touch of I114: signal is true;
	signal I116: std_logic; attribute dont_touch of I116: signal is true;
	signal I117: std_logic; attribute dont_touch of I117: signal is true;
	signal I119: std_logic; attribute dont_touch of I119: signal is true;
	signal I120: std_logic; attribute dont_touch of I120: signal is true;
	signal I123: std_logic; attribute dont_touch of I123: signal is true;
	signal I124: std_logic; attribute dont_touch of I124: signal is true;
	signal I126: std_logic; attribute dont_touch of I126: signal is true;
	signal I127: std_logic; attribute dont_touch of I127: signal is true;
	signal I128: std_logic; attribute dont_touch of I128: signal is true;
	signal I129: std_logic; attribute dont_touch of I129: signal is true;
	signal I130: std_logic; attribute dont_touch of I130: signal is true;
	signal I131: std_logic; attribute dont_touch of I131: signal is true;
	signal I133: std_logic; attribute dont_touch of I133: signal is true;
	signal I134: std_logic; attribute dont_touch of I134: signal is true;
	signal I136: std_logic; attribute dont_touch of I136: signal is true;
	signal I137: std_logic; attribute dont_touch of I137: signal is true;
	signal I140: std_logic; attribute dont_touch of I140: signal is true;
	signal I141: std_logic; attribute dont_touch of I141: signal is true;
	signal I142: std_logic; attribute dont_touch of I142: signal is true;
	signal I145: std_logic; attribute dont_touch of I145: signal is true;
	signal I146: std_logic; attribute dont_touch of I146: signal is true;
	signal I148: std_logic; attribute dont_touch of I148: signal is true;
	signal I149: std_logic; attribute dont_touch of I149: signal is true;
	signal I151: std_logic; attribute dont_touch of I151: signal is true;
	signal I152: std_logic; attribute dont_touch of I152: signal is true;
	signal I153: std_logic; attribute dont_touch of I153: signal is true;
	signal I154: std_logic; attribute dont_touch of I154: signal is true;
	signal I156: std_logic; attribute dont_touch of I156: signal is true;
	signal I157: std_logic; attribute dont_touch of I157: signal is true;
	signal I158: std_logic; attribute dont_touch of I158: signal is true;
	signal I160: std_logic; attribute dont_touch of I160: signal is true;
	signal I161: std_logic; attribute dont_touch of I161: signal is true;
	signal I163: std_logic; attribute dont_touch of I163: signal is true;
	signal I164: std_logic; attribute dont_touch of I164: signal is true;
	signal I166: std_logic; attribute dont_touch of I166: signal is true;
	signal I167: std_logic; attribute dont_touch of I167: signal is true;
	signal I169: std_logic; attribute dont_touch of I169: signal is true;
	signal I170: std_logic; attribute dont_touch of I170: signal is true;
	signal I171: std_logic; attribute dont_touch of I171: signal is true;
	signal I173: std_logic; attribute dont_touch of I173: signal is true;
	signal I174: std_logic; attribute dont_touch of I174: signal is true;
	signal I175: std_logic; attribute dont_touch of I175: signal is true;
	signal I176: std_logic; attribute dont_touch of I176: signal is true;
	signal I177: std_logic; attribute dont_touch of I177: signal is true;
	signal I179: std_logic; attribute dont_touch of I179: signal is true;
	signal I180: std_logic; attribute dont_touch of I180: signal is true;
	signal I182: std_logic; attribute dont_touch of I182: signal is true;
	signal I183: std_logic; attribute dont_touch of I183: signal is true;
	signal I185: std_logic; attribute dont_touch of I185: signal is true;
	signal I186: std_logic; attribute dont_touch of I186: signal is true;
	signal I188: std_logic; attribute dont_touch of I188: signal is true;
	signal I189: std_logic; attribute dont_touch of I189: signal is true;
	signal I191: std_logic; attribute dont_touch of I191: signal is true;
	signal I192: std_logic; attribute dont_touch of I192: signal is true;
	signal I194: std_logic; attribute dont_touch of I194: signal is true;
	signal I196: std_logic; attribute dont_touch of I196: signal is true;
	signal I197: std_logic; attribute dont_touch of I197: signal is true;
	signal I199: std_logic; attribute dont_touch of I199: signal is true;
	signal I200: std_logic; attribute dont_touch of I200: signal is true;
	signal I202: std_logic; attribute dont_touch of I202: signal is true;
	signal I203: std_logic; attribute dont_touch of I203: signal is true;
	signal I205: std_logic; attribute dont_touch of I205: signal is true;
	signal I206: std_logic; attribute dont_touch of I206: signal is true;
	signal I208: std_logic; attribute dont_touch of I208: signal is true;
	signal I209: std_logic; attribute dont_touch of I209: signal is true;
	signal I210: std_logic; attribute dont_touch of I210: signal is true;
	signal I212: std_logic; attribute dont_touch of I212: signal is true;
	signal I213: std_logic; attribute dont_touch of I213: signal is true;
	signal I215: std_logic; attribute dont_touch of I215: signal is true;
	signal I216: std_logic; attribute dont_touch of I216: signal is true;
	signal I218: std_logic; attribute dont_touch of I218: signal is true;
	signal I219: std_logic; attribute dont_touch of I219: signal is true;
	signal I220: std_logic; attribute dont_touch of I220: signal is true;
	signal I222: std_logic; attribute dont_touch of I222: signal is true;
	signal I223: std_logic; attribute dont_touch of I223: signal is true;
	signal I224: std_logic; attribute dont_touch of I224: signal is true;
	signal I226: std_logic; attribute dont_touch of I226: signal is true;
	signal I227: std_logic; attribute dont_touch of I227: signal is true;
	signal I229: std_logic; attribute dont_touch of I229: signal is true;
	signal I230: std_logic; attribute dont_touch of I230: signal is true;
	signal I232: std_logic; attribute dont_touch of I232: signal is true;
	signal I233: std_logic; attribute dont_touch of I233: signal is true;
	signal I234: std_logic; attribute dont_touch of I234: signal is true;
	signal I236: std_logic; attribute dont_touch of I236: signal is true;
	signal I237: std_logic; attribute dont_touch of I237: signal is true;
	signal I239: std_logic; attribute dont_touch of I239: signal is true;
	signal I240: std_logic; attribute dont_touch of I240: signal is true;
	signal I242: std_logic; attribute dont_touch of I242: signal is true;
	signal I243: std_logic; attribute dont_touch of I243: signal is true;
	signal I245: std_logic; attribute dont_touch of I245: signal is true;
	signal I247: std_logic; attribute dont_touch of I247: signal is true;
	signal I248: std_logic; attribute dont_touch of I248: signal is true;
	signal I250: std_logic; attribute dont_touch of I250: signal is true;
	signal I251: std_logic; attribute dont_touch of I251: signal is true;
	signal I253: std_logic; attribute dont_touch of I253: signal is true;
	signal I254: std_logic; attribute dont_touch of I254: signal is true;
	signal I256: std_logic; attribute dont_touch of I256: signal is true;
	signal I257: std_logic; attribute dont_touch of I257: signal is true;
	signal I259: std_logic; attribute dont_touch of I259: signal is true;
	signal I260: std_logic; attribute dont_touch of I260: signal is true;
	signal I262: std_logic; attribute dont_touch of I262: signal is true;
	signal I263: std_logic; attribute dont_touch of I263: signal is true;
	signal I266: std_logic; attribute dont_touch of I266: signal is true;
	signal I267: std_logic; attribute dont_touch of I267: signal is true;
	signal I269: std_logic; attribute dont_touch of I269: signal is true;
	signal I270: std_logic; attribute dont_touch of I270: signal is true;
	signal I272: std_logic; attribute dont_touch of I272: signal is true;
	signal I273: std_logic; attribute dont_touch of I273: signal is true;
	signal I275: std_logic; attribute dont_touch of I275: signal is true;
	signal I276: std_logic; attribute dont_touch of I276: signal is true;
	signal I278: std_logic; attribute dont_touch of I278: signal is true;
	signal I280: std_logic; attribute dont_touch of I280: signal is true;
	signal I281: std_logic; attribute dont_touch of I281: signal is true;
	signal I282: std_logic; attribute dont_touch of I282: signal is true;
	signal I284: std_logic; attribute dont_touch of I284: signal is true;
	signal I285: std_logic; attribute dont_touch of I285: signal is true;
	signal I287: std_logic; attribute dont_touch of I287: signal is true;
	signal I288: std_logic; attribute dont_touch of I288: signal is true;
	signal I291: std_logic; attribute dont_touch of I291: signal is true;
	signal I293: std_logic; attribute dont_touch of I293: signal is true;
	signal I294: std_logic; attribute dont_touch of I294: signal is true;
	signal I296: std_logic; attribute dont_touch of I296: signal is true;
	signal I297: std_logic; attribute dont_touch of I297: signal is true;
	signal I299: std_logic; attribute dont_touch of I299: signal is true;
	signal I300: std_logic; attribute dont_touch of I300: signal is true;
	signal I302: std_logic; attribute dont_touch of I302: signal is true;
	signal I303: std_logic; attribute dont_touch of I303: signal is true;
	signal I305: std_logic; attribute dont_touch of I305: signal is true;
	signal I306: std_logic; attribute dont_touch of I306: signal is true;
	signal I308: std_logic; attribute dont_touch of I308: signal is true;
	signal I310: std_logic; attribute dont_touch of I310: signal is true;
	signal I311: std_logic; attribute dont_touch of I311: signal is true;
	signal I314: std_logic; attribute dont_touch of I314: signal is true;
	signal I315: std_logic; attribute dont_touch of I315: signal is true;
	signal I317: std_logic; attribute dont_touch of I317: signal is true;
	signal I318: std_logic; attribute dont_touch of I318: signal is true;
	signal I320: std_logic; attribute dont_touch of I320: signal is true;
	signal I321: std_logic; attribute dont_touch of I321: signal is true;
	signal I323: std_logic; attribute dont_touch of I323: signal is true;
	signal I325: std_logic; attribute dont_touch of I325: signal is true;
	signal I326: std_logic; attribute dont_touch of I326: signal is true;
	signal I328: std_logic; attribute dont_touch of I328: signal is true;
	signal I329: std_logic; attribute dont_touch of I329: signal is true;
	signal I332: std_logic; attribute dont_touch of I332: signal is true;
	signal I333: std_logic; attribute dont_touch of I333: signal is true;
	signal I335: std_logic; attribute dont_touch of I335: signal is true;
	signal I336: std_logic; attribute dont_touch of I336: signal is true;
	signal I338: std_logic; attribute dont_touch of I338: signal is true;
	signal I339: std_logic; attribute dont_touch of I339: signal is true;
	signal I341: std_logic; attribute dont_touch of I341: signal is true;
	signal I342: std_logic; attribute dont_touch of I342: signal is true;
	signal I344: std_logic; attribute dont_touch of I344: signal is true;
	signal I346: std_logic; attribute dont_touch of I346: signal is true;
	signal I347: std_logic; attribute dont_touch of I347: signal is true;
	signal I349: std_logic; attribute dont_touch of I349: signal is true;
	signal I350: std_logic; attribute dont_touch of I350: signal is true;
	signal I352: std_logic; attribute dont_touch of I352: signal is true;
	signal I354: std_logic; attribute dont_touch of I354: signal is true;
	signal I356: std_logic; attribute dont_touch of I356: signal is true;
	signal I357: std_logic; attribute dont_touch of I357: signal is true;
	signal I359: std_logic; attribute dont_touch of I359: signal is true;
	signal I360: std_logic; attribute dont_touch of I360: signal is true;
	signal I362: std_logic; attribute dont_touch of I362: signal is true;
	signal I363: std_logic; attribute dont_touch of I363: signal is true;
	signal I365: std_logic; attribute dont_touch of I365: signal is true;
	signal I366: std_logic; attribute dont_touch of I366: signal is true;
	signal I368: std_logic; attribute dont_touch of I368: signal is true;
	signal I369: std_logic; attribute dont_touch of I369: signal is true;
	signal I371: std_logic; attribute dont_touch of I371: signal is true;
	signal I372: std_logic; attribute dont_touch of I372: signal is true;
	signal I374: std_logic; attribute dont_touch of I374: signal is true;
	signal I375: std_logic; attribute dont_touch of I375: signal is true;
	signal I377: std_logic; attribute dont_touch of I377: signal is true;
	signal I378: std_logic; attribute dont_touch of I378: signal is true;
	signal I380: std_logic; attribute dont_touch of I380: signal is true;
	signal I381: std_logic; attribute dont_touch of I381: signal is true;
	signal I383: std_logic; attribute dont_touch of I383: signal is true;
	signal I384: std_logic; attribute dont_touch of I384: signal is true;
	signal I386: std_logic; attribute dont_touch of I386: signal is true;
	signal I387: std_logic; attribute dont_touch of I387: signal is true;
	signal I389: std_logic; attribute dont_touch of I389: signal is true;
	signal I390: std_logic; attribute dont_touch of I390: signal is true;
	signal I392: std_logic; attribute dont_touch of I392: signal is true;
	signal I393: std_logic; attribute dont_touch of I393: signal is true;
	signal I395: std_logic; attribute dont_touch of I395: signal is true;
	signal I396: std_logic; attribute dont_touch of I396: signal is true;
	signal I398: std_logic; attribute dont_touch of I398: signal is true;
	signal I399: std_logic; attribute dont_touch of I399: signal is true;
	signal I402: std_logic; attribute dont_touch of I402: signal is true;
	signal I403: std_logic; attribute dont_touch of I403: signal is true;
	signal I405: std_logic; attribute dont_touch of I405: signal is true;
	signal I406: std_logic; attribute dont_touch of I406: signal is true;
	signal I409: std_logic; attribute dont_touch of I409: signal is true;
	signal I412: std_logic; attribute dont_touch of I412: signal is true;
	signal I414: std_logic; attribute dont_touch of I414: signal is true;
	signal I415: std_logic; attribute dont_touch of I415: signal is true;
	signal I417: std_logic; attribute dont_touch of I417: signal is true;
	signal I419: std_logic; attribute dont_touch of I419: signal is true;
	signal I420: std_logic; attribute dont_touch of I420: signal is true;
	signal I423: std_logic; attribute dont_touch of I423: signal is true;
	signal I425: std_logic; attribute dont_touch of I425: signal is true;
	signal I427: std_logic; attribute dont_touch of I427: signal is true;
	signal I429: std_logic; attribute dont_touch of I429: signal is true;
	signal I430: std_logic; attribute dont_touch of I430: signal is true;
	signal I432: std_logic; attribute dont_touch of I432: signal is true;
	signal I433: std_logic; attribute dont_touch of I433: signal is true;
	signal I435: std_logic; attribute dont_touch of I435: signal is true;
	signal I436: std_logic; attribute dont_touch of I436: signal is true;
	signal I438: std_logic; attribute dont_touch of I438: signal is true;
	signal I439: std_logic; attribute dont_touch of I439: signal is true;
	signal I441: std_logic; attribute dont_touch of I441: signal is true;
	signal I442: std_logic; attribute dont_touch of I442: signal is true;
	signal I444: std_logic; attribute dont_touch of I444: signal is true;
	signal I446: std_logic; attribute dont_touch of I446: signal is true;
	signal I447: std_logic; attribute dont_touch of I447: signal is true;
	signal I449: std_logic; attribute dont_touch of I449: signal is true;
	signal I450: std_logic; attribute dont_touch of I450: signal is true;
	signal I452: std_logic; attribute dont_touch of I452: signal is true;
	signal I453: std_logic; attribute dont_touch of I453: signal is true;
	signal I456: std_logic; attribute dont_touch of I456: signal is true;
	signal I457: std_logic; attribute dont_touch of I457: signal is true;
	signal I460: std_logic; attribute dont_touch of I460: signal is true;
	signal I461: std_logic; attribute dont_touch of I461: signal is true;
	signal I463: std_logic; attribute dont_touch of I463: signal is true;
	signal I464: std_logic; attribute dont_touch of I464: signal is true;
	signal I466: std_logic; attribute dont_touch of I466: signal is true;
	signal I468: std_logic; attribute dont_touch of I468: signal is true;
	signal I470: std_logic; attribute dont_touch of I470: signal is true;
	signal I471: std_logic; attribute dont_touch of I471: signal is true;
	signal I473: std_logic; attribute dont_touch of I473: signal is true;
	signal I475: std_logic; attribute dont_touch of I475: signal is true;
	signal I476: std_logic; attribute dont_touch of I476: signal is true;
	signal I478: std_logic; attribute dont_touch of I478: signal is true;
	signal I479: std_logic; attribute dont_touch of I479: signal is true;
	signal I482: std_logic; attribute dont_touch of I482: signal is true;
	signal I483: std_logic; attribute dont_touch of I483: signal is true;
	signal I485: std_logic; attribute dont_touch of I485: signal is true;
	signal I486: std_logic; attribute dont_touch of I486: signal is true;
	signal I489: std_logic; attribute dont_touch of I489: signal is true;
	signal I491: std_logic; attribute dont_touch of I491: signal is true;
	signal I492: std_logic; attribute dont_touch of I492: signal is true;
	signal I494: std_logic; attribute dont_touch of I494: signal is true;
	signal I495: std_logic; attribute dont_touch of I495: signal is true;
	signal I497: std_logic; attribute dont_touch of I497: signal is true;
	signal I498: std_logic; attribute dont_touch of I498: signal is true;
	signal I500: std_logic; attribute dont_touch of I500: signal is true;
	signal I501: std_logic; attribute dont_touch of I501: signal is true;
	signal I503: std_logic; attribute dont_touch of I503: signal is true;
	signal I505: std_logic; attribute dont_touch of I505: signal is true;
	signal I506: std_logic; attribute dont_touch of I506: signal is true;
	signal I508: std_logic; attribute dont_touch of I508: signal is true;
	signal I510: std_logic; attribute dont_touch of I510: signal is true;
	signal I513: std_logic; attribute dont_touch of I513: signal is true;
	signal I514: std_logic; attribute dont_touch of I514: signal is true;
	signal I516: std_logic; attribute dont_touch of I516: signal is true;
	signal I518: std_logic; attribute dont_touch of I518: signal is true;
	signal I520: std_logic; attribute dont_touch of I520: signal is true;
	signal I524: std_logic; attribute dont_touch of I524: signal is true;
	signal I528: std_logic; attribute dont_touch of I528: signal is true;
	signal I533: std_logic; attribute dont_touch of I533: signal is true;
	signal I534: std_logic; attribute dont_touch of I534: signal is true;
	signal I537: std_logic; attribute dont_touch of I537: signal is true;
	signal I538: std_logic; attribute dont_touch of I538: signal is true;
	signal I542: std_logic; attribute dont_touch of I542: signal is true;
	signal I546: std_logic; attribute dont_touch of I546: signal is true;
	signal I547: std_logic; attribute dont_touch of I547: signal is true;
	signal I548: std_logic; attribute dont_touch of I548: signal is true;
	signal I554: std_logic; attribute dont_touch of I554: signal is true;
	signal I555: std_logic; attribute dont_touch of I555: signal is true;
	signal I559: std_logic; attribute dont_touch of I559: signal is true;
	signal I560: std_logic; attribute dont_touch of I560: signal is true;
	signal I610: std_logic; attribute dont_touch of I610: signal is true;
	signal I642: std_logic; attribute dont_touch of I642: signal is true;
	signal I650: std_logic; attribute dont_touch of I650: signal is true;
	signal I653: std_logic; attribute dont_touch of I653: signal is true;
	signal I656: std_logic; attribute dont_touch of I656: signal is true;
	signal I659: std_logic; attribute dont_touch of I659: signal is true;
	signal I662: std_logic; attribute dont_touch of I662: signal is true;
	signal I665: std_logic; attribute dont_touch of I665: signal is true;
	signal I668: std_logic; attribute dont_touch of I668: signal is true;
	signal I671: std_logic; attribute dont_touch of I671: signal is true;
	signal I674: std_logic; attribute dont_touch of I674: signal is true;
	signal I677: std_logic; attribute dont_touch of I677: signal is true;
	signal I680: std_logic; attribute dont_touch of I680: signal is true;
	signal I683: std_logic; attribute dont_touch of I683: signal is true;
	signal I686: std_logic; attribute dont_touch of I686: signal is true;
	signal I689: std_logic; attribute dont_touch of I689: signal is true;
	signal I692: std_logic; attribute dont_touch of I692: signal is true;
	signal I695: std_logic; attribute dont_touch of I695: signal is true;
	signal I698: std_logic; attribute dont_touch of I698: signal is true;
	signal I701: std_logic; attribute dont_touch of I701: signal is true;
	signal I704: std_logic; attribute dont_touch of I704: signal is true;
	signal I707: std_logic; attribute dont_touch of I707: signal is true;
	signal I710: std_logic; attribute dont_touch of I710: signal is true;
	signal I713: std_logic; attribute dont_touch of I713: signal is true;
	signal I716: std_logic; attribute dont_touch of I716: signal is true;
	signal I719: std_logic; attribute dont_touch of I719: signal is true;
	signal I722: std_logic; attribute dont_touch of I722: signal is true;
	signal II142: std_logic; attribute dont_touch of II142: signal is true;
	signal II254: std_logic; attribute dont_touch of II254: signal is true;
	signal II329: std_logic; attribute dont_touch of II329: signal is true;
	signal II368: std_logic; attribute dont_touch of II368: signal is true;
	signal II491: std_logic; attribute dont_touch of II491: signal is true;
	signal II497: std_logic; attribute dont_touch of II497: signal is true;
	signal V0E: std_logic; attribute dont_touch of V0E: signal is true;
	signal V1E: std_logic; attribute dont_touch of V1E: signal is true;
	signal V2E: std_logic; attribute dont_touch of V2E: signal is true;
	signal V3E: std_logic; attribute dont_touch of V3E: signal is true;
	signal V4E: std_logic; attribute dont_touch of V4E: signal is true;
	signal V5E: std_logic; attribute dont_touch of V5E: signal is true;
	signal V6E: std_logic; attribute dont_touch of V6E: signal is true;
	signal V7: std_logic; attribute dont_touch of V7: signal is true;
	signal V7E: std_logic; attribute dont_touch of V7E: signal is true;
	signal V8: std_logic; attribute dont_touch of V8: signal is true;
	signal V8E: std_logic; attribute dont_touch of V8E: signal is true;
	signal V9: std_logic; attribute dont_touch of V9: signal is true;
	signal V9E: std_logic; attribute dont_touch of V9E: signal is true;
	signal V10: std_logic; attribute dont_touch of V10: signal is true;
	signal V10E: std_logic; attribute dont_touch of V10E: signal is true;
	signal V11: std_logic; attribute dont_touch of V11: signal is true;
	signal V11E: std_logic; attribute dont_touch of V11E: signal is true;
	signal V12: std_logic; attribute dont_touch of V12: signal is true;
	signal V12E: std_logic; attribute dont_touch of V12E: signal is true;
	signal V13_D_0: std_logic; attribute dont_touch of V13_D_0: signal is true;
	signal V13_D_0C: std_logic; attribute dont_touch of V13_D_0C: signal is true;
	signal V13_D_1: std_logic; attribute dont_touch of V13_D_1: signal is true;
	signal V13_D_1C: std_logic; attribute dont_touch of V13_D_1C: signal is true;
	signal V13_D_2: std_logic; attribute dont_touch of V13_D_2: signal is true;
	signal V13_D_2C: std_logic; attribute dont_touch of V13_D_2C: signal is true;
	signal V13_D_3: std_logic; attribute dont_touch of V13_D_3: signal is true;
	signal V13_D_3C: std_logic; attribute dont_touch of V13_D_3C: signal is true;
	signal V13_D_4: std_logic; attribute dont_touch of V13_D_4: signal is true;
	signal V13_D_4C: std_logic; attribute dont_touch of V13_D_4C: signal is true;
	signal V13_D_5: std_logic; attribute dont_touch of V13_D_5: signal is true;
	signal V13_D_5C: std_logic; attribute dont_touch of V13_D_5C: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			V7<=V13_D_0C;
			V8<=V13_D_1C;
			V9<=V13_D_2C;
			V10<=V13_D_3C;
			V11<=V13_D_4C;
			V12<=V13_D_5C;
		end if;
	end process;
	C30DE<= not C30D;
	C49DE<= not C49D;
	C70DE<= not C70D;
	C81DE<= not C81D;
	C83DE<= not C83D;
	C90DE<= not C90D;
	C104DE<= not C104D;
	C108DE<= not C108D;
	C117DE<= not C117D;
	C118DE<= not C118D;
	C124DE<= not C124D;
	C129DE<= not C129D;
	C131DE<= not C131D;
	C138DE<= not C138D;
	C141DE<= not C141D;
	C144DE<= not C144D;
	C157DE<= not C157D;
	C165DE<= not C165D;
	C166DE<= not C166D;
	C180DE<= not C180D;
	C191DE<= not C191D;
	C194DE<= not C194D;
	C195DE<= not C195D;
	C208DE<= not C208D;
	C218DE<= not C218D;
	C220DE<= not C220D;
	I650<= not AV13_D_24B;
	I653<= not AV13_D_23B;
	I656<= not AV13_D_22B;
	I659<= not AV13_D_21B;
	I662<= not AV13_D_20B;
	I665<= not AV13_D_19B;
	I668<= not AV13_D_18B;
	I671<= not AV13_D_17B;
	I674<= not AV13_D_16B;
	I677<= not AV13_D_15B;
	I680<= not AV13_D_14B;
	I683<= not AV13_D_13B;
	I686<= not AV13_D_12B;
	I689<= not AV13_D_11B;
	I692<= not AV13_D_10B;
	I695<= not AV13_D_9B;
	I698<= not AV13_D_8B;
	I701<= not AV13_D_7B;
	I704<= not AV13_D_6B;
	I707<= not AV13_D_5B;
	I710<= not AV13_D_4B;
	I713<= not AV13_D_3B;
	I716<= not AV13_D_2B;
	I719<= not AV13_D_1B;
	I722<= not AV13_D_0B;
	V0E<= not V0;
	V1E<= not V1;
	V2E<= not V2;
	V3E<= not V3;
	V4E<= not V4;
	V5E<= not V5;
	V6E<= not V6;
	V7E<= not V7;
	V8E<= not V8;
	V9E<= not V9;
	V10E<= not V10;
	V11E<= not V11;
	V12E<= not V12;
	V13_D_0<= not I722;
	V13_D_1<= not I719;
	V13_D_2<= not I716;
	V13_D_3<= not I713;
	V13_D_4<= not I710;
	V13_D_5<= not I707;
	V13_D_6<= not I704;
	V13_D_7<= not I701;
	V13_D_8<= not I698;
	V13_D_9<= not I695;
	V13_D_10<= not I692;
	V13_D_11<= not I689;
	V13_D_12<= not I686;
	V13_D_13<= not I683;
	V13_D_14<= not I680;
	V13_D_15<= not I677;
	V13_D_16<= not I674;
	V13_D_17<= not I671;
	V13_D_18<= not I668;
	V13_D_19<= not I665;
	V13_D_20<= not I662;
	V13_D_21<= not I659;
	V13_D_22<= not I656;
	V13_D_23<= not I653;
	V13_D_24<= not I650;
	AV13_D_9B<=C153D and V12E;
	AV13_D_15B<=V7E and V12E and I548;
	AV13_D_16B<=C200D and V8 and V10;
	AV13_D_18B<=C210D and V7E and V12E;
	AV13_D_20B<=C138DE and C220DE and C104D and I329;
	AV13_D_21B<=C213D and V7E and V10E and V12E;
	AV13_D_23B<=C216D and V7E and V8E;
	I27<=C184D and V7;
	I28<=V7E and C188D;
	I29<=C190D and V10;
	I31<=C108DE and C83DE and I642;
	I32<=C207D and V2;
	I34<=C91D and C165DE;
	I35<=C79D and V7 and V9 and V12E;
	I36<=V7E and C89D;
	I38<=C102D and V7E;
	I39<=C103D and V10E;
	I40<=V2 and C92D;
	I41<=V7 and V12E and C96D;
	I43<=V8 and V10 and C108DE;
	I44<=V2E and C106D;
	I45<=C116D and V7E;
	I46<=V7 and C110D;
	I48<=C177D and V8E;
	I49<=V8 and C176D;
	I51<=C132D and V7;
	I52<=C135D and V7E;
	I54<=C186D and V9E;
	I55<=C187D and V12E;
	I58<=C75D and C129DE;
	I59<=V7 and C67D;
	I60<=V7E and C74D;
	I62<=V6E and C95D;
	I63<=V8 and C99D;
	I64<=V11E and C157DE;
	I65<=V9 and C185D;
	I66<=V8E and V12E and C100D;
	I68<=C206D and V12E;
	I69<=V7 and C202D;
	I71<=V2E and C28D;
	I72<=C38D and V7E;
	I73<=V7 and C31D and V8;
	I75<=C129DE and C144DE;
	I76<=V7E and C174D;
	I78<=V7E and C196D;
	I79<=V8 and C170D;
	I80<=V7 and V12E and C192D;
	I82<=V0E and C217D and C108DE;
	I83<=C225D and V11;
	I84<=V7E and C224D;
	I86<=C54D and C165DE;
	I87<=C53D and V7E;
	I88<=V2E and C43D;
	I89<=V7 and C48D;
	I91<=C148D and C131DE;
	I92<=V7 and C140D;
	I93<=V7E and C147D;
	I95<=C76D and C81DE;
	I96<=V8 and C85D;
	I97<=C88D and V11E;
	I98<=V8E and V12 and C87D;
	I100<=C134D and V9E;
	I101<=C127D and C128D and V12E;
	I103<=C115D and V10;
	I104<=V3 and C107D and V12;
	I105<=V8 and C113D;
	I106<=V8E and C114D;
	I108<=C181D and C83DE;
	I109<=C179D and V2 and V8 and V11;
	I111<=C98D and V10E;
	I112<=V11E and V12;
	I113<=V2E and V12E and C93D;
	I114<=V9 and C97D;
	I116<=C37D and V9;
	I117<=V8E and C35D;
	I119<=C126D and V8;
	I120<=V7E and C123D;
	I123<=V8 and C162D;
	I124<=C164D and V12E;
	I126<=V2 and C58D;
	I127<=C73D and V10E;
	I128<=V8 and C69D;
	I129<=V8E and C72D;
	I130<=C60D and C83D;
	I131<=V9 and V11E and C157DE;
	I133<=C152D and V9;
	I134<=V7E and V10 and C151D;
	I136<=C47D and C144DE;
	I137<=V8 and C46D;
	I140<=V8E and V10E and C144DE;
	I141<=C170D and V8;
	I142<=V7E and V9 and V11E;
	I145<=C49DE and C166DE and C220DE;
	I146<=C223D and V8E and V9E;
	I148<=V9 and V10E and C144DE;
	I149<=C112D and V10;
	I151<=V9 and C138DE;
	I152<=V8 and V12E and C129DE;
	I153<=C52D and V8E;
	I154<=V2 and C40D;
	I156<=C80D and V9;
	I157<=C82D and V9E;
	I158<=C84D and V10E;
	I160<=V8 and C65D;
	I161<=C144DE and C191D;
	I163<=V11E and V12E and C118DE;
	I164<=C133D and V8E;
	I166<=C205D and V10;
	I167<=V8 and V11 and C129D;
	I169<=C195D and V8E;
	I170<=V10 and V11E;
	I171<=V8 and C193D;
	I173<=C146D and V11E;
	I174<=V8E and C143D;
	I175<=V9 and C144D;
	I176<=V10E and C145D;
	I177<=C137D and C127D;
	I179<=V9 and V10 and C144DE;
	I180<=C173D and V9E;
	I182<=V8E and V10E and C144DE;
	I183<=C183D and V8;
	I185<=V8E and C195DE;
	I186<=V8 and V11 and C117DE;
	I188<=C175D and V11;
	I189<=V7 and V12E;
	I191<=V8 and V11 and C117DE;
	I192<=V8E and V9E and C44D;
	I194<=V3 and V12 and C77D;
	I196<=C161D and V11;
	I197<=C158D and V7 and V11E;
	I199<=V9E and C63D;
	I200<=V12E and C124D;
	I202<=V9E and C144DE and C83DE and C194DE;
	I203<=C34D and V9;
	I205<=V8E and C30DE;
	I206<=V7 and C150D;
	I208<=C122D and V11E;
	I209<=V8 and C119D;
	I210<=V9 and C120D;
	I212<=V9E and C49DE;
	I213<=C57D and V10E;
	I215<=V1 and V9 and C144DE;
	I216<=C189D and V9E;
	I218<=V12E and C44D and C83DE;
	I219<=C49D and V9;
	I220<=C51D and V12;
	I222<=C156D and C83DE;
	I223<=V7E and C160D and V9E;
	I224<=C163D and V8E and V11;
	I226<=V8E and V10E and C144DE;
	I227<=C139D and V8 and V10;
	I229<=V9 and V10 and C144DE;
	I230<=C109D and V10E;
	I232<=C165D and C83DE;
	I233<=C168D and V8E;
	I234<=V8 and C167D;
	I236<=V2E and V8 and C219D;
	I237<=V7 and V12E and C221D;
	I239<=V9 and V12 and C124DE;
	I240<=C125D and V9E;
	I242<=C130D and C165DE;
	I243<=C131D and V9 and C144DE;
	I245<=C185D and V8E;
	I247<=V10 and C144DE;
	I248<=C45D and V10E;
	I250<=C77D and V3 and C138DE;
	I251<=V6E and V11E and V12E;
	I253<=V1E and V10E and C138DE;
	I254<=V1 and V6 and V7E and V8E;
	I256<=V9 and V10 and C138DE;
	I257<=C215D and V9E;
	I259<=V12E and C129DE and C83DE;
	I260<=V3E and C78D;
	I262<=C42D and V8;
	I263<=V7E and V11 and C41D;
	I266<=V7 and C49DE and C220DE;
	I267<=C214D and V7E and V10E;
	I269<=V11E and C108DE and C83DE;
	I270<=V1E and C55D;
	I272<=V10E and C144DE;
	I273<=C201D and V8;
	I275<=V7 and V8 and C90DE;
	I276<=C27D and V7E and V9 and V12E;
	I278<=V10E and C138DE;
	I280<=V1E and C26D;
	I281<=V3E and C29D;
	I282<=C36D and V12;
	I284<=V11E and C157DE;
	I285<=C222D and V10E;
	I287<=V9 and V11;
	I288<=V7E and C203D;
	I291<=C142D and V11;
	I293<=C138DE and C118DE and I368;
	I294<=C211D and V3 and V7E and V11E;
	I296<=V8E and V9E and C124DE and C83DE;
	I297<=C209D and C208D and V11;
	I299<=V11E and C108DE;
	I300<=V0E and C105D;
	I302<=V11E and C157DE;
	I303<=C172D and V12E;
	I305<=V9 and C49DE;
	I306<=C129DE and C138D;
	I308<=C111D and C144DE;
	I310<=V6E and V9 and V12E and C124DE;
	I311<=C71D and V9E;
	I314<=V10 and C90DE;
	I315<=C155D and V12E and C129D;
	I317<=V10 and V11E;
	I318<=V11 and C118D;
	I320<=V11 and C141D;
	I321<=C33D and V11E and V12E;
	I323<=V10E and C127D;
	I325<=V10 and C90DE;
	I326<=C81DE and C129D;
	I328<=V3 and V12E and C124DE;
	I329<=V3 and V7E and V10;
	I332<=C138D and V9E;
	I333<=V11E and V12E;
	I335<=V12E and C218DE;
	I336<=C124D and V12;
	I338<=C108D and C165DE;
	I339<=V8E and C144DE;
	I341<=V11E and C118DE;
	I342<=C159D and V8E;
	I344<=C83D and V12E;
	I346<=V12 and C191DE;
	I347<=C90D and V10E;
	I349<=C118D and V11E;
	I350<=V11 and C117D;
	I352<=V8 and C124D;
	I354<=C191D and V11;
	I356<=C50D and V10E;
	I357<=V10 and V11E;
	I359<=V12E and C165DE;
	I360<=V3E and C59D;
	I362<=V8 and C138DE;
	I363<=V1E and C178D;
	I365<=C56D and V8 and V11;
	I366<=V8E and V9 and V11E and V12E;
	I368<=V7 and V8 and V9E;
	I369<=V9 and C124DE;
	I371<=V10E and C90DE;
	I372<=C129D and V12E;
	I374<=V9E and C30DE;
	I375<=C86D and V10E;
	I377<=V7 and V10 and C90DE;
	I378<=C218D and V5E and V9 and V12E;
	I380<=V2 and V11;
	I381<=C166D and V11E;
	I383<=C70D and C141DE;
	I384<=V10E and C138DE;
	I386<=V0 and C104D and V8 and C30DE;
	I387<=V8E and V9E and C124DE;
	I389<=V8 and V9 and V10;
	I390<=C220D and V10E;
	I392<=C81D and V11E;
	I393<=V10E and V12E;
	I395<=C157D and V9E;
	I396<=V10E and V12E;
	I398<=V12E and C118DE;
	I399<=V8 and C141D;
	I402<=V8 and V9E and C30DE;
	I403<=V9 and V12E and C124DE and I254;
	I405<=V8E and V9E and C194DE;
	I406<=V8 and V11 and C117DE;
	I409<=V9 and V11E;
	I412<=V3 and V10E and V12E;
	I414<=V6 and C138DE;
	I415<=V8E and V11E and V12E;
	I417<=V5E and V11E and V12E;
	I419<=V5E and V7E and V8E and C30DE;
	I420<=V2E and V7 and C131DE;
	I423<=V3E and C157DE;
	I425<=V8E and V10E;
	I427<=V8E and V9 and V10;
	I429<=V9E and C30DE;
	I430<=V1E and V9 and V10E;
	I432<=V7 and C90DE;
	I433<=V10 and C144DE;
	I435<=V12 and C165DE;
	I436<=V8E and V9 and C144DE;
	I438<=V0 and V10 and C144DE;
	I439<=V6 and V12 and C124DE;
	I441<=V11 and C220DE;
	I442<=V7E and V8E and V9E;
	I444<=V3E and V9E;
	I446<=V11E and C90DE;
	I447<=V8E and V9 and V10E and V12E;
	I449<=C108DE and C83DE;
	I450<=V3 and V8 and C138DE and C104DE;
	I452<=V12E and C220DE;
	I453<=V8E and V10E and V12;
	I456<=V9 and C30DE;
	I457<=V6 and C124DE and C90DE;
	I460<=V2E and V12E and C165DE;
	I461<=V8E and V9 and V12;
	I463<=C165DE and C191DE;
	I464<=V8E and V10E and V11;
	I466<=V8E and V11E and V12E;
	I468<=V9 and C83DE;
	I470<=V8 and V12E and C83DE;
	I471<=V1 and V10E and V12;
	I473<=V0E and C30DE;
	I475<=V2E and V8 and C138DE;
	I476<=V8E and V9 and V11E and V12E;
	I478<=V10E and C83DE;
	I479<=V0 and V11;
	I482<=V2 and C220DE;
	I483<=V8E and V9E and V11E and C83DE;
	I485<=V6 and C141DE and C220DE;
	I486<=V6E and V8E and V12 and C129DE;
	I489<=V8E and V11;
	I492<=V10 and V11E;
	I494<=V8E and V10 and C108DE;
	I495<=V9 and V11 and C131DE;
	I498<=V8 and C117DE;
	I500<=V8 and V11 and C83DE;
	I501<=V8E and V11E;
	I503<=V9E and C30DE;
	I505<=V7 and V8 and C138DE and C191DE;
	I506<=V7E and V9 and V10E and V12E;
	I508<=V9E and V11E;
	I510<=V9 and V10;
	I513<=V12E and C166DE and I142;
	I514<=V2 and V7 and V9E and C138DE;
	I516<=V1 and V12;
	I518<=V9 and V10E;
	I520<=V3E and V6E;
	I524<=V6 and V11E;
	I528<=V9E and V11;
	I533<=V9 and V10;
	I534<=V8E and V10E;
	I537<=V6E and V7E and V8E and V12;
	I538<=V8 and V12E;
	I546<=V0 and V11;
	I547<=V10 and V11E;
	I548<=C199D and V4 and V5E;
	I554<=V2E and V8 and V9E;
	I555<=V0 and V8E and V11;
	I559<=V8 and V11;
	I560<=V7E and V12E;
	I642<=V7E and V8E and C124DE;
	II142<=V7E and C169D;
	II254<=C39D and V8E;
	II329<=V9 and V12 and C30D;
	II368<=C30D and C90DE;
	II491<=V10E and C138DE;
	II497<=V8E and V9E and C194DE;
	V13_D_0C<=V13_D_0 and CLR;
	V13_D_1C<=V13_D_1 and CLR;
	V13_D_2C<=V13_D_2 and CLR;
	V13_D_3C<=V13_D_3 and CLR;
	V13_D_4C<=V13_D_4 and CLR;
	V13_D_5C<=V13_D_5 and CLR;
	AV13_D_0B<=I71 or I72 or I73;
	AV13_D_1B<=I86 or I87 or I88 or I89;
	AV13_D_2B<=I58 or I59 or I60;
	AV13_D_3B<=I34 or I35 or I36;
	AV13_D_4B<=I38 or I39 or I40 or I41;
	AV13_D_5B<=I43 or I44 or I45 or I46;
	AV13_D_6B<=I119 or I120;
	AV13_D_7B<=I51 or I52;
	AV13_D_8B<=I91 or I92 or I93;
	AV13_D_10B<=I123 or I124;
	AV13_D_11B<=I140 or I141 or II142;
	AV13_D_12B<=I48 or I49;
	AV13_D_13B<=I27 or I28 or I29;
	AV13_D_14B<=I78 or I79 or I80;
	AV13_D_17B<=I31 or I32;
	AV13_D_19B<=I293 or I294;
	AV13_D_22B<=I266 or I267;
	AV13_D_24B<=I82 or I83 or I84;
	C26D<=I414 or I415;
	C27D<=I500 or I501;
	C28D<=I275 or I276;
	C29D<=C138DE or I466;
	C30D<=V10E or V11E;
	C31D<=II368 or I369;
	C33D<=V6E or V10;
	C34D<=I320 or I321;
	C35D<=I202 or I203;
	C36D<=C165DE or V10E;
	C37D<=I280 or I281 or I282;
	C38D<=I116 or I117;
	C39D<=I423 or V9;
	C40D<=I253 or II254;
	C41D<=I470 or I471;
	C42D<=I432 or I433;
	C43D<=I262 or I263;
	C44D<=I473 or C124DE;
	C45D<=C90DE or V11E;
	C46D<=I247 or I248;
	C47D<=I533 or I534;
	C48D<=I136 or I137;
	C49D<=C141D or V11;
	C50D<=I520 or V11;
	C51D<=I356 or I357;
	C52D<=I218 or I219 or I220;
	C53D<=I151 or I152 or I153 or I154;
	C54D<=C90DE or I412;
	C55D<=I475 or I476;
	C56D<=V9 or I516;
	C57D<=I365 or I366;
	C58D<=I212 or I213;
	C59D<=I537 or I538;
	C60D<=I494 or I495;
	C63D<=V12E or I317 or I318;
	C65D<=I199 or I200;
	C67D<=I160 or I161;
	C69D<=I328 or II329;
	C70D<=V0 or V11E;
	C71D<=I383 or I384;
	C72D<=I310 or I311;
	C73D<=I269 or I270;
	C74D<=I129 or I130 or I131 or I542;
	C75D<=I359 or I360;
	C76D<=C131DE or I427;
	C77D<=C104D or V0E;
	C78D<=I452 or I453;
	C79D<=C131DE or V11;
	C80D<=I250 or I251;
	C81D<=V2E or V12;
	C82D<=I392 or I393;
	C83D<=V4E or V5E;
	C84D<=C138DE or I344;
	C85D<=I156 or I157 or I158;
	C86D<=V9 or I524;
	C87D<=I374 or I375;
	C88D<=I259 or I260;
	C89D<=I95 or I96 or I97 or I98;
	C90D<=V9 or V12E;
	C91D<=I346 or I347;
	C92D<=I505 or I506;
	C93D<=C191DE or I468;
	C95D<=I446 or I447;
	C96D<=I463 or I464;
	C97D<=V11E or I194;
	C98D<=C144D or I444;
	C99D<=I111 or I112 or I113 or I114;
	C100D<=I429 or I430;
	C102D<=I65 or I66 or I610;
	C103D<=I435 or I436;
	C104D<=V1 or V6E;
	C105D<=I449 or I450;
	C106D<=I402 or I403;
	C107D<=I386 or I387;
	C108D<=V9 or V12;
	C109D<=I338 or I339;
	C110D<=I229 or I230;
	C111D<=C83DE or V2;
	C112D<=I308 or V9E;
	C113D<=I148 or I149;
	C114D<=I456 or I457;
	C115D<=I299 or I300;
	C116D<=I103 or I104 or I105 or I106;
	C117D<=V9E or V2;
	C118D<=V2E or V10E;
	C119D<=I349 or V12 or I350;
	C120D<=C144D or I425;
	C122D<=V12 or I323;
	C123D<=C157DE or I208 or I209 or I210;
	C124D<=V10 or V11;
	C125D<=I335 or I336;
	C126D<=I239 or I240;
	C127D<=V5E or V4;
	C128D<=I405 or I406;
	C129D<=V9 or V10;
	C130D<=I371 or I372;
	C131D<=V8E or V10;
	C132D<=I242 or I243;
	C133D<=C49DE or I278;
	C134D<=I163 or I164;
	C135D<=I100 or I101;
	C137D<=C117DE or I489;
	C138D<=V11E or V12E;
	C139D<=I332 or I333;
	C140D<=I226 or I227;
	C141D<=V10E or V12;
	C142D<=V0 or V12;
	C143D<=C49DE or V9 or I291;
	C144D<=V11E or V12;
	C145D<=I528 or V12;
	C146D<=I398 or I399;
	C147D<=I176 or I177 or I491;
	C148D<=C90DE or I409;
	C150D<=C30DE or I352;
	C151D<=I554 or I555;
	C152D<=I205 or I206;
	C153D<=I133 or I134;
	C155D<=V2 or V7;
	C156D<=I441 or I442;
	C157D<=V10E or V12E;
	C158D<=I395 or I396;
	C159D<=I546 or I547;
	C160D<=I341 or I342;
	C161D<=I314 or I315;
	C162D<=I196 or I197;
	C163D<=C129DE or I510;
	C164D<=I222 or I223 or I224;
	C165D<=V8E or V11;
	C166D<=V3E or V6E;
	C167D<=I380 or I381;
	C168D<=C159D or V9;
	C169D<=I232 or I233 or V12 or I234;
	C170D<=C124DE or V9E;
	C172D<=I478 or I479;
	C173D<=I302 or I303;
	C174D<=I179 or I180;
	C175D<=I325 or I326;
	C176D<=I188 or I189;
	C177D<=I75 or I76;
	C178D<=I559 or I560;
	C179D<=V10 or I518;
	C180D<=C194DE or V11E;
	C181D<=I185 or I186;
	C183D<=I305 or I306;
	C184D<=I182 or I183;
	C185D<=II491 or I492;
	C186D<=C49DE or I245;
	C187D<=I108 or I109;
	C188D<=I54 or I55;
	C189D<=I362 or I363;
	C190D<=I215 or I216;
	C191D<=V10E or V9;
	C192D<=V8 or I354;
	C193D<=V2 or V11E;
	C194D<=V0 or V10E;
	C195D<=C180DE or V9;
	C196D<=I170 or V12 or I171 or I497;
	C199D<=I191 or I192;
	C200D<=I513 or I514;
	C201D<=I503 or V12E;
	C202D<=I272 or I273;
	C203D<=C70DE or I508;
	C205D<=I287 or I288;
	C206D<=I166 or I167;
	C207D<=I68 or I69;
	C208D<=V5 or V4;
	C209D<=II497 or I498;
	C210D<=I296 or I297;
	C211D<=I485 or I486;
	C213D<=I482 or I483;
	C214D<=I460 or I461;
	C215D<=I438 or I439;
	C216D<=I256 or I257;
	C217D<=I419 or I420;
	C218D<=V7E or V10;
	C219D<=I377 or I378;
	C220D<=V8E or V9E;
	C221D<=I389 or I390;
	C222D<=C138DE or I417;
	C223D<=I284 or I285;
	C224D<=I145 or I146;
	C225D<=I236 or I237;
	I491<=I173 or I174 or I175;
	I497<=C208DE or C83DE or I169;
	I542<=I126 or I127 or I128;
	I610<=I62 or I63 or I64;
end RTL;
