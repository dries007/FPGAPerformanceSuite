-- File created by Bench2VHDL
-- Name: s38584
-- File: bench/s38584.bench
-- Timestamp: 2019-05-21T22:08:28.667278
--
-- Original File
-- =============
--	# s38584.1
--	# 38 inputs
--	# 304 outputs
--	# 1426 D-type flipflops
--	# 7805 inverters
--	# 11448 gates (5516 ANDs + 2126 NANDs + 2621 ORs + 1185 NORs)
--	
--	INPUT(g35)
--	INPUT(g36)
--	INPUT(g6744)
--	INPUT(g6745)
--	INPUT(g6746)
--	INPUT(g6747)
--	INPUT(g6748)
--	INPUT(g6749)
--	INPUT(g6750)
--	INPUT(g6751)
--	INPUT(g6752)
--	INPUT(g6753)
--	INPUT(g84)
--	INPUT(g120)
--	INPUT(g5)
--	INPUT(g113)
--	INPUT(g126)
--	INPUT(g99)
--	INPUT(g53)
--	INPUT(g116)
--	INPUT(g92)
--	INPUT(g56)
--	INPUT(g91)
--	INPUT(g44)
--	INPUT(g57)
--	INPUT(g100)
--	INPUT(g54)
--	INPUT(g124)
--	INPUT(g125)
--	INPUT(g114)
--	INPUT(g134)
--	INPUT(g72)
--	INPUT(g115)
--	INPUT(g135)
--	INPUT(g90)
--	INPUT(g127)
--	INPUT(g64)
--	INPUT(g73)
--	
--	OUTPUT(g7243)
--	OUTPUT(g7245)
--	OUTPUT(g7257)
--	OUTPUT(g7260)
--	OUTPUT(g7540)
--	OUTPUT(g7916)
--	OUTPUT(g7946)
--	OUTPUT(g8132)
--	OUTPUT(g8178)
--	OUTPUT(g8215)
--	OUTPUT(g8235)
--	OUTPUT(g8277)
--	OUTPUT(g8279)
--	OUTPUT(g8283)
--	OUTPUT(g8291)
--	OUTPUT(g8342)
--	OUTPUT(g8344)
--	OUTPUT(g8353)
--	OUTPUT(g8358)
--	OUTPUT(g8398)
--	OUTPUT(g8403)
--	OUTPUT(g8416)
--	OUTPUT(g8475)
--	OUTPUT(g8719)
--	OUTPUT(g8783)
--	OUTPUT(g8784)
--	OUTPUT(g8785)
--	OUTPUT(g8786)
--	OUTPUT(g8787)
--	OUTPUT(g8788)
--	OUTPUT(g8789)
--	OUTPUT(g8839)
--	OUTPUT(g8870)
--	OUTPUT(g8915)
--	OUTPUT(g8916)
--	OUTPUT(g8917)
--	OUTPUT(g8918)
--	OUTPUT(g8919)
--	OUTPUT(g8920)
--	OUTPUT(g9019)
--	OUTPUT(g9048)
--	OUTPUT(g9251)
--	OUTPUT(g9497)
--	OUTPUT(g9553)
--	OUTPUT(g9555)
--	OUTPUT(g9615)
--	OUTPUT(g9617)
--	OUTPUT(g9680)
--	OUTPUT(g9682)
--	OUTPUT(g9741)
--	OUTPUT(g9743)
--	OUTPUT(g9817)
--	OUTPUT(g10122)
--	OUTPUT(g10306)
--	OUTPUT(g10500)
--	OUTPUT(g10527)
--	OUTPUT(g11349)
--	OUTPUT(g11388)
--	OUTPUT(g11418)
--	OUTPUT(g11447)
--	OUTPUT(g11678)
--	OUTPUT(g11770)
--	OUTPUT(g12184)
--	OUTPUT(g12238)
--	OUTPUT(g12300)
--	OUTPUT(g12350)
--	OUTPUT(g12368)
--	OUTPUT(g12422)
--	OUTPUT(g12470)
--	OUTPUT(g12832)
--	OUTPUT(g12919)
--	OUTPUT(g12923)
--	OUTPUT(g13039)
--	OUTPUT(g13049)
--	OUTPUT(g13068)
--	OUTPUT(g13085)
--	OUTPUT(g13099)
--	OUTPUT(g13259)
--	OUTPUT(g13272)
--	OUTPUT(g13865)
--	OUTPUT(g13881)
--	OUTPUT(g13895)
--	OUTPUT(g13906)
--	OUTPUT(g13926)
--	OUTPUT(g13966)
--	OUTPUT(g14096)
--	OUTPUT(g14125)
--	OUTPUT(g14147)
--	OUTPUT(g14167)
--	OUTPUT(g14189)
--	OUTPUT(g14201)
--	OUTPUT(g14217)
--	OUTPUT(g14421)
--	OUTPUT(g14451)
--	OUTPUT(g14518)
--	OUTPUT(g14597)
--	OUTPUT(g14635)
--	OUTPUT(g14662)
--	OUTPUT(g14673)
--	OUTPUT(g14694)
--	OUTPUT(g14705)
--	OUTPUT(g14738)
--	OUTPUT(g14749)
--	OUTPUT(g14779)
--	OUTPUT(g14828)
--	OUTPUT(g16603)
--	OUTPUT(g16624)
--	OUTPUT(g16627)
--	OUTPUT(g16656)
--	OUTPUT(g16659)
--	OUTPUT(g16686)
--	OUTPUT(g16693)
--	OUTPUT(g16718)
--	OUTPUT(g16722)
--	OUTPUT(g16744)
--	OUTPUT(g16748)
--	OUTPUT(g16775)
--	OUTPUT(g16874)
--	OUTPUT(g16924)
--	OUTPUT(g16955)
--	OUTPUT(g17291)
--	OUTPUT(g17316)
--	OUTPUT(g17320)
--	OUTPUT(g17400)
--	OUTPUT(g17404)
--	OUTPUT(g17423)
--	OUTPUT(g17519)
--	OUTPUT(g17577)
--	OUTPUT(g17580)
--	OUTPUT(g17604)
--	OUTPUT(g17607)
--	OUTPUT(g17639)
--	OUTPUT(g17646)
--	OUTPUT(g17649)
--	OUTPUT(g17674)
--	OUTPUT(g17678)
--	OUTPUT(g17685)
--	OUTPUT(g17688)
--	OUTPUT(g17711)
--	OUTPUT(g17715)
--	OUTPUT(g17722)
--	OUTPUT(g17739)
--	OUTPUT(g17743)
--	OUTPUT(g17760)
--	OUTPUT(g17764)
--	OUTPUT(g17778)
--	OUTPUT(g17787)
--	OUTPUT(g17813)
--	OUTPUT(g17819)
--	OUTPUT(g17845)
--	OUTPUT(g17871)
--	OUTPUT(g18092)
--	OUTPUT(g18094)
--	OUTPUT(g18095)
--	OUTPUT(g18096)
--	OUTPUT(g18097)
--	OUTPUT(g18098)
--	OUTPUT(g18099)
--	OUTPUT(g18100)
--	OUTPUT(g18101)
--	OUTPUT(g18881)
--	OUTPUT(g19334)
--	OUTPUT(g19357)
--	OUTPUT(g20049)
--	OUTPUT(g20557)
--	OUTPUT(g20652)
--	OUTPUT(g20654)
--	OUTPUT(g20763)
--	OUTPUT(g20899)
--	OUTPUT(g20901)
--	OUTPUT(g21176)
--	OUTPUT(g21245)
--	OUTPUT(g21270)
--	OUTPUT(g21292)
--	OUTPUT(g21698)
--	OUTPUT(g21727)
--	OUTPUT(g23002)
--	OUTPUT(g23190)
--	OUTPUT(g23612)
--	OUTPUT(g23652)
--	OUTPUT(g23683)
--	OUTPUT(g23759)
--	OUTPUT(g24151)
--	OUTPUT(g25114)
--	OUTPUT(g25167)
--	OUTPUT(g25219)
--	OUTPUT(g25259)
--	OUTPUT(g25582)
--	OUTPUT(g25583)
--	OUTPUT(g25584)
--	OUTPUT(g25585)
--	OUTPUT(g25586)
--	OUTPUT(g25587)
--	OUTPUT(g25588)
--	OUTPUT(g25589)
--	OUTPUT(g25590)
--	OUTPUT(g26801)
--	OUTPUT(g26875)
--	OUTPUT(g26876)
--	OUTPUT(g26877)
--	OUTPUT(g27831)
--	OUTPUT(g28030)
--	OUTPUT(g28041)
--	OUTPUT(g28042)
--	OUTPUT(g28753)
--	OUTPUT(g29210)
--	OUTPUT(g29211)
--	OUTPUT(g29212)
--	OUTPUT(g29213)
--	OUTPUT(g29214)
--	OUTPUT(g29215)
--	OUTPUT(g29216)
--	OUTPUT(g29217)
--	OUTPUT(g29218)
--	OUTPUT(g29219)
--	OUTPUT(g29220)
--	OUTPUT(g29221)
--	OUTPUT(g30327)
--	OUTPUT(g30329)
--	OUTPUT(g30330)
--	OUTPUT(g30331)
--	OUTPUT(g30332)
--	OUTPUT(g31521)
--	OUTPUT(g31656)
--	OUTPUT(g31665)
--	OUTPUT(g31793)
--	OUTPUT(g31860)
--	OUTPUT(g31861)
--	OUTPUT(g31862)
--	OUTPUT(g31863)
--	OUTPUT(g32185)
--	OUTPUT(g32429)
--	OUTPUT(g32454)
--	OUTPUT(g32975)
--	OUTPUT(g33079)
--	OUTPUT(g33435)
--	OUTPUT(g33533)
--	OUTPUT(g33636)
--	OUTPUT(g33659)
--	OUTPUT(g33874)
--	OUTPUT(g33894)
--	OUTPUT(g33935)
--	OUTPUT(g33945)
--	OUTPUT(g33946)
--	OUTPUT(g33947)
--	OUTPUT(g33948)
--	OUTPUT(g33949)
--	OUTPUT(g33950)
--	OUTPUT(g33959)
--	OUTPUT(g34201)
--	OUTPUT(g34221)
--	OUTPUT(g34232)
--	OUTPUT(g34233)
--	OUTPUT(g34234)
--	OUTPUT(g34235)
--	OUTPUT(g34236)
--	OUTPUT(g34237)
--	OUTPUT(g34238)
--	OUTPUT(g34239)
--	OUTPUT(g34240)
--	OUTPUT(g34383)
--	OUTPUT(g34425)
--	OUTPUT(g34435)
--	OUTPUT(g34436)
--	OUTPUT(g34437)
--	OUTPUT(g34597)
--	OUTPUT(g34788)
--	OUTPUT(g34839)
--	OUTPUT(g34913)
--	OUTPUT(g34915)
--	OUTPUT(g34917)
--	OUTPUT(g34919)
--	OUTPUT(g34921)
--	OUTPUT(g34923)
--	OUTPUT(g34925)
--	OUTPUT(g34927)
--	OUTPUT(g34956)
--	OUTPUT(g34972)
--	OUTPUT(g24168)
--	OUTPUT(g24178)
--	OUTPUT(g12833)
--	OUTPUT(g24174)
--	OUTPUT(g24181)
--	OUTPUT(g24172)
--	OUTPUT(g24161)
--	OUTPUT(g24177)
--	OUTPUT(g24171)
--	OUTPUT(g24163)
--	OUTPUT(g24170)
--	OUTPUT(g24185)
--	OUTPUT(g24164)
--	OUTPUT(g24173)
--	OUTPUT(g24162)
--	OUTPUT(g24179)
--	OUTPUT(g24180)
--	OUTPUT(g24175)
--	OUTPUT(g24183)
--	OUTPUT(g24166)
--	OUTPUT(g24176)
--	OUTPUT(g24184)
--	OUTPUT(g24169)
--	OUTPUT(g24182)
--	OUTPUT(g24165)
--	OUTPUT(g24167)
--	
--	g5057 = DFF(g33046)
--	g2771 = DFF(g34441)
--	g1882 = DFF(g33982)
--	g6462 = DFF(g25751)
--	g2299 = DFF(g34007)
--	g4040 = DFF(g24276)
--	g2547 = DFF(g30381)
--	g559 = DFF(g640)
--	g3017 = DFF(g31877)
--	g3243 = DFF(g30405)
--	g452 = DFF(g25604)
--	g464 = DFF(g25607)
--	g3542 = DFF(g30416)
--	g5232 = DFF(g30466)
--	g5813 = DFF(g25736)
--	g2907 = DFF(g34617)
--	g1744 = DFF(g33974)
--	g5909 = DFF(g30505)
--	g1802 = DFF(g33554)
--	g3554 = DFF(g30432)
--	g6219 = DFF(g33064)
--	g807 = DFF(g34881)
--	g6031 = DFF(g6027)
--	g847 = DFF(g24216)
--	g976 = DFF(g24232)
--	g4172 = DFF(g34733)
--	g4372 = DFF(g34882)
--	g3512 = DFF(g33026)
--	g749 = DFF(g31867)
--	g3490 = DFF(g25668)
--	g6005 = DFF(g24344)
--	g4235 = DFF(g4232)
--	g1600 = DFF(g33966)
--	g1714 = DFF(g33550)
--	g3649 = DFF(g3625)
--	g3155 = DFF(g30393)
--	g3355 = DFF(g31880)
--	g2236 = DFF(g29248)
--	g4555 = DFF(g4571)
--	g3698 = DFF(g24274)
--	g6073 = DFF(g31920)
--	g1736 = DFF(g33973)
--	g1968 = DFF(g30360)
--	g4621 = DFF(g34460)
--	g5607 = DFF(g30494)
--	g2657 = DFF(g30384)
--	g5659 = DFF(g24340)
--	g490 = DFF(g29223)
--	g311 = DFF(g26881)
--	g6069 = DFF(g31925)
--	g772 = DFF(g34252)
--	g5587 = DFF(g30489)
--	g6177 = DFF(g29301)
--	g6377 = DFF(g6373)
--	g3167 = DFF(g33022)
--	g5615 = DFF(g30496)
--	g4567 = DFF(g33043)
--	g3057 = DFF(g28062)
--	g3457 = DFF(g29263)
--	g6287 = DFF(g30533)
--	g1500 = DFF(g24256)
--	g2563 = DFF(g34015)
--	g4776 = DFF(g34031)
--	g4593 = DFF(g34452)
--	g6199 = DFF(g34646)
--	g2295 = DFF(g34001)
--	g1384 = DFF(g25633)
--	g1339 = DFF(g24259)
--	g5180 = DFF(g33049)
--	g2844 = DFF(g34609)
--	g1024 = DFF(g31869)
--	g5591 = DFF(g30490)
--	g3598 = DFF(g30427)
--	g4264 = DFF(g21894)
--	g767 = DFF(g33965)
--	g5853 = DFF(g34645)
--	g3321 = DFF(g3317)
--	g2089 = DFF(g33571)
--	g4933 = DFF(g34267)
--	g4521 = DFF(g26971)
--	g5507 = DFF(g34644)
--	g3625 = DFF(g3618)
--	g6291 = DFF(g30534)
--	g294 = DFF(g33535)
--	g5559 = DFF(g30498)
--	g5794 = DFF(g25728)
--	g6144 = DFF(g25743)
--	g3813 = DFF(g25684)
--	g562 = DFF(g25613)
--	g608 = DFF(g34438)
--	g1205 = DFF(g24244)
--	g3909 = DFF(g30439)
--	g6259 = DFF(g30541)
--	g5905 = DFF(g30519)
--	g921 = DFF(g25621)
--	g2955 = DFF(g34807)
--	g203 = DFF(g25599)
--	g6088 = DFF(g31924)
--	g1099 = DFF(g24235)
--	g4878 = DFF(g34036)
--	g5204 = DFF(g30476)
--	g5630 = DFF(g5623)
--	g3606 = DFF(g30429)
--	g1926 = DFF(g32997)
--	g6215 = DFF(g33063)
--	g3586 = DFF(g30424)
--	g291 = DFF(g32977)
--	g4674 = DFF(g34026)
--	g3570 = DFF(g30420)
--	g640 = DFF(g637)
--	g5969 = DFF(g6012)
--	g1862 = DFF(g33560)
--	g676 = DFF(g29226)
--	g843 = DFF(g25619)
--	g4132 = DFF(g28076)
--	g4332 = DFF(g34455)
--	g4153 = DFF(g30457)
--	g5666 = DFF(g5637)
--	g6336 = DFF(g33625)
--	g622 = DFF(g34790)
--	g3506 = DFF(g30414)
--	g4558 = DFF(g26966)
--	g6065 = DFF(g31923)
--	g6322 = DFF(g6315)
--	g3111 = DFF(g25656)
--	g117 = DFF(g30390)
--	g2837 = DFF(g26935)
--	g939 = DFF(g34727)
--	g278 = DFF(g25594)
--	g4492 = DFF(g26963)
--	g4864 = DFF(g34034)
--	g1036 = DFF(g33541)
--	g128 = DFF(g28093)
--	g1178 = DFF(g24236)
--	g3239 = DFF(g30404)
--	g718 = DFF(g28051)
--	g6195 = DFF(g29303)
--	g1135 = DFF(g26917)
--	g6137 = DFF(g25741)
--	g6395 = DFF(g33624)
--	g3380 = DFF(g31882)
--	g5343 = DFF(g24337)
--	g554 = DFF(g34911)
--	g496 = DFF(g33963)
--	g3853 = DFF(g34627)
--	g5134 = DFF(g29282)
--	g1422 = DFF(g1418)
--	g3794 = DFF(g25676)
--	g2485 = DFF(g33013)
--	g925 = DFF(g32981)
--	g48 = DFF(g34993)
--	g5555 = DFF(g30483)
--	g878 = DFF(g875)
--	g1798 = DFF(g32994)
--	g4076 = DFF(g28070)
--	g2941 = DFF(g34806)
--	g3905 = DFF(g30453)
--	g763 = DFF(g33539)
--	g6255 = DFF(g30526)
--	g4375 = DFF(g26951)
--	g4871 = DFF(g34035)
--	g4722 = DFF(g34636)
--	g590 = DFF(g32978)
--	g6692 = DFF(g6668)
--	g1632 = DFF(g30348)
--	g5313 = DFF(g24336)
--	g3100 = DFF(g3092)
--	g1495 = DFF(g24250)
--	g6497 = DFF(g6490)
--	g1437 = DFF(g29236)
--	g6154 = DFF(g29298)
--	g1579 = DFF(g1576)
--	g5567 = DFF(g30499)
--	g1752 = DFF(g33976)
--	g1917 = DFF(g32996)
--	g744 = DFF(g30335)
--	g3040 = DFF(g31878)
--	g4737 = DFF(g34637)
--	g4809 = DFF(g25693)
--	g6267 = DFF(g30528)
--	g3440 = DFF(g25661)
--	g3969 = DFF(g4012)
--	g1442 = DFF(g24251)
--	g5965 = DFF(g30521)
--	g4477 = DFF(g26960)
--	g1233 = DFF(g24239)
--	g4643 = DFF(g34259)
--	g5264 = DFF(g30474)
--	g6329 = DFF(g6351)
--	g2610 = DFF(g33016)
--	g5160 = DFF(g34643)
--	g5360 = DFF(g31905)
--	g5933 = DFF(g30510)
--	g1454 = DFF(g29239)
--	g753 = DFF(g26897)
--	g1296 = DFF(g34729)
--	g3151 = DFF(g34625)
--	g2980 = DFF(g34800)
--	g6727 = DFF(g24353)
--	g3530 = DFF(g33029)
--	g4742 = DFF(g21903)
--	g4104 = DFF(g33615)
--	g1532 = DFF(g24253)
--	g4304 = DFF(g24281)
--	g2177 = DFF(g33997)
--	g3010 = DFF(g25651)
--	g52 = DFF(g34997)
--	g4754 = DFF(g34263)
--	g1189 = DFF(g24237)
--	g2287 = DFF(g33584)
--	g4273 = DFF(g24280)
--	g1389 = DFF(g26920)
--	g1706 = DFF(g33548)
--	g5835 = DFF(g29296)
--	g1171 = DFF(g30338)
--	g4269 = DFF(g21895)
--	g2399 = DFF(g33588)
--	g3372 = DFF(g31886)
--	g4983 = DFF(g34041)
--	g5611 = DFF(g30495)
--	g3618 = DFF(g3661)
--	g4572 = DFF(g29279)
--	g3143 = DFF(g25655)
--	g2898 = DFF(g34795)
--	g3343 = DFF(g24269)
--	g3235 = DFF(g30403)
--	g4543 = DFF(g33042)
--	g3566 = DFF(g30419)
--	g4534 = DFF(g34023)
--	g4961 = DFF(g28090)
--	g6398 = DFF(g31926)
--	g4927 = DFF(g34642)
--	g2259 = DFF(g30370)
--	g2819 = DFF(g34448)
--	g4414 = DFF(g26946)
--	g5802 = DFF(g5794)
--	g2852 = DFF(g34610)
--	g417 = DFF(g24209)
--	g681 = DFF(g28047)
--	g437 = DFF(g24206)
--	g351 = DFF(g26891)
--	g5901 = DFF(g30504)
--	g2886 = DFF(g34798)
--	g3494 = DFF(g25669)
--	g5511 = DFF(g30480)
--	g3518 = DFF(g33027)
--	g1604 = DFF(g33972)
--	g4135 = DFF(g28077)
--	g5092 = DFF(g25697)
--	g4831 = DFF(g28099)
--	g4382 = DFF(g26947)
--	g6386 = DFF(g24350)
--	g479 = DFF(g24210)
--	g3965 = DFF(g30455)
--	g4749 = DFF(g28084)
--	g2008 = DFF(g33993)
--	g736 = DFF(g802)
--	g3933 = DFF(g30444)
--	g222 = DFF(g33537)
--	g3050 = DFF(g25650)
--	g5736 = DFF(g31915)
--	g1052 = DFF(g25625)
--	g58 = DFF(g30328)
--	g5623 = DFF(g5666)
--	g2122 = DFF(g30366)
--	g2465 = DFF(g33593)
--	g6483 = DFF(g25755)
--	g5889 = DFF(g30502)
--	g4495 = DFF(g33036)
--	g365 = DFF(g25595)
--	g4653 = DFF(g34462)
--	g3179 = DFF(g33024)
--	g1728 = DFF(g33552)
--	g2433 = DFF(g34014)
--	g3835 = DFF(g29273)
--	g6187 = DFF(g25748)
--	g4917 = DFF(g34638)
--	g1070 = DFF(g30341)
--	g822 = DFF(g26899)
--	g6027 = DFF(g6023)
--	g914 = DFF(g30336)
--	g5339 = DFF(g5335)
--	g4164 = DFF(g26940)
--	g969 = DFF(g25622)
--	g2807 = DFF(g34447)
--	g5424 = DFF(g25709)
--	g4054 = DFF(g33613)
--	g6191 = DFF(g25749)
--	g5077 = DFF(g25704)
--	g5523 = DFF(g33053)
--	g3680 = DFF(g3676)
--	g6637 = DFF(g30555)
--	g174 = DFF(g25601)
--	g1682 = DFF(g33971)
--	g355 = DFF(g26892)
--	g1087 = DFF(g1083)
--	g1105 = DFF(g26915)
--	g2342 = DFF(g33008)
--	g6307 = DFF(g30538)
--	g3802 = DFF(g3794)
--	g6159 = DFF(g25750)
--	g2255 = DFF(g30369)
--	g2815 = DFF(g34446)
--	g911 = DFF(g29230)
--	g43 = DFF(g34789)
--	g4012 = DFF(g3983)
--	g1748 = DFF(g33975)
--	g5551 = DFF(g30497)
--	g5742 = DFF(g31917)
--	g3558 = DFF(g30418)
--	g5499 = DFF(g25721)
--	g2960 = DFF(g34622)
--	g3901 = DFF(g30438)
--	g4888 = DFF(g34266)
--	g6251 = DFF(g30540)
--	g6315 = DFF(g6358)
--	g1373 = DFF(g32986)
--	g3092 = DFF(g25648)
--	g157 = DFF(g33960)
--	g2783 = DFF(g34442)
--	g4281 = DFF(g4277)
--	g3574 = DFF(g30421)
--	g2112 = DFF(g33573)
--	g1283 = DFF(g34730)
--	g433 = DFF(g24205)
--	g4297 = DFF(g4294)
--	g5983 = DFF(g6005)
--	g1459 = DFF(g1399)
--	g758 = DFF(g32979)
--	g5712 = DFF(g25731)
--	g4138 = DFF(g28078)
--	g4639 = DFF(g34025)
--	g6537 = DFF(g25763)
--	g5543 = DFF(g30481)
--	g1582 = DFF(g1500)
--	g3736 = DFF(g31890)
--	g5961 = DFF(g30517)
--	g6243 = DFF(g30539)
--	g632 = DFF(g34880)
--	g1227 = DFF(g24242)
--	g3889 = DFF(g30436)
--	g3476 = DFF(g29265)
--	g1664 = DFF(g32990)
--	g1246 = DFF(g24245)
--	g6128 = DFF(g25739)
--	g6629 = DFF(g30553)
--	g246 = DFF(g26907)
--	g4049 = DFF(g24278)
--	g4449 = DFF(g26955)
--	g2932 = DFF(g24282)
--	g4575 = DFF(g29276)
--	g4098 = DFF(g31894)
--	g4498 = DFF(g33037)
--	g528 = DFF(g26894)
--	g5436 = DFF(g25711)
--	g16 = DFF(g34593)
--	g3139 = DFF(g25654)
--	g102 = DFF(g33962)
--	g4584 = DFF(g34451)
--	g142 = DFF(g34250)
--	g5335 = DFF(g5331)
--	g5831 = DFF(g29295)
--	g239 = DFF(g26905)
--	g1216 = DFF(g25629)
--	g2848 = DFF(g34792)
--	g5805 = DFF(g5798)
--	g5022 = DFF(g25703)
--	g4019 = DFF(g4000)
--	g1030 = DFF(g32983)
--	g3672 = DFF(g3668)
--	g3231 = DFF(g30402)
--	g6490 = DFF(g25757)
--	g1430 = DFF(g1426)
--	g4452 = DFF(g4446)
--	g2241 = DFF(g33999)
--	g1564 = DFF(g24262)
--	g5798 = DFF(g25729)
--	g6148 = DFF(g6140)
--	g6649 = DFF(g30558)
--	g110 = DFF(g34848)
--	g884 = DFF(g881)
--	g3742 = DFF(g31892)
--	g225 = DFF(g26901)
--	g4486 = DFF(g26961)
--	g4504 = DFF(g33039)
--	g5873 = DFF(g33059)
--	g5037 = DFF(g31899)
--	g2319 = DFF(g33007)
--	g5495 = DFF(g25720)
--	g4185 = DFF(g21891)
--	g5208 = DFF(g30462)
--	g2152 = DFF(g18422)
--	g5579 = DFF(g30487)
--	g5869 = DFF(g33058)
--	g5719 = DFF(g31916)
--	g1589 = DFF(g24261)
--	g5752 = DFF(g25730)
--	g6279 = DFF(g30531)
--	g5917 = DFF(g30506)
--	g2975 = DFF(g34804)
--	g6167 = DFF(g25747)
--	g3983 = DFF(g4005)
--	g2599 = DFF(g33601)
--	g1448 = DFF(g26922)
--	g881 = DFF(g878)
--	g3712 = DFF(g25679)
--	g2370 = DFF(g29250)
--	g5164 = DFF(g30459)
--	g1333 = DFF(g1582)
--	g153 = DFF(g33534)
--	g6549 = DFF(g30543)
--	g4087 = DFF(g29275)
--	g4801 = DFF(g34030)
--	g2984 = DFF(g34980)
--	g3961 = DFF(g30451)
--	g5770 = DFF(g25723)
--	g962 = DFF(g25627)
--	g101 = DFF(g34787)
--	g4226 = DFF(g4222)
--	g6625 = DFF(g30552)
--	g51 = DFF(g34996)
--	g1018 = DFF(g30337)
--	g1418 = DFF(g24254)
--	g4045 = DFF(g24277)
--	g1467 = DFF(g29237)
--	g2461 = DFF(g30378)
--	g5706 = DFF(g31912)
--	g457 = DFF(g25603)
--	g2756 = DFF(g33019)
--	g5990 = DFF(g33623)
--	g471 = DFF(g25608)
--	g1256 = DFF(g29235)
--	g5029 = DFF(g31902)
--	g6519 = DFF(g29306)
--	g4169 = DFF(g28080)
--	g1816 = DFF(g33978)
--	g4369 = DFF(g26970)
--	g3436 = DFF(g25660)
--	g5787 = DFF(g25726)
--	g4578 = DFF(g29278)
--	g4459 = DFF(g34253)
--	g3831 = DFF(g29272)
--	g2514 = DFF(g33595)
--	g3288 = DFF(g33610)
--	g2403 = DFF(g33589)
--	g2145 = DFF(g34605)
--	g1700 = DFF(g30350)
--	g513 = DFF(g25611)
--	g2841 = DFF(g26936)
--	g5297 = DFF(g33619)
--	g3805 = DFF(g3798)
--	g2763 = DFF(g34022)
--	g4793 = DFF(g34033)
--	g952 = DFF(g34726)
--	g1263 = DFF(g31870)
--	g1950 = DFF(g33985)
--	g5138 = DFF(g29283)
--	g2307 = DFF(g34003)
--	g5109 = DFF(g5101)
--	g5791 = DFF(g25727)
--	g3798 = DFF(g25677)
--	g4664 = DFF(g34463)
--	g2223 = DFF(g33006)
--	g5808 = DFF(g29292)
--	g6645 = DFF(g30557)
--	g2016 = DFF(g33989)
--	g5759 = DFF(g28098)
--	g3873 = DFF(g33033)
--	g3632 = DFF(g3654)
--	g2315 = DFF(g34005)
--	g2811 = DFF(g26932)
--	g5957 = DFF(g30516)
--	g2047 = DFF(g33575)
--	g3869 = DFF(g33032)
--	g6358 = DFF(g6329)
--	g3719 = DFF(g31891)
--	g5575 = DFF(g30486)
--	g46 = DFF(g34991)
--	g3752 = DFF(g25678)
--	g3917 = DFF(g30440)
--	g4188 = DFF(g4191)
--	g1585 = DFF(g1570)
--	g4388 = DFF(g26949)
--	g6275 = DFF(g30530)
--	g6311 = DFF(g30542)
--	g4216 = DFF(g4213)
--	g1041 = DFF(g25624)
--	g2595 = DFF(g30383)
--	g2537 = DFF(g33597)
--	g136 = DFF(g34598)
--	g4430 = DFF(g26957)
--	g4564 = DFF(g26967)
--	g3454 = DFF(g3447)
--	g4826 = DFF(g28102)
--	g6239 = DFF(g30524)
--	g3770 = DFF(g25671)
--	g232 = DFF(g26903)
--	g5268 = DFF(g30475)
--	g6545 = DFF(g34647)
--	g2417 = DFF(g30377)
--	g1772 = DFF(g33553)
--	g4741 = DFF(g21902)
--	g5052 = DFF(g31903)
--	g5452 = DFF(g25715)
--	g1890 = DFF(g33984)
--	g2629 = DFF(g33602)
--	g572 = DFF(g28045)
--	g2130 = DFF(g34603)
--	g4108 = DFF(g33035)
--	g4308 = DFF(g4304)
--	g475 = DFF(g24208)
--	g990 = DFF(g1239)
--	g31 = DFF(g34596)
--	g3412 = DFF(g28064)
--	g45 = DFF(g34990)
--	g799 = DFF(g24213)
--	g3706 = DFF(g31887)
--	g3990 = DFF(g33614)
--	g5385 = DFF(g31907)
--	g5881 = DFF(g33060)
--	g1992 = DFF(g30362)
--	g3029 = DFF(g31875)
--	g3171 = DFF(g33023)
--	g3787 = DFF(g25674)
--	g812 = DFF(g26898)
--	g832 = DFF(g25618)
--	g5897 = DFF(g30518)
--	g4165 = DFF(g28079)
--	g4571 = DFF(g6974)
--	g3281 = DFF(g3303)
--	g4455 = DFF(g26959)
--	g2902 = DFF(g34801)
--	g333 = DFF(g26884)
--	g168 = DFF(g25600)
--	g2823 = DFF(g26933)
--	g3684 = DFF(g28066)
--	g3639 = DFF(g33612)
--	g5331 = DFF(g5327)
--	g3338 = DFF(g24268)
--	g5406 = DFF(g25716)
--	g3791 = DFF(g25675)
--	g269 = DFF(g26906)
--	g401 = DFF(g24203)
--	g6040 = DFF(g24346)
--	g441 = DFF(g24207)
--	g5105 = DFF(g25701)
--	g3808 = DFF(g29269)
--	g9 = DFF(g34592)
--	g3759 = DFF(g28068)
--	g4467 = DFF(g34255)
--	g3957 = DFF(g30450)
--	g4093 = DFF(g30456)
--	g1760 = DFF(g32991)
--	g6151 = DFF(g6144)
--	g6351 = DFF(g24348)
--	g160 = DFF(g34249)
--	g5445 = DFF(g25713)
--	g5373 = DFF(g31909)
--	g2279 = DFF(g30371)
--	g3498 = DFF(g29268)
--	g586 = DFF(g29224)
--	g869 = DFF(g859)
--	g2619 = DFF(g33017)
--	g1183 = DFF(g30339)
--	g1608 = DFF(g33967)
--	g4197 = DFF(g4194)
--	g5283 = DFF(g5276)
--	g1779 = DFF(g33559)
--	g2652 = DFF(g29255)
--	g5459 = DFF(g5452)
--	g2193 = DFF(g30368)
--	g2393 = DFF(g30375)
--	g5767 = DFF(g25732)
--	g661 = DFF(g28052)
--	g4950 = DFF(g28089)
--	g5535 = DFF(g33055)
--	g2834 = DFF(g30392)
--	g1361 = DFF(g30343)
--	g3419 = DFF(g25657)
--	g6235 = DFF(g30523)
--	g1146 = DFF(g24233)
--	g2625 = DFF(g33018)
--	g150 = DFF(g32976)
--	g1696 = DFF(g30349)
--	g6555 = DFF(g33067)
--	g859 = DFF(g26900)
--	g3385 = DFF(g31883)
--	g3881 = DFF(g33034)
--	g6621 = DFF(g30551)
--	g3470 = DFF(g25667)
--	g3897 = DFF(g30452)
--	g518 = DFF(g25612)
--	g3025 = DFF(g31874)
--	g538 = DFF(g34719)
--	g2606 = DFF(g33607)
--	g1472 = DFF(g26923)
--	g6113 = DFF(g25746)
--	g542 = DFF(g24211)
--	g5188 = DFF(g33050)
--	g5689 = DFF(g24341)
--	g1116 = DFF(g1056)
--	g405 = DFF(g24201)
--	g5216 = DFF(g30463)
--	g6494 = DFF(g6486)
--	g4669 = DFF(g34464)
--	g5428 = DFF(g25710)
--	g996 = DFF(g24243)
--	g4531 = DFF(g24335)
--	g2860 = DFF(g34611)
--	g4743 = DFF(g34262)
--	g6593 = DFF(g30546)
--	g2710 = DFF(g18527)
--	g215 = DFF(g25591)
--	g4411 = DFF(g4414)
--	g1413 = DFF(g30347)
--	g4474 = DFF(g10384)
--	g5308 = DFF(g5283)
--	g6641 = DFF(g30556)
--	g3045 = DFF(g33020)
--	g6 = DFF(g34589)
--	g1936 = DFF(g33562)
--	g55 = DFF(g35002)
--	g504 = DFF(g25610)
--	g2587 = DFF(g33015)
--	g4480 = DFF(g31896)
--	g2311 = DFF(g34004)
--	g3602 = DFF(g30428)
--	g5571 = DFF(g30485)
--	g3578 = DFF(g30422)
--	g468 = DFF(g25606)
--	g5448 = DFF(g25714)
--	g3767 = DFF(g25680)
--	g5827 = DFF(g29294)
--	g3582 = DFF(g30423)
--	g6271 = DFF(g30529)
--	g4688 = DFF(g34028)
--	g5774 = DFF(g25724)
--	g2380 = DFF(g33587)
--	g5196 = DFF(g30460)
--	g5396 = DFF(g31910)
--	g3227 = DFF(g30401)
--	g2020 = DFF(g33990)
--	g4000 = DFF(g3976)
--	g1079 = DFF(g1075)
--	g6541 = DFF(g29309)
--	g3203 = DFF(g30411)
--	g1668 = DFF(g33546)
--	g4760 = DFF(g28085)
--	g262 = DFF(g26904)
--	g1840 = DFF(g33556)
--	g70 = DFF(g18093)
--	g5467 = DFF(g25722)
--	g460 = DFF(g25605)
--	g6209 = DFF(g33062)
--	g74 = DFF(g26893)
--	g5290 = DFF(g5313)
--	g655 = DFF(g28050)
--	g3502 = DFF(g34626)
--	g2204 = DFF(g33583)
--	g5256 = DFF(g30472)
--	g4608 = DFF(g34454)
--	g794 = DFF(g34850)
--	g4023 = DFF(g4019)
--	g4423 = DFF(g4537)
--	g3689 = DFF(g24272)
--	g5381 = DFF(g31906)
--	g5685 = DFF(g5681)
--	g703 = DFF(g24214)
--	g5421 = DFF(g25718)
--	g862 = DFF(g26909)
--	g3247 = DFF(g30406)
--	g2040 = DFF(g33569)
--	g4999 = DFF(g25694)
--	g4146 = DFF(g34628)
--	g4633 = DFF(g34458)
--	g1157 = DFF(g24240)
--	g5723 = DFF(g31918)
--	g4732 = DFF(g34634)
--	g5101 = DFF(g25700)
--	g5817 = DFF(g29293)
--	g2151 = DFF(g18421)
--	g2351 = DFF(g33009)
--	g2648 = DFF(g33603)
--	g6736 = DFF(g24355)
--	g4944 = DFF(g34268)
--	g4072 = DFF(g25691)
--	g344 = DFF(g26890)
--	g4443 = DFF(g4449)
--	g3466 = DFF(g29264)
--	g4116 = DFF(g28072)
--	g5041 = DFF(g31900)
--	g5441 = DFF(g25712)
--	g4434 = DFF(g26956)
--	g3827 = DFF(g29271)
--	g6500 = DFF(g29304)
--	g5673 = DFF(g5654)
--	g3133 = DFF(g29261)
--	g3333 = DFF(g28063)
--	g979 = DFF(g1116)
--	g4681 = DFF(g34027)
--	g298 = DFF(g33961)
--	g3774 = DFF(g25672)
--	g2667 = DFF(g33604)
--	g3396 = DFF(g33025)
--	g4210 = DFF(g4207)
--	g1894 = DFF(g32995)
--	g2988 = DFF(g34624)
--	g3538 = DFF(g30415)
--	g301 = DFF(g33536)
--	g341 = DFF(g26888)
--	g827 = DFF(g28055)
--	g1075 = DFF(g24238)
--	g6077 = DFF(g31921)
--	g2555 = DFF(g33600)
--	g5011 = DFF(g28105)
--	g199 = DFF(g34721)
--	g6523 = DFF(g29307)
--	g1526 = DFF(g30345)
--	g4601 = DFF(g34453)
--	g854 = DFF(g32980)
--	g1484 = DFF(g29238)
--	g4922 = DFF(g34639)
--	g5080 = DFF(g25695)
--	g5863 = DFF(g33057)
--	g4581 = DFF(g26969)
--	g3021 = DFF(g31879)
--	g2518 = DFF(g29253)
--	g2567 = DFF(g34021)
--	g568 = DFF(g26895)
--	g3263 = DFF(g30413)
--	g6613 = DFF(g30549)
--	g6044 = DFF(g24347)
--	g6444 = DFF(g25758)
--	g2965 = DFF(g34808)
--	g5857 = DFF(g30501)
--	g1616 = DFF(g33969)
--	g890 = DFF(g34440)
--	g5976 = DFF(g5969)
--	g3562 = DFF(g30433)
--	g4294 = DFF(g21900)
--	g1404 = DFF(g26921)
--	g3723 = DFF(g31893)
--	g3817 = DFF(g29270)
--	g93 = DFF(g34878)
--	g4501 = DFF(g33038)
--	g287 = DFF(g31865)
--	g2724 = DFF(g26926)
--	g4704 = DFF(g28083)
--	g22 = DFF(g29209)
--	g2878 = DFF(g34797)
--	g5220 = DFF(g30478)
--	g617 = DFF(g34724)
--	g637 = DFF(g24212)
--	g316 = DFF(g26883)
--	g1277 = DFF(g32985)
--	g6513 = DFF(g25761)
--	g336 = DFF(g26886)
--	g2882 = DFF(g34796)
--	g933 = DFF(g32982)
--	g1906 = DFF(g33561)
--	g305 = DFF(g26880)
--	g8 = DFF(g34591)
--	g3368 = DFF(g31884)
--	g2799 = DFF(g26931)
--	g887 = DFF(g884)
--	g5327 = DFF(g5308)
--	g4912 = DFF(g34641)
--	g4157 = DFF(g34629)
--	g2541 = DFF(g33598)
--	g2153 = DFF(g33576)
--	g550 = DFF(g34720)
--	g255 = DFF(g26902)
--	g1945 = DFF(g29244)
--	g5240 = DFF(g30468)
--	g1478 = DFF(g26924)
--	g3080 = DFF(g25645)
--	g3863 = DFF(g33031)
--	g1959 = DFF(g29245)
--	g3480 = DFF(g29266)
--	g6653 = DFF(g30559)
--	g6719 = DFF(g6715)
--	g2864 = DFF(g34794)
--	g4894 = DFF(g28087)
--	g5681 = DFF(g5677)
--	g3857 = DFF(g30435)
--	g3976 = DFF(g3969)
--	g499 = DFF(g25609)
--	g5413 = DFF(g28095)
--	g1002 = DFF(g28057)
--	g776 = DFF(g34439)
--	g28 = DFF(g34595)
--	g1236 = DFF(g1233)
--	g4646 = DFF(g34260)
--	g2476 = DFF(g33012)
--	g1657 = DFF(g32989)
--	g2375 = DFF(g34006)
--	g63 = DFF(g34847)
--	g6012 = DFF(g5983)
--	g358 = DFF(g365)
--	g896 = DFF(g26910)
--	g967 = DFF(g21722)
--	g3423 = DFF(g25658)
--	g283 = DFF(g28043)
--	g3161 = DFF(g33021)
--	g2384 = DFF(g29251)
--	g3361 = DFF(g25665)
--	g6675 = DFF(g6697)
--	g4616 = DFF(g34456)
--	g4561 = DFF(g26968)
--	g2024 = DFF(g33991)
--	g3451 = DFF(g3443)
--	g2795 = DFF(g26930)
--	g613 = DFF(g34599)
--	g4527 = DFF(g28082)
--	g1844 = DFF(g33557)
--	g5937 = DFF(g30511)
--	g4546 = DFF(g33045)
--	g3103 = DFF(g3096)
--	g2523 = DFF(g30379)
--	g3303 = DFF(g24267)
--	g2643 = DFF(g34020)
--	g6109 = DFF(g28100)
--	g1489 = DFF(g24249)
--	g5390 = DFF(g31908)
--	g194 = DFF(g25592)
--	g2551 = DFF(g30382)
--	g5156 = DFF(g29285)
--	g3072 = DFF(g25644)
--	g1242 = DFF(g1227)
--	g47 = DFF(g34992)
--	g3443 = DFF(g25662)
--	g4277 = DFF(g21896)
--	g1955 = DFF(g33563)
--	g6049 = DFF(g33622)
--	g3034 = DFF(g31876)
--	g2273 = DFF(g33582)
--	g6715 = DFF(g6711)
--	g4771 = DFF(g28086)
--	g6098 = DFF(g25744)
--	g3147 = DFF(g29262)
--	g3347 = DFF(g24270)
--	g2269 = DFF(g33581)
--	g191 = DFF(g194)
--	g2712 = DFF(g26937)
--	g626 = DFF(g34849)
--	g2729 = DFF(g28060)
--	g5357 = DFF(g33618)
--	g4991 = DFF(g34038)
--	g6019 = DFF(g6000)
--	g4709 = DFF(g34032)
--	g6419 = DFF(g31927)
--	g6052 = DFF(g31919)
--	g2927 = DFF(g34803)
--	g4340 = DFF(g34459)
--	g5929 = DFF(g30509)
--	g4907 = DFF(g34640)
--	g3317 = DFF(g3298)
--	g4035 = DFF(g28069)
--	g2946 = DFF(g21899)
--	g918 = DFF(g31868)
--	g4082 = DFF(g26938)
--	g6486 = DFF(g25756)
--	g2036 = DFF(g30363)
--	g577 = DFF(g30334)
--	g1620 = DFF(g33970)
--	g2831 = DFF(g30391)
--	g667 = DFF(g25615)
--	g930 = DFF(g33540)
--	g3937 = DFF(g30445)
--	g5782 = DFF(g25725)
--	g817 = DFF(g25617)
--	g1249 = DFF(g24247)
--	g837 = DFF(g24215)
--	g3668 = DFF(g3649)
--	g599 = DFF(g33964)
--	g5475 = DFF(g25719)
--	g739 = DFF(g29228)
--	g5949 = DFF(g30514)
--	g6682 = DFF(g33627)
--	g6105 = DFF(g28101)
--	g904 = DFF(g24231)
--	g2873 = DFF(g34615)
--	g1854 = DFF(g30356)
--	g5084 = DFF(g25696)
--	g5603 = DFF(g30493)
--	g4222 = DFF(g4219)
--	g2495 = DFF(g33594)
--	g2437 = DFF(g34009)
--	g2102 = DFF(g30365)
--	g2208 = DFF(g33004)
--	g2579 = DFF(g34018)
--	g4064 = DFF(g25685)
--	g4899 = DFF(g34040)
--	g2719 = DFF(g25639)
--	g4785 = DFF(g34029)
--	g5583 = DFF(g30488)
--	g781 = DFF(g34600)
--	g6173 = DFF(g29300)
--	g6373 = DFF(g6369)
--	g2917 = DFF(g34802)
--	g686 = DFF(g25614)
--	g1252 = DFF(g28058)
--	g671 = DFF(g29225)
--	g2265 = DFF(g33580)
--	g6283 = DFF(g30532)
--	g6369 = DFF(g6365)
--	g5276 = DFF(g5320)
--	g6459 = DFF(g25760)
--	g901 = DFF(g25620)
--	g4194 = DFF(g4188)
--	g5527 = DFF(g33054)
--	g4489 = DFF(g26962)
--	g1974 = DFF(g33564)
--	g1270 = DFF(g32984)
--	g4966 = DFF(g34039)
--	g6415 = DFF(g31932)
--	g6227 = DFF(g33065)
--	g3929 = DFF(g30443)
--	g5503 = DFF(g29291)
--	g4242 = DFF(g24279)
--	g5925 = DFF(g30508)
--	g1124 = DFF(g29232)
--	g4955 = DFF(g34269)
--	g5224 = DFF(g30464)
--	g2012 = DFF(g33988)
--	g6203 = DFF(g30522)
--	g5120 = DFF(g25708)
--	g5320 = DFF(g5290)
--	g2389 = DFF(g30374)
--	g4438 = DFF(g26953)
--	g2429 = DFF(g34008)
--	g2787 = DFF(g34444)
--	g1287 = DFF(g34731)
--	g2675 = DFF(g33606)
--	g66 = DFF(g24334)
--	g4836 = DFF(g34265)
--	g1199 = DFF(g30340)
--	g1399 = DFF(g24257)
--	g5547 = DFF(g30482)
--	g3782 = DFF(g25673)
--	g6428 = DFF(g31929)
--	g2138 = DFF(g34604)
--	g3661 = DFF(g3632)
--	g2338 = DFF(g33591)
--	g4229 = DFF(g4226)
--	g6247 = DFF(g30525)
--	g2791 = DFF(g26929)
--	g3949 = DFF(g30448)
--	g1291 = DFF(g34602)
--	g5945 = DFF(g30513)
--	g5244 = DFF(g30469)
--	g2759 = DFF(g33608)
--	g6741 = DFF(g33626)
--	g785 = DFF(g34725)
--	g1259 = DFF(g30342)
--	g3484 = DFF(g29267)
--	g209 = DFF(g25593)
--	g6609 = DFF(g30548)
--	g5517 = DFF(g33052)
--	g2449 = DFF(g34012)
--	g2575 = DFF(g34017)
--	g65 = DFF(g34785)
--	g2715 = DFF(g24263)
--	g936 = DFF(g26912)
--	g2098 = DFF(g30364)
--	g4462 = DFF(g34254)
--	g604 = DFF(g34251)
--	g6589 = DFF(g30560)
--	g1886 = DFF(g33983)
--	g6466 = DFF(g25752)
--	g6365 = DFF(g6346)
--	g6711 = DFF(g6692)
--	g429 = DFF(g24204)
--	g1870 = DFF(g33980)
--	g4249 = DFF(g34631)
--	g6455 = DFF(g28103)
--	g3004 = DFF(g31873)
--	g1825 = DFF(g29243)
--	g6133 = DFF(g25740)
--	g1008 = DFF(g25623)
--	g4392 = DFF(g26950)
--	g5002 = DFF(g4999)
--	g3546 = DFF(g30431)
--	g5236 = DFF(g30467)
--	g1768 = DFF(g30353)
--	g4854 = DFF(g34467)
--	g3925 = DFF(g30442)
--	g6509 = DFF(g29305)
--	g732 = DFF(g25616)
--	g2504 = DFF(g29252)
--	g1322 = DFF(g1459)
--	g4520 = DFF(g6972)
--	g4219 = DFF(g4216)
--	g2185 = DFF(g33003)
--	g37 = DFF(g34613)
--	g4031 = DFF(g4027)
--	g2070 = DFF(g33570)
--	g4812 = DFF(g4809)
--	g6093 = DFF(g33061)
--	g968 = DFF(g21723)
--	g4176 = DFF(g34734)
--	g4005 = DFF(g24275)
--	g4405 = DFF(g4408)
--	g872 = DFF(g887)
--	g6181 = DFF(g29302)
--	g6381 = DFF(g24349)
--	g4765 = DFF(g34264)
--	g5563 = DFF(g30484)
--	g1395 = DFF(g25634)
--	g1913 = DFF(g33567)
--	g2331 = DFF(g33585)
--	g6263 = DFF(g30527)
--	g50 = DFF(g34995)
--	g3945 = DFF(g30447)
--	g347 = DFF(g344)
--	g5731 = DFF(g31914)
--	g4473 = DFF(g34256)
--	g1266 = DFF(g25630)
--	g5489 = DFF(g29290)
--	g714 = DFF(g29227)
--	g2748 = DFF(g31872)
--	g5471 = DFF(g29287)
--	g4540 = DFF(g31897)
--	g6723 = DFF(g6719)
--	g6605 = DFF(g30562)
--	g2445 = DFF(g34011)
--	g2173 = DFF(g33996)
--	g4287 = DFF(g21898)
--	g2491 = DFF(g33014)
--	g4849 = DFF(g34465)
--	g2169 = DFF(g33995)
--	g2283 = DFF(g30372)
--	g6585 = DFF(g30545)
--	g121 = DFF(g30389)
--	g2407 = DFF(g33590)
--	g2868 = DFF(g34616)
--	g2767 = DFF(g26927)
--	g1783 = DFF(g32992)
--	g3310 = DFF(g3281)
--	g1312 = DFF(g25631)
--	g5212 = DFF(g30477)
--	g4245 = DFF(g34632)
--	g645 = DFF(g28046)
--	g4291 = DFF(g4287)
--	g79 = DFF(g26896)
--	g182 = DFF(g25602)
--	g1129 = DFF(g26916)
--	g2227 = DFF(g33578)
--	g6058 = DFF(g25745)
--	g4207 = DFF(g4204)
--	g2246 = DFF(g33579)
--	g1830 = DFF(g30354)
--	g3590 = DFF(g30425)
--	g392 = DFF(g24200)
--	g1592 = DFF(g33544)
--	g6505 = DFF(g25764)
--	g6411 = DFF(g31930)
--	g1221 = DFF(g24246)
--	g5921 = DFF(g30507)
--	g106 = DFF(g26889)
--	g146 = DFF(g30333)
--	g218 = DFF(g215)
--	g6474 = DFF(g25753)
--	g1932 = DFF(g32998)
--	g1624 = DFF(g32987)
--	g5062 = DFF(g25702)
--	g5462 = DFF(g29286)
--	g2689 = DFF(g34606)
--	g6573 = DFF(g33070)
--	g1677 = DFF(g29240)
--	g2028 = DFF(g32999)
--	g2671 = DFF(g33605)
--	g1576 = DFF(g24255)
--	g4408 = DFF(g26945)
--	g34 = DFF(g34877)
--	g1848 = DFF(g33558)
--	g3089 = DFF(g25647)
--	g3731 = DFF(g31889)
--	g86 = DFF(g25699)
--	g5485 = DFF(g29289)
--	g2741 = DFF(g30388)
--	g802 = DFF(g799)
--	g2638 = DFF(g29254)
--	g4122 = DFF(g28074)
--	g4322 = DFF(g34450)
--	g5941 = DFF(g30512)
--	g2108 = DFF(g33572)
--	g6000 = DFF(g5976)
--	g25 = DFF(g15048)
--	g1644 = DFF(g33551)
--	g595 = DFF(g33538)
--	g2217 = DFF(g33005)
--	g1319 = DFF(g24248)
--	g2066 = DFF(g33002)
--	g1152 = DFF(g24234)
--	g5252 = DFF(g30471)
--	g2165 = DFF(g34000)
--	g2571 = DFF(g34016)
--	g5176 = DFF(g33048)
--	g391 = DFF(g26911)
--	g5005 = DFF(g5002)
--	g2711 = DFF(g18528)
--	g6023 = DFF(g6019)
--	g1211 = DFF(g25628)
--	g2827 = DFF(g26934)
--	g6423 = DFF(g31928)
--	g875 = DFF(g869)
--	g4859 = DFF(g34468)
--	g424 = DFF(g24202)
--	g1274 = DFF(g33542)
--	g1426 = DFF(g1422)
--	g85 = DFF(g34717)
--	g2803 = DFF(g34445)
--	g6451 = DFF(g28104)
--	g1821 = DFF(g33555)
--	g2509 = DFF(g34013)
--	g5073 = DFF(g28091)
--	g1280 = DFF(g26919)
--	g4815 = DFF(g4812)
--	g6346 = DFF(g6322)
--	g6633 = DFF(g30554)
--	g5124 = DFF(g29281)
--	g1083 = DFF(g1079)
--	g6303 = DFF(g30537)
--	g5069 = DFF(g28092)
--	g2994 = DFF(g34732)
--	g650 = DFF(g28049)
--	g1636 = DFF(g33545)
--	g3921 = DFF(g30441)
--	g2093 = DFF(g29247)
--	g6732 = DFF(g24354)
--	g1306 = DFF(g25636)
--	g5377 = DFF(g31911)
--	g1061 = DFF(g26914)
--	g3462 = DFF(g25670)
--	g2181 = DFF(g33998)
--	g956 = DFF(g25626)
--	g1756 = DFF(g33977)
--	g5849 = DFF(g29297)
--	g4112 = DFF(g28071)
--	g2685 = DFF(g30387)
--	g2197 = DFF(g33577)
--	g6116 = DFF(g25737)
--	g2421 = DFF(g33592)
--	g1046 = DFF(g26913)
--	g482 = DFF(g28044)
--	g4401 = DFF(g26948)
--	g6434 = DFF(g31931)
--	g1514 = DFF(g30344)
--	g329 = DFF(g26885)
--	g6565 = DFF(g33069)
--	g2950 = DFF(g34621)
--	g4129 = DFF(g28075)
--	g1345 = DFF(g28059)
--	g6533 = DFF(g25762)
--	g3298 = DFF(g3274)
--	g3085 = DFF(g25646)
--	g4727 = DFF(g34633)
--	g6697 = DFF(g24352)
--	g1536 = DFF(g26925)
--	g3941 = DFF(g30446)
--	g370 = DFF(g25597)
--	g5694 = DFF(g24342)
--	g1858 = DFF(g30357)
--	g446 = DFF(g26908)
--	g4932 = DFF(g21905)
--	g3219 = DFF(g30399)
--	g1811 = DFF(g29242)
--	g3431 = DFF(g25659)
--	g6601 = DFF(g30547)
--	g3376 = DFF(g31881)
--	g2441 = DFF(g34010)
--	g1874 = DFF(g33986)
--	g4349 = DFF(g34257)
--	g6581 = DFF(g30544)
--	g6597 = DFF(g30561)
--	g5008 = DFF(g5005)
--	g3610 = DFF(g30430)
--	g2890 = DFF(g34799)
--	g1978 = DFF(g33565)
--	g1612 = DFF(g33968)
--	g112 = DFF(g34879)
--	g2856 = DFF(g34793)
--	g6479 = DFF(g25754)
--	g1982 = DFF(g33566)
--	g6668 = DFF(g6661)
--	g5228 = DFF(g30465)
--	g4119 = DFF(g28073)
--	g6390 = DFF(g24351)
--	g1542 = DFF(g30346)
--	g4258 = DFF(g21893)
--	g4818 = DFF(g4815)
--	g5033 = DFF(g31904)
--	g4717 = DFF(g34635)
--	g1554 = DFF(g25637)
--	g3849 = DFF(g29274)
--	g6704 = DFF(g6675)
--	g3199 = DFF(g30396)
--	g5845 = DFF(g25735)
--	g4975 = DFF(g34037)
--	g790 = DFF(g34791)
--	g5913 = DFF(g30520)
--	g1902 = DFF(g30358)
--	g6163 = DFF(g29299)
--	g4125 = DFF(g28081)
--	g4821 = DFF(g28096)
--	g4939 = DFF(g28088)
--	g1056 = DFF(g24241)
--	g3207 = DFF(g30397)
--	g4483 = DFF(g4520)
--	g3259 = DFF(g30409)
--	g5142 = DFF(g29284)
--	g5248 = DFF(g30470)
--	g2126 = DFF(g30367)
--	g3694 = DFF(g24273)
--	g5481 = DFF(g29288)
--	g1964 = DFF(g30359)
--	g5097 = DFF(g25698)
--	g3215 = DFF(g30398)
--	g4027 = DFF(g4023)
--	g111 = DFF(g34718)
--	g4427 = DFF(g26952)
--	g7 = DFF(g34590)
--	g2779 = DFF(g26928)
--	g4200 = DFF(g4197)
--	g4446 = DFF(g26954)
--	g1720 = DFF(g30351)
--	g1367 = DFF(g31871)
--	g5112 = DFF(g5105)
--	g19 = DFF(g34594)
--	g4145 = DFF(g26939)
--	g2161 = DFF(g33994)
--	g376 = DFF(g25596)
--	g2361 = DFF(g33586)
--	g4191 = DFF(g21901)
--	g582 = DFF(g31866)
--	g2051 = DFF(g33000)
--	g1193 = DFF(g26918)
--	g5401 = DFF(g33051)
--	g3408 = DFF(g28065)
--	g2327 = DFF(g30373)
--	g907 = DFF(g28056)
--	g947 = DFF(g34601)
--	g1834 = DFF(g30355)
--	g3594 = DFF(g30426)
--	g2999 = DFF(g34805)
--	g5727 = DFF(g31913)
--	g2303 = DFF(g34002)
--	g6661 = DFF(g6704)
--	g3065 = DFF(g25652)
--	g699 = DFF(g28053)
--	g723 = DFF(g29229)
--	g5703 = DFF(g33620)
--	g546 = DFF(g34722)
--	g2472 = DFF(g33599)
--	g5953 = DFF(g30515)
--	g3096 = DFF(g25649)
--	g6439 = DFF(g33066)
--	g1740 = DFF(g33979)
--	g3550 = DFF(g30417)
--	g3845 = DFF(g25683)
--	g2116 = DFF(g33574)
--	g5677 = DFF(g5673)
--	g3195 = DFF(g30410)
--	g3913 = DFF(g30454)
--	g4537 = DFF(g34024)
--	g1687 = DFF(g33547)
--	g2681 = DFF(g30386)
--	g2533 = DFF(g33596)
--	g324 = DFF(g26887)
--	g2697 = DFF(g34607)
--	g5747 = DFF(g33056)
--	g4417 = DFF(g31895)
--	g6561 = DFF(g33068)
--	g1141 = DFF(g29233)
--	g1570 = DFF(g24258)
--	g2413 = DFF(g30376)
--	g1710 = DFF(g33549)
--	g6527 = DFF(g29308)
--	g6404 = DFF(g25759)
--	g3255 = DFF(g30408)
--	g1691 = DFF(g29241)
--	g2936 = DFF(g34620)
--	g5644 = DFF(g33621)
--	g5152 = DFF(g25707)
--	g5352 = DFF(g24339)
--	g4213 = DFF(g4185)
--	g6120 = DFF(g25738)
--	g2775 = DFF(g34443)
--	g2922 = DFF(g34619)
--	g1111 = DFF(g29234)
--	g5893 = DFF(g30503)
--	g1311 = DFF(g21724)
--	g3267 = DFF(g3310)
--	g6617 = DFF(g30550)
--	g2060 = DFF(g33001)
--	g4512 = DFF(g33040)
--	g5599 = DFF(g30492)
--	g3401 = DFF(g25664)
--	g4366 = DFF(g26944)
--	g3676 = DFF(g3672)
--	g94 = DFF(g34614)
--	g3129 = DFF(g29260)
--	g3329 = DFF(g3325)
--	g5170 = DFF(g33047)
--	g4456 = DFF(g25692)
--	g5821 = DFF(g25733)
--	g6299 = DFF(g30536)
--	g1239 = DFF(g1157)
--	g3727 = DFF(g31888)
--	g2079 = DFF(g29246)
--	g4698 = DFF(g34261)
--	g3703 = DFF(g33611)
--	g1559 = DFF(g25638)
--	g943 = DFF(g34728)
--	g411 = DFF(g29222)
--	g6140 = DFF(g25742)
--	g3953 = DFF(g30449)
--	g3068 = DFF(g25643)
--	g2704 = DFF(g34608)
--	g6035 = DFF(g24345)
--	g6082 = DFF(g31922)
--	g49 = DFF(g34994)
--	g1300 = DFF(g25635)
--	g4057 = DFF(g25686)
--	g5200 = DFF(g30461)
--	g4843 = DFF(g34466)
--	g5046 = DFF(g31901)
--	g2250 = DFF(g29249)
--	g319 = DFF(g26882)
--	g4549 = DFF(g33041)
--	g2453 = DFF(g33011)
--	g5841 = DFF(g25734)
--	g5763 = DFF(g28097)
--	g3747 = DFF(g33030)
--	g5637 = DFF(g5659)
--	g2912 = DFF(g34618)
--	g2357 = DFF(g33010)
--	g4232 = DFF(g4229)
--	g164 = DFF(g31864)
--	g4253 = DFF(g34630)
--	g5016 = DFF(g31898)
--	g3119 = DFF(g25653)
--	g1351 = DFF(g25632)
--	g1648 = DFF(g32988)
--	g4519 = DFF(g33616)
--	g5115 = DFF(g29280)
--	g3352 = DFF(g33609)
--	g6657 = DFF(g30563)
--	g4552 = DFF(g33044)
--	g3893 = DFF(g30437)
--	g3211 = DFF(g30412)
--	g5654 = DFF(g5630)
--	g929 = DFF(g21725)
--	g3274 = DFF(g3267)
--	g5595 = DFF(g30491)
--	g3614 = DFF(g30434)
--	g2894 = DFF(g34612)
--	g3125 = DFF(g29259)
--	g3325 = DFF(g3321)
--	g3821 = DFF(g25681)
--	g4141 = DFF(g25687)
--	g4570 = DFF(g33617)
--	g5272 = DFF(g30479)
--	g2735 = DFF(g29256)
--	g728 = DFF(g28054)
--	g6295 = DFF(g30535)
--	g5417 = DFF(g28094)
--	g2661 = DFF(g30385)
--	g1988 = DFF(g30361)
--	g5128 = DFF(g25705)
--	g1548 = DFF(g24260)
--	g3106 = DFF(g29257)
--	g4659 = DFF(g34461)
--	g4358 = DFF(g34258)
--	g1792 = DFF(g32993)
--	g2084 = DFF(g33992)
--	g3061 = DFF(g28061)
--	g3187 = DFF(g30394)
--	g4311 = DFF(g34449)
--	g2583 = DFF(g34019)
--	g3003 = DFF(g21726)
--	g1094 = DFF(g29231)
--	g3841 = DFF(g25682)
--	g4284 = DFF(g21897)
--	g3763 = DFF(g28067)
--	g3191 = DFF(g30395)
--	g4239 = DFF(g21892)
--	g3391 = DFF(g31885)
--	g4180 = DFF(g4210)
--	g691 = DFF(g28048)
--	g534 = DFF(g34723)
--	g5366 = DFF(g25717)
--	g385 = DFF(g25598)
--	g2004 = DFF(g33987)
--	g2527 = DFF(g30380)
--	g5456 = DFF(g5448)
--	g4420 = DFF(g26965)
--	g5148 = DFF(g25706)
--	g4507 = DFF(g30458)
--	g5348 = DFF(g24338)
--	g3223 = DFF(g30400)
--	g4931 = DFF(g21904)
--	g2970 = DFF(g34623)
--	g5698 = DFF(g24343)
--	g3416 = DFF(g25666)
--	g5260 = DFF(g30473)
--	g1521 = DFF(g24252)
--	g3522 = DFF(g33028)
--	g3115 = DFF(g29258)
--	g3251 = DFF(g30407)
--	g1 = DFF(g26958)
--	g4628 = DFF(g34457)
--	g1996 = DFF(g33568)
--	g3447 = DFF(g25663)
--	g4515 = DFF(g26964)
--	g4204 = DFF(g4200)
--	g4300 = DFF(g34735)
--	g1724 = DFF(g30352)
--	g1379 = DFF(g33543)
--	g3654 = DFF(g24271)
--	g12 = DFF(g30326)
--	g1878 = DFF(g33981)
--	g5619 = DFF(g30500)
--	g71 = DFF(g34786)
--	g59 = DFF(g29277)
--	
--	I28349 = NOT(g28367)
--	g19408 = NOT(g16066)
--	I21294 = NOT(g18274)
--	g13297 = NOT(g10831)
--	g19635 = NOT(g16349)
--	g32394 = NOT(g30601)
--	I19778 = NOT(g17781)
--	g9900 = NOT(g6)
--	g11889 = NOT(g9954)
--	g13103 = NOT(g10905)
--	g17470 = NOT(g14454)
--	g23499 = NOT(g20785)
--	g6895 = NOT(g3288)
--	g9797 = NOT(g5441)
--	g31804 = NOT(g29385)
--	g6837 = NOT(g968)
--	I15824 = NOT(g1116)
--	g20066 = NOT(g17433)
--	g33804 = NOT(g33250)
--	g20231 = NOT(g17821)
--	I19786 = NOT(g17844)
--	g24066 = NOT(g21127)
--	g11888 = NOT(g10160)
--	g9510 = NOT(g5835)
--	I22692 = NOT(g21308)
--	g12884 = NOT(g10392)
--	g22494 = NOT(g19801)
--	g9245 = NOT(I13031)
--	g8925 = NOT(I12910)
--	g34248 = NOT(I32243)
--	g10289 = NOT(g1319)
--	g11181 = NOT(g8134)
--	I20116 = NOT(g15737)
--	g7888 = NOT(g1536)
--	g9291 = NOT(g3021)
--	g28559 = NOT(g27700)
--	g21056 = NOT(g15426)
--	I33246 = NOT(g34970)
--	g10288 = NOT(I13718)
--	g8224 = NOT(g3774)
--	g21611 = NOT(I21210)
--	g16718 = NOT(I17932)
--	g21722 = NOT(I21285)
--	I12530 = NOT(g4815)
--	g16521 = NOT(g13543)
--	I22400 = NOT(g19620)
--	g23611 = NOT(g18833)
--	g10571 = NOT(g10233)
--	g17467 = NOT(g14339)
--	g17494 = NOT(g14339)
--	g10308 = NOT(g4459)
--	g27015 = NOT(g26869)
--	g23988 = NOT(g19277)
--	g23924 = NOT(g18997)
--	g12217 = NOT(I15070)
--	g14571 = NOT(I16688)
--	g32318 = NOT(g31596)
--	g32446 = NOT(g31596)
--	g14308 = NOT(I16471)
--	I24041 = NOT(g22182)
--	I14935 = NOT(g9902)
--	g34778 = NOT(I32976)
--	g20511 = NOT(g17929)
--	g26672 = NOT(g25275)
--	g11931 = NOT(I14749)
--	g20763 = NOT(I20816)
--	g23432 = NOT(g21514)
--	I18165 = NOT(g13177)
--	I18523 = NOT(g14443)
--	g21271 = NOT(I21002)
--	I31776 = NOT(g33204)
--	g23271 = NOT(g20785)
--	g22155 = NOT(g19074)
--	I22539 = NOT(g19606)
--	I32231 = NOT(g34123)
--	g34786 = NOT(I32988)
--	g9259 = NOT(g5176)
--	I15190 = NOT(g6005)
--	g17782 = NOT(I18788)
--	g8277 = NOT(I12483)
--	g9819 = NOT(g92)
--	I16969 = NOT(g13943)
--	g32540 = NOT(g30614)
--	g25027 = NOT(I24191)
--	g19711 = NOT(g17062)
--	g22170 = NOT(g19210)
--	g13190 = NOT(g10939)
--	g7297 = NOT(g6069)
--	g17419 = NOT(g14965)
--	g20660 = NOT(g17873)
--	g16861 = NOT(I18051)
--	g21461 = NOT(g15348)
--	g10816 = NOT(I14054)
--	g28713 = NOT(g27907)
--	g15755 = NOT(g13134)
--	g23461 = NOT(g18833)
--	I24237 = NOT(g23823)
--	g34945 = NOT(g34933)
--	g8789 = NOT(I12779)
--	g31833 = NOT(g29385)
--	I18006 = NOT(g13638)
--	I20035 = NOT(g15706)
--	I17207 = NOT(g13835)
--	g30999 = NOT(g29722)
--	g25249 = NOT(g22228)
--	g9488 = NOT(g1878)
--	g19537 = NOT(g15938)
--	g17155 = NOT(I18205)
--	I16855 = NOT(g10473)
--	g15563 = NOT(I17140)
--	g23031 = NOT(g19801)
--	g30090 = NOT(g29134)
--	g30998 = NOT(g29719)
--	g25248 = NOT(g22228)
--	g23650 = NOT(g20653)
--	g7138 = NOT(g5360)
--	g16099 = NOT(g13437)
--	g34998 = NOT(g34981)
--	g23887 = NOT(g18997)
--	g25552 = NOT(g22594)
--	g20916 = NOT(g18008)
--	g27084 = NOT(g26673)
--	g30182 = NOT(I28419)
--	g7963 = NOT(g4146)
--	g10374 = NOT(g6903)
--	I32763 = NOT(g34511)
--	g19606 = NOT(g17614)
--	g19492 = NOT(g16349)
--	g22167 = NOT(g19074)
--	g22194 = NOT(I21776)
--	g7109 = NOT(g5011)
--	g7791 = NOT(I12199)
--	g34672 = NOT(I32800)
--	g16777 = NOT(I18003)
--	g20550 = NOT(g15864)
--	g23529 = NOT(g20558)
--	g6854 = NOT(g2685)
--	g18930 = NOT(g15789)
--	g13024 = NOT(g11900)
--	g32902 = NOT(g30673)
--	g6941 = NOT(g3990)
--	g12110 = NOT(I14970)
--	g32957 = NOT(g31672)
--	g9951 = NOT(g6133)
--	g32377 = NOT(g30984)
--	g12922 = NOT(g12297)
--	g23528 = NOT(g18833)
--	g12321 = NOT(g9637)
--	g28678 = NOT(g27800)
--	g32739 = NOT(g30735)
--	g21393 = NOT(g17264)
--	g23843 = NOT(g19147)
--	g26026 = NOT(I25105)
--	g25081 = NOT(g22342)
--	g20085 = NOT(g16187)
--	g23393 = NOT(g20739)
--	g19750 = NOT(g16326)
--	g30331 = NOT(I28594)
--	g24076 = NOT(g19984)
--	g24085 = NOT(g20857)
--	g17589 = NOT(g14981)
--	g20596 = NOT(I20690)
--	g34932 = NOT(g34914)
--	g23764 = NOT(g21308)
--	g25786 = NOT(g24518)
--	I25869 = NOT(g25851)
--	g32738 = NOT(g31376)
--	g32562 = NOT(g30673)
--	g32645 = NOT(g30825)
--	g14669 = NOT(g12301)
--	g20054 = NOT(g17328)
--	I26337 = NOT(g26835)
--	g24054 = NOT(g19919)
--	I20130 = NOT(g15748)
--	g17588 = NOT(g14782)
--	g17524 = NOT(g14933)
--	I18600 = NOT(g5335)
--	g23869 = NOT(g19277)
--	g32699 = NOT(g31528)
--	g10392 = NOT(g6989)
--	I28576 = NOT(g28431)
--	I28585 = NOT(g30217)
--	I15987 = NOT(g12381)
--	g14668 = NOT(g12450)
--	g25356 = NOT(g22763)
--	g24431 = NOT(g22722)
--	g29725 = NOT(g28349)
--	I15250 = NOT(g9152)
--	g28294 = NOT(g27295)
--	g8945 = NOT(g608)
--	g10489 = NOT(g9259)
--	g11987 = NOT(I14833)
--	g13625 = NOT(g10971)
--	I25161 = NOT(g24920)
--	g17477 = NOT(g14848)
--	g23868 = NOT(g19277)
--	g32698 = NOT(g30614)
--	g31812 = NOT(g29385)
--	g11250 = NOT(g7502)
--	g25380 = NOT(g23776)
--	I32550 = NOT(g34398)
--	g7957 = NOT(g1252)
--	g13250 = NOT(I15811)
--	g20269 = NOT(g15844)
--	g34505 = NOT(g34409)
--	g7049 = NOT(g5853)
--	g20773 = NOT(I20830)
--	g25090 = NOT(g23630)
--	g6958 = NOT(g4372)
--	g20268 = NOT(g18008)
--	g14424 = NOT(g11136)
--	g34717 = NOT(I32881)
--	g12417 = NOT(g7175)
--	g25182 = NOT(g22763)
--	g12936 = NOT(g12601)
--	g20655 = NOT(I20753)
--	g8340 = NOT(g3050)
--	g13943 = NOT(I16231)
--	g21225 = NOT(g17428)
--	g24156 = NOT(I23312)
--	g23259 = NOT(g21070)
--	g24655 = NOT(g23067)
--	I12109 = NOT(g749)
--	I18063 = NOT(g14357)
--	g7715 = NOT(g1178)
--	g29744 = NOT(g28431)
--	g8478 = NOT(g3103)
--	g20180 = NOT(g17533)
--	g17616 = NOT(g14309)
--	g20670 = NOT(g15426)
--	I29447 = NOT(g30729)
--	g10830 = NOT(g10087)
--	I32243 = NOT(g34134)
--	g22305 = NOT(g19801)
--	g24180 = NOT(I23384)
--	g32632 = NOT(g31070)
--	g31795 = NOT(I29371)
--	g9594 = NOT(g2307)
--	g6829 = NOT(g1319)
--	g7498 = NOT(g6675)
--	g23258 = NOT(g20924)
--	g26811 = NOT(g25206)
--	I16590 = NOT(g11966)
--	g10544 = NOT(I13906)
--	g15573 = NOT(I17154)
--	I27492 = NOT(g27511)
--	g9806 = NOT(g5782)
--	g14544 = NOT(I16663)
--	I14653 = NOT(g9417)
--	I33044 = NOT(g34775)
--	I16741 = NOT(g5677)
--	g25513 = NOT(g23870)
--	g32661 = NOT(g31070)
--	g20993 = NOT(g15615)
--	g32547 = NOT(g30614)
--	g32895 = NOT(g30673)
--	g8876 = NOT(I12855)
--	g24839 = NOT(g23436)
--	g23244 = NOT(I22343)
--	g24993 = NOT(g22384)
--	g22177 = NOT(g19074)
--	g16162 = NOT(g13437)
--	g11855 = NOT(I14671)
--	g20667 = NOT(g15224)
--	g17466 = NOT(g12983)
--	g9887 = NOT(g5802)
--	g6974 = NOT(I11746)
--	g24667 = NOT(g23112)
--	g9934 = NOT(g5849)
--	g21069 = NOT(g15277)
--	g25505 = NOT(g22228)
--	g34433 = NOT(I32470)
--	g34387 = NOT(g34188)
--	g10042 = NOT(g2671)
--	g24131 = NOT(g21209)
--	g32481 = NOT(g31194)
--	g14705 = NOT(I16803)
--	I13321 = NOT(g6486)
--	g18975 = NOT(g15938)
--	g19553 = NOT(g16782)
--	g19862 = NOT(I20233)
--	g30097 = NOT(g29118)
--	g8915 = NOT(I12884)
--	g16629 = NOT(g13990)
--	I16150 = NOT(g10430)
--	g21657 = NOT(g17657)
--	g16472 = NOT(g14098)
--	I20781 = NOT(g17155)
--	g21068 = NOT(g15277)
--	g14255 = NOT(g12381)
--	I21477 = NOT(g18695)
--	g14189 = NOT(I16391)
--	g32551 = NOT(g30735)
--	g32572 = NOT(g30735)
--	g23375 = NOT(g20924)
--	I24781 = NOT(g24264)
--	I33146 = NOT(g34903)
--	g7162 = NOT(g4521)
--	g25212 = NOT(g22763)
--	g7268 = NOT(g1636)
--	I11740 = NOT(g4519)
--	g7362 = NOT(g1906)
--	g12909 = NOT(g10412)
--	g9433 = NOT(g5148)
--	g26850 = NOT(I25576)
--	g12543 = NOT(g9417)
--	g17642 = NOT(g14691)
--	g20502 = NOT(g15373)
--	g10678 = NOT(I13990)
--	I22725 = NOT(g21250)
--	I13740 = NOT(g85)
--	g23879 = NOT(g19210)
--	g20557 = NOT(I20647)
--	g23970 = NOT(g19277)
--	g34343 = NOT(g34089)
--	g20210 = NOT(g16897)
--	I22114 = NOT(g19935)
--	g12908 = NOT(g10414)
--	g20618 = NOT(g15277)
--	g11867 = NOT(I14679)
--	g11894 = NOT(I14702)
--	I11685 = NOT(g117)
--	g8310 = NOT(g2051)
--	g23878 = NOT(g19147)
--	g21337 = NOT(g15758)
--	g20443 = NOT(g15171)
--	g10383 = NOT(g6978)
--	g23337 = NOT(g20924)
--	g19757 = NOT(g17224)
--	g9496 = NOT(g3303)
--	g14383 = NOT(I16535)
--	g17733 = NOT(g14238)
--	I16526 = NOT(g10430)
--	g8663 = NOT(g3343)
--	g10030 = NOT(g116)
--	g23886 = NOT(g21468)
--	I18614 = NOT(g6315)
--	g32490 = NOT(g30673)
--	g10093 = NOT(g5703)
--	g18884 = NOT(g15938)
--	g27242 = NOT(g26183)
--	I14576 = NOT(g8791)
--	g11714 = NOT(g8107)
--	g22166 = NOT(g18997)
--	g11450 = NOT(I14455)
--	I17114 = NOT(g14358)
--	I27192 = NOT(g27662)
--	g23792 = NOT(g19074)
--	g23967 = NOT(g19210)
--	g23994 = NOT(g19277)
--	g32784 = NOT(g31672)
--	g9891 = NOT(g6173)
--	I18320 = NOT(g13605)
--	g28037 = NOT(g26365)
--	g8002 = NOT(g1389)
--	g9337 = NOT(g1608)
--	g9913 = NOT(g2403)
--	g32956 = NOT(g30825)
--	I21285 = NOT(g18215)
--	g11819 = NOT(g7717)
--	g11910 = NOT(g10185)
--	g14065 = NOT(g11048)
--	g7086 = NOT(g4826)
--	g13707 = NOT(g11360)
--	g31829 = NOT(g29385)
--	g32889 = NOT(g31376)
--	g11202 = NOT(I14267)
--	g8236 = NOT(g4812)
--	g33920 = NOT(I31786)
--	I21254 = NOT(g16540)
--	g24039 = NOT(g21256)
--	g25620 = NOT(I24759)
--	g21425 = NOT(g15509)
--	g29221 = NOT(I27579)
--	I17744 = NOT(g14912)
--	g23459 = NOT(g21611)
--	I16917 = NOT(g10582)
--	g20038 = NOT(g17328)
--	g23425 = NOT(g20751)
--	g31828 = NOT(g29385)
--	g32888 = NOT(g30673)
--	I15070 = NOT(g10108)
--	g25097 = NOT(g22342)
--	g32824 = NOT(g31376)
--	g10219 = NOT(g2697)
--	g13055 = NOT(I15682)
--	g9807 = NOT(g5712)
--	I30901 = NOT(g32407)
--	g19673 = NOT(g16931)
--	g24038 = NOT(g21193)
--	g14219 = NOT(g12381)
--	g19397 = NOT(g16449)
--	g21458 = NOT(g15758)
--	g6849 = NOT(g2551)
--	I15590 = NOT(g11988)
--	g28155 = NOT(I26664)
--	I13762 = NOT(g6755)
--	g13070 = NOT(g11984)
--	g23458 = NOT(I22583)
--	g32671 = NOT(g31528)
--	I21036 = NOT(g17221)
--	g34229 = NOT(g33936)
--	g10218 = NOT(g2527)
--	I18034 = NOT(g13680)
--	g16172 = NOT(g13584)
--	g20601 = NOT(g17433)
--	g21010 = NOT(g15634)
--	g11986 = NOT(I14830)
--	g7470 = NOT(g5623)
--	I12483 = NOT(g3096)
--	g17476 = NOT(g14665)
--	g17485 = NOT(I18408)
--	I16077 = NOT(g10430)
--	I14745 = NOT(g10029)
--	g11741 = NOT(g10033)
--	g22907 = NOT(g20453)
--	g23545 = NOT(g21562)
--	g23444 = NOT(I22561)
--	g25369 = NOT(g22228)
--	g32931 = NOT(g30937)
--	g33682 = NOT(I31515)
--	g6900 = NOT(g3440)
--	g19634 = NOT(g16349)
--	g19872 = NOT(g17015)
--	g34716 = NOT(I32878)
--	I20542 = NOT(g16508)
--	I25598 = NOT(g25424)
--	g8928 = NOT(g4340)
--	g29812 = NOT(g28381)
--	I28241 = NOT(g28709)
--	g12841 = NOT(g10357)
--	g22594 = NOT(I21934)
--	I16688 = NOT(g10981)
--	g9815 = NOT(g6098)
--	g8064 = NOT(g3376)
--	I18408 = NOT(g13017)
--	I20913 = NOT(g16964)
--	g23086 = NOT(g20283)
--	I32815 = NOT(g34470)
--	g30310 = NOT(g28830)
--	g8899 = NOT(g807)
--	g11735 = NOT(g8534)
--	g29371 = NOT(I27735)
--	I11908 = NOT(g4449)
--	g9692 = NOT(g1756)
--	g13877 = NOT(g11350)
--	I32601 = NOT(g34319)
--	g8785 = NOT(I12767)
--	g24169 = NOT(I23351)
--	g24791 = NOT(g23850)
--	g9497 = NOT(I13166)
--	I16102 = NOT(g10430)
--	g26681 = NOT(g25396)
--	g20168 = NOT(g17533)
--	g9154 = NOT(I12994)
--	g25133 = NOT(g23733)
--	g34925 = NOT(I33167)
--	I26309 = NOT(g26825)
--	g9354 = NOT(g2719)
--	g27014 = NOT(g25888)
--	I27564 = NOT(g28166)
--	g24168 = NOT(I23348)
--	g23322 = NOT(I22425)
--	g32546 = NOT(g31170)
--	g9960 = NOT(g6474)
--	g22519 = NOT(g19801)
--	g22176 = NOT(g18997)
--	g14201 = NOT(I16401)
--	g26802 = NOT(I25514)
--	g28119 = NOT(g27008)
--	g12835 = NOT(g10352)
--	g7635 = NOT(g1002)
--	g14277 = NOT(I16455)
--	g20666 = NOT(g15224)
--	g13018 = NOT(I15636)
--	I16231 = NOT(g10520)
--	g32024 = NOT(I29582)
--	g25228 = NOT(g23828)
--	I19802 = NOT(g15727)
--	g19574 = NOT(g16826)
--	g7766 = NOT(I12189)
--	g19452 = NOT(g16326)
--	g6819 = NOT(g1046)
--	g16540 = NOT(I17744)
--	I19857 = NOT(g16640)
--	g22154 = NOT(g19074)
--	g7087 = NOT(g6336)
--	I33297 = NOT(g35000)
--	g25011 = NOT(g22763)
--	g32860 = NOT(g30673)
--	I18891 = NOT(g16676)
--	g7487 = NOT(g1259)
--	I33103 = NOT(g34846)
--	g8237 = NOT(g255)
--	g18953 = NOT(g16077)
--	I14761 = NOT(g7753)
--	g19912 = NOT(g17328)
--	g17519 = NOT(I18460)
--	g21561 = NOT(g15595)
--	I12183 = NOT(g2719)
--	g21656 = NOT(g17700)
--	g6923 = NOT(g3791)
--	g26765 = NOT(g25309)
--	I25680 = NOT(g25641)
--	g22935 = NOT(g20283)
--	g17092 = NOT(g14011)
--	g34944 = NOT(g34932)
--	g10037 = NOT(g1848)
--	I32791 = NOT(g34578)
--	g32497 = NOT(g30673)
--	g21295 = NOT(g17533)
--	g23353 = NOT(g20924)
--	g29507 = NOT(g28353)
--	I32884 = NOT(g34690)
--	g8844 = NOT(I12826)
--	g11402 = NOT(g7594)
--	g17518 = NOT(g14918)
--	g26549 = NOT(I25391)
--	g17154 = NOT(g14348)
--	g22883 = NOT(g20391)
--	g20556 = NOT(g15483)
--	g23823 = NOT(I22989)
--	g17637 = NOT(g12933)
--	g20580 = NOT(g17328)
--	g26548 = NOT(g25255)
--	g10419 = NOT(g8821)
--	g11866 = NOT(g9883)
--	g11917 = NOT(I14727)
--	g32700 = NOT(g31579)
--	I26687 = NOT(g27880)
--	g32659 = NOT(g30735)
--	g21336 = NOT(g17367)
--	g32625 = NOT(g31070)
--	g10352 = NOT(g6804)
--	g23336 = NOT(g20924)
--	I32479 = NOT(g34302)
--	g19592 = NOT(I20035)
--	g34429 = NOT(I32458)
--	g10155 = NOT(g2643)
--	g10418 = NOT(g8818)
--	g12041 = NOT(I14905)
--	g32658 = NOT(g31579)
--	g19780 = NOT(g16449)
--	g16739 = NOT(g13223)
--	g12430 = NOT(I15250)
--	I16660 = NOT(g10981)
--	g34428 = NOT(I32455)
--	I21074 = NOT(g17766)
--	g23966 = NOT(g19210)
--	g22215 = NOT(g19277)
--	g28036 = NOT(g26365)
--	g27237 = NOT(g26162)
--	g32943 = NOT(g31710)
--	g20110 = NOT(g16897)
--	g11706 = NOT(I14579)
--	g24084 = NOT(g20720)
--	g16738 = NOT(I17956)
--	g9761 = NOT(g2445)
--	g13706 = NOT(g11280)
--	g16645 = NOT(g13756)
--	g12465 = NOT(g7192)
--	I11992 = NOT(g763)
--	g24110 = NOT(g21209)
--	g20922 = NOT(I20891)
--	g27983 = NOT(g26725)
--	g20321 = NOT(g17821)
--	g23017 = NOT(g20453)
--	g32644 = NOT(g30735)
--	g33648 = NOT(I31482)
--	I21238 = NOT(g16540)
--	g34690 = NOT(I32840)
--	g6870 = NOT(g3089)
--	g9828 = NOT(g2024)
--	g20179 = NOT(g17249)
--	g34549 = NOT(I32617)
--	g8948 = NOT(g785)
--	g20531 = NOT(g15907)
--	g12983 = NOT(I15600)
--	g24179 = NOT(I23381)
--	g16290 = NOT(g13260)
--	g32969 = NOT(g30735)
--	g13280 = NOT(I15846)
--	g6825 = NOT(g979)
--	g33755 = NOT(I31610)
--	g17501 = NOT(I18434)
--	g7369 = NOT(g1996)
--	g27142 = NOT(g26105)
--	g8955 = NOT(g1418)
--	g20178 = NOT(g16971)
--	g10194 = NOT(g6741)
--	g19396 = NOT(g16431)
--	g17577 = NOT(I18504)
--	g13624 = NOT(g10951)
--	I14241 = NOT(g8356)
--	I21941 = NOT(g18918)
--	g24178 = NOT(I23378)
--	g14167 = NOT(I16371)
--	g32968 = NOT(g31376)
--	g19731 = NOT(g17093)
--	g29920 = NOT(g28824)
--	g34504 = NOT(g34408)
--	g29358 = NOT(I27718)
--	g7868 = NOT(g1099)
--	I15102 = NOT(g5313)
--	I26195 = NOT(g26260)
--	I11835 = NOT(g101)
--	I20891 = NOT(g17700)
--	g9746 = NOT(I13326)
--	g20373 = NOT(g17929)
--	g32855 = NOT(g30825)
--	g23289 = NOT(g20924)
--	g24685 = NOT(g23139)
--	g24373 = NOT(g22908)
--	I33024 = NOT(g34783)
--	g8150 = NOT(g2185)
--	g10401 = NOT(g7041)
--	g22906 = NOT(g20453)
--	g20654 = NOT(I20750)
--	I16596 = NOT(g12640)
--	g34317 = NOT(g34115)
--	g8350 = NOT(g4646)
--	g18908 = NOT(g16100)
--	g32870 = NOT(g31021)
--	g7535 = NOT(g1500)
--	g32527 = NOT(g30673)
--	I13007 = NOT(g65)
--	g8038 = NOT(I12360)
--	g10119 = NOT(g2841)
--	I24474 = NOT(g22546)
--	g16632 = NOT(g14454)
--	g21308 = NOT(g17485)
--	g8438 = NOT(g3100)
--	g23571 = NOT(g18833)
--	g28693 = NOT(g27837)
--	g23308 = NOT(g21024)
--	g31794 = NOT(I29368)
--	g6972 = NOT(I11740)
--	g31845 = NOT(g29385)
--	g8009 = NOT(g3106)
--	I31497 = NOT(g33187)
--	g7261 = NOT(g4449)
--	g24417 = NOT(g22171)
--	g33845 = NOT(I31694)
--	g10118 = NOT(g2541)
--	I19775 = NOT(g17780)
--	g9932 = NOT(g5805)
--	g28166 = NOT(I26687)
--	g28009 = NOT(I26516)
--	g16661 = NOT(g14454)
--	I17507 = NOT(g13416)
--	g25549 = NOT(g22763)
--	g13876 = NOT(g11432)
--	g13885 = NOT(g10862)
--	g32503 = NOT(g31194)
--	g23495 = NOT(I22622)
--	I31659 = NOT(g33219)
--	g14749 = NOT(I16829)
--	g32867 = NOT(g30673)
--	g32894 = NOT(g30614)
--	I31625 = NOT(g33197)
--	g14616 = NOT(I16733)
--	g34245 = NOT(I32234)
--	I32953 = NOT(g34656)
--	g8836 = NOT(g736)
--	g30299 = NOT(g28765)
--	g6887 = NOT(g3333)
--	g23816 = NOT(g21308)
--	g25548 = NOT(g22550)
--	g34323 = NOT(g34105)
--	g34299 = NOT(g34080)
--	I32654 = NOT(g34378)
--	g22139 = NOT(I21722)
--	g8918 = NOT(I12893)
--	g24964 = NOT(I24128)
--	g7246 = NOT(g4446)
--	I11746 = NOT(g4570)
--	g26856 = NOT(I25586)
--	g13763 = NOT(g10971)
--	g14276 = NOT(I16452)
--	g31521 = NOT(I29182)
--	I32800 = NOT(g34582)
--	g32581 = NOT(g31070)
--	g32714 = NOT(g31528)
--	g32450 = NOT(g31591)
--	g10053 = NOT(g6381)
--	g23985 = NOT(g19210)
--	g22138 = NOT(g21370)
--	g15739 = NOT(g13284)
--	I26705 = NOT(g27967)
--	g34775 = NOT(I32967)
--	I20750 = NOT(g16677)
--	g20587 = NOT(g15373)
--	g32707 = NOT(g31579)
--	g32819 = NOT(g30825)
--	g9576 = NOT(g6565)
--	g31832 = NOT(g29385)
--	I20982 = NOT(g16300)
--	g23954 = NOT(I23099)
--	g24587 = NOT(g23112)
--	g8229 = NOT(g3881)
--	g9716 = NOT(g5057)
--	I22788 = NOT(g18940)
--	I26679 = NOT(g27773)
--	g12863 = NOT(g10371)
--	g8993 = NOT(g385)
--	g15562 = NOT(g14943)
--	g32818 = NOT(g30735)
--	g10036 = NOT(g1816)
--	g32496 = NOT(g30614)
--	g19787 = NOT(g17096)
--	g16127 = NOT(g13437)
--	g8822 = NOT(g4975)
--	g10177 = NOT(g1834)
--	g20909 = NOT(g17955)
--	g20543 = NOT(g17955)
--	I13684 = NOT(g128)
--	g31861 = NOT(I29441)
--	g9848 = NOT(g4462)
--	g21669 = NOT(I21230)
--	g19357 = NOT(I19837)
--	g17415 = NOT(g14797)
--	g6845 = NOT(g2126)
--	g7502 = NOT(I11992)
--	I15550 = NOT(g10430)
--	g32590 = NOT(g31154)
--	g9699 = NOT(g2311)
--	g9747 = NOT(I13329)
--	g24117 = NOT(g21209)
--	g24000 = NOT(g19277)
--	I33197 = NOT(g34930)
--	g23260 = NOT(g21070)
--	g19743 = NOT(g17125)
--	I14584 = NOT(g9766)
--	g33926 = NOT(I31796)
--	g25245 = NOT(g22763)
--	g34697 = NOT(g34545)
--	g26831 = NOT(g24836)
--	g20569 = NOT(g15277)
--	I20840 = NOT(g17727)
--	g34995 = NOT(I33285)
--	g23842 = NOT(g19147)
--	g32741 = NOT(g31710)
--	g13314 = NOT(g10893)
--	I23348 = NOT(g23384)
--	g25299 = NOT(g22763)
--	g32384 = NOT(g31666)
--	I19831 = NOT(g16533)
--	g33388 = NOT(g32382)
--	I18252 = NOT(g13177)
--	I16502 = NOT(g10430)
--	g20568 = NOT(g15509)
--	g23489 = NOT(g21468)
--	g25533 = NOT(g22550)
--	g13085 = NOT(I15717)
--	g19769 = NOT(g16987)
--	g24568 = NOT(g22942)
--	g20242 = NOT(g16308)
--	g25298 = NOT(g23760)
--	g11721 = NOT(g10074)
--	g7689 = NOT(I12159)
--	g29927 = NOT(g28861)
--	I17121 = NOT(g14366)
--	g34512 = NOT(g34420)
--	g21424 = NOT(g15426)
--	g23559 = NOT(g21070)
--	g13596 = NOT(g10971)
--	g23525 = NOT(g21562)
--	g23488 = NOT(g21468)
--	g28675 = NOT(g27779)
--	g23016 = NOT(g20453)
--	I32909 = NOT(g34712)
--	g7216 = NOT(g822)
--	g11431 = NOT(g7618)
--	g12952 = NOT(I15572)
--	g23558 = NOT(g20924)
--	g13431 = NOT(I15932)
--	g32801 = NOT(g30937)
--	g14630 = NOT(g12402)
--	g32735 = NOT(g31021)
--	g24123 = NOT(g21143)
--	g32877 = NOT(g30825)
--	g7028 = NOT(I11785)
--	I30686 = NOT(g32381)
--	g8895 = NOT(g599)
--	g10166 = NOT(g6040)
--	g17576 = NOT(g14953)
--	g17585 = NOT(g14974)
--	g20772 = NOT(g15171)
--	g9644 = NOT(g2016)
--	g22200 = NOT(g19277)
--	g23893 = NOT(g19074)
--	I15773 = NOT(g10430)
--	g11269 = NOT(g7516)
--	I15942 = NOT(g12381)
--	g14166 = NOT(g11048)
--	g8620 = NOT(g3065)
--	g19881 = NOT(g15915)
--	g8462 = NOT(g1183)
--	g25232 = NOT(g22228)
--	g29491 = NOT(I27777)
--	g7247 = NOT(g5377)
--	g20639 = NOT(g15224)
--	I17173 = NOT(g13716)
--	g16931 = NOT(I18101)
--	I16468 = NOT(g12760)
--	g23544 = NOT(g21562)
--	g23865 = NOT(g21308)
--	I12046 = NOT(g613)
--	g32695 = NOT(g30735)
--	I31581 = NOT(g33164)
--	g11268 = NOT(g7515)
--	g20230 = NOT(I20499)
--	g12790 = NOT(g7097)
--	g17609 = NOT(g14817)
--	g29755 = NOT(I28002)
--	g7564 = NOT(g336)
--	g9152 = NOT(g2834)
--	g20638 = NOT(g15224)
--	I18509 = NOT(g5623)
--	g9818 = NOT(g6490)
--	g13655 = NOT(g10573)
--	g34316 = NOT(g34093)
--	g17200 = NOT(I18238)
--	g32526 = NOT(g30614)
--	g20265 = NOT(g17821)
--	g29981 = NOT(g28942)
--	g6815 = NOT(g929)
--	I12787 = NOT(g4311)
--	g12873 = NOT(g10380)
--	I22028 = NOT(g20204)
--	I29211 = NOT(g30298)
--	g8788 = NOT(I12776)
--	I18872 = NOT(g13745)
--	I23333 = NOT(g22683)
--	g30989 = NOT(g29672)
--	g33766 = NOT(I31619)
--	g19662 = NOT(g17432)
--	g21610 = NOT(g15615)
--	g14454 = NOT(I16613)
--	g23610 = NOT(g18833)
--	g10570 = NOT(g9021)
--	g34989 = NOT(I33267)
--	g8249 = NOT(g1917)
--	g20391 = NOT(I20562)
--	g32457 = NOT(g30735)
--	g21189 = NOT(g15634)
--	g24992 = NOT(g22417)
--	I33070 = NOT(g34810)
--	g20510 = NOT(g17226)
--	g23189 = NOT(g20060)
--	g11930 = NOT(g9281)
--	g12422 = NOT(I15238)
--	g26736 = NOT(g25349)
--	g9186 = NOT(I13010)
--	g17745 = NOT(g14978)
--	g34988 = NOT(I33264)
--	g22973 = NOT(g20330)
--	g34924 = NOT(I33164)
--	g6960 = NOT(g1)
--	g9386 = NOT(g5727)
--	I15667 = NOT(g12143)
--	I32639 = NOT(g34345)
--	g21270 = NOT(I20999)
--	g32866 = NOT(g30614)
--	g32917 = NOT(g30937)
--	g23270 = NOT(g20785)
--	g19482 = NOT(g16349)
--	g21678 = NOT(g16540)
--	g17813 = NOT(I18813)
--	g12834 = NOT(g10349)
--	g20579 = NOT(g17249)
--	g34432 = NOT(I32467)
--	g7308 = NOT(g1668)
--	g11965 = NOT(I14797)
--	g8085 = NOT(I12382)
--	g9599 = NOT(g3310)
--	g10074 = NOT(g718)
--	g19710 = NOT(g17059)
--	g18983 = NOT(g16077)
--	g24579 = NOT(g23067)
--	g34271 = NOT(g34160)
--	g19552 = NOT(g16856)
--	g21460 = NOT(g15628)
--	g21686 = NOT(g16540)
--	g9274 = NOT(g5857)
--	g20578 = NOT(g15563)
--	g26843 = NOT(I25567)
--	g23460 = NOT(g21611)
--	g23939 = NOT(g19074)
--	g21383 = NOT(g17367)
--	g19779 = NOT(g16431)
--	I19843 = NOT(g16594)
--	g9614 = NOT(g5128)
--	I33067 = NOT(g34812)
--	g17674 = NOT(I18647)
--	g12021 = NOT(g9543)
--	g14238 = NOT(g10823)
--	g20586 = NOT(g15171)
--	g23030 = NOT(g20453)
--	g32706 = NOT(g30673)
--	g23938 = NOT(g18997)
--	g32597 = NOT(g31154)
--	I18574 = NOT(g13075)
--	g25316 = NOT(g22763)
--	g8854 = NOT(g613)
--	g21267 = NOT(g15680)
--	g24586 = NOT(g23067)
--	I32391 = NOT(g34153)
--	g23267 = NOT(g20097)
--	g9821 = NOT(g115)
--	I13236 = NOT(g5452)
--	I18205 = NOT(g14563)
--	g34145 = NOT(I32096)
--	I16168 = NOT(g3321)
--	g26869 = NOT(g24842)
--	g32689 = NOT(g30825)
--	g15824 = NOT(I17324)
--	g20442 = NOT(g15171)
--	g10382 = NOT(g6958)
--	I18912 = NOT(g15050)
--	I22240 = NOT(g20086)
--	g32923 = NOT(g31021)
--	g33451 = NOT(g32132)
--	g19786 = NOT(g17062)
--	I14833 = NOT(g10142)
--	g16659 = NOT(I17857)
--	g12614 = NOT(g9935)
--	g22761 = NOT(g21024)
--	g9280 = NOT(I13054)
--	g10519 = NOT(g9326)
--	g34736 = NOT(I32904)
--	g10176 = NOT(g44)
--	I16479 = NOT(g10430)
--	g27320 = NOT(I26004)
--	g16987 = NOT(I18135)
--	g32688 = NOT(g30735)
--	g32624 = NOT(g30825)
--	I23312 = NOT(g21681)
--	g13279 = NOT(I15843)
--	I16217 = NOT(g3632)
--	I21115 = NOT(g15714)
--	g16658 = NOT(g14157)
--	I22604 = NOT(g21143)
--	g10518 = NOT(g9311)
--	g10154 = NOT(g2547)
--	g12905 = NOT(g10408)
--	g20615 = NOT(g15509)
--	g33246 = NOT(g32212)
--	g9083 = NOT(g626)
--	g23875 = NOT(g18997)
--	g25080 = NOT(g23742)
--	g24116 = NOT(g21143)
--	g14518 = NOT(I16639)
--	g23219 = NOT(I22316)
--	I18051 = NOT(g13680)
--	g30330 = NOT(I28591)
--	g13278 = NOT(g10738)
--	g26709 = NOT(g25435)
--	I29969 = NOT(g30991)
--	g8219 = NOT(g3731)
--	g27565 = NOT(g26645)
--	I17491 = NOT(g13416)
--	I16486 = NOT(g11204)
--	g20041 = NOT(g15569)
--	g9636 = NOT(g72)
--	g22214 = NOT(g19210)
--	g7827 = NOT(g4688)
--	g12122 = NOT(g9705)
--	g20275 = NOT(g17929)
--	g24041 = NOT(g19968)
--	g19998 = NOT(g15915)
--	g8431 = NOT(g3085)
--	g11468 = NOT(g7624)
--	g16644 = NOT(I17842)
--	g13039 = NOT(I15663)
--	g8812 = NOT(I12805)
--	g15426 = NOT(I17121)
--	g22207 = NOT(I21787)
--	g6828 = NOT(g1300)
--	g19672 = NOT(g16931)
--	g34132 = NOT(g33831)
--	g17400 = NOT(I18333)
--	I12890 = NOT(g4219)
--	g29045 = NOT(g27779)
--	g34960 = NOT(I33218)
--	g11038 = NOT(g8632)
--	g16969 = NOT(g14262)
--	g6830 = NOT(g1389)
--	g17013 = NOT(g14262)
--	I18350 = NOT(g13716)
--	g8005 = NOT(g3025)
--	g20237 = NOT(g17213)
--	g21160 = NOT(g17508)
--	g7196 = NOT(I11860)
--	g11815 = NOT(g7582)
--	g8405 = NOT(I12572)
--	g9187 = NOT(g518)
--	g16968 = NOT(g14238)
--	I27552 = NOT(g28162)
--	I15677 = NOT(g5654)
--	g31859 = NOT(g29385)
--	I32116 = NOT(g33937)
--	g20035 = NOT(g16430)
--	g31825 = NOT(g29385)
--	g32876 = NOT(g30735)
--	g32885 = NOT(g31021)
--	g34161 = NOT(g33851)
--	g16197 = NOT(g13861)
--	g24035 = NOT(g20841)
--	g11677 = NOT(g7689)
--	g21455 = NOT(g15426)
--	I12003 = NOT(g767)
--	g8286 = NOT(g53)
--	g8765 = NOT(g3333)
--	g17328 = NOT(I18313)
--	g31858 = NOT(g29385)
--	g13975 = NOT(g11048)
--	g32854 = NOT(g30735)
--	g7780 = NOT(g2878)
--	I12779 = NOT(g4210)
--	g16527 = NOT(g14048)
--	g25198 = NOT(g22228)
--	g30259 = NOT(g28463)
--	g25529 = NOT(g22763)
--	g14215 = NOT(g12198)
--	g32511 = NOT(g30614)
--	g23915 = NOT(g19277)
--	g32763 = NOT(g31710)
--	I15937 = NOT(g11676)
--	I17395 = NOT(g12952)
--	I28434 = NOT(g28114)
--	g30087 = NOT(g29121)
--	g11143 = NOT(g8032)
--	g19961 = NOT(g17328)
--	g26810 = NOT(g25220)
--	I29894 = NOT(g31771)
--	I14033 = NOT(g8912)
--	g34471 = NOT(g34423)
--	g9200 = NOT(g1548)
--	g25528 = NOT(g22594)
--	I21934 = NOT(g21273)
--	g31844 = NOT(g29385)
--	I31597 = NOT(g33187)
--	g8733 = NOT(g3698)
--	g19505 = NOT(g16349)
--	g23277 = NOT(I22380)
--	g7018 = NOT(g5297)
--	g8974 = NOT(I12930)
--	I11726 = NOT(g4273)
--	I32237 = NOT(g34130)
--	I17633 = NOT(g13258)
--	g32660 = NOT(g30825)
--	g7418 = NOT(g2361)
--	I13726 = NOT(g4537)
--	g9003 = NOT(g790)
--	g6953 = NOT(g4157)
--	g7994 = NOT(I12336)
--	g29997 = NOT(g29060)
--	g11884 = NOT(g8125)
--	g21467 = NOT(g15758)
--	I16676 = NOT(g10588)
--	g25869 = NOT(g25250)
--	g10349 = NOT(g6956)
--	g23494 = NOT(I22619)
--	g26337 = NOT(g24818)
--	I32806 = NOT(g34585)
--	g8796 = NOT(g4785)
--	I32684 = NOT(g34430)
--	g32456 = NOT(g31376)
--	g34244 = NOT(I32231)
--	I33300 = NOT(g35001)
--	g20130 = NOT(g17328)
--	g22683 = NOT(I22000)
--	g13410 = NOT(I15921)
--	I12826 = NOT(g4349)
--	g21037 = NOT(I20913)
--	g24130 = NOT(g20998)
--	g32480 = NOT(g31070)
--	g10083 = NOT(g2407)
--	g10348 = NOT(I13762)
--	g32916 = NOT(g31021)
--	g14348 = NOT(g10887)
--	g12891 = NOT(g10399)
--	g8324 = NOT(g2476)
--	g26792 = NOT(g25439)
--	g20523 = NOT(g17821)
--	I16417 = NOT(g875)
--	I21013 = NOT(g15806)
--	g32550 = NOT(g31376)
--	g9637 = NOT(I13252)
--	g23984 = NOT(g19210)
--	g18952 = NOT(g16053)
--	g24165 = NOT(I23339)
--	g30068 = NOT(g29157)
--	g34810 = NOT(I33020)
--	g31227 = NOT(g29744)
--	g17683 = NOT(g15027)
--	g23419 = NOT(g21468)
--	g34068 = NOT(g33728)
--	g21352 = NOT(g16322)
--	g13015 = NOT(g11875)
--	g8540 = NOT(g3408)
--	g23352 = NOT(g20924)
--	g25259 = NOT(I24445)
--	g25225 = NOT(g23802)
--	g21155 = NOT(g15656)
--	g34879 = NOT(I33109)
--	g21418 = NOT(g17821)
--	g22882 = NOT(g20391)
--	g28608 = NOT(g27670)
--	g23418 = NOT(g21468)
--	g32721 = NOT(g31021)
--	g20006 = NOT(g17328)
--	I26466 = NOT(g26870)
--	I15556 = NOT(g11928)
--	g32596 = NOT(g31070)
--	g9223 = NOT(g1216)
--	g12109 = NOT(I14967)
--	g19433 = NOT(g15915)
--	g23170 = NOT(g20046)
--	g7197 = NOT(g812)
--	g22407 = NOT(g19455)
--	g34878 = NOT(I33106)
--	g19387 = NOT(g16431)
--	I16762 = NOT(g5290)
--	g6848 = NOT(g2417)
--	g7397 = NOT(g890)
--	I27449 = NOT(g27737)
--	g15969 = NOT(I17416)
--	I20846 = NOT(g16923)
--	g19620 = NOT(g17296)
--	g12108 = NOT(I14964)
--	g10139 = NOT(g136)
--	I15223 = NOT(g10119)
--	I17612 = NOT(g13250)
--	I24396 = NOT(g23453)
--	g6855 = NOT(g2711)
--	g17414 = NOT(g14627)
--	g27492 = NOT(g26598)
--	g8287 = NOT(g160)
--	I17324 = NOT(g14119)
--	g9416 = NOT(g2429)
--	g13223 = NOT(I15800)
--	g24437 = NOT(g22654)
--	g25244 = NOT(g23802)
--	g19343 = NOT(g16136)
--	g34994 = NOT(I33282)
--	I17098 = NOT(g14336)
--	g32773 = NOT(g31376)
--	g32942 = NOT(g30825)
--	g9251 = NOT(I13037)
--	g20703 = NOT(g15373)
--	g29220 = NOT(I27576)
--	I11635 = NOT(g9)
--	g23589 = NOT(g21468)
--	g10415 = NOT(g7109)
--	g18422 = NOT(I19238)
--	g32655 = NOT(g30614)
--	g8399 = NOT(g3798)
--	g11110 = NOT(g8728)
--	g29911 = NOT(g28780)
--	g19369 = NOT(g15995)
--	g33377 = NOT(I30901)
--	g34425 = NOT(I32446)
--	g12381 = NOT(I15223)
--	g23524 = NOT(g21562)
--	g27091 = NOT(g26725)
--	g28184 = NOT(I26705)
--	g32670 = NOT(g30673)
--	g33120 = NOT(I30686)
--	I12026 = NOT(g344)
--	I21100 = NOT(g16284)
--	g8898 = NOT(g676)
--	g20600 = NOT(g15348)
--	I16117 = NOT(g10430)
--	g34919 = NOT(I33149)
--	g19368 = NOT(g16326)
--	I32222 = NOT(g34118)
--	g20781 = NOT(I20840)
--	g16877 = NOT(I18071)
--	g23477 = NOT(g21468)
--	g32734 = NOT(g31710)
--	g33645 = NOT(I31477)
--	g22759 = NOT(g19857)
--	I17140 = NOT(g13835)
--	g26817 = NOT(g25242)
--	g7631 = NOT(g74)
--	g34918 = NOT(I33146)
--	g17584 = NOT(g14773)
--	I26693 = NOT(g27930)
--	g10664 = NOT(g8928)
--	I20929 = NOT(g17663)
--	g32839 = NOT(g30735)
--	g32930 = NOT(g31021)
--	g20372 = NOT(g17847)
--	g30079 = NOT(g29097)
--	g19412 = NOT(g16489)
--	g7257 = NOT(I11903)
--	g22758 = NOT(g20330)
--	g24372 = NOT(g22885)
--	g16695 = NOT(g14454)
--	g25171 = NOT(g22228)
--	g20175 = NOT(I20433)
--	g7301 = NOT(g925)
--	I16747 = NOT(g12729)
--	g8291 = NOT(I12503)
--	g11373 = NOT(g7566)
--	g23864 = NOT(g19210)
--	g25886 = NOT(g24537)
--	g23022 = NOT(g20283)
--	g32667 = NOT(g30825)
--	g32694 = NOT(g31376)
--	g32838 = NOT(g31376)
--	I31550 = NOT(g33204)
--	g33698 = NOT(I31539)
--	g24175 = NOT(I23369)
--	g29147 = NOT(I27449)
--	g32965 = NOT(g31710)
--	g12840 = NOT(g10356)
--	g6818 = NOT(g976)
--	g17759 = NOT(g14864)
--	g6867 = NOT(I11685)
--	g16526 = NOT(g13898)
--	g23749 = NOT(g18997)
--	I15800 = NOT(g11607)
--	g15714 = NOT(I17228)
--	g9880 = NOT(g5787)
--	g23313 = NOT(g21070)
--	g25994 = NOT(g24575)
--	g8344 = NOT(I12523)
--	g9537 = NOT(g1748)
--	g29950 = NOT(g28896)
--	g24063 = NOT(g20014)
--	g17758 = NOT(g14861)
--	g26656 = NOT(g25495)
--	g20516 = NOT(I20609)
--	g10554 = NOT(g8974)
--	g18905 = NOT(g16077)
--	g24137 = NOT(g20998)
--	g32487 = NOT(g30825)
--	g24516 = NOT(g22670)
--	g7751 = NOT(g1521)
--	g23285 = NOT(g20887)
--	g26680 = NOT(g25300)
--	g32619 = NOT(g30614)
--	g8259 = NOT(g2217)
--	g21305 = NOT(g15758)
--	g21053 = NOT(g15373)
--	g32502 = NOT(g31070)
--	g14609 = NOT(I16724)
--	g15979 = NOT(I17420)
--	g10200 = NOT(g2138)
--	g23305 = NOT(g20391)
--	g32557 = NOT(g31376)
--	g13334 = NOT(g11048)
--	g29151 = NOT(g27858)
--	g29172 = NOT(g27020)
--	I24787 = NOT(g24266)
--	g9978 = NOT(g2756)
--	g30322 = NOT(g28431)
--	g10608 = NOT(g9155)
--	g29996 = NOT(g28962)
--	I12811 = NOT(g4340)
--	g10115 = NOT(g2283)
--	I16639 = NOT(g4000)
--	g21466 = NOT(g15509)
--	g32618 = NOT(g31154)
--	I18662 = NOT(g6322)
--	g8088 = NOT(g1554)
--	g6975 = NOT(g4507)
--	g9417 = NOT(I13124)
--	g34159 = NOT(I32116)
--	g11762 = NOT(g7964)
--	g7041 = NOT(g5644)
--	g9935 = NOT(I13483)
--	I13606 = NOT(g74)
--	g11964 = NOT(g9154)
--	g21036 = NOT(I20910)
--	g7441 = NOT(g862)
--	g20209 = NOT(g17821)
--	g33661 = NOT(I31497)
--	g33895 = NOT(I31751)
--	g9982 = NOT(g3976)
--	g21177 = NOT(I20957)
--	g21560 = NOT(g17873)
--	g16077 = NOT(I17456)
--	g9234 = NOT(g5170)
--	I15587 = NOT(g11985)
--	g32469 = NOT(g30673)
--	I27368 = NOT(g27881)
--	I18482 = NOT(g13350)
--	g20208 = NOT(g17533)
--	g14745 = NOT(g12423)
--	g13216 = NOT(g10939)
--	g17141 = NOT(I18191)
--	I11750 = NOT(g4474)
--	I18248 = NOT(g12938)
--	g19379 = NOT(g17327)
--	g26631 = NOT(g25467)
--	g12862 = NOT(g10370)
--	g17652 = NOT(g15033)
--	g34656 = NOT(I32770)
--	g8215 = NOT(I12451)
--	g30295 = NOT(I28540)
--	g22332 = NOT(I21838)
--	g9542 = NOT(g2173)
--	I16391 = NOT(g859)
--	g26364 = NOT(I25327)
--	g32468 = NOT(g30614)
--	g6821 = NOT(I11655)
--	I18003 = NOT(g13638)
--	g19050 = NOT(I19759)
--	g34680 = NOT(I32820)
--	g8951 = NOT(g554)
--	g16689 = NOT(g13923)
--	g34144 = NOT(I32093)
--	g34823 = NOT(I33037)
--	g20542 = NOT(g17873)
--	g16923 = NOT(I18089)
--	g20453 = NOT(I20584)
--	g16280 = NOT(g13330)
--	g6984 = NOT(g4709)
--	g32038 = NOT(g30934)
--	g24021 = NOT(g20841)
--	g28241 = NOT(g27064)
--	g29318 = NOT(g29029)
--	g16688 = NOT(g14045)
--	g16624 = NOT(I17814)
--	g22406 = NOT(g19506)
--	g8114 = NOT(g3522)
--	g10184 = NOT(g4486)
--	g12040 = NOT(I14902)
--	I16579 = NOT(g10981)
--	g16300 = NOT(I17626)
--	g19386 = NOT(g16431)
--	g10805 = NOT(I14046)
--	I22785 = NOT(g18940)
--	g20913 = NOT(g15373)
--	I18778 = NOT(g6704)
--	g34336 = NOT(g34112)
--	g32815 = NOT(g30937)
--	g14184 = NOT(g12381)
--	g19603 = NOT(g16349)
--	g19742 = NOT(g17096)
--	g13117 = NOT(g10981)
--	g17135 = NOT(g14297)
--	g12904 = NOT(g10410)
--	g20614 = NOT(g15426)
--	g32601 = NOT(g31376)
--	I15569 = NOT(g11965)
--	g9554 = NOT(g5105)
--	g20436 = NOT(I20569)
--	g23874 = NOT(g18997)
--	g8870 = NOT(I12837)
--	g32677 = NOT(g30673)
--	g33127 = NOT(g31950)
--	g25322 = NOT(I24497)
--	I31694 = NOT(g33176)
--	I32834 = NOT(g34472)
--	g32975 = NOT(I30537)
--	g21693 = NOT(I21254)
--	g20607 = NOT(g17955)
--	g13569 = NOT(g10951)
--	g8650 = NOT(g4664)
--	I12896 = NOT(g4229)
--	g20320 = NOT(g17015)
--	I18647 = NOT(g5320)
--	g20073 = NOT(g16540)
--	I28832 = NOT(g30301)
--	I33131 = NOT(g34906)
--	g30017 = NOT(g29085)
--	g20274 = NOT(g17847)
--	g9213 = NOT(I13020)
--	g24073 = NOT(g21127)
--	g20530 = NOT(g15509)
--	g21665 = NOT(I21226)
--	g25158 = NOT(g22228)
--	I21744 = NOT(g19338)
--	g20593 = NOT(g15277)
--	I17754 = NOT(g13494)
--	g23665 = NOT(g21562)
--	g25783 = NOT(g25250)
--	I17355 = NOT(g14591)
--	g32937 = NOT(g31021)
--	g19429 = NOT(g16489)
--	I23345 = NOT(g23320)
--	g33385 = NOT(g32038)
--	I21849 = NOT(g19620)
--	g29044 = NOT(g27742)
--	g10761 = NOT(g8411)
--	g7411 = NOT(g2040)
--	g25561 = NOT(g22550)
--	g18891 = NOT(g16053)
--	g20565 = NOT(g18008)
--	I31619 = NOT(g33212)
--	I15814 = NOT(g11129)
--	g24122 = NOT(g20857)
--	I23399 = NOT(g23450)
--	g8136 = NOT(g269)
--	g19730 = NOT(g17062)
--	g19428 = NOT(g16090)
--	g12183 = NOT(I15033)
--	g9902 = NOT(g100)
--	I18233 = NOT(g14639)
--	g33354 = NOT(g32329)
--	I33210 = NOT(g34943)
--	g32791 = NOT(g31672)
--	g23476 = NOT(g21468)
--	g23485 = NOT(g20785)
--	I25555 = NOT(g25241)
--	g31824 = NOT(g29385)
--	g32884 = NOT(g30825)
--	g33888 = NOT(g33346)
--	g8594 = NOT(g3849)
--	g19765 = NOT(g16897)
--	g6756 = NOT(I11623)
--	g24034 = NOT(g19968)
--	g7074 = NOT(I11801)
--	g11772 = NOT(I14623)
--	g10400 = NOT(g7002)
--	g20641 = NOT(g15509)
--	g26816 = NOT(g25260)
--	g21454 = NOT(g15373)
--	I33279 = NOT(g34986)
--	g23555 = NOT(I22692)
--	I32607 = NOT(g34358)
--	g7474 = NOT(I11980)
--	g17221 = NOT(I18245)
--	g19690 = NOT(g16826)
--	g30309 = NOT(g28959)
--	g7992 = NOT(g5008)
--	g9490 = NOT(g2563)
--	I14563 = NOT(g802)
--	g16511 = NOT(g14130)
--	g9166 = NOT(g837)
--	g20153 = NOT(g16782)
--	g23570 = NOT(g18833)
--	I32274 = NOT(g34195)
--	g23914 = NOT(g19210)
--	g32479 = NOT(g30735)
--	g32666 = NOT(g31376)
--	I13483 = NOT(g6035)
--	g11293 = NOT(g7527)
--	g24153 = NOT(I23303)
--	I31469 = NOT(g33388)
--	g6904 = NOT(g3494)
--	g32363 = NOT(I29891)
--	I12112 = NOT(g794)
--	g12872 = NOT(g10379)
--	g13638 = NOT(I16057)
--	g34308 = NOT(g34088)
--	g9056 = NOT(g3017)
--	g23907 = NOT(g19074)
--	g32478 = NOT(g31376)
--	g32015 = NOT(I29571)
--	g19504 = NOT(g16349)
--	g9456 = NOT(g6073)
--	g33931 = NOT(I31807)
--	I32464 = NOT(g34245)
--	g8228 = NOT(g3835)
--	g9529 = NOT(g6561)
--	g7863 = NOT(g1249)
--	g20136 = NOT(I20399)
--	g20635 = NOT(g18008)
--	I27742 = NOT(g28819)
--	g13416 = NOT(I15929)
--	g25017 = NOT(g23699)
--	I25567 = NOT(g25272)
--	I25594 = NOT(g25531)
--	I18897 = NOT(g16738)
--	g24136 = NOT(g20857)
--	g32486 = NOT(g30735)
--	I13326 = NOT(g66)
--	g23239 = NOT(g21308)
--	g33426 = NOT(g32017)
--	g11841 = NOT(g9800)
--	g9155 = NOT(I12997)
--	I14395 = NOT(g3654)
--	g6841 = NOT(g2145)
--	I17420 = NOT(g13394)
--	g23567 = NOT(g21562)
--	g32556 = NOT(g31554)
--	I32797 = NOT(g34581)
--	I14899 = NOT(g10198)
--	g8033 = NOT(g157)
--	g23238 = NOT(g20924)
--	g11510 = NOT(g7633)
--	g13510 = NOT(I15981)
--	g17812 = NOT(I18810)
--	g34816 = NOT(I33030)
--	I20647 = NOT(g17010)
--	g32580 = NOT(g30825)
--	g9698 = NOT(g2181)
--	g28441 = NOT(g27629)
--	g26260 = NOT(g24759)
--	I14633 = NOT(g9340)
--	g9964 = NOT(g126)
--	I13252 = NOT(g6751)
--	g20164 = NOT(g16826)
--	g34985 = NOT(I33255)
--	I20999 = NOT(g16709)
--	g23941 = NOT(g19074)
--	g18091 = NOT(I18879)
--	g19128 = NOT(I19778)
--	g23382 = NOT(g20682)
--	g24164 = NOT(I23336)
--	g25289 = NOT(g22228)
--	g21176 = NOT(I20954)
--	g21185 = NOT(g15277)
--	g23519 = NOT(g21468)
--	I27730 = NOT(g28752)
--	g12047 = NOT(g9591)
--	g16307 = NOT(I17633)
--	g13835 = NOT(I16150)
--	g34954 = NOT(I33210)
--	g13014 = NOT(g11872)
--	g25023 = NOT(g22457)
--	g24891 = NOT(g23231)
--	I33143 = NOT(g34903)
--	g19626 = NOT(g17409)
--	g25288 = NOT(g22228)
--	g25224 = NOT(g22763)
--	I20233 = NOT(g17487)
--	g16721 = NOT(g14072)
--	I12793 = NOT(g4578)
--	g23518 = NOT(g21070)
--	g23154 = NOT(I22264)
--	g26488 = NOT(I25366)
--	g26424 = NOT(I25356)
--	g20575 = NOT(g17929)
--	g31860 = NOT(I29438)
--	g13007 = NOT(g11852)
--	g25308 = NOT(g22763)
--	g8195 = NOT(g1783)
--	g8137 = NOT(g411)
--	g32922 = NOT(g31710)
--	g8891 = NOT(g582)
--	g19533 = NOT(g16261)
--	g24474 = NOT(g23620)
--	g20711 = NOT(g15509)
--	I16193 = NOT(g3281)
--	g16431 = NOT(I17675)
--	I27549 = NOT(g28161)
--	g27051 = NOT(I25779)
--	g32531 = NOT(g31070)
--	I13847 = NOT(g7266)
--	I31791 = NOT(g33354)
--	g20327 = NOT(g15224)
--	g23935 = NOT(g19210)
--	g24711 = NOT(g23139)
--	g34669 = NOT(I32791)
--	g26830 = NOT(g24411)
--	g27592 = NOT(g26715)
--	g12051 = NOT(g9595)
--	g20537 = NOT(g15345)
--	g24109 = NOT(g21143)
--	g32740 = NOT(g31672)
--	g15885 = NOT(I17374)
--	g8807 = NOT(g79)
--	g11615 = NOT(g6875)
--	g9619 = NOT(g5845)
--	g17507 = NOT(g15030)
--	I24331 = NOT(g22976)
--	g34668 = NOT(I32788)
--	g13116 = NOT(g10935)
--	g16773 = NOT(g14021)
--	I18148 = NOT(g13526)
--	g24108 = NOT(g20998)
--	I28162 = NOT(g28803)
--	g32186 = NOT(I29720)
--	g34392 = NOT(g34202)
--	g32676 = NOT(g30614)
--	g32685 = NOT(g31528)
--	g33659 = NOT(I31491)
--	g28399 = NOT(g27074)
--	g30195 = NOT(I28434)
--	g7400 = NOT(g911)
--	g8859 = NOT(g772)
--	g32953 = NOT(g31327)
--	g19737 = NOT(g17015)
--	g11720 = NOT(I14589)
--	g20283 = NOT(I20529)
--	g6811 = NOT(g714)
--	g34195 = NOT(I32150)
--	g20606 = NOT(g17955)
--	g33250 = NOT(g32186)
--	g16655 = NOT(g14151)
--	g10882 = NOT(g7601)
--	I18104 = NOT(g13177)
--	g10414 = NOT(g7092)
--	I13634 = NOT(g79)
--	g31658 = NOT(I29242)
--	I13872 = NOT(g7474)
--	g13041 = NOT(I15667)
--	g32654 = NOT(g31070)
--	g9843 = NOT(g4311)
--	g33658 = NOT(g33080)
--	g16180 = NOT(g13437)
--	g30016 = NOT(g29049)
--	g9989 = NOT(g5077)
--	I24448 = NOT(g22923)
--	g11430 = NOT(g7617)
--	g22541 = NOT(I21911)
--	g34559 = NOT(g34384)
--	g12350 = NOT(I15190)
--	g10407 = NOT(g7063)
--	g32800 = NOT(g31021)
--	g32936 = NOT(g31710)
--	g19697 = NOT(g16886)
--	I31486 = NOT(g33197)
--	g23215 = NOT(g20785)
--	g12820 = NOT(g10233)
--	I17699 = NOT(g13416)
--	g23501 = NOT(g20924)
--	g6874 = NOT(g3143)
--	I29965 = NOT(g31189)
--	I32109 = NOT(g33631)
--	I21033 = NOT(g17221)
--	g20381 = NOT(g17955)
--	g8342 = NOT(I12519)
--	g11237 = NOT(I14305)
--	g9834 = NOT(g2579)
--	g9971 = NOT(g2093)
--	I21234 = NOT(g16540)
--	g24982 = NOT(g22763)
--	g26679 = NOT(g25385)
--	g34830 = NOT(I33044)
--	g34893 = NOT(I33119)
--	g9686 = NOT(g73)
--	g22359 = NOT(g19495)
--	g8255 = NOT(g2028)
--	g17473 = NOT(g14841)
--	g20091 = NOT(g17328)
--	I22366 = NOT(g19757)
--	g24091 = NOT(g20720)
--	g7183 = NOT(g4608)
--	g8481 = NOT(I12618)
--	I12128 = NOT(g4253)
--	g17789 = NOT(g14321)
--	g29956 = NOT(I28185)
--	g29385 = NOT(g28180)
--	g34544 = NOT(I32613)
--	g15480 = NOT(I17125)
--	I26664 = NOT(g27708)
--	g22358 = NOT(g19801)
--	g32762 = NOT(g31672)
--	g9598 = NOT(g2571)
--	g24174 = NOT(I23366)
--	g8097 = NOT(g3029)
--	g25260 = NOT(I24448)
--	g32964 = NOT(g31672)
--	g29980 = NOT(g28935)
--	g7779 = NOT(g1413)
--	g34713 = NOT(I32871)
--	g8497 = NOT(g3436)
--	g13142 = NOT(g10632)
--	g21349 = NOT(g15758)
--	g8154 = NOT(g3139)
--	I28591 = NOT(g29371)
--	g17325 = NOT(I18304)
--	g8354 = NOT(g4815)
--	g18948 = NOT(g15800)
--	g7023 = NOT(g5445)
--	g31855 = NOT(g29385)
--	g10206 = NOT(g4489)
--	g14441 = NOT(I16590)
--	g14584 = NOT(g11048)
--	g9321 = NOT(g5863)
--	g7423 = NOT(g2433)
--	g9670 = NOT(g5022)
--	I22547 = NOT(g20720)
--	g25195 = NOT(g22763)
--	g16487 = NOT(I17695)
--	g23906 = NOT(g19074)
--	g26093 = NOT(g24814)
--	g30610 = NOT(I28872)
--	g18904 = NOT(g16053)
--	g32587 = NOT(g30735)
--	g15085 = NOT(I17008)
--	I32982 = NOT(g34749)
--	g23284 = NOT(g20785)
--	g19445 = NOT(g15915)
--	g10725 = NOT(g7846)
--	g21304 = NOT(g17367)
--	g25525 = NOT(g22550)
--	g34042 = NOT(g33674)
--	g25424 = NOT(g23800)
--	I20433 = NOT(g16234)
--	g23304 = NOT(g20785)
--	g25016 = NOT(g23666)
--	g6978 = NOT(g4616)
--	I33179 = NOT(g34893)
--	g7161 = NOT(I11843)
--	g19499 = NOT(g16782)
--	g17121 = NOT(g14321)
--	g7361 = NOT(g1874)
--	g22682 = NOT(g19379)
--	g10114 = NOT(g2116)
--	g20192 = NOT(g17268)
--	g9253 = NOT(g5037)
--	I16821 = NOT(g5983)
--	I17661 = NOT(g13329)
--	g27929 = NOT(I26448)
--	g25558 = NOT(g22594)
--	g23566 = NOT(g21562)
--	g32909 = NOT(g30614)
--	g10082 = NOT(g2375)
--	g32543 = NOT(g31376)
--	g34270 = NOT(g34159)
--	I27232 = NOT(g27993)
--	g19498 = NOT(g16752)
--	g34188 = NOT(g33875)
--	g7051 = NOT(I11793)
--	g10107 = NOT(I13606)
--	g22173 = NOT(I21757)
--	g34124 = NOT(g33819)
--	g9909 = NOT(g1978)
--	g12929 = NOT(g12550)
--	g25830 = NOT(g24485)
--	g27583 = NOT(g26686)
--	g20663 = NOT(g15373)
--	g27928 = NOT(g26810)
--	g25893 = NOT(g24541)
--	g8783 = NOT(I12761)
--	g7451 = NOT(g2070)
--	g32908 = NOT(g31327)
--	g6982 = NOT(g4531)
--	g7327 = NOT(g2165)
--	g24522 = NOT(g22689)
--	g33894 = NOT(I31748)
--	g11165 = NOT(I14222)
--	g8112 = NOT(g3419)
--	g8218 = NOT(g3490)
--	g34939 = NOT(g34922)
--	g9740 = NOT(g5821)
--	g8267 = NOT(g2342)
--	g25544 = NOT(g22594)
--	g32569 = NOT(g30673)
--	g34383 = NOT(I32388)
--	g29190 = NOT(g27046)
--	I32840 = NOT(g34480)
--	g17291 = NOT(I18276)
--	g14744 = NOT(g12578)
--	g16286 = NOT(I17615)
--	g21139 = NOT(g15634)
--	g21653 = NOT(g17663)
--	g26837 = NOT(g24869)
--	g7633 = NOT(I12120)
--	g34938 = NOT(g34920)
--	g23653 = NOT(I22788)
--	g9552 = NOT(g3654)
--	g15655 = NOT(g13202)
--	I31800 = NOT(g33164)
--	g10399 = NOT(g7017)
--	g32568 = NOT(g31170)
--	g32747 = NOT(g30825)
--	I18310 = NOT(g12978)
--	I20369 = NOT(g17690)
--	g18062 = NOT(I18872)
--	g21138 = NOT(g15634)
--	g24483 = NOT(I23688)
--	g19432 = NOT(g15885)
--	I19837 = NOT(g1399)
--	g30065 = NOT(g29049)
--	I11820 = NOT(g3869)
--	g23138 = NOT(g20453)
--	I26799 = NOT(g27660)
--	g20553 = NOT(g17929)
--	g31819 = NOT(g29385)
--	g8676 = NOT(g4821)
--	I15727 = NOT(g10981)
--	I32192 = NOT(g33628)
--	g10398 = NOT(g6999)
--	I18379 = NOT(g13012)
--	g14398 = NOT(I16555)
--	g10141 = NOT(I13634)
--	g29211 = NOT(I27549)
--	g10652 = NOT(g7601)
--	g10804 = NOT(g9772)
--	g6800 = NOT(g203)
--	I13152 = NOT(g6746)
--	g9687 = NOT(I13287)
--	g31818 = NOT(g29385)
--	g32814 = NOT(g31021)
--	g20326 = NOT(g18008)
--	g23333 = NOT(g20785)
--	g13222 = NOT(g10590)
--	g19753 = NOT(g16987)
--	g16601 = NOT(I17783)
--	g17760 = NOT(I18752)
--	g16677 = NOT(I17879)
--	I22889 = NOT(g18926)
--	g20536 = NOT(g18065)
--	g20040 = NOT(g17271)
--	g13437 = NOT(I15937)
--	I20412 = NOT(g16213)
--	g32751 = NOT(g31327)
--	g32807 = NOT(g31021)
--	g32772 = NOT(g31327)
--	g28463 = NOT(I26952)
--	g32974 = NOT(g30937)
--	g8830 = NOT(g767)
--	g24040 = NOT(g19919)
--	g7753 = NOT(I12183)
--	g20702 = NOT(g17955)
--	g30218 = NOT(g28918)
--	g25188 = NOT(g23909)
--	g32639 = NOT(g31070)
--	g20904 = NOT(g17433)
--	I17956 = NOT(g14562)
--	g23963 = NOT(g19147)
--	g19650 = NOT(g16971)
--	g28033 = NOT(g26365)
--	g8592 = NOT(g3805)
--	g7072 = NOT(g6199)
--	g14332 = NOT(I16492)
--	I11691 = NOT(g36)
--	I28540 = NOT(g28954)
--	g32638 = NOT(g30825)
--	g7472 = NOT(g6329)
--	g19529 = NOT(g16349)
--	g12640 = NOT(I15382)
--	I15600 = NOT(g10430)
--	g22927 = NOT(I22128)
--	g9860 = NOT(g5417)
--	g10406 = NOT(g7046)
--	I24228 = NOT(g22409)
--	g20564 = NOT(g15373)
--	g10361 = NOT(g6841)
--	I25576 = NOT(g25296)
--	g7443 = NOT(g914)
--	g8703 = NOT(I12709)
--	g14406 = NOT(g12249)
--	g19528 = NOT(g16349)
--	g19696 = NOT(g17015)
--	g34160 = NOT(I32119)
--	g25267 = NOT(g22228)
--	g19330 = NOT(g17326)
--	I17181 = NOT(g13745)
--	I17671 = NOT(g13280)
--	I29363 = NOT(g30218)
--	g23585 = NOT(g21070)
--	g32841 = NOT(g31672)
--	g11236 = NOT(g8357)
--	I21291 = NOT(g18273)
--	g7116 = NOT(g22)
--	g22649 = NOT(g19063)
--	g10500 = NOT(I13875)
--	g27881 = NOT(I26430)
--	g19365 = NOT(g16249)
--	g20673 = NOT(g15277)
--	g32510 = NOT(g31194)
--	g9691 = NOT(g1706)
--	g31801 = NOT(g29385)
--	I15821 = NOT(g11143)
--	I12056 = NOT(g2748)
--	g24183 = NOT(I23393)
--	I32904 = NOT(g34708)
--	g14833 = NOT(g11405)
--	g19869 = NOT(g16540)
--	g21609 = NOT(g18008)
--	g19960 = NOT(g17433)
--	g23609 = NOT(g21611)
--	g24397 = NOT(g22908)
--	g29339 = NOT(g28274)
--	g12881 = NOT(g10388)
--	g7565 = NOT(I12046)
--	g22903 = NOT(g20330)
--	g13175 = NOT(g10909)
--	g34915 = NOT(I33137)
--	I16593 = NOT(g10498)
--	I25115 = NOT(g25322)
--	g32579 = NOT(g30735)
--	g8068 = NOT(g3457)
--	I13020 = NOT(g6750)
--	I32621 = NOT(g34335)
--	g23312 = NOT(g21070)
--	I31569 = NOT(g33197)
--	I28301 = NOT(g29042)
--	g25219 = NOT(I24393)
--	I27271 = NOT(g27998)
--	g21608 = NOT(g17955)
--	g24062 = NOT(g19968)
--	g17649 = NOT(I18614)
--	g20509 = NOT(g15277)
--	g23608 = NOT(g21611)
--	g34201 = NOT(I32158)
--	g9607 = NOT(g5046)
--	g24509 = NOT(g22689)
--	g32578 = NOT(g31376)
--	g32835 = NOT(g31710)
--	g33695 = NOT(g33187)
--	g34277 = NOT(I32274)
--	g25218 = NOT(g23949)
--	g9962 = NOT(g6519)
--	g11790 = NOT(I14630)
--	g14004 = NOT(g11149)
--	g17648 = NOT(g15024)
--	g20508 = NOT(g15277)
--	g9158 = NOT(g513)
--	g27662 = NOT(I26296)
--	g17491 = NOT(g12983)
--	g22981 = NOT(g20283)
--	g20634 = NOT(g15373)
--	I21029 = NOT(g15816)
--	g21052 = NOT(g15373)
--	g28163 = NOT(I26682)
--	g8677 = NOT(g4854)
--	g25837 = NOT(g25064)
--	g7533 = NOT(g1306)
--	g19709 = NOT(g16987)
--	g32586 = NOT(g31376)
--	I22211 = NOT(g21463)
--	g9506 = NOT(g5774)
--	g17604 = NOT(I18555)
--	g34595 = NOT(I32693)
--	g7697 = NOT(g4087)
--	g10613 = NOT(g10233)
--	g23745 = NOT(g20900)
--	I18504 = NOT(g5283)
--	I22024 = NOT(g19350)
--	g32442 = NOT(g31213)
--	I31814 = NOT(g33149)
--	g19471 = NOT(g16449)
--	g30037 = NOT(g29121)
--	g12890 = NOT(g10397)
--	g16580 = NOT(I17754)
--	g23813 = NOT(g18997)
--	g7596 = NOT(I12070)
--	I31751 = NOT(g33228)
--	I31807 = NOT(g33149)
--	g16223 = NOT(g13437)
--	g10273 = NOT(I13708)
--	g33457 = NOT(I30989)
--	I32062 = NOT(g33653)
--	I12199 = NOT(g6215)
--	g10106 = NOT(g16)
--	g9311 = NOT(g5523)
--	I11743 = NOT(g4564)
--	g22845 = NOT(g20682)
--	I12887 = NOT(g4216)
--	g34984 = NOT(I33252)
--	g32615 = NOT(g31376)
--	I15834 = NOT(g11164)
--	g13209 = NOT(g10632)
--	g8848 = NOT(g358)
--	g20213 = NOT(g17062)
--	I15208 = NOT(g637)
--	g33917 = NOT(I31779)
--	g21184 = NOT(g15509)
--	g34419 = NOT(g34151)
--	g9615 = NOT(I13236)
--	g21674 = NOT(g16540)
--	g10812 = NOT(I14050)
--	g32720 = NOT(g31710)
--	g30155 = NOT(I28390)
--	g8398 = NOT(I12563)
--	g28325 = NOT(g27463)
--	g12779 = NOT(g9444)
--	g22898 = NOT(g20283)
--	g9174 = NOT(g1205)
--	g34418 = NOT(g34150)
--	g17794 = NOT(g13350)
--	g26836 = NOT(g24866)
--	g17845 = NOT(I18835)
--	g9374 = NOT(g5188)
--	g20574 = NOT(g17847)
--	g20452 = NOT(g17200)
--	I15542 = NOT(g1570)
--	g32430 = NOT(g30984)
--	g10033 = NOT(g655)
--	g10371 = NOT(g6918)
--	g32746 = NOT(g30735)
--	g32493 = NOT(g30735)
--	g22719 = NOT(I22024)
--	g24452 = NOT(g22722)
--	I26100 = NOT(g26365)
--	g7936 = NOT(g1061)
--	g9985 = NOT(g4332)
--	g24047 = NOT(g19919)
--	g12778 = NOT(g9856)
--	I18245 = NOT(g14676)
--	I12764 = NOT(g4194)
--	g23732 = NOT(g18833)
--	g8241 = NOT(g1792)
--	I20793 = NOT(g17694)
--	g20912 = NOT(g15171)
--	g19602 = NOT(g16349)
--	g32465 = NOT(g30825)
--	g7117 = NOT(I11816)
--	I18323 = NOT(g13680)
--	g19657 = NOT(g16349)
--	g22718 = NOT(g20887)
--	g16740 = NOT(g13980)
--	I12132 = NOT(g577)
--	g19068 = NOT(g16031)
--	g15169 = NOT(I17094)
--	g28121 = NOT(g27093)
--	g9284 = NOT(g2161)
--	g19375 = NOT(I19863)
--	g10795 = NOT(g7202)
--	I25692 = NOT(g25689)
--	g9239 = NOT(g5511)
--	g33923 = NOT(I31791)
--	g9180 = NOT(g3719)
--	g16186 = NOT(g13555)
--	g16676 = NOT(I17876)
--	g16685 = NOT(g14038)
--	I20690 = NOT(g15733)
--	I29936 = NOT(g30606)
--	I17658 = NOT(g13394)
--	g9380 = NOT(g5471)
--	g12945 = NOT(g12467)
--	g31624 = NOT(I29218)
--	g32806 = NOT(g31710)
--	g20072 = NOT(g17384)
--	g32684 = NOT(g30673)
--	g33688 = NOT(I31523)
--	g29707 = NOT(g28504)
--	g9832 = NOT(g2399)
--	I15073 = NOT(g10109)
--	g19878 = NOT(g17271)
--	g24051 = NOT(g21127)
--	g24072 = NOT(g20982)
--	g34589 = NOT(I32675)
--	g17718 = NOT(g14776)
--	g17521 = NOT(g14727)
--	g16654 = NOT(g14136)
--	g20592 = NOT(g15277)
--	g27998 = NOT(I26512)
--	I16575 = NOT(g3298)
--	g15479 = NOT(g14895)
--	g9853 = NOT(g5297)
--	I15593 = NOT(g11989)
--	g8644 = NOT(g3352)
--	g6989 = NOT(g4575)
--	g9020 = NOT(g4287)
--	g24756 = NOT(g22763)
--	I32452 = NOT(g34241)
--	I12709 = NOT(g4284)
--	g21400 = NOT(g17847)
--	g20780 = NOT(g15509)
--	g7922 = NOT(g1312)
--	g8119 = NOT(g3727)
--	g13530 = NOT(g12641)
--	g23400 = NOT(g20676)
--	g12998 = NOT(g11829)
--	g34836 = NOT(I33050)
--	g13593 = NOT(g10556)
--	g28173 = NOT(I26693)
--	g18929 = NOT(g16100)
--	g32517 = NOT(g31194)
--	g23013 = NOT(g20330)
--	I28572 = NOT(g28274)
--	g12233 = NOT(g10338)
--	I31586 = NOT(g33149)
--	g23214 = NOT(g20785)
--	g11122 = NOT(g8751)
--	I14902 = NOT(g9821)
--	I14301 = NOT(g8571)
--	g12182 = NOT(I15030)
--	g29978 = NOT(g28927)
--	g12672 = NOT(g10003)
--	g7581 = NOT(g1379)
--	g21329 = NOT(g16577)
--	g22926 = NOT(g20391)
--	g25155 = NOT(g22472)
--	g9559 = NOT(g6077)
--	g13565 = NOT(g11006)
--	g6971 = NOT(I11737)
--	g8818 = NOT(I12808)
--	I25005 = NOT(g24417)
--	g14421 = NOT(I16575)
--	I19704 = NOT(g17653)
--	g25266 = NOT(g22228)
--	g25170 = NOT(g22498)
--	g9931 = NOT(g5763)
--	g23539 = NOT(g21070)
--	g17573 = NOT(g12911)
--	g7597 = NOT(g952)
--	g11034 = NOT(g7611)
--	g23005 = NOT(g20283)
--	g13034 = NOT(g11920)
--	g17247 = NOT(I18259)
--	I32051 = NOT(g33631)
--	g30022 = NOT(g29001)
--	g34118 = NOT(I32051)
--	I16606 = NOT(g3649)
--	g15580 = NOT(g13242)
--	g12932 = NOT(I15550)
--	g23538 = NOT(g20924)
--	g34864 = NOT(g34840)
--	I16492 = NOT(g12430)
--	g17389 = NOT(g14915)
--	g17926 = NOT(I18852)
--	g16964 = NOT(I18120)
--	g24152 = NOT(I23300)
--	g19458 = NOT(I19927)
--	g30313 = NOT(g28843)
--	g34749 = NOT(I32921)
--	g17612 = NOT(g15014)
--	g24396 = NOT(g22885)
--	g8211 = NOT(g2319)
--	g29067 = NOT(I27401)
--	g9905 = NOT(g802)
--	g10541 = NOT(g9407)
--	g16423 = NOT(g14066)
--	g27961 = NOT(g26816)
--	g8186 = NOT(g990)
--	g34313 = NOT(g34086)
--	I13552 = NOT(g121)
--	g10473 = NOT(I13857)
--	g17324 = NOT(I18301)
--	g32523 = NOT(g30825)
--	I24128 = NOT(g23009)
--	g31854 = NOT(g29385)
--	g14541 = NOT(g11405)
--	g16216 = NOT(I17557)
--	I29909 = NOT(g31791)
--	I33041 = NOT(g34772)
--	g12897 = NOT(g10400)
--	g13409 = NOT(I15918)
--	g16587 = NOT(I17763)
--	g17777 = NOT(g14908)
--	g25167 = NOT(I24331)
--	g25194 = NOT(g22763)
--	I13779 = NOT(g6868)
--	I26584 = NOT(g26943)
--	g9630 = NOT(g6527)
--	g29150 = NOT(g27886)
--	g34276 = NOT(g34058)
--	g34285 = NOT(I32284)
--	g7995 = NOT(g153)
--	g30305 = NOT(g28939)
--	g11136 = NOT(I14192)
--	g30053 = NOT(g29121)
--	g8026 = NOT(g3857)
--	g25524 = NOT(g22228)
--	I27970 = NOT(g28803)
--	g18827 = NOT(g16000)
--	g34053 = NOT(g33683)
--	g7479 = NOT(g1008)
--	g9300 = NOT(g5180)
--	g10359 = NOT(g6830)
--	I32820 = NOT(g34474)
--	g8426 = NOT(g3045)
--	g32475 = NOT(g30614)
--	g14359 = NOT(I16515)
--	g8170 = NOT(g3770)
--	g7840 = NOT(g4878)
--	g22997 = NOT(g20391)
--	g32727 = NOT(g31710)
--	g10358 = NOT(g6827)
--	g33660 = NOT(I31494)
--	g32863 = NOT(g31021)
--	g29196 = NOT(g27059)
--	I32846 = NOT(g34502)
--	g14535 = NOT(g12318)
--	g24405 = NOT(g22722)
--	g8125 = NOT(g3869)
--	g30036 = NOT(g29085)
--	g14358 = NOT(I16512)
--	g25119 = NOT(g22384)
--	I22819 = NOT(g19862)
--	g8821 = NOT(I12811)
--	g16000 = NOT(I17425)
--	g15740 = NOT(g13342)
--	I25683 = NOT(g25642)
--	I29242 = NOT(g29313)
--	g32437 = NOT(I29965)
--	g14828 = NOT(I16875)
--	g23235 = NOT(g20785)
--	g33456 = NOT(I30986)
--	g10121 = NOT(g2327)
--	g11164 = NOT(g8085)
--	g25118 = NOT(g22417)
--	g26693 = NOT(g25300)
--	g8280 = NOT(g3443)
--	g23683 = NOT(I22816)
--	g15373 = NOT(I17118)
--	g9973 = NOT(g2112)
--	g33916 = NOT(I31776)
--	I22111 = NOT(g19919)
--	g7356 = NOT(g1802)
--	I17819 = NOT(g3618)
--	g16747 = NOT(g14113)
--	g20583 = NOT(g17873)
--	g32703 = NOT(g30825)
--	I12994 = NOT(g6748)
--	I15474 = NOT(g10364)
--	g24020 = NOT(g20014)
--	g19532 = NOT(g16821)
--	g22360 = NOT(I21849)
--	g9040 = NOT(g499)
--	g28648 = NOT(g27693)
--	g18881 = NOT(I19671)
--	I13672 = NOT(g106)
--	g13474 = NOT(g11048)
--	I25882 = NOT(g25776)
--	g20046 = NOT(g16540)
--	g9969 = NOT(g1682)
--	g19783 = NOT(g16931)
--	I17111 = NOT(g13809)
--	g16123 = NOT(g13530)
--	g24046 = NOT(g21256)
--	g17871 = NOT(I18845)
--	g16814 = NOT(g14058)
--	g21414 = NOT(g17929)
--	g32600 = NOT(g31542)
--	g7704 = NOT(I12167)
--	I16663 = NOT(g10981)
--	g23515 = NOT(g20785)
--	g28604 = NOT(g27759)
--	g23882 = NOT(g19277)
--	g23414 = NOT(I22525)
--	g32781 = NOT(g31376)
--	I23099 = NOT(g20682)
--	g31596 = NOT(I29204)
--	g8106 = NOT(g3133)
--	g14173 = NOT(g12076)
--	I23324 = NOT(g21697)
--	g20113 = NOT(g16826)
--	g21407 = NOT(g15171)
--	g31243 = NOT(g29933)
--	I17590 = NOT(g14591)
--	g19353 = NOT(I19831)
--	g24113 = NOT(g19984)
--	I32929 = NOT(g34649)
--	g32952 = NOT(g30937)
--	g19144 = NOT(g16031)
--	g12811 = NOT(g10319)
--	g27971 = NOT(g26673)
--	g8187 = NOT(g1657)
--	g32821 = NOT(g31021)
--	g8387 = NOT(g3080)
--	g25036 = NOT(g23733)
--	I31523 = NOT(g33187)
--	g7163 = NOT(g4593)
--	g29597 = NOT(g28444)
--	g25101 = NOT(g22384)
--	g20105 = NOT(g17433)
--	g24357 = NOT(g22325)
--	g25560 = NOT(g22550)
--	g10029 = NOT(I13548)
--	g8756 = NOT(g4049)
--	g22220 = NOT(I21802)
--	g13303 = NOT(I15869)
--	g24105 = NOT(g19935)
--	I17094 = NOT(g14331)
--	I18031 = NOT(g13680)
--	g29689 = NOT(I27954)
--	g14029 = NOT(g11283)
--	g29923 = NOT(g28874)
--	g25642 = NOT(I24787)
--	g32790 = NOT(g30825)
--	g9648 = NOT(g2177)
--	g32137 = NOT(g31134)
--	g10028 = NOT(g8)
--	g9875 = NOT(g5747)
--	g32516 = NOT(g31070)
--	g31655 = NOT(I29233)
--	I29579 = NOT(g30565)
--	g28262 = NOT(I26785)
--	I24445 = NOT(g22923)
--	g20640 = NOT(g15426)
--	I17801 = NOT(g14936)
--	g20769 = NOT(g17955)
--	g17472 = NOT(g14656)
--	I26406 = NOT(g26187)
--	g12368 = NOT(I15208)
--	I16040 = NOT(g10430)
--	I20499 = NOT(g16224)
--	I12086 = NOT(g622)
--	g33670 = NOT(I31504)
--	I31727 = NOT(g33076)
--	g32873 = NOT(g30614)
--	g8046 = NOT(g528)
--	g25064 = NOT(I24228)
--	g16510 = NOT(g14008)
--	g19364 = NOT(g15825)
--	g20768 = NOT(g17955)
--	g28633 = NOT(g27687)
--	g8514 = NOT(g4258)
--	I19238 = NOT(g15079)
--	g34570 = NOT(g34392)
--	g34712 = NOT(I32868)
--	g21725 = NOT(I21294)
--	g11796 = NOT(g7985)
--	g16579 = NOT(g13267)
--	g33335 = NOT(I30861)
--	g8403 = NOT(I12568)
--	g23759 = NOT(I22886)
--	g13174 = NOT(g10741)
--	I21766 = NOT(g19620)
--	I17695 = NOT(g14330)
--	g26941 = NOT(I25689)
--	g34914 = NOT(I33134)
--	g31839 = NOT(g29385)
--	g33839 = NOT(I31686)
--	I32827 = NOT(g34477)
--	g8345 = NOT(g3794)
--	g8841 = NOT(I12823)
--	I14671 = NOT(g7717)
--	g7157 = NOT(g5706)
--	I12159 = NOT(g608)
--	g22147 = NOT(g18997)
--	g26519 = NOT(I25380)
--	g16578 = NOT(I17750)
--	g15569 = NOT(I17148)
--	g8763 = NOT(I12749)
--	I16564 = NOT(g10429)
--	g23435 = NOT(g18833)
--	g31667 = NOT(g30142)
--	g31838 = NOT(g29385)
--	g23082 = NOT(g21024)
--	g32834 = NOT(g31672)
--	g9839 = NOT(g2724)
--	g30074 = NOT(g29046)
--	g26518 = NOT(g25233)
--	g17591 = NOT(I18526)
--	g12896 = NOT(g10402)
--	g17776 = NOT(g14905)
--	g27011 = NOT(g25917)
--	I27561 = NOT(g28163)
--	g15568 = NOT(g14984)
--	g15747 = NOT(g13307)
--	g25009 = NOT(g22472)
--	I13723 = NOT(g3167)
--	I26004 = NOT(g26818)
--	I18868 = NOT(g14315)
--	I23360 = NOT(g23360)
--	g18945 = NOT(g16100)
--	g30567 = NOT(g29930)
--	I30962 = NOT(g32021)
--	g17147 = NOT(g14321)
--	g22858 = NOT(g20751)
--	g34594 = NOT(I32690)
--	I13149 = NOT(g6745)
--	g17754 = NOT(g14262)
--	I16847 = NOT(g6329)
--	g26935 = NOT(I25677)
--	g25008 = NOT(g22432)
--	g32542 = NOT(g31554)
--	g8107 = NOT(g3179)
--	I32803 = NOT(g34584)
--	I25399 = NOT(g24489)
--	g31487 = NOT(I29149)
--	g32021 = NOT(I29579)
--	g32453 = NOT(I29981)
--	I29720 = NOT(g30931)
--	g11192 = NOT(g8038)
--	g22151 = NOT(I21734)
--	I11620 = NOT(g1)
--	I21162 = NOT(g17292)
--	I12144 = NOT(g554)
--	I12823 = NOT(g4311)
--	I18709 = NOT(g6668)
--	g20662 = NOT(g15171)
--	g21399 = NOT(g15224)
--	g23849 = NOT(g19277)
--	g22996 = NOT(g20330)
--	g23940 = NOT(g19074)
--	g25892 = NOT(g24528)
--	I20753 = NOT(g16677)
--	I15663 = NOT(g5308)
--	g23399 = NOT(g21514)
--	g32726 = NOT(g31672)
--	g32913 = NOT(g30825)
--	g24027 = NOT(g20014)
--	I18259 = NOT(g12946)
--	g9618 = NOT(g5794)
--	g11663 = NOT(g6905)
--	g16615 = NOT(I17801)
--	g22844 = NOT(g21163)
--	g13522 = NOT(g10981)
--	g34941 = NOT(g34926)
--	g13663 = NOT(g10971)
--	g21398 = NOT(g18008)
--	g23848 = NOT(g19210)
--	g25555 = NOT(g22550)
--	g32614 = NOT(g31542)
--	g7626 = NOT(I12112)
--	I12336 = NOT(g52)
--	g23398 = NOT(g21468)
--	I32881 = NOT(g34688)
--	g8858 = NOT(g671)
--	g33443 = NOT(I30971)
--	g16720 = NOT(g14234)
--	g9282 = NOT(g723)
--	g34675 = NOT(I32809)
--	I20650 = NOT(g17010)
--	g23652 = NOT(I22785)
--	g32607 = NOT(g31542)
--	g8016 = NOT(g3391)
--	g10981 = NOT(I14119)
--	g8757 = NOT(I12746)
--	g32905 = NOT(g30825)
--	g14563 = NOT(I16676)
--	g8416 = NOT(I12580)
--	g27112 = NOT(g26793)
--	g20710 = NOT(g15509)
--	g16746 = NOT(g14258)
--	I20529 = NOT(g16309)
--	I21911 = NOT(g21278)
--	g17844 = NOT(I18832)
--	g20552 = NOT(g17847)
--	g32530 = NOT(g30825)
--	g9693 = NOT(g1886)
--	g13483 = NOT(g11270)
--	I33264 = NOT(g34978)
--	I15862 = NOT(g11215)
--	g17367 = NOT(I18320)
--	g32593 = NOT(g31542)
--	g18932 = NOT(g16136)
--	g6985 = NOT(g4669)
--	I33137 = NOT(g34884)
--	g20204 = NOT(g16578)
--	g19687 = NOT(g17096)
--	I21246 = NOT(g16540)
--	g24003 = NOT(g21514)
--	g23263 = NOT(I22366)
--	I12631 = NOT(g1242)
--	g8522 = NOT(g298)
--	g20779 = NOT(g15509)
--	g22319 = NOT(I21831)
--	g12378 = NOT(g9417)
--	g34935 = NOT(I33189)
--	g23332 = NOT(g20785)
--	g32565 = NOT(g30735)
--	g32464 = NOT(g30735)
--	g25239 = NOT(g23972)
--	g19954 = NOT(g16540)
--	g11949 = NOT(I14773)
--	I24393 = NOT(g23453)
--	g19374 = NOT(g16047)
--	g20778 = NOT(g15224)
--	g34883 = NOT(g34852)
--	g10794 = NOT(g8470)
--	g9555 = NOT(I13206)
--	g18897 = NOT(g15509)
--	I15536 = NOT(g1227)
--	g10395 = NOT(g6995)
--	g22227 = NOT(g19801)
--	g24778 = NOT(g23286)
--	g9804 = NOT(g5456)
--	g10262 = NOT(g586)
--	g24081 = NOT(g21209)
--	g21406 = NOT(g17955)
--	g16684 = NOT(g14223)
--	g11948 = NOT(g10224)
--	I21776 = NOT(g21308)
--	I15702 = NOT(g12217)
--	g14262 = NOT(g10838)
--	g12944 = NOT(g12659)
--	I18810 = NOT(g13716)
--	g23406 = NOT(g20330)
--	g9792 = NOT(g5401)
--	g32641 = NOT(g30614)
--	g6832 = NOT(I11665)
--	g32797 = NOT(g30825)
--	g23962 = NOT(g19147)
--	g31815 = NOT(g29385)
--	g23361 = NOT(I22464)
--	g28032 = NOT(g26365)
--	I32482 = NOT(g34304)
--	g11702 = NOT(g6928)
--	g7778 = NOT(g1339)
--	g15579 = NOT(I17159)
--	g31601 = NOT(I29207)
--	g8654 = NOT(g1087)
--	I16452 = NOT(g11182)
--	I18879 = NOT(g13267)
--	g9621 = NOT(g6423)
--	g10191 = NOT(g6386)
--	g23500 = NOT(g20924)
--	g24356 = NOT(g22594)
--	g13621 = NOT(g10573)
--	g21049 = NOT(g17433)
--	I11896 = NOT(g4446)
--	g25185 = NOT(g22228)
--	g17059 = NOT(I18151)
--	g20380 = NOT(g17955)
--	g26083 = NOT(g24809)
--	g14191 = NOT(g12381)
--	g30729 = NOT(I28883)
--	I15564 = NOT(g11949)
--	g25092 = NOT(g23666)
--	g24999 = NOT(g23626)
--	g26284 = NOT(g24875)
--	I18337 = NOT(g1422)
--	g34501 = NOT(g34400)
--	g27730 = NOT(g26424)
--	g10521 = NOT(I13889)
--	g12857 = NOT(I15474)
--	I19348 = NOT(g15084)
--	g21048 = NOT(g17533)
--	g25154 = NOT(g22457)
--	g20090 = NOT(g17433)
--	g17058 = NOT(I18148)
--	g32635 = NOT(g31542)
--	g8880 = NOT(I12861)
--	g31937 = NOT(g30991)
--	g8595 = NOT(I12666)
--	g24090 = NOT(g19935)
--	g19489 = NOT(g16449)
--	g20233 = NOT(g17873)
--	g33937 = NOT(I31823)
--	g12793 = NOT(g10287)
--	I11716 = NOT(g4054)
--	g20182 = NOT(g16897)
--	g20651 = NOT(g15483)
--	g20672 = NOT(g15277)
--	I17876 = NOT(g13070)
--	g23004 = NOT(g20283)
--	I27495 = NOT(g27961)
--	g7475 = NOT(g896)
--	g21221 = NOT(g15680)
--	g24182 = NOT(I23390)
--	g19559 = NOT(g16129)
--	g23221 = NOT(g20785)
--	I14644 = NOT(g7717)
--	g11183 = NOT(g8135)
--	g29942 = NOT(g28867)
--	g22957 = NOT(I22143)
--	g31791 = NOT(I29363)
--	g7627 = NOT(g4311)
--	g19558 = NOT(g15938)
--	g6905 = NOT(I11708)
--	g16523 = NOT(g14041)
--	g8612 = NOT(g2775)
--	g23613 = NOT(I22748)
--	g9518 = NOT(g6219)
--	g15615 = NOT(I17181)
--	I17763 = NOT(g13191)
--	I31607 = NOT(g33164)
--	g13062 = NOT(g10981)
--	g7526 = NOT(I12013)
--	g7998 = NOT(g392)
--	g11509 = NOT(g7632)
--	g22146 = NOT(g18997)
--	g26653 = NOT(g25337)
--	g20513 = NOT(g18065)
--	g17301 = NOT(g14454)
--	g20449 = NOT(g15277)
--	g28162 = NOT(I26679)
--	g10389 = NOT(g6986)
--	g32891 = NOT(g30825)
--	I15872 = NOT(g11236)
--	g13933 = NOT(g11419)
--	g23947 = NOT(g19210)
--	g31479 = NOT(I29139)
--	g31666 = NOT(I29248)
--	I27954 = NOT(g28803)
--	g18097 = NOT(I18897)
--	g21273 = NOT(I21006)
--	g17120 = NOT(g14262)
--	g19544 = NOT(g16349)
--	g23273 = NOT(g21070)
--	g19865 = NOT(g15885)
--	g17739 = NOT(I18728)
--	g10612 = NOT(g10233)
--	g11872 = NOT(I14684)
--	g23605 = NOT(g20739)
--	g9776 = NOT(g5073)
--	g10099 = NOT(g6682)
--	g15746 = NOT(g13121)
--	g16475 = NOT(g14107)
--	g20448 = NOT(g15509)
--	g34304 = NOT(I32309)
--	I12954 = NOT(g4358)
--	g10388 = NOT(g6983)
--	I32651 = NOT(g34375)
--	g32575 = NOT(g31170)
--	g32474 = NOT(g31194)
--	g19713 = NOT(g16816)
--	g7439 = NOT(g6351)
--	g29930 = NOT(I28162)
--	g22698 = NOT(I22009)
--	g29993 = NOT(g29018)
--	g16727 = NOT(g14454)
--	g17738 = NOT(g14813)
--	g17645 = NOT(g15018)
--	g20505 = NOT(g15426)
--	g21463 = NOT(g15588)
--	g23812 = NOT(g18997)
--	g32711 = NOT(g31070)
--	g8130 = NOT(g4515)
--	g14701 = NOT(g12351)
--	I17456 = NOT(g13680)
--	I23318 = NOT(g21689)
--	g8542 = NOT(I12644)
--	g24505 = NOT(g22689)
--	g8330 = NOT(g2587)
--	g24404 = NOT(g22908)
--	g10272 = NOT(I13705)
--	g9965 = NOT(g127)
--	g29965 = NOT(g28903)
--	I33034 = NOT(g34769)
--	g14251 = NOT(g12308)
--	I17916 = NOT(g13087)
--	g20026 = NOT(g17271)
--	g32537 = NOT(g30825)
--	I18078 = NOT(g13350)
--	g20212 = NOT(g17194)
--	g23234 = NOT(g20375)
--	g24026 = NOT(g19919)
--	g9264 = NOT(g5396)
--	g15806 = NOT(I17302)
--	I21058 = NOT(g17747)
--	g25438 = NOT(g22763)
--	g6973 = NOT(I11743)
--	I17314 = NOT(g14078)
--	I32449 = NOT(g34127)
--	g19679 = NOT(g16782)
--	I18086 = NOT(g13856)
--	g27245 = NOT(g26209)
--	g34653 = NOT(I32763)
--	g9360 = NOT(g3372)
--	g9933 = NOT(g5759)
--	g32606 = NOT(g30673)
--	g10032 = NOT(g562)
--	I29236 = NOT(g29498)
--	g32492 = NOT(g31376)
--	g19678 = NOT(g16752)
--	I15205 = NOT(g10139)
--	g14032 = NOT(g11048)
--	g10140 = NOT(g19)
--	g29210 = NOT(I27546)
--	g9050 = NOT(g1087)
--	g17427 = NOT(I18364)
--	I13802 = NOT(g6971)
--	g13574 = NOT(I16024)
--	I25514 = NOT(g25073)
--	I13857 = NOT(g9780)
--	g17366 = NOT(g14454)
--	g7952 = NOT(g3774)
--	g25083 = NOT(g23782)
--	g25348 = NOT(g22763)
--	g9450 = NOT(g5817)
--	I14450 = NOT(g4191)
--	g16600 = NOT(I17780)
--	g19686 = NOT(g17062)
--	g25284 = NOT(I24474)
--	g21514 = NOT(I21189)
--	I11793 = NOT(g6049)
--	g11912 = NOT(g8989)
--	g26576 = NOT(I25399)
--	I26682 = NOT(g27774)
--	g28147 = NOT(I26654)
--	I27558 = NOT(g28155)
--	g32750 = NOT(g30937)
--	I12016 = NOT(g772)
--	I18125 = NOT(g13191)
--	g10061 = NOT(I13581)
--	g13311 = NOT(I15878)
--	g28754 = NOT(I27238)
--	g32381 = NOT(I29909)
--	g7616 = NOT(I12086)
--	I19484 = NOT(g15122)
--	g23507 = NOT(g21562)
--	g34852 = NOT(g34845)
--	g20433 = NOT(g17929)
--	g25566 = NOT(g22550)
--	g18896 = NOT(g16031)
--	g24149 = NOT(g19338)
--	g20387 = NOT(g15426)
--	g28370 = NOT(g27528)
--	I28866 = NOT(g29730)
--	I22180 = NOT(g21366)
--	g16821 = NOT(I18031)
--	g21421 = NOT(g15171)
--	g27737 = NOT(g26718)
--	I12893 = NOT(g4226)
--	g7004 = NOT(I11777)
--	g9379 = NOT(g5424)
--	g23421 = NOT(g21562)
--	g13051 = NOT(g11964)
--	g20097 = NOT(g17691)
--	g32796 = NOT(g31376)
--	g7527 = NOT(I12016)
--	I33164 = NOT(g34894)
--	g24097 = NOT(g19935)
--	g26608 = NOT(g25334)
--	g11592 = NOT(I14537)
--	g20104 = NOT(g17433)
--	g7647 = NOT(I12132)
--	g34664 = NOT(I32782)
--	I27713 = NOT(g28224)
--	I13548 = NOT(g94)
--	g10360 = NOT(g6836)
--	g23012 = NOT(g20330)
--	g24104 = NOT(g19890)
--	g17226 = NOT(I18252)
--	g25139 = NOT(g22472)
--	g17715 = NOT(I18700)
--	g6875 = NOT(I11697)
--	g9777 = NOT(g5112)
--	g17481 = NOT(g15005)
--	I25541 = NOT(g25180)
--	g32840 = NOT(g30825)
--	I28597 = NOT(g29374)
--	g28367 = NOT(I26880)
--	I31474 = NOT(g33212)
--	g24971 = NOT(g23590)
--	g27880 = NOT(I26427)
--	g25138 = NOT(g22472)
--	g34576 = NOT(I32654)
--	g16873 = NOT(I18063)
--	g23541 = NOT(g21514)
--	g31800 = NOT(g29385)
--	g12995 = NOT(g11820)
--	g7503 = NOT(g1351)
--	g7970 = NOT(g4688)
--	g13350 = NOT(I15906)
--	g23473 = NOT(g20785)
--	g33800 = NOT(I31642)
--	g8056 = NOT(g1246)
--	I13317 = NOT(g6144)
--	g11820 = NOT(I14644)
--	g33936 = NOT(I31820)
--	g8456 = NOT(g56)
--	g12880 = NOT(g10387)
--	I22131 = NOT(g19984)
--	I24078 = NOT(g22360)
--	g23789 = NOT(g21308)
--	I17839 = NOT(g13412)
--	g32192 = NOT(g31262)
--	I33109 = NOT(g34851)
--	I15846 = NOT(g11183)
--	I16357 = NOT(g884)
--	I25359 = NOT(g24715)
--	I19799 = NOT(g17817)
--	g30312 = NOT(g28970)
--	I12189 = NOT(g5869)
--	I19813 = NOT(g17952)
--	g24368 = NOT(g22228)
--	g21724 = NOT(I21291)
--	g23788 = NOT(g18997)
--	g8155 = NOT(g3380)
--	g34312 = NOT(g34098)
--	g26973 = NOT(g26105)
--	g34200 = NOT(g33895)
--	g7224 = NOT(g4601)
--	g32522 = NOT(g30735)
--	g23359 = NOT(I22458)
--	g32663 = NOT(g30673)
--	g8355 = NOT(I12534)
--	g8851 = NOT(g590)
--	I13057 = NOT(g112)
--	g14451 = NOT(I16606)
--	I23366 = NOT(g23321)
--	I18364 = NOT(g13009)
--	I22619 = NOT(g21193)
--	I17131 = NOT(g14384)
--	I22502 = NOT(g19376)
--	g22980 = NOT(I22153)
--	g21434 = NOT(g17248)
--	I22557 = NOT(g20695)
--	g21358 = NOT(g16307)
--	g6839 = NOT(g1858)
--	g23434 = NOT(g21611)
--	g24850 = NOT(I24022)
--	g30052 = NOT(g29018)
--	I19674 = NOT(g15932)
--	g8964 = NOT(g4269)
--	I29913 = NOT(g30605)
--	g27831 = NOT(I26406)
--	I11626 = NOT(g31)
--	g11413 = NOT(g9100)
--	g34921 = NOT(I33155)
--	g13413 = NOT(g11737)
--	g34052 = NOT(g33635)
--	g23946 = NOT(g19210)
--	g24133 = NOT(g19935)
--	g29169 = NOT(g27886)
--	g18096 = NOT(I18894)
--	g18944 = NOT(g15938)
--	g20229 = NOT(g17015)
--	g32483 = NOT(g30673)
--	g19617 = NOT(g16349)
--	g19470 = NOT(g16000)
--	g22181 = NOT(g19277)
--	g11691 = NOT(I14570)
--	g19915 = NOT(g16349)
--	g12831 = NOT(g9569)
--	g26732 = NOT(g25389)
--	I16803 = NOT(g6369)
--	I12030 = NOT(g595)
--	I17557 = NOT(g14510)
--	g9541 = NOT(g2012)
--	g32553 = NOT(g31170)
--	g32862 = NOT(g30825)
--	g7617 = NOT(I12089)
--	g16726 = NOT(g14454)
--	I26649 = NOT(g27675)
--	g34813 = NOT(I33027)
--	g10776 = NOT(I14033)
--	g19277 = NOT(I19813)
--	g32949 = NOT(g30825)
--	g9332 = NOT(g64)
--	g14591 = NOT(I16709)
--	g14785 = NOT(g12629)
--	I21226 = NOT(g16540)
--	I22286 = NOT(g19446)
--	g7516 = NOT(I12003)
--	g21682 = NOT(g16540)
--	I18224 = NOT(g13793)
--	g9680 = NOT(I13276)
--	g9153 = NOT(I12991)
--	g10147 = NOT(g728)
--	g20716 = NOT(g15277)
--	g27989 = NOT(g26759)
--	g29217 = NOT(I27567)
--	g34973 = NOT(I33235)
--	g25554 = NOT(g22550)
--	I15929 = NOT(g10430)
--	I18571 = NOT(g13074)
--	g21291 = NOT(g16620)
--	g32536 = NOT(g31376)
--	g14147 = NOT(I16357)
--	g30184 = NOT(g28144)
--	I31796 = NOT(g33176)
--	g10355 = NOT(g6816)
--	g32948 = NOT(g30735)
--	g23291 = NOT(g21070)
--	g16607 = NOT(g13960)
--	g19494 = NOT(g16349)
--	g11929 = NOT(I14745)
--	I11737 = NOT(g4467)
--	g34674 = NOT(I32806)
--	g8279 = NOT(I12487)
--	g16320 = NOT(g14454)
--	g20582 = NOT(g17873)
--	g32702 = NOT(g30735)
--	g9744 = NOT(g6486)
--	g10370 = NOT(g7095)
--	g31000 = NOT(g29737)
--	g32757 = NOT(g30937)
--	g32904 = NOT(g30735)
--	g6988 = NOT(g4765)
--	I14866 = NOT(g9748)
--	g16530 = NOT(g14454)
--	g26400 = NOT(I25351)
--	g11928 = NOT(I14742)
--	g25115 = NOT(I24281)
--	g13583 = NOT(I16028)
--	g32621 = NOT(g31542)
--	g8872 = NOT(g4258)
--	g22520 = NOT(g19801)
--	I22601 = NOT(g21127)
--	g10151 = NOT(g1992)
--	g28120 = NOT(g27108)
--	I32228 = NOT(g34122)
--	I11697 = NOT(g3352)
--	g10172 = NOT(g6459)
--	g20627 = NOT(g17433)
--	I12837 = NOT(g4222)
--	g7892 = NOT(g4801)
--	g34934 = NOT(g34918)
--	g9558 = NOT(g5841)
--	g20379 = NOT(g17821)
--	g8057 = NOT(g3068)
--	g32564 = NOT(g31376)
--	I13995 = NOT(g8744)
--	g24379 = NOT(g22550)
--	g8457 = NOT(g225)
--	g8989 = NOT(I12935)
--	g19352 = NOT(g15758)
--	g22546 = NOT(I21918)
--	g23760 = NOT(I22889)
--	g20050 = NOT(I20321)
--	g23029 = NOT(g20453)
--	g6804 = NOT(g490)
--	g24112 = NOT(g19935)
--	g10367 = NOT(g6870)
--	g10394 = NOT(g6994)
--	I25028 = NOT(g24484)
--	g24050 = NOT(g20841)
--	g9901 = NOT(g84)
--	g34692 = NOT(I32846)
--	I22143 = NOT(g20189)
--	I21784 = NOT(g19638)
--	g23506 = NOT(g21514)
--	g23028 = NOT(g20391)
--	I18752 = NOT(g6358)
--	I28480 = NOT(g28652)
--	g31814 = NOT(g29385)
--	g32673 = NOT(g31376)
--	g32847 = NOT(g30735)
--	g20386 = NOT(g15224)
--	I21297 = NOT(g18597)
--	g8971 = NOT(I12927)
--	g22860 = NOT(g20000)
--	g24386 = NOT(g22594)
--	g20603 = NOT(g17873)
--	g9511 = NOT(g5881)
--	g27736 = NOT(I26356)
--	g7738 = NOT(I12176)
--	g31807 = NOT(g29385)
--	g8686 = NOT(g2819)
--	g13302 = NOT(g12321)
--	g20096 = NOT(g16782)
--	g24603 = NOT(g23108)
--	g33772 = NOT(I31622)
--	g7991 = NOT(g4878)
--	I23354 = NOT(g23277)
--	g24096 = NOT(g19890)
--	g29922 = NOT(g28837)
--	g34400 = NOT(g34142)
--	g7244 = NOT(g4408)
--	g12887 = NOT(g10394)
--	g10420 = NOT(g9239)
--	I17143 = NOT(g14412)
--	g22497 = NOT(g19513)
--	g25184 = NOT(g22763)
--	g32509 = NOT(g31070)
--	g31639 = NOT(I29225)
--	g10319 = NOT(I13740)
--	g17088 = NOT(I18160)
--	g32933 = NOT(g31376)
--	g30329 = NOT(I28588)
--	g9492 = NOT(g2759)
--	I21181 = NOT(g17413)
--	g16136 = NOT(I17491)
--	g7340 = NOT(g4443)
--	g20681 = NOT(g15483)
--	g9600 = NOT(g3632)
--	I23671 = NOT(g23202)
--	g32508 = NOT(g30825)
--	g9574 = NOT(g6462)
--	g31638 = NOT(g29689)
--	g9864 = NOT(I13424)
--	g32634 = NOT(g30673)
--	g32851 = NOT(g31327)
--	g32872 = NOT(g31327)
--	g33638 = NOT(I31469)
--	g35001 = NOT(I33297)
--	g30328 = NOT(I28585)
--	g7907 = NOT(g3072)
--	g11640 = NOT(I14550)
--	g11769 = NOT(g8626)
--	g34539 = NOT(g34354)
--	g9714 = NOT(g4012)
--	g12843 = NOT(g10359)
--	g17497 = NOT(g14879)
--	g22987 = NOT(g20391)
--	g34328 = NOT(g34096)
--	g10059 = NOT(g6451)
--	g23927 = NOT(g19074)
--	I18842 = NOT(g13809)
--	g24429 = NOT(g22722)
--	g19524 = NOT(g15695)
--	I29891 = NOT(g31578)
--	g7517 = NOT(g962)
--	g22658 = NOT(I21969)
--	g29953 = NOT(g28907)
--	g10540 = NOT(g9392)
--	g10058 = NOT(g6497)
--	g31841 = NOT(g29385)
--	g24428 = NOT(g22722)
--	I32096 = NOT(g33641)
--	g33391 = NOT(g32384)
--	g19477 = NOT(g16431)
--	g12869 = NOT(g10376)
--	g16164 = NOT(I17507)
--	g23649 = NOT(g18833)
--	g26683 = NOT(g25514)
--	g7876 = NOT(g1495)
--	g25692 = NOT(I24839)
--	g15614 = NOT(g14914)
--	g22339 = NOT(g19801)
--	g20765 = NOT(g17748)
--	g8938 = NOT(g4899)
--	I19235 = NOT(g15078)
--	I20495 = NOT(g16283)
--	g29800 = NOT(g28363)
--	g10203 = NOT(g2393)
--	g12868 = NOT(g10377)
--	g21903 = NOT(I21480)
--	g14203 = NOT(g12381)
--	g20549 = NOT(g15277)
--	g23648 = NOT(g18833)
--	g13881 = NOT(I16181)
--	I16090 = NOT(g10430)
--	g22338 = NOT(g19801)
--	g23491 = NOT(g21514)
--	I20816 = NOT(g17088)
--	g23903 = NOT(g18997)
--	I33252 = NOT(g34974)
--	I32681 = NOT(g34429)
--	g10044 = NOT(g5357)
--	g34241 = NOT(I32222)
--	g27709 = NOT(I26337)
--	g21604 = NOT(g15938)
--	I22580 = NOT(g20982)
--	I16651 = NOT(g10542)
--	g20548 = NOT(g15426)
--	g8519 = NOT(g287)
--	g8740 = NOT(I12735)
--	g31578 = NOT(I29199)
--	g25013 = NOT(g23599)
--	g31835 = NOT(g29385)
--	g32574 = NOT(g31070)
--	I20985 = NOT(g16300)
--	g24548 = NOT(g22942)
--	I31564 = NOT(g33204)
--	g17296 = NOT(I18280)
--	g25214 = NOT(g22228)
--	g27708 = NOT(I26334)
--	I12418 = NOT(g55)
--	g17644 = NOT(g15002)
--	g20504 = NOT(g18008)
--	g30100 = NOT(g29131)
--	g23563 = NOT(g20682)
--	g10377 = NOT(g6940)
--	g32912 = NOT(g30735)
--	g8606 = NOT(g4653)
--	I18865 = NOT(g14314)
--	I20954 = NOT(g16228)
--	g19748 = NOT(g17015)
--	g10120 = NOT(g1902)
--	g22197 = NOT(g19074)
--	g14377 = NOT(g12201)
--	I11753 = NOT(g4492)
--	g22855 = NOT(g20391)
--	g19276 = NOT(g17367)
--	g9889 = NOT(g6128)
--	g13027 = NOT(I15647)
--	g7110 = NOT(g6682)
--	I14660 = NOT(g9746)
--	g33442 = NOT(g31937)
--	g22870 = NOT(g20887)
--	g22527 = NOT(g19546)
--	I21860 = NOT(g19638)
--	g34683 = NOT(I32827)
--	g28127 = NOT(g27102)
--	g25538 = NOT(g22594)
--	g29216 = NOT(I27564)
--	I32690 = NOT(g34432)
--	g11249 = NOT(g8405)
--	I28838 = NOT(g29372)
--	I13031 = NOT(g6747)
--	g14738 = NOT(I16821)
--	g13249 = NOT(g10590)
--	g14562 = NOT(g12036)
--	g14645 = NOT(I16755)
--	I30861 = NOT(g32383)
--	g20129 = NOT(g17328)
--	g16606 = NOT(g14110)
--	g17197 = NOT(I18233)
--	g18880 = NOT(g15656)
--	g23767 = NOT(g18997)
--	g23794 = NOT(g19147)
--	g21395 = NOT(g17873)
--	g24129 = NOT(g20857)
--	g32592 = NOT(g30673)
--	g20057 = NOT(g16349)
--	g32756 = NOT(g31021)
--	g23395 = NOT(I22502)
--	g24057 = NOT(g20841)
--	g20128 = NOT(g17533)
--	I12167 = NOT(g5176)
--	g14290 = NOT(I16460)
--	g17870 = NOT(I18842)
--	g17411 = NOT(g14454)
--	g17527 = NOT(g14741)
--	g23899 = NOT(g19277)
--	g7002 = NOT(g5160)
--	g13003 = NOT(I15609)
--	g24128 = NOT(g20720)
--	g11204 = NOT(I14271)
--	I14550 = NOT(g10072)
--	g7824 = NOT(g4169)
--	g30991 = NOT(I28925)
--	g6996 = NOT(g4955)
--	g25241 = NOT(g23651)
--	g11779 = NOT(g9602)
--	I18270 = NOT(g13191)
--	g16750 = NOT(g14454)
--	g22867 = NOT(g20391)
--	g34991 = NOT(I33273)
--	g7236 = NOT(g4608)
--	g9285 = NOT(g2715)
--	g20626 = NOT(g15483)
--	g27774 = NOT(I26381)
--	I27401 = NOT(g27051)
--	I11843 = NOT(g111)
--	g23898 = NOT(g19277)
--	g9500 = NOT(g5495)
--	g20323 = NOT(g17873)
--	I21250 = NOT(g16540)
--	g29117 = NOT(g27886)
--	g24626 = NOT(g23139)
--	g33430 = NOT(g32421)
--	g23191 = NOT(I22289)
--	g20533 = NOT(g17271)
--	g10427 = NOT(g10053)
--	g12955 = NOT(I15577)
--	g32820 = NOT(g31672)
--	I18460 = NOT(g5276)
--	g8341 = NOT(g3119)
--	g10366 = NOT(g6895)
--	g24533 = NOT(g22876)
--	g25100 = NOT(g22384)
--	g12879 = NOT(g10381)
--	g22714 = NOT(g20436)
--	g11786 = NOT(g7549)
--	g14366 = NOT(I16526)
--	g17503 = NOT(g14892)
--	I14054 = NOT(g10028)
--	g9184 = NOT(g6120)
--	g23521 = NOT(g21468)
--	g28181 = NOT(I26700)
--	g25771 = NOT(I24920)
--	g20775 = NOT(g18008)
--	g18831 = NOT(g15224)
--	I15647 = NOT(g12109)
--	I23339 = NOT(g23232)
--	g32846 = NOT(g31376)
--	g9339 = NOT(g2295)
--	I19759 = NOT(g17767)
--	g19733 = NOT(g16856)
--	I24558 = NOT(g23777)
--	g12878 = NOT(g10386)
--	g26758 = NOT(g25389)
--	I27749 = NOT(g28917)
--	I20830 = NOT(g17657)
--	g12337 = NOT(g9340)
--	g32731 = NOT(g31376)
--	g31806 = NOT(g29385)
--	g22202 = NOT(I21784)
--	g33806 = NOT(I31650)
--	g9024 = NOT(g4358)
--	I12749 = NOT(g4575)
--	g11826 = NOT(I14650)
--	g17714 = NOT(g14930)
--	g12886 = NOT(g10393)
--	g22979 = NOT(g20453)
--	g20737 = NOT(g15656)
--	g22496 = NOT(g19510)
--	g10403 = NOT(g7040)
--	I21969 = NOT(g21370)
--	g23440 = NOT(I22557)
--	g13999 = NOT(g11048)
--	g7222 = NOT(g4427)
--	g27967 = NOT(I26479)
--	g27994 = NOT(g26793)
--	g33142 = NOT(g32072)
--	g19630 = NOT(g16897)
--	g9809 = NOT(g6082)
--	g20232 = NOT(g16931)
--	I14773 = NOT(g9581)
--	g29814 = NOT(I28062)
--	g17819 = NOT(I18825)
--	g17707 = NOT(g14758)
--	I33047 = NOT(g34776)
--	g30206 = NOT(g28436)
--	g7928 = NOT(g4776)
--	g26744 = NOT(g25400)
--	g12967 = NOT(g11790)
--	g23861 = NOT(g19147)
--	g23573 = NOT(g20248)
--	g32691 = NOT(g30673)
--	g18989 = NOT(g16000)
--	g8879 = NOT(I12858)
--	g8607 = NOT(g37)
--	g11233 = NOT(g9664)
--	I18875 = NOT(g13782)
--	g21247 = NOT(g15171)
--	g23247 = NOT(g20924)
--	g11182 = NOT(I14241)
--	I11708 = NOT(g3703)
--	g7064 = NOT(g5990)
--	g17818 = NOT(I18822)
--	g9672 = NOT(g5390)
--	I13708 = NOT(g136)
--	g20697 = NOT(g17433)
--	g14226 = NOT(g11618)
--	g9077 = NOT(g504)
--	g17496 = NOT(g14683)
--	I19345 = NOT(g15083)
--	g22986 = NOT(g20330)
--	g8659 = NOT(g2815)
--	g25882 = NOT(g25026)
--	g23926 = NOT(g19074)
--	g8358 = NOT(I12541)
--	g18988 = NOT(g15979)
--	I32775 = NOT(g34512)
--	g9477 = NOT(I13149)
--	g8506 = NOT(g3782)
--	I30766 = NOT(g32363)
--	g9523 = NOT(g6419)
--	g24995 = NOT(g22763)
--	g34759 = NOT(I32935)
--	g7785 = NOT(g4621)
--	g16522 = NOT(g13889)
--	g23612 = NOT(I22745)
--	g10572 = NOT(g10233)
--	I25534 = NOT(g25448)
--	I17964 = NOT(g3661)
--	g23388 = NOT(g21070)
--	I15932 = NOT(g12381)
--	g17590 = NOT(I18523)
--	g19476 = NOT(g16326)
--	g12919 = NOT(I15536)
--	I12808 = NOT(g4322)
--	g6799 = NOT(g199)
--	g26804 = NOT(g25400)
--	g20512 = NOT(g18062)
--	g34435 = NOT(I32476)
--	g23777 = NOT(I22918)
--	g23534 = NOT(I22665)
--	I26451 = NOT(g26862)
--	g13932 = NOT(g11534)
--	g32929 = NOT(g31710)
--	g8587 = NOT(g3689)
--	I14839 = NOT(g9689)
--	g23272 = NOT(g20924)
--	g11513 = NOT(g7948)
--	g19454 = NOT(g16349)
--	g7563 = NOT(g6322)
--	g17741 = NOT(g12972)
--	g12918 = NOT(I15533)
--	I18160 = NOT(g14441)
--	I15448 = NOT(g10877)
--	g17384 = NOT(I18323)
--	g32583 = NOT(g30614)
--	g32928 = NOT(g31672)
--	g19570 = NOT(g16349)
--	g19712 = NOT(g17096)
--	g6997 = NOT(g4578)
--	g22150 = NOT(g21280)
--	g11897 = NOT(I14705)
--	I22000 = NOT(g20277)
--	g10490 = NOT(g9274)
--	g9551 = NOT(g3281)
--	g9742 = NOT(g6144)
--	g9104 = NOT(I12987)
--	g23462 = NOT(I22589)
--	g9099 = NOT(g3706)
--	g34345 = NOT(I32352)
--	g9499 = NOT(g5152)
--	g11404 = NOT(g7596)
--	g15750 = NOT(g13291)
--	g34940 = NOT(g34924)
--	g13505 = NOT(g10981)
--	I15717 = NOT(g6346)
--	g16326 = NOT(I17658)
--	g18887 = NOT(g15373)
--	g20445 = NOT(g15224)
--	I31820 = NOT(g33323)
--	I12064 = NOT(g617)
--	g23032 = NOT(I22211)
--	g10376 = NOT(g6923)
--	g10385 = NOT(I13805)
--	g25206 = NOT(g23613)
--	g12598 = NOT(g7004)
--	g14376 = NOT(g12126)
--	g14385 = NOT(I16541)
--	g34848 = NOT(I33070)
--	g19074 = NOT(I19772)
--	g17735 = NOT(g14807)
--	g14297 = NOT(g10869)
--	g20499 = NOT(g15483)
--	g7394 = NOT(g5637)
--	g10980 = NOT(g9051)
--	g11026 = NOT(g8434)
--	I26785 = NOT(g27013)
--	g12086 = NOT(g9654)
--	g32787 = NOT(g30937)
--	g13026 = NOT(g11018)
--	g31863 = NOT(I29447)
--	I14619 = NOT(g4185)
--	g10354 = NOT(g6811)
--	I23315 = NOT(g21685)
--	I33152 = NOT(g34900)
--	g19567 = NOT(g16164)
--	g14095 = NOT(g11326)
--	g29014 = NOT(g27742)
--	g22526 = NOT(g19801)
--	I17569 = NOT(g14564)
--	g9754 = NOT(g2020)
--	g21061 = NOT(I20929)
--	g28126 = NOT(g27122)
--	g18528 = NOT(I19348)
--	g20498 = NOT(g15348)
--	g6802 = NOT(g468)
--	g8284 = NOT(g5002)
--	g23061 = NOT(g20283)
--	g8239 = NOT(g1056)
--	g28250 = NOT(g27074)
--	g10181 = NOT(g2551)
--	g25114 = NOT(I24278)
--	g7557 = NOT(g1500)
--	g8180 = NOT(g262)
--	I17747 = NOT(g13298)
--	g12322 = NOT(I15162)
--	g27977 = NOT(g26105)
--	g32743 = NOT(g30937)
--	g32827 = NOT(g31672)
--	g25082 = NOT(g22342)
--	g8591 = NOT(g3763)
--	g30332 = NOT(I28597)
--	g24056 = NOT(g20014)
--	g9613 = NOT(g5062)
--	g12901 = NOT(g10404)
--	g20611 = NOT(g18008)
--	g17526 = NOT(I18469)
--	g12977 = NOT(I15590)
--	g20080 = NOT(g17328)
--	g7471 = NOT(g6012)
--	g9044 = NOT(g604)
--	g20924 = NOT(I20895)
--	g19519 = NOT(g16795)
--	g24080 = NOT(g21143)
--	g19675 = NOT(g16987)
--	g9444 = NOT(g5535)
--	g9269 = NOT(g5517)
--	g22866 = NOT(g20330)
--	I17814 = NOT(g3274)
--	g32640 = NOT(g31154)
--	g20432 = NOT(g17847)
--	g32769 = NOT(g31672)
--	g23360 = NOT(I22461)
--	g29116 = NOT(g27837)
--	g19518 = NOT(g16239)
--	g8507 = NOT(g3712)
--	g9983 = NOT(g4239)
--	g12656 = NOT(g7028)
--	I15620 = NOT(g12038)
--	I17772 = NOT(g14888)
--	g25849 = NOT(g24491)
--	g9862 = NOT(g5413)
--	I27555 = NOT(g28142)
--	g23447 = NOT(g21562)
--	g32768 = NOT(g30825)
--	g32803 = NOT(g31376)
--	g25399 = NOT(g22763)
--	g12295 = NOT(g7139)
--	I23384 = NOT(g23362)
--	g10190 = NOT(g6044)
--	g29041 = NOT(I27385)
--	g13620 = NOT(g10556)
--	g12823 = NOT(g9206)
--	I17639 = NOT(g13350)
--	I27570 = NOT(g28262)
--	I15811 = NOT(g11128)
--	I21067 = NOT(g15573)
--	I18822 = NOT(g13745)
--	g16509 = NOT(g13873)
--	I32056 = NOT(g33641)
--	g11811 = NOT(g9724)
--	I12712 = NOT(g59)
--	g20145 = NOT(g17533)
--	g34833 = NOT(I33047)
--	g34049 = NOT(g33678)
--	I13010 = NOT(g6749)
--	g31821 = NOT(g29385)
--	g32881 = NOT(g30673)
--	I32988 = NOT(g34755)
--	g24031 = NOT(g21193)
--	I33020 = NOT(g34781)
--	g16508 = NOT(I17704)
--	I24455 = NOT(g22541)
--	g26605 = NOT(g25293)
--	g20650 = NOT(g15348)
--	g23629 = NOT(g21514)
--	g21451 = NOT(I21162)
--	g16872 = NOT(I18060)
--	I12907 = NOT(g4322)
--	g22923 = NOT(I22124)
--	I17416 = NOT(g13806)
--	g23472 = NOT(g21062)
--	g15483 = NOT(I17128)
--	g9534 = NOT(g90)
--	g9729 = NOT(g5138)
--	g9961 = NOT(g6404)
--	g7438 = NOT(g5983)
--	g25263 = NOT(g22763)
--	g29983 = NOT(g28977)
--	g20529 = NOT(g15509)
--	g22300 = NOT(I21815)
--	g26812 = NOT(g25439)
--	I21019 = NOT(g17325)
--	g27017 = NOT(g25895)
--	I27567 = NOT(g28181)
--	g15862 = NOT(I17355)
--	g8515 = NOT(I12631)
--	g34221 = NOT(I32192)
--	g8630 = NOT(g4843)
--	g21246 = NOT(I20985)
--	I27238 = NOT(g27320)
--	g23246 = NOT(g20785)
--	g20528 = NOT(g15224)
--	g20696 = NOT(g17533)
--	g25135 = NOT(g22457)
--	g20330 = NOT(I20542)
--	g9927 = NOT(g5689)
--	g32662 = NOT(g30614)
--	g8300 = NOT(g1242)
--	g32027 = NOT(I29585)
--	I32461 = NOT(g34244)
--	g19577 = NOT(g16129)
--	g17688 = NOT(I18667)
--	g9014 = NOT(g3004)
--	g20764 = NOT(I20819)
--	g10497 = NOT(g10102)
--	I25591 = NOT(g25380)
--	g32890 = NOT(g30735)
--	I33282 = NOT(g34987)
--	I27941 = NOT(g28803)
--	g9414 = NOT(g2004)
--	g7212 = NOT(g6411)
--	g19439 = NOT(g15885)
--	g9660 = NOT(g3267)
--	g9946 = NOT(g6093)
--	g20132 = NOT(g16931)
--	g24365 = NOT(g22594)
--	g20869 = NOT(g15615)
--	g13412 = NOT(g11963)
--	g23776 = NOT(g21177)
--	g34947 = NOT(g34938)
--	I12382 = NOT(g47)
--	g24132 = NOT(g19890)
--	g32482 = NOT(g30614)
--	g24869 = NOT(I24041)
--	g24960 = NOT(g23716)
--	g19438 = NOT(g16249)
--	I12519 = NOT(g3447)
--	g17157 = NOT(g13350)
--	I12176 = NOT(g5523)
--	g9903 = NOT(g681)
--	g13133 = NOT(g11330)
--	g32710 = NOT(g30825)
--	I12092 = NOT(g790)
--	g14700 = NOT(g12512)
--	g21355 = NOT(g17821)
--	g32552 = NOT(g30825)
--	g31834 = NOT(g29385)
--	g23355 = NOT(g21070)
--	g34812 = NOT(I33024)
--	g10658 = NOT(I13979)
--	g21370 = NOT(g16323)
--	g23859 = NOT(g19074)
--	g28819 = NOT(I27271)
--	g16311 = NOT(g13273)
--	g32779 = NOT(g30937)
--	I17442 = NOT(g13638)
--	g18878 = NOT(g15426)
--	g24161 = NOT(I23327)
--	g29130 = NOT(g27907)
--	I32696 = NOT(g34434)
--	I32843 = NOT(g34499)
--	g7993 = NOT(I12333)
--	g20709 = NOT(g15426)
--	g11011 = NOT(g10274)
--	g22854 = NOT(g20330)
--	g34951 = NOT(g34941)
--	g34972 = NOT(I33232)
--	g23858 = NOT(g18997)
--	g13011 = NOT(I15623)
--	I12935 = NOT(g6753)
--	g32778 = NOT(g31021)
--	g18886 = NOT(g16000)
--	I31803 = NOT(g33176)
--	g9036 = NOT(g5084)
--	I18313 = NOT(g13350)
--	g25221 = NOT(g23653)
--	I22275 = NOT(g20127)
--	g8440 = NOT(g3431)
--	g20708 = NOT(g15426)
--	g22763 = NOT(I22046)
--	g9679 = NOT(g5475)
--	g23172 = NOT(I22275)
--	g13716 = NOT(I16090)
--	I17615 = NOT(g13251)
--	g20087 = NOT(g17249)
--	g32786 = NOT(g31021)
--	g33726 = NOT(I31581)
--	I32960 = NOT(g34653)
--	g8123 = NOT(g3808)
--	g19566 = NOT(g16136)
--	g14338 = NOT(I16502)
--	g24087 = NOT(g21143)
--	I18276 = NOT(g1075)
--	I18285 = NOT(g13638)
--	g28590 = NOT(g27724)
--	g23844 = NOT(g21308)
--	g32647 = NOT(g31154)
--	g23394 = NOT(I22499)
--	I32868 = NOT(g34579)
--	g9831 = NOT(g2269)
--	g32945 = NOT(g30937)
--	g33436 = NOT(I30962)
--	g22660 = NOT(g19140)
--	g15509 = NOT(I17136)
--	I19012 = NOT(g15060)
--	g17763 = NOT(g15011)
--	g8666 = NOT(g3703)
--	g10060 = NOT(g6541)
--	I18900 = NOT(g16767)
--	g27976 = NOT(g26703)
--	g27985 = NOT(g26131)
--	I32161 = NOT(g33791)
--	g32826 = NOT(g30825)
--	g25273 = NOT(g23978)
--	g29863 = NOT(g28410)
--	g24043 = NOT(g20982)
--	g10197 = NOT(g31)
--	I21300 = NOT(g18598)
--	g22456 = NOT(g19801)
--	g12976 = NOT(I15587)
--	g15634 = NOT(I17188)
--	I23688 = NOT(g23244)
--	I23300 = NOT(g21665)
--	g14197 = NOT(g12160)
--	g32090 = NOT(g31003)
--	g9805 = NOT(g5485)
--	g9916 = NOT(g3625)
--	g19653 = NOT(g16897)
--	g33346 = NOT(g32132)
--	I18101 = NOT(g13416)
--	I32225 = NOT(g34121)
--	g10527 = NOT(I13892)
--	I12577 = NOT(g1227)
--	g10411 = NOT(g7086)
--	g23420 = NOT(g21514)
--	g9749 = NOT(g1691)
--	I18177 = NOT(g13191)
--	I18560 = NOT(g5969)
--	g32651 = NOT(g31376)
--	g18918 = NOT(I19704)
--	g32672 = NOT(g31579)
--	I19789 = NOT(g17793)
--	g24069 = NOT(g19968)
--	g22550 = NOT(I21922)
--	I33027 = NOT(g34767)
--	g26788 = NOT(g25349)
--	g26724 = NOT(g25341)
--	g20657 = NOT(g17433)
--	g20774 = NOT(g18008)
--	I26427 = NOT(g26859)
--	g8655 = NOT(g2787)
--	g23446 = NOT(g21562)
--	I16057 = NOT(g10430)
--	I28908 = NOT(g30182)
--	g19636 = NOT(g16987)
--	g23227 = NOT(g20924)
--	g30012 = NOT(I28241)
--	g19415 = NOT(g15758)
--	g24068 = NOT(g19919)
--	g24375 = NOT(g22722)
--	g21059 = NOT(g15509)
--	I33249 = NOT(g34971)
--	g7462 = NOT(g2599)
--	g23059 = NOT(g20453)
--	g31797 = NOT(g29385)
--	g6838 = NOT(g1724)
--	g13096 = NOT(I15727)
--	g33641 = NOT(I31474)
--	g32932 = NOT(g31327)
--	g33797 = NOT(g33306)
--	I31482 = NOT(g33204)
--	g19852 = NOT(g17015)
--	g22721 = NOT(I22028)
--	g10503 = NOT(g8879)
--	I16626 = NOT(g11986)
--	g21058 = NOT(g15426)
--	g6809 = NOT(g341)
--	g32513 = NOT(g31376)
--	I20864 = NOT(g16960)
--	g23058 = NOT(g20453)
--	g32449 = NOT(I29977)
--	g14503 = NOT(g12256)
--	g16691 = NOT(g14160)
--	I24022 = NOT(g22182)
--	g19963 = NOT(g16326)
--	g12842 = NOT(g10355)
--	g34473 = NOT(g34426)
--	I12083 = NOT(g568)
--	g17085 = NOT(g14238)
--	I31779 = NOT(g33212)
--	g24171 = NOT(I23357)
--	g32897 = NOT(g30735)
--	g32961 = NOT(g31376)
--	g23203 = NOT(g20073)
--	g8839 = NOT(I12819)
--	g34789 = NOT(I32997)
--	g7788 = NOT(g4674)
--	g11429 = NOT(g7616)
--	g17721 = NOT(g12915)
--	g29372 = NOT(I27738)
--	g10581 = NOT(g9529)
--	I16775 = NOT(g12183)
--	g13857 = NOT(I16163)
--	g32505 = NOT(g31566)
--	g20994 = NOT(g15615)
--	g9095 = NOT(g3368)
--	g32404 = NOT(I29936)
--	I14800 = NOT(g10107)
--	g33136 = NOT(g32057)
--	g9037 = NOT(g164)
--	g14714 = NOT(g11405)
--	g33635 = NOT(g33436)
--	g24994 = NOT(g22432)
--	g14315 = NOT(I16479)
--	g30325 = NOT(I28576)
--	g34788 = NOT(I32994)
--	g11793 = NOT(I14633)
--	g11428 = NOT(g7615)
--	g26682 = NOT(g25309)
--	g9653 = NOT(g2441)
--	g17431 = NOT(I18376)
--	g13793 = NOT(I16120)
--	g22341 = NOT(g19801)
--	g32717 = NOT(g30735)
--	g34325 = NOT(g34092)
--	I15765 = NOT(g10823)
--	I18009 = NOT(g13680)
--	g21281 = NOT(g16286)
--	g18977 = NOT(g16100)
--	I31786 = NOT(g33197)
--	I32970 = NOT(g34716)
--	g22156 = NOT(g19147)
--	g27830 = NOT(g26802)
--	g21902 = NOT(I21477)
--	g34920 = NOT(I33152)
--	g8172 = NOT(g3873)
--	g8278 = NOT(g3096)
--	g34434 = NOT(I32473)
--	g23902 = NOT(g21468)
--	g23301 = NOT(g21037)
--	g34358 = NOT(I32364)
--	g28917 = NOT(I27314)
--	g23377 = NOT(g21070)
--	I32878 = NOT(g34501)
--	g22180 = NOT(g19210)
--	g24425 = NOT(g22722)
--	g19554 = NOT(g16861)
--	g10111 = NOT(g1858)
--	g12830 = NOT(g9995)
--	g12893 = NOT(g10391)
--	I11816 = NOT(g93)
--	g16583 = NOT(g14069)
--	g7392 = NOT(g4438)
--	g20919 = NOT(g15224)
--	g15756 = NOT(g13315)
--	I25146 = NOT(g24911)
--	g34946 = NOT(g34934)
--	I25562 = NOT(g25250)
--	g19609 = NOT(g16264)
--	g8235 = NOT(I12463)
--	g8343 = NOT(g3447)
--	I18476 = NOT(g14031)
--	g34121 = NOT(I32056)
--	I14964 = NOT(g10230)
--	g19200 = NOT(I19789)
--	g21562 = NOT(I21199)
--	g9752 = NOT(g1840)
--	g12865 = NOT(g10372)
--	g20010 = NOT(g17226)
--	g8282 = NOT(g3841)
--	g20918 = NOT(g15224)
--	g23645 = NOT(g20875)
--	g8566 = NOT(g3831)
--	I18555 = NOT(g5630)
--	g24010 = NOT(g21562)
--	g9917 = NOT(I13473)
--	I32967 = NOT(g34648)
--	I32994 = NOT(g34739)
--	g10741 = NOT(g8411)
--	I21480 = NOT(g18696)
--	g7854 = NOT(g1152)
--	g13504 = NOT(g11303)
--	g25541 = NOT(g22763)
--	g20545 = NOT(g15373)
--	g20079 = NOT(g17328)
--	g20444 = NOT(g15373)
--	g21290 = NOT(I21029)
--	g32723 = NOT(g31327)
--	I31672 = NOT(g33149)
--	g10384 = NOT(I13802)
--	g8134 = NOT(I12415)
--	g23290 = NOT(g20924)
--	I33182 = NOT(g34910)
--	I13374 = NOT(g6490)
--	g8334 = NOT(g3034)
--	g24079 = NOT(g20998)
--	g21698 = NOT(g18562)
--	g14384 = NOT(I16538)
--	g22667 = NOT(g21156)
--	g34682 = NOT(I32824)
--	g29209 = NOT(I27543)
--	g20599 = NOT(g18065)
--	g6926 = NOT(g3853)
--	I16512 = NOT(g12811)
--	g23698 = NOT(g21611)
--	I12415 = NOT(g48)
--	g11317 = NOT(I14346)
--	g20078 = NOT(g16846)
--	I12333 = NOT(g45)
--	g32433 = NOT(I29961)
--	g19745 = NOT(g16877)
--	g24078 = NOT(g20857)
--	g6754 = NOT(I11617)
--	g12705 = NOT(g7051)
--	g20598 = NOT(g17929)
--	g32620 = NOT(g30673)
--	I28579 = NOT(g29474)
--	g20086 = NOT(I20355)
--	g19799 = NOT(g17062)
--	g25325 = NOT(g22228)
--	I32458 = NOT(g34243)
--	g11129 = NOT(g7994)
--	I25366 = NOT(g24477)
--	g8804 = NOT(g4035)
--	g10150 = NOT(g1700)
--	g24086 = NOT(g20998)
--	g16743 = NOT(g13986)
--	g21427 = NOT(g17367)
--	g15731 = NOT(g13326)
--	g9364 = NOT(g5041)
--	g10877 = NOT(I14079)
--	g23427 = NOT(I22542)
--	g25535 = NOT(g22763)
--	g32811 = NOT(g30735)
--	I12963 = NOT(g640)
--	g14150 = NOT(g12381)
--	g21366 = NOT(I21100)
--	g32646 = NOT(g31070)
--	g8792 = NOT(I12790)
--	g7219 = NOT(g4405)
--	g19798 = NOT(g17200)
--	I28014 = NOT(g28158)
--	g11128 = NOT(g7993)
--	g7640 = NOT(I12128)
--	I18238 = NOT(g13144)
--	g10019 = NOT(g6479)
--	g28157 = NOT(I26670)
--	I15626 = NOT(g12041)
--	g22210 = NOT(I21792)
--	g20322 = NOT(g17873)
--	g32971 = NOT(g31672)
--	g7431 = NOT(g2555)
--	I32079 = NOT(g33937)
--	g7252 = NOT(g1592)
--	g16640 = NOT(I17834)
--	g29913 = NOT(g28840)
--	g34760 = NOT(I32938)
--	g7812 = NOT(I12214)
--	g16769 = NOT(g13530)
--	g20159 = NOT(g17533)
--	g34134 = NOT(I32079)
--	g25121 = NOT(g22432)
--	g20901 = NOT(I20867)
--	g13626 = NOT(g11273)
--	g20532 = NOT(g15277)
--	g17487 = NOT(I18414)
--	I27576 = NOT(g28173)
--	I15533 = NOT(g11867)
--	g24159 = NOT(I23321)
--	g13323 = NOT(g11048)
--	g24125 = NOT(g19890)
--	g6983 = NOT(g4698)
--	I18382 = NOT(g13350)
--	g21661 = NOT(I21222)
--	g17502 = NOT(g14697)
--	g16768 = NOT(g13223)
--	I19927 = NOT(g17408)
--	g20158 = NOT(g16971)
--	g8113 = NOT(g3466)
--	g12938 = NOT(I15556)
--	I16498 = NOT(g10430)
--	g23403 = NOT(I22512)
--	g23547 = NOT(g21611)
--	g23895 = NOT(g19147)
--	I13424 = NOT(g5689)
--	g24158 = NOT(I23318)
--	g33750 = NOT(I31607)
--	I18092 = NOT(g3668)
--	g7405 = NOT(g1936)
--	g13298 = NOT(I15862)
--	g19732 = NOT(g17096)
--	I22264 = NOT(g20100)
--	I30980 = NOT(g32132)
--	I24008 = NOT(g22182)
--	g29905 = NOT(g28783)
--	g20561 = NOT(g17873)
--	g20656 = NOT(g17249)
--	g9553 = NOT(I13202)
--	I18518 = NOT(g13835)
--	I18154 = NOT(g13177)
--	g23226 = NOT(g20924)
--	g7765 = NOT(g4165)
--	g20680 = NOT(g15348)
--	g26648 = NOT(g25115)
--	g20144 = NOT(g17533)
--	g10402 = NOT(g7023)
--	g23715 = NOT(g20764)
--	g23481 = NOT(I22604)
--	g32850 = NOT(g30937)
--	g31796 = NOT(g29385)
--	g19761 = NOT(g17015)
--	I12608 = NOT(g1582)
--	g12875 = NOT(I15494)
--	I21734 = NOT(g19268)
--	g6961 = NOT(I11734)
--	g8567 = NOT(g4082)
--	I21930 = NOT(g21297)
--	g34927 = NOT(I33173)
--	g7733 = NOT(g4093)
--	I22422 = NOT(g19330)
--	I15697 = NOT(g6000)
--	I17873 = NOT(g15017)
--	g31840 = NOT(g29385)
--	I32158 = NOT(g33791)
--	g12218 = NOT(I15073)
--	g32896 = NOT(g31376)
--	g12837 = NOT(g10354)
--	g23127 = NOT(g21163)
--	g6927 = NOT(g3845)
--	I21838 = NOT(g19263)
--	g25134 = NOT(g22417)
--	g10001 = NOT(g6105)
--	g22975 = NOT(g20391)
--	g13856 = NOT(I16160)
--	I23694 = NOT(g23252)
--	I29248 = NOT(g29491)
--	g9888 = NOT(g5831)
--	g10077 = NOT(g1724)
--	g13995 = NOT(g11261)
--	I33149 = NOT(g34900)
--	g8593 = NOT(g3759)
--	g29153 = NOT(g27937)
--	g24966 = NOT(g22763)
--	g7073 = NOT(g6191)
--	I12799 = NOT(g59)
--	g20631 = NOT(g15171)
--	g17815 = NOT(g14348)
--	g10597 = NOT(g10233)
--	g23490 = NOT(g21514)
--	g25506 = NOT(g22228)
--	g9429 = NOT(g3723)
--	I13705 = NOT(g63)
--	I29204 = NOT(g29505)
--	g32716 = NOT(g31376)
--	g7473 = NOT(g6697)
--	g16249 = NOT(I17590)
--	g18976 = NOT(g16100)
--	g14597 = NOT(I16713)
--	g19539 = NOT(g16129)
--	g6946 = NOT(I11721)
--	g24017 = NOT(g18833)
--	g11512 = NOT(g7634)
--	g34648 = NOT(I32752)
--	g24364 = NOT(g22722)
--	g17677 = NOT(g14882)
--	g34491 = NOT(I32550)
--	I22542 = NOT(g19773)
--	g16482 = NOT(g13464)
--	I17834 = NOT(g14977)
--	g31522 = NOT(I29185)
--	g32582 = NOT(g31170)
--	g7980 = NOT(g3161)
--	g21297 = NOT(I21042)
--	g18954 = NOT(g17427)
--	g23376 = NOT(g21070)
--	g23385 = NOT(I22488)
--	I25095 = NOT(g25265)
--	g19538 = NOT(g16100)
--	g6903 = NOT(g3502)
--	g7069 = NOT(g6137)
--	g9281 = NOT(I13057)
--	I12805 = NOT(g4098)
--	g26990 = NOT(g26105)
--	g34755 = NOT(I32929)
--	g23889 = NOT(g20682)
--	I13124 = NOT(g2729)
--	I18728 = NOT(g6012)
--	I21210 = NOT(g17526)
--	g23354 = NOT(g20453)
--	I14579 = NOT(g8792)
--	g22169 = NOT(g19147)
--	I26700 = NOT(g27956)
--	g34770 = NOT(I32956)
--	g12470 = NOT(I15284)
--	g7540 = NOT(I12026)
--	g8160 = NOT(g3423)
--	g22884 = NOT(g20453)
--	g34981 = NOT(g34973)
--	g23888 = NOT(g18997)
--	g23824 = NOT(g21271)
--	I15831 = NOT(g10416)
--	g32627 = NOT(g30673)
--	g28307 = NOT(g27306)
--	g32959 = NOT(g30937)
--	g32925 = NOT(g31327)
--	g21181 = NOT(g15426)
--	g22168 = NOT(g19147)
--	g10102 = NOT(g6727)
--	g10157 = NOT(g2036)
--	g31862 = NOT(I29444)
--	g32958 = NOT(g31710)
--	I15316 = NOT(g10087)
--	I19719 = NOT(g17431)
--	g8450 = NOT(g3821)
--	g24023 = NOT(g21127)
--	g26718 = NOT(g25168)
--	I32364 = NOT(g34208)
--	g17791 = NOT(g14950)
--	g20571 = NOT(g15277)
--	g9684 = NOT(g6191)
--	g11316 = NOT(g8967)
--	g9745 = NOT(g6537)
--	g12075 = NOT(I14935)
--	I17436 = NOT(g13416)
--	g28431 = NOT(I26925)
--	g9639 = NOT(g1752)
--	I18906 = NOT(g16963)
--	g9338 = NOT(g1870)
--	g24571 = NOT(g22942)
--	g10231 = NOT(g2661)
--	I18083 = NOT(g13394)
--	g9963 = NOT(g7)
--	I26296 = NOT(g26820)
--	g33326 = NOT(g32318)
--	g17410 = NOT(g12955)
--	I12761 = NOT(g4188)
--	g11498 = NOT(I14475)
--	g34767 = NOT(I32947)
--	g14231 = NOT(g12246)
--	g26832 = NOT(g24850)
--	g34845 = NOT(g34773)
--	g32603 = NOT(g31070)
--	g6831 = NOT(g1413)
--	I22464 = NOT(g21222)
--	g23931 = NOT(g20875)
--	g32742 = NOT(g31021)
--	I29233 = NOT(g30295)
--	g9309 = NOT(g5462)
--	I23306 = NOT(g21673)
--	g30990 = NOT(g29676)
--	I18304 = NOT(g14790)
--	g19771 = NOT(g17096)
--	g25240 = NOT(g23650)
--	g32944 = NOT(g31021)
--	I29182 = NOT(g30012)
--	g29474 = NOT(I27758)
--	g34990 = NOT(I33270)
--	g11989 = NOT(I14839)
--	I25190 = NOT(g25423)
--	g16826 = NOT(I18034)
--	g17479 = NOT(g14855)
--	g21426 = NOT(g15277)
--	g8179 = NOT(g4999)
--	g12037 = NOT(I14893)
--	g20495 = NOT(g17926)
--	g23426 = NOT(I22539)
--	g25903 = NOT(I25005)
--	g27984 = NOT(g26737)
--	I13875 = NOT(g1233)
--	g33702 = NOT(I31545)
--	g9808 = NOT(g5827)
--	g19683 = NOT(g16931)
--	g23190 = NOT(I22286)
--	I16709 = NOT(g10430)
--	g11988 = NOT(I14836)
--	I21815 = NOT(g21308)
--	g17478 = NOT(g14996)
--	g28156 = NOT(I26667)
--	I12013 = NOT(g590)
--	g17015 = NOT(I18143)
--	g32681 = NOT(g30735)
--	I32309 = NOT(g34210)
--	I12214 = NOT(g6561)
--	g16182 = NOT(g13846)
--	g16651 = NOT(g14005)
--	I22153 = NOT(g20014)
--	g23520 = NOT(g21468)
--	g27155 = NOT(g26131)
--	g9759 = NOT(g2265)
--	g18830 = NOT(g18008)
--	I16471 = NOT(g12367)
--	g17486 = NOT(I18411)
--	g7898 = NOT(g4991)
--	g25563 = NOT(g22594)
--	g32802 = NOT(g31327)
--	g32857 = NOT(g30937)
--	g22223 = NOT(g19210)
--	g13271 = NOT(I15834)
--	g34718 = NOT(I32884)
--	g24985 = NOT(g23586)
--	g34521 = NOT(g34270)
--	g32730 = NOT(g31327)
--	g23546 = NOT(g21611)
--	I24215 = NOT(g22360)
--	g32793 = NOT(g31021)
--	I18653 = NOT(g5681)
--	g20374 = NOT(g18065)
--	g23211 = NOT(g21308)
--	I30644 = NOT(g32024)
--	g19882 = NOT(g16540)
--	g19414 = NOT(g16349)
--	g26701 = NOT(g25341)
--	g7245 = NOT(I11896)
--	g17580 = NOT(I18509)
--	g11753 = NOT(g8587)
--	I29961 = NOT(g30984)
--	I12538 = NOT(g58)
--	g26777 = NOT(g25439)
--	g20643 = NOT(g15962)
--	I18138 = NOT(g14277)
--	g9049 = NOT(g640)
--	g23088 = NOT(I22240)
--	g31847 = NOT(g29385)
--	g32765 = NOT(g31327)
--	g19407 = NOT(g16268)
--	g9449 = NOT(g5770)
--	g16449 = NOT(I17679)
--	g11031 = NOT(g8609)
--	g22922 = NOT(g20330)
--	g23860 = NOT(g19074)
--	I15650 = NOT(g12110)
--	g32690 = NOT(g31070)
--	g9575 = NOT(g6509)
--	g32549 = NOT(g31554)
--	I15736 = NOT(g12322)
--	I14684 = NOT(g7717)
--	I18333 = NOT(g1083)
--	g22179 = NOT(g19210)
--	I29717 = NOT(g30931)
--	g25262 = NOT(g22763)
--	I11617 = NOT(g1)
--	g11736 = NOT(g8165)
--	g20669 = NOT(g15426)
--	I17136 = NOT(g14398)
--	g16897 = NOT(I18083)
--	I26503 = NOT(g26811)
--	g34573 = NOT(I32645)
--	g7344 = NOT(g5659)
--	g25899 = NOT(g24997)
--	g13736 = NOT(g11313)
--	g32548 = NOT(g30673)
--	I18852 = NOT(g13716)
--	I32687 = NOT(g34431)
--	g34247 = NOT(I32240)
--	I32976 = NOT(g34699)
--	I32985 = NOT(g34736)
--	g22178 = NOT(g19147)
--	g9498 = NOT(g5101)
--	g6873 = NOT(g3151)
--	g20668 = NOT(g15426)
--	g34926 = NOT(I33170)
--	g32504 = NOT(g30673)
--	g31851 = NOT(g29385)
--	I15843 = NOT(g11181)
--	I32752 = NOT(g34510)
--	g9833 = NOT(g2449)
--	g10287 = NOT(I13715)
--	g7259 = NOT(g4375)
--	g21659 = NOT(g17727)
--	I33050 = NOT(g34777)
--	g14314 = NOT(I16476)
--	g16717 = NOT(g13951)
--	g17531 = NOT(I18476)
--	g12836 = NOT(g10351)
--	g20195 = NOT(g16931)
--	I26581 = NOT(g26942)
--	g8997 = NOT(g577)
--	g23987 = NOT(g19277)
--	g10085 = NOT(g1768)
--	g8541 = NOT(g3498)
--	g23250 = NOT(g21070)
--	g24489 = NOT(I23694)
--	I23363 = NOT(g23385)
--	g14307 = NOT(I16468)
--	I27235 = NOT(g27320)
--	g17178 = NOT(I18214)
--	g6869 = NOT(I11691)
--	g34777 = NOT(I32973)
--	g12477 = NOT(I15295)
--	g20525 = NOT(g17955)
--	I15869 = NOT(g11234)
--	g18939 = NOT(g16077)
--	g8132 = NOT(I12411)
--	g28443 = NOT(I26936)
--	g34272 = NOT(g34229)
--	g24525 = NOT(g22670)
--	g24424 = NOT(g22722)
--	I11623 = NOT(g28)
--	g13132 = NOT(g10632)
--	g17685 = NOT(I18662)
--	g17676 = NOT(g12941)
--	g13869 = NOT(g10831)
--	g20558 = NOT(I20650)
--	g8680 = NOT(g686)
--	g22936 = NOT(g20283)
--	I13623 = NOT(g4294)
--	I21486 = NOT(g18727)
--	g17953 = NOT(I18861)
--	I22327 = NOT(g19367)
--	g23339 = NOT(g21070)
--	g8353 = NOT(I12530)
--	g18938 = NOT(g16053)
--	g23943 = NOT(g19147)
--	g18093 = NOT(I18885)
--	I13037 = NOT(g4304)
--	I29149 = NOT(g29384)
--	g14431 = NOT(g12208)
--	g31213 = NOT(I29013)
--	g11868 = NOT(g9185)
--	g12864 = NOT(g10373)
--	g13868 = NOT(g11493)
--	g6917 = NOT(g3684)
--	g8744 = NOT(g691)
--	g23338 = NOT(g20453)
--	g18065 = NOT(I18875)
--	g24893 = NOT(I24060)
--	g12749 = NOT(g7074)
--	g19435 = NOT(g16449)
--	g9162 = NOT(g622)
--	g9019 = NOT(I12950)
--	g17417 = NOT(g14804)
--	I18609 = NOT(g5976)
--	g7886 = NOT(g1442)
--	g20544 = NOT(g15171)
--	g23969 = NOT(g19277)
--	g32626 = NOT(g30614)
--	g28039 = NOT(g26365)
--	I32195 = NOT(g33628)
--	I13352 = NOT(g4146)
--	g11709 = NOT(I14584)
--	g30997 = NOT(g29702)
--	g10156 = NOT(g2675)
--	g20713 = NOT(g15277)
--	g21060 = NOT(g15509)
--	g34997 = NOT(I33291)
--	I12991 = NOT(g6752)
--	g23060 = NOT(g19908)
--	g23968 = NOT(g18833)
--	g18875 = NOT(g15171)
--	g32533 = NOT(g30614)
--	g8558 = NOT(g3787)
--	g28038 = NOT(g26365)
--	I32525 = NOT(g34285)
--	g13259 = NOT(I15824)
--	g33912 = NOT(I31770)
--	g19744 = NOT(g15885)
--	g16620 = NOT(I17808)
--	g7314 = NOT(g1740)
--	g10180 = NOT(g2259)
--	I14006 = NOT(g9104)
--	I17108 = NOT(g13782)
--	I14475 = NOT(g10175)
--	g11471 = NOT(g7626)
--	g19345 = NOT(g17591)
--	g25099 = NOT(g22369)
--	g13087 = NOT(g12012)
--	g32775 = NOT(g30825)
--	g25388 = NOT(g22763)
--	g25324 = NOT(g22228)
--	I14727 = NOT(g7753)
--	g13258 = NOT(I15821)
--	g12900 = NOT(g10406)
--	g19399 = NOT(g16489)
--	g20610 = NOT(g18008)
--	g7870 = NOT(g1193)
--	g21411 = NOT(g15426)
--	g17762 = NOT(g13000)
--	g20705 = NOT(I20793)
--	g34766 = NOT(g34703)
--	g23870 = NOT(g21293)
--	I16010 = NOT(g11148)
--	g23411 = NOT(g20734)
--	g23527 = NOT(g21611)
--	g28187 = NOT(I26710)
--	I14222 = NOT(g8286)
--	I21922 = NOT(g21335)
--	g25534 = NOT(g22763)
--	g15932 = NOT(I17395)
--	g25098 = NOT(g22369)
--	g10335 = NOT(g4483)
--	I23321 = NOT(g21693)
--	g7650 = NOT(g4064)
--	g27101 = NOT(g26770)
--	g25272 = NOT(g23715)
--	g29862 = NOT(g28406)
--	g24042 = NOT(g20014)
--	g33072 = NOT(g31945)
--	g20189 = NOT(I20447)
--	g19398 = NOT(g16489)
--	g20679 = NOT(g15634)
--	I29368 = NOT(g30321)
--	g17423 = NOT(I18360)
--	g16971 = NOT(I18131)
--	g11043 = NOT(g8561)
--	g12036 = NOT(g9245)
--	g9086 = NOT(g847)
--	g32737 = NOT(g31327)
--	I18813 = NOT(g5673)
--	g17216 = NOT(g14454)
--	g20270 = NOT(g15277)
--	g9728 = NOT(g5109)
--	g19652 = NOT(g16897)
--	I30986 = NOT(g32437)
--	I17750 = NOT(g14383)
--	g22543 = NOT(g19801)
--	g17587 = NOT(I18518)
--	g9730 = NOT(g5436)
--	I31504 = NOT(g33164)
--	g24124 = NOT(g21209)
--	g8092 = NOT(g1589)
--	g14694 = NOT(I16795)
--	g29948 = NOT(g28853)
--	g8492 = NOT(g3396)
--	g9185 = NOT(I13007)
--	g23503 = NOT(g21468)
--	g23894 = NOT(g19074)
--	g19263 = NOT(I19799)
--	g32697 = NOT(g31070)
--	g27064 = NOT(I25786)
--	I18674 = NOT(g13101)
--	g25032 = NOT(g23639)
--	g20383 = NOT(g15373)
--	g32856 = NOT(g31021)
--	I28913 = NOT(g30322)
--	g11810 = NOT(g9664)
--	g25140 = NOT(g22228)
--	g9070 = NOT(g5428)
--	g8714 = NOT(g4859)
--	g7594 = NOT(I12064)
--	g31820 = NOT(g29385)
--	g10487 = NOT(g10233)
--	g32880 = NOT(g30614)
--	g13068 = NOT(I15697)
--	g25997 = NOT(I25095)
--	g7972 = NOT(g1046)
--	g24030 = NOT(g21127)
--	g20267 = NOT(g17955)
--	g24093 = NOT(g20998)
--	g10502 = NOT(g8876)
--	g26776 = NOT(g25498)
--	g23714 = NOT(g20751)
--	I27758 = NOT(g28119)
--	g23450 = NOT(I22571)
--	I29228 = NOT(g30314)
--	g32512 = NOT(g31566)
--	g7806 = NOT(g4681)
--	I15878 = NOT(g11249)
--	g20065 = NOT(g16846)
--	g31846 = NOT(g29385)
--	g7943 = NOT(g1395)
--	g24065 = NOT(g20982)
--	g11878 = NOT(I14690)
--	g19361 = NOT(I19843)
--	I20609 = NOT(g16539)
--	I12758 = NOT(g4093)
--	g23819 = NOT(g19147)
--	g12874 = NOT(g10383)
--	g26754 = NOT(g25300)
--	g34472 = NOT(I32525)
--	g25766 = NOT(g24439)
--	g28479 = NOT(g27654)
--	I32678 = NOT(g34428)
--	g23202 = NOT(I22302)
--	g14443 = NOT(I16596)
--	g23257 = NOT(g20924)
--	g26859 = NOT(I25591)
--	g27009 = NOT(g25911)
--	g26825 = NOT(I25541)
--	g21055 = NOT(g15224)
--	g23496 = NOT(g20248)
--	g7322 = NOT(g1862)
--	g16228 = NOT(I17569)
--	g20219 = NOT(I20495)
--	g23055 = NOT(g20887)
--	g6990 = NOT(g4742)
--	g17242 = NOT(g14454)
--	g34246 = NOT(I32237)
--	g10278 = NOT(g4628)
--	g33413 = NOT(g31971)
--	g29847 = NOT(g28395)
--	I29582 = NOT(g30591)
--	g23111 = NOT(g20391)
--	g12009 = NOT(I14862)
--	g21070 = NOT(I20937)
--	g6888 = NOT(I11701)
--	g22974 = NOT(g20330)
--	g32831 = NOT(g31376)
--	g33691 = NOT(I31528)
--	g32445 = NOT(I29973)
--	I32938 = NOT(g34663)
--	I32093 = NOT(g33670)
--	I13276 = NOT(g5798)
--	g16716 = NOT(g13948)
--	g9678 = NOT(g5406)
--	g10039 = NOT(g2273)
--	g10306 = NOT(I13726)
--	g32499 = NOT(g31376)
--	g23986 = NOT(g18833)
--	g30591 = NOT(I28851)
--	g6956 = NOT(g4242)
--	g18984 = NOT(g17486)
--	g8623 = NOT(g3990)
--	I11809 = NOT(g6741)
--	g34591 = NOT(I32681)
--	I18214 = NOT(g12918)
--	g12892 = NOT(g10398)
--	g34785 = NOT(I32985)
--	g16582 = NOT(g13915)
--	g17772 = NOT(g14297)
--	g34776 = NOT(I32970)
--	g11425 = NOT(g7640)
--	g10038 = NOT(g2241)
--	g32498 = NOT(g31566)
--	g23384 = NOT(I22485)
--	g17639 = NOT(I18600)
--	I12141 = NOT(g599)
--	g34147 = NOT(g33823)
--	g9682 = NOT(I13280)
--	g9766 = NOT(g2748)
--	g15811 = NOT(g13125)
--	g16310 = NOT(g13223)
--	g7096 = NOT(g6537)
--	g10815 = NOT(g9917)
--	g13458 = NOT(g11048)
--	g24160 = NOT(I23324)
--	I15918 = NOT(g12381)
--	g9305 = NOT(g5381)
--	g7496 = NOT(g5969)
--	g33929 = NOT(I31803)
--	g16627 = NOT(I17819)
--	g17638 = NOT(g14838)
--	g22841 = NOT(g20391)
--	g34950 = NOT(g34940)
--	g12914 = NOT(g12235)
--	g13010 = NOT(I15620)
--	g32611 = NOT(g31154)
--	g7845 = NOT(g1146)
--	I33232 = NOT(g34957)
--	g25451 = NOT(g22228)
--	g32722 = NOT(g30937)
--	g25220 = NOT(I24396)
--	g32924 = NOT(g30937)
--	g33928 = NOT(I31800)
--	g19947 = NOT(g17226)
--	g7195 = NOT(g25)
--	g12907 = NOT(g10415)
--	g20617 = NOT(g15277)
--	g17416 = NOT(g14956)
--	g7395 = NOT(g6005)
--	g7891 = NOT(g2994)
--	g8651 = NOT(g758)
--	g16958 = NOT(g14238)
--	g9748 = NOT(g114)
--	g13545 = NOT(I16010)
--	g23877 = NOT(g19147)
--	g19273 = NOT(g16100)
--	g20915 = NOT(I20882)
--	g7913 = NOT(g1052)
--	g27074 = NOT(I25790)
--	g28321 = NOT(g27317)
--	I32837 = NOT(g34498)
--	g30996 = NOT(g29694)
--	g25246 = NOT(g23828)
--	g34151 = NOT(I32106)
--	I12135 = NOT(g807)
--	g10143 = NOT(g568)
--	g29213 = NOT(I27555)
--	g34996 = NOT(I33288)
--	g23019 = NOT(g19866)
--	I33261 = NOT(g34977)
--	g8285 = NOT(I12497)
--	g12074 = NOT(I14932)
--	I25695 = NOT(g25690)
--	g9226 = NOT(g1564)
--	g20277 = NOT(g16487)
--	g16603 = NOT(I17787)
--	g16742 = NOT(g13983)
--	g23196 = NOT(g20785)
--	g34844 = NOT(g34737)
--	I22564 = NOT(g20857)
--	g16096 = NOT(g13530)
--	g23018 = NOT(g19801)
--	g32753 = NOT(g30735)
--	g12238 = NOT(I15102)
--	g32461 = NOT(g30614)
--	I21242 = NOT(g16540)
--	g10169 = NOT(g6395)
--	g24075 = NOT(g19935)
--	g17579 = NOT(g14959)
--	g19371 = NOT(I19857)
--	g20595 = NOT(g15877)
--	g23526 = NOT(g21611)
--	g6808 = NOT(g554)
--	g20494 = NOT(g17847)
--	g14169 = NOT(g12381)
--	g8139 = NOT(g1648)
--	I16289 = NOT(g12107)
--	I32455 = NOT(g34242)
--	g7266 = NOT(g35)
--	g29912 = NOT(g28827)
--	g29311 = NOT(g28998)
--	g10410 = NOT(g7069)
--	g20623 = NOT(g17929)
--	g27675 = NOT(I26309)
--	I12049 = NOT(g781)
--	g9373 = NOT(g5142)
--	g17014 = NOT(g14297)
--	g27092 = NOT(g26737)
--	g9091 = NOT(g1430)
--	g20037 = NOT(g17328)
--	g31827 = NOT(g29385)
--	g32736 = NOT(g30937)
--	I32617 = NOT(g34333)
--	g13322 = NOT(g10918)
--	g32887 = NOT(g30614)
--	I32470 = NOT(g34247)
--	g24623 = NOT(g23076)
--	g33827 = NOT(I31672)
--	g9491 = NOT(g2729)
--	I14905 = NOT(g9822)
--	g24037 = NOT(g21127)
--	g34420 = NOT(g34152)
--	g16429 = NOT(I17671)
--	I11665 = NOT(g1589)
--	g20782 = NOT(g15853)
--	g21457 = NOT(g17367)
--	g13901 = NOT(g11480)
--	g23402 = NOT(g20875)
--	I13166 = NOT(g5101)
--	g32529 = NOT(g30735)
--	g23457 = NOT(I22580)
--	g25370 = NOT(g22228)
--	g8795 = NOT(I12793)
--	g10363 = NOT(I13779)
--	I24400 = NOT(g23954)
--	g10217 = NOT(g2102)
--	I14593 = NOT(g9978)
--	g30318 = NOT(g28274)
--	g14363 = NOT(I16521)
--	g14217 = NOT(I16417)
--	g9283 = NOT(g1736)
--	I14346 = NOT(g10233)
--	g16428 = NOT(I17668)
--	g9369 = NOT(g5084)
--	g32528 = NOT(g31554)
--	g32696 = NOT(g30825)
--	g9007 = NOT(g1083)
--	I21230 = NOT(g16540)
--	g32843 = NOT(g31021)
--	g6957 = NOT(g2932)
--	g24419 = NOT(g22722)
--	g32393 = NOT(g30922)
--	g9407 = NOT(g6549)
--	I15295 = NOT(g8515)
--	I11892 = NOT(g4408)
--	g34059 = NOT(g33658)
--	g8672 = NOT(g4669)
--	g9920 = NOT(g4322)
--	I15144 = NOT(g5659)
--	I13892 = NOT(g1576)
--	g31803 = NOT(g29385)
--	g32764 = NOT(g30937)
--	g24155 = NOT(I23309)
--	g24418 = NOT(g22722)
--	I32467 = NOT(g34246)
--	g20266 = NOT(g17873)
--	g8477 = NOT(g3061)
--	g34540 = NOT(I32607)
--	g11823 = NOT(I14647)
--	g13680 = NOT(I16077)
--	g17615 = NOT(I18574)
--	g12883 = NOT(g10390)
--	g13144 = NOT(I15773)
--	g22493 = NOT(g19801)
--	g7097 = NOT(I11809)
--	g23001 = NOT(g19801)
--	g34058 = NOT(g33660)
--	g24170 = NOT(I23354)
--	g32869 = NOT(g30735)
--	I18882 = NOT(g16580)
--	g32960 = NOT(g31327)
--	I18414 = NOT(g14359)
--	g7497 = NOT(g6358)
--	I14797 = NOT(g9636)
--	g19421 = NOT(g16326)
--	g17720 = NOT(g15045)
--	I33056 = NOT(g34778)
--	I25689 = NOT(g25688)
--	g9582 = NOT(g703)
--	g11336 = NOT(g7620)
--	g7960 = NOT(g1404)
--	g32868 = NOT(g31376)
--	g8205 = NOT(g2208)
--	I32782 = NOT(g34571)
--	g10223 = NOT(g4561)
--	g21689 = NOT(I21250)
--	g23256 = NOT(g20785)
--	I12106 = NOT(g626)
--	I12605 = NOT(g1570)
--	g17430 = NOT(I18373)
--	g17746 = NOT(g14825)
--	g20853 = NOT(g15595)
--	g34044 = NOT(g33675)
--	g21280 = NOT(g16601)
--	g23923 = NOT(g18997)
--	I14409 = NOT(g8364)
--	g29152 = NOT(g27907)
--	g29846 = NOT(g28391)
--	I32352 = NOT(g34169)
--	I29002 = NOT(g29675)
--	g21300 = NOT(I21047)
--	g20167 = NOT(g16971)
--	g20194 = NOT(g16897)
--	g20589 = NOT(g15224)
--	g32709 = NOT(g30735)
--	g11966 = NOT(I14800)
--	g23300 = NOT(g20283)
--	I12463 = NOT(g4812)
--	g17465 = NOT(g12955)
--	g8742 = NOT(g4035)
--	g13966 = NOT(I16246)
--	g10084 = NOT(g2837)
--	g24167 = NOT(I23345)
--	g9415 = NOT(g2169)
--	g19541 = NOT(g16136)
--	g30301 = NOT(I28548)
--	g10110 = NOT(g661)
--	g11631 = NOT(g8595)
--	g19473 = NOT(g16349)
--	g18101 = NOT(I18909)
--	g11017 = NOT(g10289)
--	g20588 = NOT(g18008)
--	g20524 = NOT(g17873)
--	g32708 = NOT(g31376)
--	I32170 = NOT(g33638)
--	I12033 = NOT(g776)
--	g13017 = NOT(I15633)
--	I28174 = NOT(g28803)
--	I29245 = NOT(g29491)
--	g32471 = NOT(g31376)
--	g19789 = NOT(g17015)
--	g24524 = NOT(g22876)
--	g24836 = NOT(I24008)
--	g16129 = NOT(I17488)
--	g25227 = NOT(g22763)
--	g14321 = NOT(g10874)
--	g34739 = NOT(I32909)
--	g10531 = NOT(g8925)
--	g17684 = NOT(g15036)
--	g27438 = NOT(I26130)
--	g14179 = NOT(g11048)
--	g25025 = NOT(g22498)
--	g7267 = NOT(g1604)
--	g24477 = NOT(I23680)
--	g10178 = NOT(g2126)
--	g26632 = NOT(g25473)
--	g24119 = NOT(g19935)
--	g27349 = NOT(g26352)
--	I31650 = NOT(g33212)
--	g23066 = NOT(g20330)
--	I28390 = NOT(g29185)
--	g9721 = NOT(g5097)
--	g23231 = NOT(g20050)
--	g34699 = NOT(I32855)
--	g19434 = NOT(g16326)
--	g16626 = NOT(g14133)
--	g8273 = NOT(g2453)
--	g10685 = NOT(I13995)
--	I16489 = NOT(g12793)
--	g16323 = NOT(I17653)
--	g24118 = NOT(g19890)
--	g10373 = NOT(g6917)
--	g14186 = NOT(g11346)
--	g14676 = NOT(I16775)
--	g24022 = NOT(g20982)
--	g34698 = NOT(g34550)
--	g7293 = NOT(g4452)
--	g12906 = NOT(g10413)
--	g16533 = NOT(I17733)
--	g20616 = NOT(g15277)
--	I18114 = NOT(g14509)
--	g23876 = NOT(g19074)
--	I18758 = NOT(g6719)
--	g13023 = NOT(g11897)
--	g18874 = NOT(g15938)
--	I31528 = NOT(g33219)
--	g25044 = NOT(g23675)
--	I19661 = NOT(g17587)
--	g29929 = NOT(g28914)
--	g16775 = NOT(I17999)
--	I18107 = NOT(g4019)
--	g10417 = NOT(g7117)
--	I25511 = NOT(g25073)
--	g32602 = NOT(g30825)
--	g32810 = NOT(g31376)
--	I13637 = NOT(g102)
--	I20882 = NOT(g17619)
--	g32657 = NOT(g31528)
--	g32774 = NOT(g30735)
--	g33778 = NOT(I31625)
--	g7828 = NOT(g4871)
--	g32955 = NOT(g30735)
--	g21511 = NOT(g15483)
--	g29928 = NOT(g28871)
--	I26670 = NOT(g27709)
--	g20704 = NOT(g15373)
--	g23511 = NOT(I22640)
--	g34427 = NOT(I32452)
--	I32119 = NOT(g33648)
--	g32879 = NOT(g31327)
--	g8572 = NOT(I12654)
--	g20053 = NOT(g17328)
--	g32970 = NOT(g30825)
--	g10334 = NOT(g4420)
--	g19682 = NOT(g17015)
--	I14537 = NOT(g10106)
--	g24053 = NOT(g21256)
--	g25120 = NOT(g22432)
--	I17780 = NOT(g13303)
--	g17523 = NOT(g14732)
--	g20900 = NOT(I20864)
--	g8712 = NOT(I12712)
--	g7592 = NOT(g347)
--	I16544 = NOT(g11931)
--	I18849 = NOT(g14290)
--	g18008 = NOT(I18868)
--	g32878 = NOT(g30937)
--	g31945 = NOT(g31189)
--	g21660 = NOT(g17694)
--	g24466 = NOT(I23671)
--	I16713 = NOT(g5331)
--	g9689 = NOT(g124)
--	g10762 = NOT(g8470)
--	g25562 = NOT(g22763)
--	g18892 = NOT(g15680)
--	g20036 = NOT(g17433)
--	g31826 = NOT(g29385)
--	g32886 = NOT(g31327)
--	I33161 = NOT(g34894)
--	I18398 = NOT(g13745)
--	g20101 = NOT(g17533)
--	g24036 = NOT(g20982)
--	I12541 = NOT(g194)
--	g20560 = NOT(g17328)
--	g16856 = NOT(I18048)
--	g21456 = NOT(g15509)
--	I26667 = NOT(g27585)
--	g11985 = NOT(I14827)
--	g17475 = NOT(I18398)
--	g24101 = NOT(g20998)
--	I23684 = NOT(g23230)
--	g32792 = NOT(g31710)
--	g23456 = NOT(g21514)
--	g13976 = NOT(g11130)
--	g24177 = NOT(I23375)
--	g24560 = NOT(g22942)
--	I15954 = NOT(g12381)
--	g32967 = NOT(g31327)
--	g10216 = NOT(I13684)
--	g14423 = NOT(I16579)
--	g8534 = NOT(g3338)
--	I16610 = NOT(g10981)
--	g9671 = NOT(g5134)
--	g20642 = NOT(g15277)
--	g23480 = NOT(I22601)
--	g27415 = NOT(g26382)
--	I20584 = NOT(g16587)
--	g23916 = NOT(g19277)
--	g9030 = NOT(g4793)
--	g19760 = NOT(g17015)
--	I32305 = NOT(g34209)
--	I14381 = NOT(g8300)
--	g16512 = NOT(g14015)
--	I16679 = NOT(g12039)
--	g23550 = NOT(g20248)
--	g26784 = NOT(g25341)
--	g9247 = NOT(g1559)
--	I33258 = NOT(g34976)
--	I32809 = NOT(g34586)
--	g18907 = NOT(g15979)
--	g7624 = NOT(I12106)
--	g32459 = NOT(g31070)
--	g20064 = NOT(g17533)
--	g7953 = NOT(g4966)
--	g30572 = NOT(g29945)
--	g24064 = NOT(g20841)
--	g28579 = NOT(g27714)
--	g9564 = NOT(g6120)
--	I18135 = NOT(g13144)
--	g23307 = NOT(g20924)
--	g32919 = NOT(g30735)
--	g23085 = NOT(g19957)
--	g32458 = NOT(g30825)
--	I24759 = NOT(g24229)
--	g14543 = NOT(I16660)
--	g33932 = NOT(I31810)
--	g9826 = NOT(g1844)
--	g10117 = NOT(g2509)
--	g10000 = NOT(g6151)
--	g26824 = NOT(g25298)
--	I16460 = NOT(g10430)
--	g20874 = NOT(g15680)
--	g21054 = NOT(g15373)
--	g32918 = NOT(g31327)
--	g23243 = NOT(g21070)
--	g20630 = NOT(g17955)
--	g11842 = NOT(I14660)
--	g21431 = NOT(g18065)
--	g9741 = NOT(I13317)
--	g8903 = NOT(g1075)
--	g23431 = NOT(g21514)
--	I13906 = NOT(g7620)
--	g32545 = NOT(g31070)
--	g9910 = NOT(g2108)
--	g17600 = NOT(g14659)
--	I19671 = NOT(g15932)
--	g34490 = NOT(I32547)
--	g20166 = NOT(g16886)
--	g20009 = NOT(g16349)
--	I22583 = NOT(g20998)
--	g27576 = NOT(g26081)
--	g27585 = NOT(g25994)
--	g20665 = NOT(g15373)
--	g25547 = NOT(g22550)
--	g32599 = NOT(g30673)
--	I20744 = NOT(g17141)
--	I31810 = NOT(g33164)
--	g9638 = NOT(g1620)
--	g21269 = NOT(g15506)
--	g24166 = NOT(I23342)
--	g24665 = NOT(g23067)
--	g7716 = NOT(g1199)
--	g7149 = NOT(g4564)
--	g34784 = NOT(I32982)
--	g7349 = NOT(g1270)
--	g30297 = NOT(g28758)
--	g27554 = NOT(g26625)
--	g20008 = NOT(g16449)
--	g34956 = NOT(I33214)
--	g17952 = NOT(I18858)
--	g32598 = NOT(g30614)
--	g13016 = NOT(g11878)
--	I22046 = NOT(g19330)
--	g23942 = NOT(g21562)
--	I20399 = NOT(g16205)
--	g23341 = NOT(g21163)
--	g18092 = NOT(I18882)
--	g21268 = NOT(g15680)
--	I14192 = NOT(g10233)
--	I18048 = NOT(g13638)
--	I28062 = NOT(g29194)
--	g25226 = NOT(g22763)
--	g22137 = NOT(g21370)
--	g21156 = NOT(g17247)
--	g17821 = NOT(I18829)
--	g8178 = NOT(I12437)
--	g6801 = NOT(g391)
--	I21006 = NOT(g15579)
--	g28615 = NOT(g27817)
--	I16875 = NOT(g6675)
--	g25481 = NOT(g22228)
--	I15893 = NOT(g10430)
--	I31878 = NOT(g33696)
--	g19649 = NOT(g17015)
--	I32874 = NOT(g34504)
--	g21180 = NOT(g18008)
--	I14663 = NOT(g9747)
--	g21670 = NOT(g16540)
--	I18221 = NOT(g13605)
--	g16722 = NOT(I17938)
--	g16924 = NOT(I18092)
--	g20555 = NOT(g15480)
--	g32817 = NOT(g31376)
--	I28851 = NOT(g29317)
--	I28872 = NOT(g30072)
--	I32693 = NOT(g34433)
--	g8135 = NOT(I12418)
--	I21222 = NOT(g18091)
--	g19491 = NOT(g16349)
--	g34181 = NOT(g33913)
--	g34671 = NOT(I32797)
--	g20570 = NOT(g15277)
--	g20712 = NOT(g15509)
--	g11865 = NOT(g10124)
--	I22302 = NOT(g19353)
--	g13865 = NOT(I16168)
--	g20914 = NOT(g15373)
--	g21335 = NOT(I21067)
--	g18883 = NOT(g15938)
--	g32532 = NOT(g31170)
--	g32901 = NOT(g31327)
--	g14639 = NOT(I16747)
--	g10230 = NOT(I13694)
--	g23335 = NOT(g20391)
--	I32665 = NOT(g34386)
--	g19755 = NOT(g15915)
--	g6755 = NOT(I11620)
--	g12921 = NOT(g12228)
--	g23839 = NOT(g18997)
--	I17787 = NOT(g3267)
--	g17873 = NOT(I18849)
--	g23930 = NOT(g19147)
--	g23993 = NOT(g19277)
--	g32783 = NOT(g30825)
--	g19770 = NOT(g17062)
--	I29199 = NOT(g30237)
--	g30931 = NOT(I28913)
--	g8805 = NOT(I12799)
--	I14862 = NOT(g8092)
--	g8916 = NOT(I12887)
--	I16160 = NOT(g11237)
--	g21694 = NOT(g16540)
--	g23838 = NOT(g18997)
--	g9861 = NOT(g5459)
--	g10416 = NOT(g10318)
--	I15705 = NOT(g12218)
--	g9048 = NOT(I12963)
--	I17302 = NOT(g14044)
--	g32561 = NOT(g30614)
--	g32656 = NOT(g30673)
--	g23965 = NOT(g21611)
--	I31459 = NOT(g33219)
--	g20239 = NOT(g17128)
--	I32476 = NOT(g34277)
--	g11705 = NOT(I14576)
--	I22640 = NOT(g21256)
--	g24074 = NOT(g21193)
--	I22769 = NOT(g21277)
--	g26860 = NOT(I25594)
--	I14326 = NOT(g8607)
--	g34426 = NOT(I32449)
--	g11042 = NOT(g8691)
--	g16031 = NOT(I17436)
--	g20567 = NOT(g15426)
--	g20594 = NOT(g15277)
--	g32680 = NOT(g31376)
--	g10391 = NOT(g6988)
--	I16455 = NOT(g11845)
--	g32823 = NOT(g31327)
--	g20238 = NOT(g17096)
--	g25297 = NOT(g23746)
--	g13255 = NOT(g10632)
--	g9827 = NOT(g1974)
--	g13189 = NOT(g10762)
--	g22542 = NOT(g19801)
--	g13679 = NOT(g10573)
--	g28142 = NOT(I26649)
--	g31811 = NOT(g29385)
--	g23487 = NOT(g20924)
--	g14510 = NOT(I16629)
--	g31646 = NOT(I29228)
--	g9333 = NOT(g417)
--	I14702 = NOT(g7717)
--	g19794 = NOT(g16489)
--	g11678 = NOT(I14563)
--	g12184 = NOT(I15036)
--	g16529 = NOT(g14055)
--	g29081 = NOT(g27837)
--	g12805 = NOT(g9511)
--	g13188 = NOT(g10909)
--	g19395 = NOT(g16431)
--	g23502 = NOT(g21070)
--	I27927 = NOT(g28803)
--	g20382 = NOT(g15171)
--	I16201 = NOT(g4023)
--	I23351 = NOT(g23263)
--	I31545 = NOT(g33219)
--	I23372 = NOT(g23361)
--	g26700 = NOT(g25429)
--	g7258 = NOT(g4414)
--	I33079 = NOT(g34809)
--	g11686 = NOT(I14567)
--	g16528 = NOT(g14154)
--	g7577 = NOT(g1263)
--	g7867 = NOT(g1489)
--	g13460 = NOT(I15942)
--	g15831 = NOT(g13385)
--	I26479 = NOT(g25771)
--	I12927 = NOT(g4332)
--	g26987 = NOT(g26131)
--	g11383 = NOT(g9061)
--	g10014 = NOT(g6439)
--	g23443 = NOT(g21468)
--	I15030 = NOT(g10073)
--	I18795 = NOT(g5327)
--	g21279 = NOT(g15680)
--	g24176 = NOT(I23372)
--	g24185 = NOT(I23399)
--	g23279 = NOT(g21037)
--	g32966 = NOT(g31021)
--	g19633 = NOT(g16931)
--	g7717 = NOT(I12172)
--	g30088 = NOT(g29094)
--	g24092 = NOT(g20857)
--	I32074 = NOT(g33670)
--	g29945 = NOT(I28174)
--	g6868 = NOT(I11688)
--	g11030 = NOT(g8292)
--	g20154 = NOT(I20412)
--	g22905 = NOT(I22114)
--	g32631 = NOT(g30825)
--	g19719 = NOT(g16897)
--	g21278 = NOT(I21013)
--	g11294 = NOT(g7598)
--	g24154 = NOT(I23306)
--	I32594 = NOT(g34298)
--	g8037 = NOT(g405)
--	g23278 = NOT(g20283)
--	g13267 = NOT(I15831)
--	g29999 = NOT(g28973)
--	g32364 = NOT(I29894)
--	g6767 = NOT(I11626)
--	g17614 = NOT(I18571)
--	g22593 = NOT(g19801)
--	g9780 = NOT(I13360)
--	g16960 = NOT(I18114)
--	g20637 = NOT(g15224)
--	g26943 = NOT(I25695)
--	g8102 = NOT(g3072)
--	g13065 = NOT(g10476)
--	g19718 = NOT(g17015)
--	g21286 = NOT(g15509)
--	g8302 = NOT(g1926)
--	g14442 = NOT(I16593)
--	g29998 = NOT(g28966)
--	g17607 = NOT(I18560)
--	g21468 = NOT(I21181)
--	g17320 = NOT(I18297)
--	g21306 = NOT(g15582)
--	g31850 = NOT(g29385)
--	g8579 = NOT(g2771)
--	g23306 = NOT(g20924)
--	I29225 = NOT(g30311)
--	I31817 = NOT(g33323)
--	g7975 = NOT(g3040)
--	g33850 = NOT(I31701)
--	g17530 = NOT(g14947)
--	g10116 = NOT(g2413)
--	g9662 = NOT(g3983)
--	g9018 = NOT(g4273)
--	g11875 = NOT(I14687)
--	g8719 = NOT(I12719)
--	g27013 = NOT(I25743)
--	g7026 = NOT(g5507)
--	I32675 = NOT(g34427)
--	g9467 = NOT(g6434)
--	g19440 = NOT(g15915)
--	g16709 = NOT(I17919)
--	g17122 = NOT(g14348)
--	g34126 = NOT(I32067)
--	g34659 = NOT(I32775)
--	I12770 = NOT(g4200)
--	I12563 = NOT(g3798)
--	g12013 = NOT(I14866)
--	g23815 = NOT(g19074)
--	g34987 = NOT(I33261)
--	I25677 = NOT(g25640)
--	I15837 = NOT(g1459)
--	I33158 = NOT(g34897)
--	g7170 = NOT(g5719)
--	g19861 = NOT(g17096)
--	g10275 = NOT(g4584)
--	g19573 = NOT(g16877)
--	g8917 = NOT(I12890)
--	g16708 = NOT(I17916)
--	g22153 = NOT(g18997)
--	g21677 = NOT(I21238)
--	g33228 = NOT(I30766)
--	g10430 = NOT(I13847)
--	g14275 = NOT(g12358)
--	g25546 = NOT(g22550)
--	g32571 = NOT(g31376)
--	I31561 = NOT(g33197)
--	I17249 = NOT(g13605)
--	g25211 = NOT(g22763)
--	I32935 = NOT(g34657)
--	g22409 = NOT(I21860)
--	g19389 = NOT(g17532)
--	g17641 = NOT(g14845)
--	g20501 = NOT(g17955)
--	g26870 = NOT(I25606)
--	g30296 = NOT(g28889)
--	g20577 = NOT(g15483)
--	g34339 = NOT(g34077)
--	g9816 = NOT(g6167)
--	g34943 = NOT(I33197)
--	I20951 = NOT(g17782)
--	g25024 = NOT(g22472)
--	g33716 = NOT(I31569)
--	I31823 = NOT(g33149)
--	g19612 = NOT(g16897)
--	g34296 = NOT(I32297)
--	g7280 = NOT(g2153)
--	g29897 = NOT(I28128)
--	g7939 = NOT(g1280)
--	g22136 = NOT(g20277)
--	g29961 = NOT(g28892)
--	g8442 = NOT(g3476)
--	g22408 = NOT(g19483)
--	g22635 = NOT(g19801)
--	I12767 = NOT(g4197)
--	g14237 = NOT(g11666)
--	g8786 = NOT(I12770)
--	g23937 = NOT(g19277)
--	g10035 = NOT(g1720)
--	g32495 = NOT(g31070)
--	g29505 = NOT(g29186)
--	g19777 = NOT(g17015)
--	g17409 = NOT(I18344)
--	I12899 = NOT(g4232)
--	g7544 = NOT(g918)
--	g8164 = NOT(g3484)
--	g9381 = NOT(g5527)
--	I15617 = NOT(g12037)
--	I13805 = NOT(g6976)
--	I18788 = NOT(g13138)
--	g8364 = NOT(g1585)
--	g32816 = NOT(g31327)
--	I15915 = NOT(g10430)
--	g24438 = NOT(g22722)
--	g11470 = NOT(g7625)
--	g17136 = NOT(g14348)
--	g10142 = NOT(I13637)
--	g17408 = NOT(I18341)
--	g34060 = NOT(g33704)
--	g29212 = NOT(I27552)
--	g7636 = NOT(g4098)
--	g9685 = NOT(g6533)
--	I26676 = NOT(g27736)
--	g9197 = NOT(g1221)
--	I18829 = NOT(g13350)
--	g32687 = NOT(g31376)
--	g9397 = NOT(g6088)
--	I18434 = NOT(g13782)
--	g33959 = NOT(I31878)
--	g9021 = NOT(I12954)
--	I12719 = NOT(g365)
--	g16602 = NOT(g14101)
--	g21410 = NOT(g15224)
--	g34197 = NOT(g33812)
--	I27718 = NOT(g28231)
--	I16401 = NOT(g869)
--	g16774 = NOT(g14024)
--	g23410 = NOT(g21562)
--	g8770 = NOT(g749)
--	I29337 = NOT(g30286)
--	g34855 = NOT(I33079)
--	I26654 = NOT(g27576)
--	I22380 = NOT(g21156)
--	g16955 = NOT(I18107)
--	g32752 = NOT(g31376)
--	g8296 = NOT(g246)
--	g25250 = NOT(I24434)
--	g27100 = NOT(g26759)
--	g32954 = NOT(g31376)
--	g8725 = NOT(g739)
--	g24083 = NOT(g19984)
--	g33378 = NOT(I30904)
--	g21666 = NOT(g16540)
--	g23479 = NOT(g21562)
--	I26936 = NOT(g27599)
--	g32643 = NOT(g31376)
--	g6940 = NOT(g4035)
--	I15494 = NOT(g10385)
--	g13075 = NOT(I15705)
--	g23363 = NOT(I22470)
--	I18344 = NOT(g13003)
--	g7187 = NOT(g6065)
--	g7387 = NOT(g2421)
--	g20622 = NOT(g15595)
--	g11467 = NOT(g7623)
--	g13595 = NOT(g10951)
--	I17999 = NOT(g4012)
--	g20566 = NOT(g15224)
--	g7461 = NOT(g2567)
--	I15623 = NOT(g12040)
--	g23478 = NOT(g21514)
--	g13494 = NOT(g11912)
--	g23015 = NOT(g20391)
--	g8553 = NOT(g3747)
--	I26334 = NOT(g26834)
--	I19707 = NOT(g17590)
--	g25296 = NOT(g23745)
--	g10130 = NOT(g5694)
--	g16171 = NOT(g13530)
--	g33944 = NOT(I31829)
--	g19061 = NOT(I19762)
--	g26818 = NOT(I25530)
--	g16886 = NOT(I18078)
--	I27573 = NOT(g28157)
--	g32669 = NOT(g30614)
--	I15782 = NOT(g10430)
--	g23486 = NOT(g20785)
--	g26055 = NOT(I25115)
--	g13037 = NOT(g10981)
--	g10362 = NOT(g6850)
--	g29149 = NOT(g27837)
--	g7027 = NOT(g5499)
--	I19818 = NOT(g1056)
--	g19766 = NOT(g16449)
--	g21556 = NOT(g15669)
--	I12861 = NOT(g4372)
--	g10165 = NOT(g5698)
--	g13782 = NOT(I16117)
--	g17575 = NOT(g14921)
--	g28137 = NOT(I26638)
--	g11984 = NOT(g9186)
--	g16967 = NOT(I18125)
--	I22331 = NOT(g19417)
--	g32668 = NOT(g31070)
--	g32842 = NOT(g31710)
--	g17711 = NOT(I18694)
--	g7046 = NOT(g5791)
--	I32284 = NOT(g34052)
--	g20653 = NOT(I20747)
--	g27991 = NOT(g25852)
--	I33288 = NOT(g34989)
--	g31802 = NOT(g29385)
--	g9631 = NOT(g6573)
--	g17327 = NOT(I18310)
--	g25060 = NOT(g23708)
--	g32489 = NOT(g30614)
--	g8389 = NOT(g3125)
--	I13329 = NOT(g86)
--	I27388 = NOT(g27698)
--	g31857 = NOT(g29385)
--	g7446 = NOT(g1256)
--	g18200 = NOT(I19012)
--	g29811 = NOT(g28376)
--	g23223 = NOT(g21308)
--	g7514 = NOT(g6704)
--	g19360 = NOT(g16249)
--	g11418 = NOT(I14424)
--	g34714 = NOT(I32874)
--	g8990 = NOT(g146)
--	g12882 = NOT(g10389)
--	g9257 = NOT(g5115)
--	g22492 = NOT(g19614)
--	g25197 = NOT(g23958)
--	g29343 = NOT(g28174)
--	g7003 = NOT(g5152)
--	I13539 = NOT(g6381)
--	g22303 = NOT(g19277)
--	I27777 = NOT(g29043)
--	g9817 = NOT(I13374)
--	g32559 = NOT(g30825)
--	g34315 = NOT(g34085)
--	g10475 = NOT(g8844)
--	I17932 = NOT(g3310)
--	g24138 = NOT(g21143)
--	g32525 = NOT(g31170)
--	g32488 = NOT(g31194)
--	g11170 = NOT(g8476)
--	g34910 = NOT(g34864)
--	I29444 = NOT(g30928)
--	g8171 = NOT(g3817)
--	g10727 = NOT(I14016)
--	g7345 = NOT(g6415)
--	g7841 = NOT(g904)
--	I12534 = NOT(g50)
--	g20636 = NOT(g18008)
--	I19384 = NOT(g15085)
--	g8787 = NOT(I12773)
--	g32558 = NOT(g30735)
--	g34202 = NOT(I32161)
--	g23084 = NOT(g19954)
--	g24636 = NOT(g23121)
--	g6826 = NOT(g218)
--	g10222 = NOT(g4492)
--	g7191 = NOT(g6398)
--	g30055 = NOT(g29157)
--	g17606 = NOT(g14999)
--	g20852 = NOT(g15595)
--	g32830 = NOT(g31327)
--	g23922 = NOT(g18997)
--	g23321 = NOT(I22422)
--	g32893 = NOT(g30937)
--	I18028 = NOT(g13638)
--	g21179 = NOT(g15373)
--	I24920 = NOT(g25513)
--	g26801 = NOT(I25511)
--	I24434 = NOT(g22763)
--	g29368 = NOT(I27730)
--	g9751 = NOT(g1710)
--	g34070 = NOT(g33725)
--	g8281 = NOT(g3494)
--	g32544 = NOT(g30735)
--	g19629 = NOT(g17015)
--	g32865 = NOT(g31327)
--	g19451 = NOT(g15938)
--	g21178 = NOT(g17955)
--	g34590 = NOT(I32678)
--	g19472 = NOT(g16349)
--	g24963 = NOT(g22342)
--	g20664 = NOT(g15373)
--	g34986 = NOT(I33258)
--	g32713 = NOT(g30673)
--	g7536 = NOT(g5976)
--	g9585 = NOT(g1616)
--	g8297 = NOT(g142)
--	g10347 = NOT(I13759)
--	g21685 = NOT(I21246)
--	I16733 = NOT(g12026)
--	I12997 = NOT(g351)
--	g28726 = NOT(g27937)
--	g34384 = NOT(I32391)
--	g23953 = NOT(g19277)
--	g30067 = NOT(g29060)
--	g11401 = NOT(g7593)
--	g22840 = NOT(g20330)
--	g21654 = NOT(g17619)
--	I29977 = NOT(g31596)
--	g7858 = NOT(g947)
--	g32610 = NOT(g31070)
--	g20576 = NOT(g18065)
--	g20585 = NOT(g17955)
--	g23654 = NOT(g20248)
--	I12061 = NOT(g562)
--	g32705 = NOT(g30614)
--	g34094 = NOT(g33772)
--	g13477 = NOT(I15954)
--	g8745 = NOT(g744)
--	g28436 = NOT(I26929)
--	g8138 = NOT(g1500)
--	g8639 = NOT(g2807)
--	g24585 = NOT(g23063)
--	I22149 = NOT(g21036)
--	g19071 = NOT(g15591)
--	g23800 = NOT(g21246)
--	I23711 = NOT(g23192)
--	g20554 = NOT(g15348)
--	g23417 = NOT(g20391)
--	g32679 = NOT(g31579)
--	g16322 = NOT(I17650)
--	g8791 = NOT(I12787)
--	g10351 = NOT(g6802)
--	g23936 = NOT(g19210)
--	g10372 = NOT(g6900)
--	I23327 = NOT(g22647)
--	g25202 = NOT(g23932)
--	g19776 = NOT(g17015)
--	g19785 = NOT(g16987)
--	g34150 = NOT(I32103)
--	I32963 = NOT(g34650)
--	g16159 = NOT(g13584)
--	g22192 = NOT(g19801)
--	g20609 = NOT(g15373)
--	g28274 = NOT(I26799)
--	g15171 = NOT(I17098)
--	g34877 = NOT(I33103)
--	g10175 = NOT(g28)
--	I17723 = NOT(g13177)
--	g12082 = NOT(g9645)
--	g17390 = NOT(g14755)
--	g28593 = NOT(g27727)
--	g32678 = NOT(g31528)
--	g13022 = NOT(g11894)
--	g7522 = NOT(g6661)
--	g23334 = NOT(g20785)
--	g25055 = NOT(g23590)
--	g19147 = NOT(I19786)
--	g30019 = NOT(g29060)
--	g7115 = NOT(g12)
--	g12107 = NOT(g9687)
--	g8808 = NOT(g595)
--	g19754 = NOT(g17062)
--	g7315 = NOT(g1772)
--	g16158 = NOT(g13555)
--	g20608 = NOT(g15171)
--	g25111 = NOT(g23699)
--	g9669 = NOT(g5092)
--	g19355 = NOT(g16027)
--	I12360 = NOT(g528)
--	g25070 = NOT(g23590)
--	g32460 = NOT(g31194)
--	g32686 = NOT(g31579)
--	I22343 = NOT(g19371)
--	g24115 = NOT(g20998)
--	g32939 = NOT(g31327)
--	I18903 = NOT(g16872)
--	g30018 = NOT(g28987)
--	g32383 = NOT(I29913)
--	g19950 = NOT(g15885)
--	g14063 = NOT(g11048)
--	g19370 = NOT(g15915)
--	I19917 = NOT(g18088)
--	I14046 = NOT(g9900)
--	I17148 = NOT(g14442)
--	g16656 = NOT(I17852)
--	g9772 = NOT(I13352)
--	I26638 = NOT(g27965)
--	g20921 = NOT(g15426)
--	g12345 = NOT(g7158)
--	I16476 = NOT(g10430)
--	g14790 = NOT(I16855)
--	g20052 = NOT(g17533)
--	g23964 = NOT(g19147)
--	I23303 = NOT(g21669)
--	g32938 = NOT(g30937)
--	g28034 = NOT(g26365)
--	g33533 = NOT(I31361)
--	g29310 = NOT(g28991)
--	g16680 = NOT(g13223)
--	g24052 = NOT(g21193)
--	I17104 = NOT(g12932)
--	g12940 = NOT(g11744)
--	g17522 = NOT(g14927)
--	g21423 = NOT(g15224)
--	g12399 = NOT(g9920)
--	g9743 = NOT(I13321)
--	I16555 = NOT(g10430)
--	g23423 = NOT(g20871)
--	g8201 = NOT(g1894)
--	g9890 = NOT(g6058)
--	g13305 = NOT(g11048)
--	g6827 = NOT(g1277)
--	g14873 = NOT(I16898)
--	g23216 = NOT(g20924)
--	g11900 = NOT(I14708)
--	g19996 = NOT(g17271)
--	g29379 = NOT(I27749)
--	g29925 = NOT(g28820)
--	g13809 = NOT(I16135)
--	I23381 = NOT(g23322)
--	I15036 = NOT(g799)
--	g8449 = NOT(g3752)
--	g12804 = NOT(g9927)
--	g9011 = NOT(g1422)
--	g19367 = NOT(I19851)
--	g19394 = NOT(g16326)
--	I12451 = NOT(g3092)
--	g6846 = NOT(g2152)
--	g9856 = NOT(g5343)
--	g8575 = NOT(g291)
--	g13036 = NOT(g10981)
--	g32875 = NOT(g31376)
--	g30917 = NOT(I28897)
--	I14827 = NOT(g9686)
--	g11560 = NOT(g7647)
--	g13101 = NOT(I15736)
--	g14209 = NOT(g11415)
--	g7880 = NOT(g1291)
--	g13177 = NOT(I15782)
--	g34917 = NOT(I33143)
--	g8715 = NOT(g4927)
--	g20674 = NOT(g15277)
--	g7595 = NOT(I12067)
--	g23543 = NOT(g21514)
--	g6803 = NOT(g496)
--	g16966 = NOT(g14291)
--	g7537 = NOT(g311)
--	g24184 = NOT(I23396)
--	I18845 = NOT(g6711)
--	I32921 = NOT(g34650)
--	g16631 = NOT(g14454)
--	g14208 = NOT(g11563)
--	I18262 = NOT(g13857)
--	g29944 = NOT(g28911)
--	g22904 = NOT(I22111)
--	g23000 = NOT(g20453)
--	I26578 = NOT(g26941)
--	g23908 = NOT(g20739)
--	g17326 = NOT(I18307)
--	g32837 = NOT(g31327)
--	g31856 = NOT(g29385)
--	I13206 = NOT(g5448)
--	g8833 = NOT(g794)
--	g30077 = NOT(g29057)
--	g9992 = NOT(g5990)
--	g20732 = NOT(g15595)
--	g23569 = NOT(g21611)
--	g25196 = NOT(g22763)
--	g10542 = NOT(g7196)
--	I31610 = NOT(g33149)
--	I23390 = NOT(g23395)
--	g13064 = NOT(g11705)
--	g24732 = NOT(g23042)
--	g14453 = NOT(I16610)
--	g7017 = NOT(g128)
--	I30992 = NOT(g32445)
--	g7243 = NOT(I11892)
--	g19446 = NOT(I19917)
--	g34597 = NOT(I32699)
--	I12776 = NOT(g4207)
--	I13759 = NOT(g6754)
--	I18191 = NOT(g14385)
--	g23568 = NOT(g21611)
--	I33255 = NOT(g34975)
--	I33189 = NOT(g34929)
--	g8584 = NOT(g3639)
--	g8539 = NOT(g3454)
--	g23242 = NOT(g21070)
--	I32973 = NOT(g34714)
--	I29571 = NOT(g31783)
--	g34689 = NOT(I32837)
--	I33270 = NOT(g34982)
--	g34923 = NOT(I33161)
--	g9863 = NOT(g5503)
--	I12355 = NOT(g46)
--	g16289 = NOT(g13223)
--	g9480 = NOT(g559)
--	I17228 = NOT(g13350)
--	g6994 = NOT(g4933)
--	g21123 = NOT(g15615)
--	g18100 = NOT(I18906)
--	g34688 = NOT(I32834)
--	g9713 = NOT(g3618)
--	g10607 = NOT(g10233)
--	g12833 = NOT(I15448)
--	g22847 = NOT(g20283)
--	g16309 = NOT(I17639)
--	I12950 = NOT(g4287)
--	g23814 = NOT(g19074)
--	g10320 = NOT(g817)
--	g32617 = NOT(g30825)
--	g28575 = NOT(g27711)
--	g32470 = NOT(g31566)
--	g10073 = NOT(g134)
--	I18832 = NOT(g13782)
--	I31686 = NOT(g33164)
--	g7328 = NOT(g2197)
--	g32915 = NOT(g31710)
--	g10274 = NOT(g976)
--	g29765 = NOT(I28014)
--	g10530 = NOT(g8922)
--	g7542 = NOT(I12030)
--	I12858 = NOT(g4340)
--	g28711 = NOT(g27886)
--	g13009 = NOT(I15617)
--	g16308 = NOT(I17636)
--	g9569 = NOT(g6227)
--	g13665 = NOT(g11306)
--	g27004 = NOT(g26131)
--	g30102 = NOT(g29157)
--	g8362 = NOT(g194)
--	I13744 = NOT(g3518)
--	g31831 = NOT(g29385)
--	g32201 = NOT(g31509)
--	g24013 = NOT(g21611)
--	I33030 = NOT(g34768)
--	I12151 = NOT(g604)
--	g10122 = NOT(I13623)
--	g6816 = NOT(g933)
--	I12172 = NOT(g2715)
--	g17183 = NOT(I18221)
--	g17673 = NOT(g14723)
--	g17847 = NOT(I18839)
--	I26430 = NOT(g26856)
--	g13008 = NOT(g11855)
--	g15656 = NOT(I17198)
--	I21483 = NOT(g18726)
--	g20329 = NOT(g15277)
--	I33267 = NOT(g34979)
--	g8052 = NOT(g1211)
--	I18861 = NOT(g14307)
--	g21293 = NOT(I21036)
--	g20207 = NOT(g17015)
--	g23230 = NOT(I22327)
--	g15680 = NOT(I17207)
--	g20539 = NOT(g15483)
--	g25001 = NOT(g23666)
--	g17062 = NOT(I18154)
--	g20005 = NOT(g17433)
--	g13485 = NOT(g10476)
--	g20328 = NOT(g15867)
--	g32595 = NOT(g30825)
--	g32467 = NOT(g31194)
--	g32494 = NOT(g30825)
--	g19902 = NOT(g17200)
--	g24005 = NOT(I23149)
--	g17509 = NOT(I18446)
--	g14034 = NOT(g11048)
--	g19957 = NOT(g16540)
--	g16816 = NOT(I18028)
--	g20538 = NOT(g15348)
--	g9688 = NOT(g113)
--	g28606 = NOT(g27762)
--	g6847 = NOT(g2283)
--	g13555 = NOT(g12692)
--	g18882 = NOT(I19674)
--	g32623 = NOT(g30735)
--	g18991 = NOT(g16136)
--	I28897 = NOT(g30155)
--	g19739 = NOT(g16931)
--	I25391 = NOT(g24483)
--	g9976 = NOT(g2537)
--	g17508 = NOT(I18443)
--	g29317 = NOT(I27677)
--	g10153 = NOT(g2417)
--	g23841 = NOT(g19074)
--	I22096 = NOT(g19890)
--	g23992 = NOT(g19210)
--	g32782 = NOT(g30735)
--	g23391 = NOT(g20645)
--	g19146 = NOT(g15574)
--	g19738 = NOT(g15992)
--	g33080 = NOT(I30644)
--	g21510 = NOT(g15647)
--	g23510 = NOT(g18833)
--	g10409 = NOT(g7087)
--	g16752 = NOT(I17976)
--	I21757 = NOT(g21308)
--	I33218 = NOT(g34955)
--	I25579 = NOT(g25297)
--	g16954 = NOT(I18104)
--	g29129 = NOT(g27858)
--	g22213 = NOT(g19147)
--	g19699 = NOT(I20116)
--	g8504 = NOT(g3451)
--	g34511 = NOT(g34419)
--	g10136 = NOT(g6113)
--	g16643 = NOT(I17839)
--	g10408 = NOT(g7049)
--	g9000 = NOT(g632)
--	g32822 = NOT(g30937)
--	g13074 = NOT(I15702)
--	I24191 = NOT(g22360)
--	g29128 = NOT(g27800)
--	g14635 = NOT(I16741)
--	I12227 = NOT(g34)
--	g13239 = NOT(g10632)
--	g19698 = NOT(g16971)
--	g9326 = NOT(g6203)
--	I15238 = NOT(g6351)
--	g12951 = NOT(I15569)
--	g25157 = NOT(g22498)
--	g23578 = NOT(I22725)
--	g8070 = NOT(g3518)
--	g13594 = NOT(g11012)
--	I16438 = NOT(g11165)
--	g23014 = NOT(g20391)
--	I25586 = NOT(g25537)
--	g8470 = NOT(I12605)
--	g20100 = NOT(I20369)
--	g7512 = NOT(g5283)
--	g34660 = NOT(g34473)
--	I30983 = NOT(g32433)
--	g9760 = NOT(g2315)
--	g20771 = NOT(g15171)
--	g22311 = NOT(g18935)
--	g24100 = NOT(g20857)
--	g26054 = NOT(g24804)
--	g7490 = NOT(g2629)
--	I15382 = NOT(g9071)
--	I14647 = NOT(g7717)
--	g25231 = NOT(g22228)
--	g7166 = NOT(g4311)
--	g20235 = NOT(g15277)
--	g19427 = NOT(g16292)
--	I26130 = NOT(g26510)
--	g11941 = NOT(I14761)
--	g19366 = NOT(g15885)
--	I17857 = NOT(g3969)
--	g32853 = NOT(g30673)
--	g24683 = NOT(g23112)
--	g33736 = NOT(I31597)
--	g11519 = NOT(g8481)
--	I14999 = NOT(g10030)
--	g16195 = NOT(g13437)
--	g34480 = NOT(I32535)
--	g16489 = NOT(I17699)
--	g34916 = NOT(I33140)
--	g13675 = NOT(g10556)
--	I20861 = NOT(g16960)
--	g32589 = NOT(g31070)
--	g7456 = NOT(g2495)
--	g15224 = NOT(I17101)
--	g7148 = NOT(I11835)
--	g6817 = NOT(g956)
--	g7649 = NOT(g1345)
--	g22592 = NOT(I21930)
--	g22756 = NOT(g20436)
--	g16525 = NOT(I17723)
--	g15571 = NOT(g13211)
--	g26942 = NOT(I25692)
--	g9924 = NOT(g5644)
--	g10474 = NOT(g8841)
--	g32588 = NOT(g30825)
--	g32524 = NOT(g31070)
--	g9220 = NOT(g843)
--	g31843 = NOT(g29385)
--	g32836 = NOT(g31021)
--	g33696 = NOT(I31535)
--	g30076 = NOT(g29085)
--	g30085 = NOT(g29082)
--	g7851 = NOT(g921)
--	I33075 = NOT(g34843)
--	g9779 = NOT(g5156)
--	g26655 = NOT(g25492)
--	g13637 = NOT(g10556)
--	g20515 = NOT(g15483)
--	g34307 = NOT(g34087)
--	g23041 = NOT(g19882)
--	I20388 = NOT(g17724)
--	g32477 = NOT(g31566)
--	I18360 = NOT(g1426)
--	g21275 = NOT(g15426)
--	g24515 = NOT(g22689)
--	I31494 = NOT(g33283)
--	g24991 = NOT(g22369)
--	I12120 = NOT(g632)
--	g10109 = NOT(g135)
--	g30054 = NOT(g29134)
--	g21430 = NOT(g15608)
--	g27163 = NOT(I25869)
--	g34596 = NOT(I32696)
--	g8406 = NOT(g232)
--	g17756 = NOT(g14858)
--	I27738 = NOT(g28140)
--	g23430 = NOT(I22547)
--	g23746 = NOT(g20902)
--	g23493 = NOT(g21611)
--	g7964 = NOT(g3155)
--	g7260 = NOT(I11908)
--	g8635 = NOT(g2783)
--	g24407 = NOT(g22594)
--	g34243 = NOT(I32228)
--	g29697 = NOT(g28336)
--	g9977 = NOT(g2667)
--	g19481 = NOT(g16349)
--	g10108 = NOT(g120)
--	I14932 = NOT(g9901)
--	g29995 = NOT(g28955)
--	I33037 = NOT(g34770)
--	g34431 = NOT(I32464)
--	g12012 = NOT(g9213)
--	g32118 = NOT(g31008)
--	g15816 = NOT(I17314)
--	g8766 = NOT(g572)
--	g18940 = NOT(I19719)
--	g8087 = NOT(g1157)
--	I31782 = NOT(g33219)
--	g32864 = NOT(g30937)
--	g23237 = NOT(g20924)
--	I19734 = NOT(g17725)
--	g7063 = NOT(g4831)
--	g10606 = NOT(g10233)
--	g21340 = NOT(I21074)
--	g32749 = NOT(g31021)
--	g32616 = NOT(g30735)
--	g23340 = NOT(g21070)
--	g23983 = NOT(g19210)
--	I22128 = NOT(g19968)
--	g34773 = NOT(I32963)
--	g9051 = NOT(g1426)
--	g23684 = NOT(I22819)
--	g25480 = NOT(g22228)
--	g34942 = NOT(g34928)
--	g32748 = NOT(g31710)
--	I15577 = NOT(g10430)
--	g8748 = NOT(g776)
--	g11215 = NOT(g8285)
--	g19127 = NOT(I19775)
--	g9451 = NOT(g5873)
--	g28326 = NOT(g27414)
--	I32991 = NOT(g34759)
--	I14505 = NOT(g10140)
--	I33155 = NOT(g34897)
--	g13215 = NOT(g10909)
--	g26131 = NOT(I25161)
--	g34156 = NOT(g33907)
--	g13729 = NOT(g10951)
--	g25550 = NOT(g22763)
--	g20441 = NOT(g17873)
--	g20584 = NOT(g17873)
--	g32704 = NOT(g31070)
--	I21047 = NOT(g17429)
--	g10381 = NOT(g6957)
--	g28040 = NOT(g26365)
--	g33708 = NOT(I31555)
--	I33170 = NOT(g34890)
--	g19490 = NOT(g16489)
--	g25287 = NOT(g22228)
--	g34670 = NOT(I32794)
--	I29939 = NOT(g31667)
--	g9999 = NOT(g6109)
--	I17128 = NOT(g13835)
--	g23517 = NOT(g21070)
--	g33258 = NOT(g32296)
--	g32809 = NOT(g31327)
--	g32900 = NOT(g30937)
--	g25307 = NOT(g22763)
--	g32466 = NOT(g31070)
--	g7118 = NOT(g832)
--	g7619 = NOT(g1296)
--	g16124 = NOT(g13555)
--	I19487 = NOT(g15125)
--	g19376 = NOT(g17509)
--	g19385 = NOT(g16326)
--	I17626 = NOT(g14582)
--	g17413 = NOT(I18350)
--	g9103 = NOT(g5774)
--	g32808 = NOT(g30937)
--	I26952 = NOT(g27972)
--	g24759 = NOT(g23003)
--	I18071 = NOT(g13680)
--	g19980 = NOT(g17226)
--	g25243 = NOT(g22763)
--	g34839 = NOT(I33053)
--	g17691 = NOT(I18674)
--	g20114 = NOT(I20385)
--	g16686 = NOT(I17892)
--	g34930 = NOT(I33182)
--	g11349 = NOT(I14365)
--	g34993 = NOT(I33279)
--	g12946 = NOT(I15564)
--	g15842 = NOT(g13469)
--	g32560 = NOT(g31070)
--	g20435 = NOT(g15348)
--	g8373 = NOT(g2485)
--	I15906 = NOT(g10430)
--	g24114 = NOT(g20720)
--	g8091 = NOT(g1579)
--	I33167 = NOT(g34890)
--	g6772 = NOT(I11629)
--	g29498 = NOT(I27784)
--	g24082 = NOT(g19890)
--	I15284 = NOT(g6697)
--	g16030 = NOT(g13570)
--	g7393 = NOT(g5320)
--	g13906 = NOT(I16201)
--	g10390 = NOT(g6987)
--	g21362 = NOT(g17873)
--	g24107 = NOT(g20857)
--	g32642 = NOT(g31542)
--	g9732 = NOT(g5481)
--	g23362 = NOT(I22467)
--	g34131 = NOT(I32074)
--	g29056 = NOT(g27800)
--	g22928 = NOT(I22131)
--	g9753 = NOT(g1890)
--	I26516 = NOT(g26824)
--	g23523 = NOT(g21514)
--	g31810 = NOT(g29385)
--	g8283 = NOT(I12493)
--	g25773 = NOT(g24453)
--	I27481 = NOT(g27928)
--	g18833 = NOT(I19661)
--	g31657 = NOT(I29239)
--	g7971 = NOT(g4818)
--	g13304 = NOT(I15872)
--	I20447 = NOT(g16244)
--	I28582 = NOT(g30116)
--	I18825 = NOT(g6019)
--	I18370 = NOT(g14873)
--	g24744 = NOT(g22202)
--	I31477 = NOT(g33391)
--	g29080 = NOT(g27779)
--	g7686 = NOT(g4659)
--	g33375 = NOT(g32377)
--	g8407 = NOT(g1171)
--	g17929 = NOT(I18855)
--	g9072 = NOT(g2994)
--	g25156 = NOT(g22498)
--	I29218 = NOT(g30304)
--	g8920 = NOT(I12899)
--	g8059 = NOT(g3171)
--	g32733 = NOT(g31672)
--	I33119 = NOT(g34852)
--	g14192 = NOT(g11385)
--	I18858 = NOT(g13835)
--	g9472 = NOT(g6555)
--	g19931 = NOT(g17200)
--	g25180 = NOT(g23529)
--	g6856 = NOT(I11682)
--	I12572 = NOT(g51)
--	g15830 = NOT(g13432)
--	g17583 = NOT(g14968)
--	g8718 = NOT(g3333)
--	I18151 = NOT(g13144)
--	g34210 = NOT(I32173)
--	g32874 = NOT(g30673)
--	I28925 = NOT(g29987)
--	g9443 = NOT(g5489)
--	g21727 = NOT(I21300)
--	I22512 = NOT(g19389)
--	g20652 = NOT(I20744)
--	g28508 = NOT(I26989)
--	g32630 = NOT(g30735)
--	g7121 = NOT(I11820)
--	g23863 = NOT(g19210)
--	g32693 = NOT(g31579)
--	I31616 = NOT(g33219)
--	g21222 = NOT(g17430)
--	I23396 = NOT(g23427)
--	g7670 = NOT(g4104)
--	g23222 = NOT(g20785)
--	I18367 = NOT(g13010)
--	g26187 = NOT(I25190)
--	g29342 = NOT(g28188)
--	g9316 = NOT(g5742)
--	g25930 = NOT(I25028)
--	g7625 = NOT(I12109)
--	g32665 = NOT(g31579)
--	I31748 = NOT(g33228)
--	I13473 = NOT(g4157)
--	g19520 = NOT(g16826)
--	g6992 = NOT(g4899)
--	g12760 = NOT(g10272)
--	g9434 = NOT(g5385)
--	g13138 = NOT(I15765)
--	g17787 = NOT(I18795)
--	g7232 = NOT(g4411)
--	g10553 = NOT(g8971)
--	g25838 = NOT(g25250)
--	I27784 = NOT(g29013)
--	I15636 = NOT(g12075)
--	I33276 = NOT(g34985)
--	I33285 = NOT(g34988)
--	g18947 = NOT(g16136)
--	I27385 = NOT(g27438)
--	g30039 = NOT(g29134)
--	g30306 = NOT(g28796)
--	g25131 = NOT(g23699)
--	I33053 = NOT(g34778)
--	g15705 = NOT(g13217)
--	g26937 = NOT(I25683)
--	g17302 = NOT(I18285)
--	g32892 = NOT(g31021)
--	g23347 = NOT(I22444)
--	g24135 = NOT(g20720)
--	g32476 = NOT(g30673)
--	g32485 = NOT(g31376)
--	g33459 = NOT(I30995)
--	I31466 = NOT(g33318)
--	g7909 = NOT(g936)
--	g30038 = NOT(g29097)
--	g23253 = NOT(g21037)
--	I12103 = NOT(g572)
--	g11852 = NOT(I14668)
--	g17743 = NOT(I18734)
--	g9681 = NOT(g5798)
--	I22499 = NOT(g21160)
--	g10040 = NOT(g2652)
--	I22316 = NOT(g19361)
--	g32555 = NOT(g30673)
--	I18446 = NOT(g13028)
--	g14536 = NOT(I16651)
--	g19860 = NOT(g17226)
--	g33458 = NOT(I30992)
--	g7519 = NOT(g1157)
--	g24361 = NOT(g22885)
--	g11963 = NOT(g9153)
--	g25557 = NOT(g22763)
--	g32570 = NOT(g31554)
--	g32712 = NOT(g30614)
--	g25210 = NOT(g23802)
--	g32914 = NOT(g31672)
--	I25351 = NOT(g24466)
--	g9914 = NOT(g2533)
--	I20355 = NOT(g17613)
--	g33918 = NOT(I31782)
--	g23236 = NOT(g20785)
--	g20500 = NOT(g17873)
--	g10621 = NOT(g7567)
--	g34677 = NOT(I32815)
--	g29365 = NOT(g29067)
--	g14252 = NOT(I16438)
--	I22989 = NOT(g21175)
--	g13664 = NOT(g11252)
--	g20049 = NOT(I20318)
--	g23952 = NOT(g19277)
--	g23351 = NOT(g20924)
--	g32907 = NOT(g30937)
--	I31642 = NOT(g33204)
--	g33079 = NOT(I30641)
--	g24049 = NOT(g20014)
--	I14896 = NOT(g9820)
--	g29960 = NOT(g28885)
--	g21175 = NOT(I20951)
--	g22881 = NOT(I22096)
--	g23821 = NOT(g19210)
--	g10564 = NOT(g9462)
--	g15938 = NOT(I17401)
--	g16075 = NOT(g13597)
--	g9413 = NOT(g1744)
--	g19659 = NOT(g17062)
--	g14564 = NOT(I16679)
--	g24048 = NOT(g19968)
--	I11682 = NOT(g2756)
--	g11576 = NOT(g8542)
--	I33064 = NOT(g34784)
--	I25790 = NOT(g26424)
--	I17989 = NOT(g14173)
--	g20004 = NOT(g17249)
--	g13484 = NOT(g10981)
--	g32567 = NOT(g31070)
--	g32594 = NOT(g30735)
--	g19658 = NOT(g16987)
--	g23264 = NOT(g21037)
--	g25286 = NOT(g22228)
--	g16623 = NOT(g14127)
--	g10183 = NOT(g2595)
--	I15609 = NOT(g12013)
--	g7586 = NOT(I12056)
--	g23516 = NOT(g20924)
--	g25039 = NOT(g22498)
--	I28548 = NOT(g28147)
--	g10397 = NOT(g7018)
--	g6976 = NOT(I11750)
--	g14183 = NOT(g12381)
--	g14673 = NOT(I16770)
--	g11609 = NOT(g7660)
--	g9820 = NOT(g99)
--	g16782 = NOT(I18006)
--	g12903 = NOT(g10411)
--	g20613 = NOT(g15224)
--	I21787 = NOT(g19422)
--	I22461 = NOT(g21225)
--	g31817 = NOT(g29385)
--	g13312 = NOT(g11048)
--	I18301 = NOT(g12976)
--	g32941 = NOT(g30735)
--	g32382 = NOT(g31657)
--	g11608 = NOT(g7659)
--	g19644 = NOT(g17953)
--	g10509 = NOT(g10233)
--	I18120 = NOT(g13350)
--	g32519 = NOT(g30673)
--	I22031 = NOT(g21387)
--	I27546 = NOT(g29041)
--	g32185 = NOT(I29717)
--	g18421 = NOT(I19235)
--	g14509 = NOT(I16626)
--	I15921 = NOT(g12381)
--	g32675 = NOT(g31070)
--	g8388 = NOT(g3010)
--	I23357 = NOT(g23359)
--	g20273 = NOT(g17128)
--	g20106 = NOT(g17328)
--	g12563 = NOT(g9864)
--	g20605 = NOT(g17955)
--	g21422 = NOT(g15373)
--	I26409 = NOT(g26187)
--	g30217 = NOT(I28458)
--	g8216 = NOT(g3092)
--	g10851 = NOT(I14069)
--	I12089 = NOT(g744)
--	g10872 = NOT(g7567)
--	g9601 = NOT(g4005)
--	g23422 = NOT(g21611)
--	g32518 = NOT(g30614)
--	I16328 = NOT(g878)
--	g24106 = NOT(g19984)
--	g24605 = NOT(g23139)
--	I14050 = NOT(g9963)
--	g29043 = NOT(I27391)
--	I16538 = NOT(g10417)
--	g13745 = NOT(I16102)
--	g32637 = NOT(g30735)
--	g31656 = NOT(I29236)
--	I20318 = NOT(g16920)
--	g17249 = NOT(I18265)
--	I28002 = NOT(g28153)
--	g32935 = NOT(g31672)
--	g24463 = NOT(g23578)
--	I21769 = NOT(g19402)
--	I17650 = NOT(g13271)
--	I28128 = NOT(g28314)
--	g20033 = NOT(g16579)
--	g31823 = NOT(g29385)
--	I32613 = NOT(g34329)
--	g32883 = NOT(g30735)
--	g17248 = NOT(I18262)
--	I30641 = NOT(g32024)
--	I31555 = NOT(g33212)
--	I14742 = NOT(g9534)
--	g19411 = NOT(g16489)
--	g19527 = NOT(g16349)
--	g17710 = NOT(g14764)
--	g24033 = NOT(g19919)
--	I17198 = NOT(g13809)
--	g12845 = NOT(g10358)
--	g27990 = NOT(g26770)
--	g16853 = NOT(g13584)
--	I12497 = NOT(g49)
--	g23542 = NOT(g21514)
--	g9581 = NOT(g91)
--	g23021 = NOT(g20283)
--	g23453 = NOT(I22576)
--	g10213 = NOT(g6732)
--	I32947 = NOT(g34659)
--	g12899 = NOT(g10407)
--	g21726 = NOT(I21297)
--	g16589 = NOT(g14082)
--	g25169 = NOT(g22763)
--	g29955 = NOT(g28950)
--	g9060 = NOT(g3355)
--	I32106 = NOT(g33653)
--	g23913 = NOT(g19147)
--	g15915 = NOT(I17392)
--	g9460 = NOT(g6154)
--	g24795 = NOT(g23342)
--	g29970 = NOT(I28199)
--	g7659 = NOT(I12141)
--	g12898 = NOT(g10405)
--	g22647 = NOT(I21959)
--	g17778 = NOT(I18778)
--	g16588 = NOT(g13929)
--	g25168 = NOT(I24334)
--	g23614 = NOT(g20248)
--	g25410 = NOT(g22228)
--	g18829 = NOT(g15171)
--	I12987 = NOT(g12)
--	I15732 = NOT(g6692)
--	g8741 = NOT(g4821)
--	g10047 = NOT(g5421)
--	I32812 = NOT(g34588)
--	g19503 = NOT(g16349)
--	g29878 = NOT(g28421)
--	g15277 = NOT(I17104)
--	g21607 = NOT(g17873)
--	g22999 = NOT(g20453)
--	g23607 = NOT(g21611)
--	g21905 = NOT(I21486)
--	g14205 = NOT(g12381)
--	g26654 = NOT(g25275)
--	g20514 = NOT(g15348)
--	I25530 = NOT(g25222)
--	g32501 = NOT(g30825)
--	g32729 = NOT(g30937)
--	g18828 = NOT(g17955)
--	g31631 = NOT(I29221)
--	g10311 = NOT(g4633)
--	g23320 = NOT(I22419)
--	g23905 = NOT(g21514)
--	g9739 = NOT(g5752)
--	g32577 = NOT(g31554)
--	g33631 = NOT(I31459)
--	I14730 = NOT(g7717)
--	g18946 = NOT(g16100)
--	g29171 = NOT(g27937)
--	g21274 = NOT(g15373)
--	g14912 = NOT(I16917)
--	g30321 = NOT(I28572)
--	g23274 = NOT(g21070)
--	g20507 = NOT(g15509)
--	g23530 = NOT(g20248)
--	g22998 = NOT(g20391)
--	g27832 = NOT(I26409)
--	I32234 = NOT(g34126)
--	g34922 = NOT(I33158)
--	I24281 = NOT(g23440)
--	g26936 = NOT(I25680)
--	g15595 = NOT(I17173)
--	g32728 = NOT(g31021)
--	g21346 = NOT(g17821)
--	g25015 = NOT(g23662)
--	g6977 = NOT(I11753)
--	I20957 = NOT(g16228)
--	g19714 = NOT(g16821)
--	I13240 = NOT(g5794)
--	g7275 = NOT(g1728)
--	g22182 = NOT(I21766)
--	g29967 = NOT(g28946)
--	g29994 = NOT(g29049)
--	g34531 = NOT(I32594)
--	g9995 = NOT(g6035)
--	I12644 = NOT(g3689)
--	I11903 = NOT(g4414)
--	g23565 = NOT(g21562)
--	g10072 = NOT(g9)
--	g32438 = NOT(g30991)
--	I14690 = NOT(g9340)
--	g8883 = NOT(g4709)
--	g7615 = NOT(I12083)
--	g12440 = NOT(g9985)
--	g27573 = NOT(g26667)
--	I20562 = NOT(g16525)
--	g25556 = NOT(g22763)
--	g24163 = NOT(I23333)
--	I33176 = NOT(g34887)
--	g7174 = NOT(g6052)
--	g19979 = NOT(g17226)
--	g16748 = NOT(I17970)
--	g7374 = NOT(g2227)
--	g12861 = NOT(g10367)
--	g17651 = NOT(g14868)
--	g17672 = NOT(g14720)
--	g34676 = NOT(I32812)
--	g8217 = NOT(g3143)
--	I16515 = NOT(g12477)
--	I17471 = NOT(g13394)
--	g9390 = NOT(g5808)
--	g21292 = NOT(I21033)
--	g11214 = NOT(g9602)
--	g32906 = NOT(g31021)
--	g7985 = NOT(g3506)
--	g16285 = NOT(I17612)
--	g8466 = NOT(g1514)
--	I19762 = NOT(g15732)
--	g22449 = NOT(g19597)
--	g34654 = NOT(I32766)
--	g20541 = NOT(g17821)
--	I12855 = NOT(g4311)
--	g16305 = NOT(g13346)
--	g10350 = NOT(g6800)
--	g13329 = NOT(I15893)
--	g16053 = NOT(I17442)
--	g9501 = NOT(g5731)
--	g6999 = NOT(g86)
--	g16809 = NOT(g14387)
--	g21409 = NOT(g18008)
--	g22897 = NOT(g21024)
--	g7239 = NOT(g5033)
--	I12411 = NOT(g4809)
--	g23409 = NOT(g21514)
--	g8165 = NOT(g3530)
--	g32622 = NOT(g31376)
--	g8571 = NOT(g57)
--	g8365 = NOT(g2060)
--	I26381 = NOT(g26851)
--	g24789 = NOT(g23309)
--	g32566 = NOT(g30825)
--	g19741 = NOT(g16987)
--	I30537 = NOT(g32027)
--	g29079 = NOT(g27742)
--	g7380 = NOT(g2331)
--	g21408 = NOT(g15373)
--	g10152 = NOT(g2122)
--	g7591 = NOT(g6668)
--	g23408 = NOT(g21468)
--	g8055 = NOT(g1236)
--	g10396 = NOT(g6997)
--	g20325 = NOT(g15171)
--	g24359 = NOT(g22550)
--	g19067 = NOT(g15979)
--	g20920 = NOT(g15426)
--	g20535 = NOT(g17847)
--	I13990 = NOT(g7636)
--	g20434 = NOT(g18065)
--	g9704 = NOT(g2575)
--	g31816 = NOT(g29385)
--	g8133 = NOT(g4809)
--	g24920 = NOT(I24089)
--	g24535 = NOT(g22942)
--	I18376 = NOT(g14332)
--	g24358 = NOT(g22550)
--	I18297 = NOT(g1418)
--	I12503 = NOT(g215)
--	g17505 = NOT(g14899)
--	g17404 = NOT(I18337)
--	g10413 = NOT(g7110)
--	g8774 = NOT(g781)
--	g32653 = NOT(g30825)
--	g19801 = NOT(I20216)
--	I32473 = NOT(g34248)
--	g17717 = NOT(g14937)
--	I17879 = NOT(g14386)
--	g34423 = NOT(g34222)
--	g15588 = NOT(I17166)
--	I22886 = NOT(g18926)
--	g32138 = NOT(g31233)
--	I17970 = NOT(g4027)
--	I20895 = NOT(g16954)
--	g24121 = NOT(g20720)
--	I18888 = NOT(g16644)
--	g8396 = NOT(g3401)
--	g9250 = NOT(g1600)
--	g34587 = NOT(I32671)
--	I13718 = NOT(g890)
--	g12997 = NOT(g11826)
--	g10405 = NOT(g7064)
--	g32636 = NOT(g31376)
--	I23998 = NOT(g22182)
--	I32788 = NOT(g34577)
--	g32415 = NOT(g31591)
--	g14405 = NOT(g12170)
--	g19695 = NOT(g17015)
--	g8538 = NOT(g3412)
--	I12819 = NOT(g4277)
--	g29977 = NOT(g28920)
--	I12910 = NOT(g4340)
--	g16874 = NOT(I18066)
--	g32852 = NOT(g30614)
--	g11235 = NOT(I14301)
--	I32535 = NOT(g34296)
--	I25327 = NOT(g24641)
--	g8509 = NOT(g4141)
--	g35002 = NOT(I33300)
--	g19526 = NOT(g16349)
--	g16630 = NOT(g14142)
--	g16693 = NOT(I17901)
--	g26814 = NOT(g25221)
--	g34543 = NOT(g34359)
--	I22425 = NOT(g19379)
--	g24173 = NOT(I23363)
--	g32963 = NOT(g30825)
--	g22148 = NOT(g19074)
--	g7515 = NOT(I12000)
--	g12871 = NOT(g10378)
--	g29353 = NOT(I27713)
--	I12070 = NOT(g785)
--	I22458 = NOT(g18954)
--	g23537 = NOT(g20785)
--	g9568 = NOT(g6181)
--	g31842 = NOT(g29385)
--	g32664 = NOT(g31528)
--	g30569 = NOT(I28838)
--	I16345 = NOT(g881)
--	g8418 = NOT(g2619)
--	I19772 = NOT(g17818)
--	g34569 = NOT(I32639)
--	g22646 = NOT(g19389)
--	I22918 = NOT(g21451)
--	g17433 = NOT(I18382)
--	I25606 = NOT(g25465)
--	g8290 = NOT(g218)
--	I17425 = NOT(g13416)
--	g18903 = NOT(g15758)
--	g30568 = NOT(g29339)
--	g23283 = NOT(g20785)
--	g19866 = NOT(g16540)
--	g11991 = NOT(g9485)
--	I17919 = NOT(g14609)
--	g13414 = NOT(g11048)
--	I22444 = NOT(g19626)
--	g23492 = NOT(g21562)
--	g25423 = NOT(I24558)
--	g23303 = NOT(g20785)
--	I31622 = NOT(g33204)
--	g32576 = NOT(g30614)
--	g24134 = NOT(g19984)
--	g8093 = NOT(g1624)
--	g32484 = NOT(g31566)
--	g34242 = NOT(I32225)
--	g24029 = NOT(g20982)
--	g33424 = NOT(g32415)
--	I11701 = NOT(g4164)
--	g10113 = NOT(g2084)
--	g17811 = NOT(g12925)
--	g17646 = NOT(I18609)
--	I11777 = NOT(g5357)
--	g20506 = NOT(g15426)
--	I28199 = NOT(g28803)
--	I25750 = NOT(g26823)
--	g20028 = NOT(g15371)
--	I12067 = NOT(g739)
--	I32173 = NOT(g33645)
--	g32554 = NOT(g30614)
--	I18089 = NOT(g13144)
--	g24506 = NOT(I23711)
--	I20385 = NOT(g16194)
--	g7750 = NOT(g1070)
--	g24028 = NOT(g20841)
--	I24784 = NOT(g24265)
--	g34123 = NOT(I32062)
--	g16712 = NOT(g13223)
--	g26841 = NOT(g24893)
--	g32609 = NOT(g30735)
--	g21381 = NOT(g18008)
--	I27735 = NOT(g28779)
--	I29239 = NOT(g29498)
--	g31830 = NOT(g29385)
--	g23982 = NOT(g19147)
--	g10357 = NOT(g6825)
--	g26510 = NOT(I25369)
--	g14357 = NOT(g12181)
--	g34772 = NOT(I32960)
--	I12735 = NOT(g4572)
--	g8181 = NOT(g424)
--	g28779 = NOT(I27253)
--	g32608 = NOT(g31376)
--	g8381 = NOT(g2610)
--	g19689 = NOT(g16795)
--	g7040 = NOT(g4821)
--	g25117 = NOT(g22417)
--	I16135 = NOT(g10430)
--	g25000 = NOT(g23630)
--	g8685 = NOT(g1430)
--	g7440 = NOT(g329)
--	g8700 = NOT(g4054)
--	g28081 = NOT(I26584)
--	g32921 = NOT(g31672)
--	g33713 = NOT(I31564)
--	g8397 = NOT(g3470)
--	g19688 = NOT(g16777)
--	g9626 = NOT(g6466)
--	g8021 = NOT(g3512)
--	g16594 = NOT(I17772)
--	g26835 = NOT(I25555)
--	g13584 = NOT(g12735)
--	g18990 = NOT(g16136)
--	g32745 = NOT(g31376)
--	I29185 = NOT(g30012)
--	g22896 = NOT(g21012)
--	I18700 = NOT(g6027)
--	g23840 = NOT(g19074)
--	g15733 = NOT(I17249)
--	g32799 = NOT(g31710)
--	g18898 = NOT(g15566)
--	g23390 = NOT(g21468)
--	g32813 = NOT(g31710)
--	g22228 = NOT(I21810)
--	g6820 = NOT(g1070)
--	g33705 = NOT(I31550)
--	g25242 = NOT(g23684)
--	g7666 = NOT(g4076)
--	I17159 = NOT(g13350)
--	g20649 = NOT(g18065)
--	I17125 = NOT(g13809)
--	I22561 = NOT(g20841)
--	I23149 = NOT(g19061)
--	g31189 = NOT(I29002)
--	g34992 = NOT(I33276)
--	I17901 = NOT(g3976)
--	g34391 = NOT(g34200)
--	g32798 = NOT(g31672)
--	I22353 = NOT(g19375)
--	g28380 = NOT(g27064)
--	g20240 = NOT(g17847)
--	I23387 = NOT(g23394)
--	g32973 = NOT(g31021)
--	I30904 = NOT(g32424)
--	g34510 = NOT(g34418)
--	g22716 = NOT(g19795)
--	g23192 = NOT(g20248)
--	g16675 = NOT(I17873)
--	g20648 = NOT(g15615)
--	g10881 = NOT(g7567)
--	I17783 = NOT(g13304)
--	g20903 = NOT(g17249)
--	g32805 = NOT(g31672)
--	g13082 = NOT(g10981)
--	g32674 = NOT(g30735)
--	g24648 = NOT(g23148)
--	g7528 = NOT(g930)
--	g12859 = NOT(g10366)
--	g13107 = NOT(g10476)
--	g34579 = NOT(I32659)
--	g7648 = NOT(I12135)
--	g26615 = NOT(g25432)
--	g12950 = NOT(g12708)
--	g20604 = NOT(g17873)
--	g9683 = NOT(g6140)
--	g23522 = NOT(g21514)
--	g18832 = NOT(g15634)
--	I13360 = NOT(g5343)
--	g24604 = NOT(g23112)
--	g30578 = NOT(g29956)
--	g33460 = NOT(I30998)
--	g33686 = NOT(g33187)
--	g19885 = NOT(g17249)
--	g26720 = NOT(g25275)
--	g7655 = NOT(g4332)
--	g11744 = NOT(I14602)
--	g20770 = NOT(g17955)
--	I26508 = NOT(g26814)
--	g9778 = NOT(g5069)
--	I14271 = NOT(g8456)
--	g20563 = NOT(g15171)
--	g27996 = NOT(I26508)
--	g32732 = NOT(g30825)
--	g24770 = NOT(g22763)
--	g8631 = NOT(g283)
--	g25230 = NOT(g23314)
--	g32934 = NOT(g30735)
--	g24981 = NOT(g22763)
--	I24089 = NOT(g22409)
--	g11849 = NOT(g7601)
--	I16613 = NOT(g10430)
--	g17582 = NOT(g14768)
--	g12996 = NOT(g11823)
--	g10027 = NOT(g6523)
--	g23483 = NOT(g18833)
--	I18060 = NOT(g14198)
--	I23369 = NOT(g23347)
--	g14662 = NOT(I16762)
--	g8301 = NOT(g1399)
--	g19763 = NOT(g16431)
--	g25265 = NOT(I24455)
--	I32240 = NOT(g34131)
--	g29976 = NOT(g29018)
--	g12844 = NOT(g10360)
--	g7410 = NOT(g2008)
--	g11398 = NOT(I14409)
--	g23862 = NOT(g19147)
--	g12367 = NOT(I15205)
--	g32692 = NOT(g31528)
--	g32761 = NOT(g30825)
--	I32648 = NOT(g34371)
--	g18926 = NOT(I19707)
--	I18855 = NOT(g13745)
--	I11629 = NOT(g19)
--	g11652 = NOT(g7674)
--	g9661 = NOT(g3661)
--	g13141 = NOT(g11374)
--	g29374 = NOT(I27742)
--	g20767 = NOT(g17873)
--	g26340 = NOT(g24953)
--	g21326 = NOT(I21058)
--	g18099 = NOT(I18903)
--	I18411 = NOT(g13018)
--	g30116 = NOT(I28349)
--	I14650 = NOT(g9340)
--	g33875 = NOT(I31727)
--	I24497 = NOT(g22592)
--	g10710 = NOT(I14006)
--	g20899 = NOT(I20861)
--	I12300 = NOT(g1157)
--	g10003 = NOT(I13539)
--	g23948 = NOT(g21012)
--	I32770 = NOT(g34505)
--	g18098 = NOT(I18900)
--	g10204 = NOT(g2685)
--	I29438 = NOT(g30610)
--	g21904 = NOT(I21483)
--	g14204 = NOT(g12155)
--	g16577 = NOT(I17747)
--	g20633 = NOT(g15171)
--	g23904 = NOT(g18997)
--	I16371 = NOT(g887)
--	g31837 = NOT(g29385)
--	g14779 = NOT(I16847)
--	g21252 = NOT(g15656)
--	I22289 = NOT(g19446)
--	g32329 = NOT(g31522)
--	g29669 = NOT(I27941)
--	g34275 = NOT(g34047)
--	g19480 = NOT(g16349)
--	g23252 = NOT(I22353)
--	g17603 = NOT(g14993)
--	g20191 = NOT(g17821)
--	g34430 = NOT(I32461)
--	g17742 = NOT(g14971)
--	g32539 = NOT(g31170)
--	g10081 = NOT(g2279)
--	g17096 = NOT(I18168)
--	I18894 = NOT(g16708)
--	g6995 = NOT(g4944)
--	g7618 = NOT(I12092)
--	g8441 = NOT(g3361)
--	g22857 = NOT(g20739)
--	I22571 = NOT(g20097)
--	I11785 = NOT(g5703)
--	g7235 = NOT(g4521)
--	g7343 = NOT(g5290)
--	I14365 = NOT(g3303)
--	g30237 = NOT(I28480)
--	I16795 = NOT(g5637)
--	g25007 = NOT(g22457)
--	g32538 = NOT(g31070)
--	g24718 = NOT(g22182)
--	I32794 = NOT(g34580)
--	g14786 = NOT(g12471)
--	g29195 = NOT(I27495)
--	g9484 = NOT(g1612)
--	g30983 = NOT(g29657)
--	g9439 = NOT(g5428)
--	g17681 = NOT(g14735)
--	g7566 = NOT(I12049)
--	g6840 = NOT(g1992)
--	g8673 = NOT(g4737)
--	g16349 = NOT(I17661)
--	g34983 = NOT(I33249)
--	g18997 = NOT(I19756)
--	g10356 = NOT(g6819)
--	g33455 = NOT(I30983)
--	g21183 = NOT(g15509)
--	g21673 = NOT(I21234)
--	g7693 = NOT(g4849)
--	g11833 = NOT(g8026)
--	g17429 = NOT(I18370)
--	g7134 = NOT(g5029)
--	g21397 = NOT(g15171)
--	g23847 = NOT(g19210)
--	g13049 = NOT(I15677)
--	g10380 = NOT(g6960)
--	g30142 = NOT(g28754)
--	g18061 = NOT(g14800)
--	g16284 = NOT(I17609)
--	g19431 = NOT(g16249)
--	g34142 = NOT(I32089)
--	g25116 = NOT(g22369)
--	g17428 = NOT(I18367)
--	I22816 = NOT(g19862)
--	g7548 = NOT(g1036)
--	g11048 = NOT(I14158)
--	g8669 = NOT(g3767)
--	g10090 = NOT(g5348)
--	g20573 = NOT(g17384)
--	g10233 = NOT(I13699)
--	g20247 = NOT(g17015)
--	g29893 = NOT(g28755)
--	I24060 = NOT(g22202)
--	g16622 = NOT(g14104)
--	g23509 = NOT(g21611)
--	g10182 = NOT(g2681)
--	g28620 = NOT(g27679)
--	I21959 = NOT(g20242)
--	g20389 = NOT(g15277)
--	g8058 = NOT(g3115)
--	I14708 = NOT(g9417)
--	I28458 = NOT(g28443)
--	I29139 = NOT(g29382)
--	g8531 = NOT(g3288)
--	g19773 = NOT(g17615)
--	g24389 = NOT(g22908)
--	g8458 = NOT(g294)
--	g24045 = NOT(g21193)
--	g12902 = NOT(g10409)
--	g20612 = NOT(g18008)
--	g23508 = NOT(g21562)
--	I16163 = NOT(g11930)
--	I20870 = NOT(g16216)
--	g32771 = NOT(g31021)
--	g8743 = NOT(g550)
--	g20388 = NOT(g17297)
--	g20324 = NOT(g17955)
--	g8890 = NOT(g376)
--	I23378 = NOT(g23426)
--	g29713 = NOT(I27970)
--	g24099 = NOT(g20720)
--	g24388 = NOT(g22885)
--	g20701 = NOT(g17955)
--	g20777 = NOT(g15224)
--	g20534 = NOT(g17183)
--	g22317 = NOT(g19801)
--	g31623 = NOT(g29669)
--	g32683 = NOT(g30614)
--	I17976 = NOT(g13638)
--	g25465 = NOT(g23824)
--	g19670 = NOT(g16897)
--	g24534 = NOT(g22670)
--	g8505 = NOT(g3480)
--	g20272 = NOT(g17239)
--	g34130 = NOT(I32071)
--	g24098 = NOT(g19984)
--	g14331 = NOT(I16489)
--	g12738 = NOT(g9374)
--	I19863 = NOT(g16675)
--	g9616 = NOT(g5452)
--	g17504 = NOT(g15021)
--	I16541 = NOT(g11929)
--	g8011 = NOT(g3167)
--	g25340 = NOT(g22763)
--	g25035 = NOT(g23699)
--	I17374 = NOT(g13638)
--	g8411 = NOT(I12577)
--	g8734 = NOT(g4045)
--	g19734 = NOT(g16861)
--	g13106 = NOT(g10981)
--	g27698 = NOT(g26648)
--	g29042 = NOT(I27388)
--	g13605 = NOT(I16040)
--	g10897 = NOT(g7601)
--	I33214 = NOT(g34954)
--	I20867 = NOT(g16216)
--	I27314 = NOT(g28009)
--	g6954 = NOT(g4138)
--	g19930 = NOT(g17200)
--	g6810 = NOT(g723)
--	g9527 = NOT(g6500)
--	I14069 = NOT(g9104)
--	g11812 = NOT(g7567)
--	g7202 = NOT(g4639)
--	I16724 = NOT(g12108)
--	g10404 = NOT(g7026)
--	I12314 = NOT(g1500)
--	g13463 = NOT(g10476)
--	g31822 = NOT(g29385)
--	g32515 = NOT(g30825)
--	I31539 = NOT(g33212)
--	g32882 = NOT(g31376)
--	I14602 = NOT(g9340)
--	I15033 = NOT(g10273)
--	g19694 = NOT(g16429)
--	g7908 = NOT(g4157)
--	I32388 = NOT(g34153)
--	g24032 = NOT(g21256)
--	g22626 = NOT(I21941)
--	I21802 = NOT(g21308)
--	I16829 = NOT(g6715)
--	g25517 = NOT(g22228)
--	g11033 = NOT(g8500)
--	g11371 = NOT(g7565)
--	I16535 = NOT(g11235)
--	g18911 = NOT(g15169)
--	g23452 = NOT(g21468)
--	g10026 = NOT(g6494)
--	g32407 = NOT(I29939)
--	g9546 = NOT(g2437)
--	g13033 = NOT(g11917)
--	g21205 = NOT(g15656)
--	g11234 = NOT(g8355)
--	g10212 = NOT(g6390)
--	I14970 = NOT(g9965)
--	g29939 = NOT(g28857)
--	g17128 = NOT(I18180)
--	g7518 = NOT(g1024)
--	I17668 = NOT(g13279)
--	I20819 = NOT(g17088)
--	I22525 = NOT(g19345)
--	I22488 = NOT(g18984)
--	I17842 = NOT(g13051)
--	I20910 = NOT(g17197)
--	g16963 = NOT(I18117)
--	g23912 = NOT(g19147)
--	I17392 = NOT(g13680)
--	g34222 = NOT(I32195)
--	g9970 = NOT(g1714)
--	g24061 = NOT(g19919)
--	I29585 = NOT(g31655)
--	g29093 = NOT(g27858)
--	g34437 = NOT(I32482)
--	g20766 = NOT(g17433)
--	I26929 = NOT(g27980)
--	g8080 = NOT(g3863)
--	I18526 = NOT(g13055)
--	g31853 = NOT(g29385)
--	g19502 = NOT(g15674)
--	g8480 = NOT(g3147)
--	g19210 = NOT(I19796)
--	g17533 = NOT(I18482)
--	g25193 = NOT(g22763)
--	g8713 = NOT(g4826)
--	g21051 = NOT(g15171)
--	g7593 = NOT(I12061)
--	I17488 = NOT(g13394)
--	g15348 = NOT(I17111)
--	g19618 = NOT(g16349)
--	g19443 = NOT(g16449)
--	I14967 = NOT(g9964)
--	g12895 = NOT(g10403)
--	I12773 = NOT(g4204)
--	g16585 = NOT(g14075)
--	g13514 = NOT(I15987)
--	g25523 = NOT(g22550)
--	g31836 = NOT(g29385)
--	g32441 = NOT(I29969)
--	g32584 = NOT(g30673)
--	I32997 = NOT(g34760)
--	g24360 = NOT(g22228)
--	g29219 = NOT(I27573)
--	g15566 = NOT(I17143)
--	g20447 = NOT(g15426)
--	g14149 = NOT(g12381)
--	g10387 = NOT(g6996)
--	g16609 = NOT(g14454)
--	g19469 = NOT(g16326)
--	I28336 = NOT(g29147)
--	g10620 = NOT(g10233)
--	g17737 = NOT(g14810)
--	g22856 = NOT(g20453)
--	g29218 = NOT(I27570)
--	g22995 = NOT(g20330)
--	g32759 = NOT(g31376)
--	g16200 = NOT(g13584)
--	I33235 = NOT(g34957)
--	g23350 = NOT(g20785)
--	g25006 = NOT(g22417)
--	g32725 = NOT(g30825)
--	g24162 = NOT(I23330)
--	I32766 = NOT(g34522)
--	g7933 = NOT(g907)
--	g16608 = NOT(g14116)
--	g19468 = NOT(g15938)
--	g9617 = NOT(I13240)
--	g23820 = NOT(g19147)
--	g34952 = NOT(g34942)
--	g34351 = NOT(g34174)
--	g13012 = NOT(I15626)
--	g32758 = NOT(g31327)
--	g7521 = NOT(g5630)
--	I32871 = NOT(g34521)
--	g25222 = NOT(I24400)
--	g7050 = NOT(g5845)
--	g20629 = NOT(g17955)
--	g23152 = NOT(g20283)
--	I12930 = NOT(g4349)
--	I13699 = NOT(g4581)
--	g9516 = NOT(g6116)
--	I21002 = NOT(g16709)
--	g20451 = NOT(g15277)
--	g21396 = NOT(g17955)
--	g31616 = NOT(I29214)
--	I14079 = NOT(g7231)
--	g30063 = NOT(g29015)
--	I22124 = NOT(g21300)
--	g9771 = NOT(g3969)
--	I29973 = NOT(g31213)
--	g26834 = NOT(I25552)
--	g20911 = NOT(g15171)
--	I16028 = NOT(g12381)
--	g10369 = NOT(g6873)
--	g32744 = NOT(g31327)
--	I31515 = NOT(g33187)
--	g24911 = NOT(I24078)
--	g19677 = NOT(g17096)
--	I18280 = NOT(g12951)
--	g12490 = NOT(I15316)
--	g17512 = NOT(g12983)
--	I17679 = NOT(g13416)
--	g21413 = NOT(g15585)
--	g9299 = NOT(g5124)
--	I15788 = NOT(g10430)
--	g23413 = NOT(g21012)
--	g27956 = NOT(I26466)
--	g32849 = NOT(g31021)
--	g9547 = NOT(g2735)
--	g10368 = NOT(g6887)
--	g32940 = NOT(g31376)
--	g7379 = NOT(g2299)
--	g8400 = NOT(g4836)
--	g11724 = NOT(I14593)
--	I17188 = NOT(g13782)
--	g31809 = NOT(g29385)
--	I12487 = NOT(g3443)
--	g11325 = NOT(g7543)
--	g20071 = NOT(g16826)
--	g32848 = NOT(g30825)
--	g9892 = NOT(g6428)
--	g24071 = NOT(g20841)
--	g11829 = NOT(I14653)
--	g12889 = NOT(g10396)
--	g11920 = NOT(I14730)
--	I11632 = NOT(g16)
--	g20591 = NOT(g15509)
--	g25781 = NOT(g24510)
--	g10412 = NOT(g7072)
--	g20776 = NOT(g18008)
--	g20785 = NOT(I20846)
--	g31808 = NOT(g29385)
--	g32652 = NOT(g30735)
--	g32804 = NOT(g30735)
--	g14412 = NOT(I16564)
--	g7289 = NOT(g4382)
--	I12618 = NOT(g3338)
--	g12888 = NOT(g10395)
--	g26614 = NOT(g25426)
--	g10133 = NOT(g6049)
--	g20147 = NOT(g17328)
--	I17938 = NOT(g3676)
--	g34209 = NOT(I32170)
--	g7835 = NOT(g4125)
--	g24147 = NOT(g19402)
--	g10229 = NOT(g6736)
--	I18066 = NOT(g3317)
--	g12181 = NOT(g9478)
--	g26607 = NOT(g25382)
--	g17499 = NOT(g14885)
--	g22989 = NOT(g20453)
--	g23929 = NOT(g19147)
--	g17316 = NOT(I18293)
--	g11344 = NOT(g9015)
--	g34208 = NOT(g33838)
--	I14158 = NOT(g8806)
--	g19410 = NOT(g16449)
--	g24825 = NOT(g23204)
--	g22722 = NOT(I22031)
--	g17498 = NOT(g14688)
--	g22988 = NOT(g20391)
--	g8183 = NOT(g482)
--	g23020 = NOT(g19869)
--	I15682 = NOT(g12182)
--	g23928 = NOT(g21562)
--	g8608 = NOT(g278)
--	I18885 = NOT(g16643)
--	g30021 = NOT(g28994)
--	I32071 = NOT(g33665)
--	g19479 = NOT(g16449)
--	g19666 = NOT(g17188)
--	g6782 = NOT(I11632)
--	g25264 = NOT(g23828)
--	g16692 = NOT(g14170)
--	g25790 = NOT(g25027)
--	I29013 = NOT(g29705)
--	g25137 = NOT(g22432)
--	g9340 = NOT(I13094)
--	I13715 = NOT(g71)
--	g17056 = NOT(g13437)
--	I29214 = NOT(g30300)
--	g11291 = NOT(g7526)
--	I32591 = NOT(g34287)
--	g24172 = NOT(I23360)
--	g23046 = NOT(g20283)
--	g32962 = NOT(g30735)
--	g9478 = NOT(I13152)
--	I14823 = NOT(g8056)
--	g19478 = NOT(g16000)
--	g24996 = NOT(g22763)
--	g17611 = NOT(g14822)
--	g17722 = NOT(I18709)
--	g9907 = NOT(g1959)
--	g13173 = NOT(g10632)
--	g34913 = NOT(I33131)
--	g10582 = NOT(g7116)
--	I16755 = NOT(g12377)
--	I29207 = NOT(g30293)
--	g14582 = NOT(I16698)
--	g33874 = NOT(I31724)
--	g9959 = NOT(g6177)
--	g7674 = NOT(I12151)
--	g8977 = NOT(g4349)
--	g24367 = NOT(g22550)
--	g24394 = NOT(g22228)
--	I16770 = NOT(g6023)
--	g32500 = NOT(g30735)
--	g34436 = NOT(I32479)
--	g9517 = NOT(g6163)
--	g9690 = NOT(g732)
--	g17432 = NOT(I18379)
--	g23787 = NOT(g18997)
--	I27677 = NOT(g28156)
--	g29170 = NOT(g27907)
--	g32833 = NOT(g30825)
--	g18957 = NOT(I19734)
--	g21282 = NOT(I21019)
--	g16214 = NOT(g13437)
--	g17271 = NOT(I18270)
--	I32950 = NOT(g34713)
--	g23282 = NOT(g20330)
--	I26710 = NOT(g27511)
--	g7541 = NOT(g344)
--	g10627 = NOT(I13968)
--	I25105 = NOT(g25284)
--	g34320 = NOT(g34119)
--	g27089 = NOT(g26703)
--	g10379 = NOT(g6953)
--	g23302 = NOT(g20330)
--	I25743 = NOT(g25903)
--	g31665 = NOT(I29245)
--	g25209 = NOT(g22763)
--	g19580 = NOT(g16164)
--	g30593 = NOT(g29970)
--	g33665 = NOT(I31500)
--	g6998 = NOT(g4932)
--	g22199 = NOT(g19210)
--	g34530 = NOT(I32591)
--	g10112 = NOT(g1988)
--	g34593 = NOT(I32687)
--	g7132 = NOT(g4558)
--	g12546 = NOT(g8740)
--	I22470 = NOT(g21326)
--	g10050 = NOT(g6336)
--	g27088 = NOT(g26694)
--	g18562 = NOT(I19384)
--	g34346 = NOT(g34162)
--	g10378 = NOT(g6926)
--	g25208 = NOT(g22763)
--	g30565 = NOT(I28832)
--	g7153 = NOT(g5373)
--	g7680 = NOT(g4108)
--	g8451 = NOT(g4057)
--	g22198 = NOT(g19147)
--	g22529 = NOT(g19549)
--	g34122 = NOT(I32059)
--	g15799 = NOT(g13110)
--	I21831 = NOT(g19127)
--	g13506 = NOT(g10808)
--	g12088 = NOT(g7701)
--	g13028 = NOT(I15650)
--	g20446 = NOT(g15224)
--	g10386 = NOT(g6982)
--	g29194 = NOT(I27492)
--	g9915 = NOT(g2583)
--	g12860 = NOT(g10368)
--	g22528 = NOT(g19801)
--	g6850 = NOT(g2704)
--	g14386 = NOT(I16544)
--	g23769 = NOT(g19074)
--	I11980 = NOT(g66)
--	g22330 = NOT(g19801)
--	I13889 = NOT(g7598)
--	g25542 = NOT(g22763)
--	g7802 = NOT(g324)
--	g20059 = NOT(g17302)
--	g32613 = NOT(g30673)
--	g8146 = NOT(g1760)
--	g10096 = NOT(g5767)
--	g20025 = NOT(g17271)
--	g8346 = NOT(g3845)
--	g24059 = NOT(g21193)
--	g33454 = NOT(I30980)
--	g14096 = NOT(I16328)
--	g24025 = NOT(g21256)
--	g9214 = NOT(g617)
--	g17529 = NOT(g15039)
--	g20540 = NOT(g16646)
--	g12497 = NOT(g9780)
--	g30292 = NOT(g28736)
--	I16898 = NOT(g10615)
--	g23768 = NOT(g18997)
--	I12884 = NOT(g4213)
--	I22467 = NOT(g19662)
--	g20058 = NOT(g16782)
--	g24540 = NOT(g22942)
--	g33712 = NOT(I31561)
--	I26356 = NOT(g26843)
--	I18307 = NOT(g12977)
--	g32947 = NOT(g31376)
--	g19531 = NOT(g16816)
--	g24058 = NOT(g20982)
--	g22869 = NOT(g20875)
--	g17528 = NOT(g14940)
--	g7558 = NOT(I12041)
--	g32605 = NOT(g30614)
--	g8696 = NOT(g3347)
--	g34409 = NOT(g34145)
--	I21722 = NOT(g19264)
--	g22868 = NOT(g20453)
--	I16521 = NOT(g10430)
--	g17764 = NOT(I18758)
--	I12666 = NOT(g4040)
--	g10429 = NOT(g7148)
--	g11927 = NOT(g10207)
--	g23881 = NOT(g19277)
--	g10857 = NOT(g8712)
--	g32812 = NOT(g30825)
--	g25073 = NOT(I24237)
--	g32463 = NOT(g31566)
--	g16100 = NOT(I17471)
--	I32446 = NOT(g34127)
--	g19676 = NOT(g17062)
--	g19685 = NOT(g16987)
--	g31239 = NOT(g29916)
--	g25274 = NOT(g22763)
--	g24044 = NOT(g21127)
--	g16771 = NOT(g14018)
--	g34408 = NOT(g34144)
--	I22419 = NOT(g19638)
--	g19373 = NOT(g16449)
--	g26575 = NOT(g25268)
--	g10428 = NOT(g9631)
--	g32951 = NOT(g31021)
--	g32972 = NOT(g31710)
--	g16235 = NOT(g13437)
--	g32033 = NOT(g30929)
--	I32059 = NOT(g33648)
--	g8508 = NOT(g3827)
--	g19654 = NOT(g16931)
--	I31361 = NOT(g33120)
--	g9402 = NOT(g6209)
--	g9824 = NOT(g1825)
--	g8944 = NOT(g370)
--	g8240 = NOT(g1333)
--	g18661 = NOT(I19487)
--	g20902 = NOT(I20870)
--	g18895 = NOT(g16000)
--	g19800 = NOT(g17096)
--	I18341 = NOT(g14308)
--	g19417 = NOT(g17178)
--	g21662 = NOT(g16540)
--	g24377 = NOT(g22594)
--	g7092 = NOT(g6483)
--	I31500 = NOT(g33176)
--	g24120 = NOT(g19984)
--	g23027 = NOT(g20391)
--	g32795 = NOT(g31327)
--	g25034 = NOT(g23695)
--	I23342 = NOT(g23299)
--	g17709 = NOT(g14761)
--	g33382 = NOT(g32033)
--	I12580 = NOT(g1239)
--	g8443 = NOT(g3736)
--	g19334 = NOT(I19818)
--	g20146 = NOT(g17533)
--	g20738 = NOT(g15483)
--	I18180 = NOT(g13605)
--	g25641 = NOT(I24784)
--	g20562 = NOT(g17955)
--	g9590 = NOT(g1882)
--	g21249 = NOT(g15509)
--	I15981 = NOT(g11290)
--	g24146 = NOT(g19422)
--	g6986 = NOT(g4743)
--	g23249 = NOT(g21070)
--	I14687 = NOT(g7753)
--	g11770 = NOT(I14619)
--	I21199 = NOT(g17501)
--	I30998 = NOT(g32453)
--	g20699 = NOT(g17873)
--	g16515 = NOT(g13486)
--	g10504 = NOT(g8763)
--	g11981 = NOT(I14823)
--	g9657 = NOT(g2763)
--	g12968 = NOT(g11793)
--	g17471 = NOT(g14454)
--	g25153 = NOT(g23733)
--	I26448 = NOT(g26860)
--	g8316 = NOT(g2351)
--	g17087 = NOT(g14321)
--	g23482 = NOT(g18833)
--	I25552 = NOT(g25240)
--	g32514 = NOT(g30735)
--	I18734 = NOT(g6373)
--	g24699 = NOT(g23047)
--	g21248 = NOT(g15224)
--	g14504 = NOT(g12361)
--	g19762 = NOT(g16326)
--	g23248 = NOT(g20924)
--	g19964 = NOT(g17200)
--	I22589 = NOT(g21340)
--	g20698 = NOT(g17873)
--	g27527 = NOT(I26195)
--	g25409 = NOT(g22228)
--	g34575 = NOT(I32651)
--	I25779 = NOT(g26424)
--	g32507 = NOT(g30735)
--	g9556 = NOT(g5448)
--	I18839 = NOT(g13716)
--	g23003 = NOT(I22180)
--	g8565 = NOT(g3802)
--	g21204 = NOT(g15656)
--	g33637 = NOT(I31466)
--	g29177 = NOT(g27937)
--	g30327 = NOT(I28582)
--	g33935 = NOT(I31817)
--	g34711 = NOT(g34559)
--	g12870 = NOT(g10374)
--	I11860 = NOT(g43)
--	g25136 = NOT(g22457)
--	g34327 = NOT(g34108)
--	I18667 = NOT(g6661)
--	I18694 = NOT(g5666)
--	g32421 = NOT(g31213)
--	I23330 = NOT(g22658)
--	I23393 = NOT(g23414)
--	g10129 = NOT(g5352)
--	I29441 = NOT(g30917)
--	g11845 = NOT(I14663)
--	g9064 = NOT(g4983)
--	I18131 = NOT(g13350)
--	g8681 = NOT(g763)
--	g10002 = NOT(g6195)
--	I25786 = NOT(g26424)
--	g10057 = NOT(g6455)
--	g9899 = NOT(g6513)
--	I32645 = NOT(g34367)
--	g7262 = NOT(g5723)
--	g24366 = NOT(g22594)
--	g20632 = NOT(g15171)
--	I15633 = NOT(g12074)
--	I32699 = NOT(g34569)
--	I33273 = NOT(g34984)
--	g30606 = NOT(I28866)
--	g8697 = NOT(g3694)
--	I33106 = NOT(g34855)
--	I14668 = NOT(g7753)
--	I25356 = NOT(g24374)
--	g19543 = NOT(g16349)
--	g30303 = NOT(g28786)
--	g8914 = NOT(g4264)
--	I19796 = NOT(g17870)
--	g17602 = NOT(g14962)
--	g12867 = NOT(g10375)
--	g12894 = NOT(g10401)
--	I17401 = NOT(g13394)
--	g16584 = NOT(g13920)
--	g17774 = NOT(g14902)
--	g23647 = NOT(g18833)
--	g18889 = NOT(g15509)
--	g17955 = NOT(I18865)
--	g18980 = NOT(g16136)
--	g32541 = NOT(g30673)
--	g7623 = NOT(I12103)
--	g10323 = NOT(I13744)
--	g23945 = NOT(g21611)
--	g16206 = NOT(g13437)
--	I25380 = NOT(g24481)
--	g18095 = NOT(I18891)
--	g23356 = NOT(g21070)
--	g32473 = NOT(g31070)
--	I31463 = NOT(g33318)
--	g19908 = NOT(g16540)
--	g22171 = NOT(g18882)
--	g13191 = NOT(I15788)
--	g26840 = NOT(I25562)
--	g20661 = NOT(g15171)
--	I12654 = NOT(g1585)
--	g21380 = NOT(g17955)
--	g10533 = NOT(g8795)
--	g20547 = NOT(g15224)
--	g23999 = NOT(g21468)
--	g32789 = NOT(g30735)
--	g18888 = NOT(g15426)
--	g23380 = NOT(g20619)
--	g33729 = NOT(I31586)
--	I18443 = NOT(g13027)
--	g19569 = NOT(g16349)
--	I14424 = NOT(g4005)
--	I14016 = NOT(g9104)
--	I17118 = NOT(g14363)
--	g16725 = NOT(g13963)
--	I22748 = NOT(g19458)
--	g13521 = NOT(g11357)
--	g22994 = NOT(g20436)
--	g34982 = NOT(I33246)
--	g32788 = NOT(g31327)
--	g32724 = NOT(g30735)
--	g19747 = NOT(g17015)
--	g23233 = NOT(g21037)
--	g21182 = NOT(g15509)
--	g6789 = NOT(I11635)
--	g11832 = NOT(g8011)
--	g23182 = NOT(g21389)
--	g20715 = NOT(g15277)
--	g23651 = NOT(g20655)
--	g32829 = NOT(g30937)
--	g28080 = NOT(I26581)
--	g32920 = NOT(g30825)
--	I18469 = NOT(g13809)
--	g32535 = NOT(g31554)
--	g25327 = NOT(g22161)
--	g32434 = NOT(g31189)
--	I14830 = NOT(g10141)
--	I21258 = NOT(g16540)
--	g24481 = NOT(I23684)
--	I14893 = NOT(g9819)
--	g25109 = NOT(g23666)
--	g12818 = NOT(g8792)
--	g20551 = NOT(g17302)
--	g20572 = NOT(g15833)
--	g9194 = NOT(g827)
--	g32828 = NOT(g31710)
--	g18931 = NOT(g16031)
--	g6987 = NOT(g4754)
--	g32946 = NOT(g31327)
--	g10232 = NOT(g4527)
--	I17276 = NOT(g13605)
--	g7285 = NOT(g4643)
--	g11861 = NOT(g8070)
--	g22919 = NOT(g21163)
--	g16744 = NOT(I17964)
--	I17704 = NOT(g13144)
--	g12978 = NOT(I15593)
--	g14232 = NOT(g11083)
--	g9731 = NOT(g5366)
--	g23331 = NOT(g20905)
--	I13968 = NOT(g7697)
--	I32547 = NOT(g34397)
--	g19751 = NOT(g16044)
--	I24839 = NOT(g24298)
--	g9489 = NOT(g2303)
--	g19772 = NOT(g17183)
--	g25283 = NOT(g22763)
--	g34840 = NOT(I33056)
--	g20127 = NOT(I20388)
--	I22177 = NOT(g21366)
--	g23449 = NOT(g18833)
--	g26483 = NOT(I25359)
--	g28753 = NOT(I27235)
--	g9557 = NOT(g5499)
--	g13926 = NOT(I16217)
--	g24127 = NOT(g19984)
--	g13045 = NOT(g11941)
--	g10261 = NOT(g4555)
--	I17808 = NOT(g13311)
--	g9071 = NOT(g2831)
--	g26862 = NOT(I25598)
--	g11388 = NOT(I14395)
--	g23897 = NOT(g19210)
--	g13099 = NOT(I15732)
--	g11324 = NOT(g7542)
--	g23448 = NOT(g21611)
--	g23961 = NOT(g19074)
--	g32682 = NOT(g30825)
--	g24490 = NOT(g22594)
--	I14705 = NOT(g7717)
--	g19638 = NOT(g17324)
--	I17101 = NOT(g14338)
--	g34192 = NOT(g33921)
--	I21810 = NOT(g20596)
--	I16629 = NOT(g11987)
--	g16652 = NOT(g13892)
--	g17010 = NOT(I18138)
--	g23505 = NOT(g21514)
--	I27543 = NOT(g28187)
--	g26326 = NOT(g24872)
--	g8922 = NOT(I12907)
--	g20385 = NOT(g18008)
--	I14679 = NOT(g9332)
--	g13251 = NOT(I15814)
--	I23375 = NOT(g23403)
--	g13272 = NOT(I15837)
--	g19416 = NOT(g15885)
--	g20103 = NOT(g17433)
--	g7424 = NOT(g2465)
--	g24376 = NOT(g22722)
--	g24385 = NOT(g22908)
--	g34522 = NOT(g34271)
--	g7809 = NOT(g4864)
--	I18143 = NOT(g13350)
--	g24103 = NOT(g21209)
--	g23026 = NOT(g20391)
--	g18088 = NOT(g13267)
--	g24980 = NOT(g22384)
--	I16246 = NOT(g3983)
--	I30971 = NOT(g32015)
--	I12117 = NOT(g586)
--	g24095 = NOT(g21209)
--	g26702 = NOT(g25309)
--	g17599 = NOT(g14794)
--	I12000 = NOT(g582)
--	g25174 = NOT(g23890)
--	g28696 = NOT(g27858)
--	g31653 = NOT(g29713)
--	g6991 = NOT(g4888)
--	g33653 = NOT(I31486)
--	I14939 = NOT(g10216)
--	g7231 = NOT(g5)
--	g20671 = NOT(g15509)
--	I17733 = NOT(g14844)
--	g27018 = NOT(I25750)
--	g31138 = NOT(g29778)
--	g32760 = NOT(g30735)
--	g17086 = NOT(g14297)
--	g24181 = NOT(I23387)
--	g7523 = NOT(g305)
--	g19579 = NOT(g16000)
--	g22159 = NOT(I21744)
--	g29941 = NOT(g28900)
--	g13140 = NOT(g10632)
--	g7643 = NOT(g4322)
--	I21792 = NOT(g21308)
--	I12568 = NOT(g5005)
--	g12018 = NOT(g9538)
--	I22009 = NOT(g21269)
--	g34553 = NOT(I32621)
--	g10499 = NOT(I13872)
--	I22665 = NOT(g21308)
--	I13581 = NOT(g6727)
--	I18168 = NOT(g13191)
--	I24278 = NOT(g23440)
--	I14267 = NOT(g7835)
--	g32506 = NOT(g31376)
--	g8784 = NOT(I12764)
--	I31724 = NOT(g33076)
--	g33636 = NOT(I31463)
--	g29185 = NOT(I27481)
--	I32956 = NOT(g34654)
--	g30326 = NOT(I28579)
--	g21723 = NOT(I21288)
--	g29092 = NOT(g27800)
--	I32297 = NOT(g34059)
--	g34949 = NOT(g34939)
--	g10498 = NOT(g7161)
--	I32103 = NOT(g33661)
--	g34326 = NOT(g34091)
--	g13061 = NOT(g10981)
--	I31829 = NOT(g33454)
--	I18479 = NOT(g13041)
--	g31852 = NOT(g29385)
--	g6959 = NOT(g4420)
--	I31535 = NOT(g33377)
--	g30040 = NOT(g29025)
--	I13202 = NOT(g5105)
--	g19586 = NOT(g16349)
--	I12123 = NOT(g758)
--	g17125 = NOT(I18177)
--	g17532 = NOT(I18479)
--	g27402 = NOT(I26100)
--	g34536 = NOT(I32601)
--	I17166 = NOT(g14536)
--	g28161 = NOT(I26676)
--	g7634 = NOT(I12123)
--	g15758 = NOT(I17276)
--	g21387 = NOT(I21115)
--	I22485 = NOT(g21308)
--	I29221 = NOT(g30307)
--	g23433 = NOT(g21562)
--	I28419 = NOT(g29195)
--	I13979 = NOT(g7733)
--	I32824 = NOT(g34475)
--	g24426 = NOT(g22722)
--	g8479 = NOT(g3057)
--	g20190 = NOT(g16971)
--	g22144 = NOT(g18997)
--	I24038 = NOT(g22202)
--	g23620 = NOT(I22769)
--	g28709 = NOT(I27192)
--	g10080 = NOT(g1982)
--	I17008 = NOT(g12857)
--	I32671 = NOT(g34388)
--	g8840 = NOT(g4277)
--	g9212 = NOT(g6466)
--	g12866 = NOT(g10369)
--	I21918 = NOT(g21290)
--	I17892 = NOT(g3325)
--	g21343 = NOT(g16428)
--	I26925 = NOT(g27015)
--	g8390 = NOT(g3385)
--	g32927 = NOT(g30825)
--	g15345 = NOT(I17108)
--	g14432 = NOT(g12311)
--	g17680 = NOT(g14889)
--	g17144 = NOT(g14085)
--	g26634 = NOT(g25317)
--	g26851 = NOT(I25579)
--	g11447 = NOT(I14450)
--	g7926 = NOT(g3423)
--	I15162 = NOT(g10176)
--	g20546 = NOT(g18008)
--	g20089 = NOT(g17533)
--	g23971 = NOT(g20751)
--	I26378 = NOT(g26850)
--	g19720 = NOT(I20130)
--	g20211 = NOT(g16931)
--	I25369 = NOT(g24891)
--	g24089 = NOT(g19890)
--	I19851 = NOT(g16615)
--	g27597 = NOT(g26745)
--	g21369 = NOT(g16285)
--	I33291 = NOT(g34983)
--	g12077 = NOT(I14939)
--	g32649 = NOT(g30673)
--	g25553 = NOT(g22550)
--	g20088 = NOT(g17533)
--	I27391 = NOT(g27929)
--	g8356 = NOT(g54)
--	I20937 = NOT(g16967)
--	g9229 = NOT(g5052)
--	I13094 = NOT(g2724)
--	g14753 = NOT(g11317)
--	I33173 = NOT(g34887)
--	g24088 = NOT(g21209)
--	g19493 = NOT(g16349)
--	g24024 = NOT(g21193)
--	g14342 = NOT(g12163)
--	g34673 = NOT(I32803)
--	g34847 = NOT(I33067)
--	g31609 = NOT(I29211)
--	g29215 = NOT(I27561)
--	g10031 = NOT(I13552)
--	g32648 = NOT(g30614)
--	g32491 = NOT(g31566)
--	g32903 = NOT(g31376)
--	g25326 = NOT(g22228)
--	g14031 = NOT(I16289)
--	g9822 = NOT(g125)
--	g10199 = NOT(g1968)
--	I11801 = NOT(g6395)
--	I14455 = NOT(g10197)
--	g16605 = NOT(g13955)
--	g11472 = NOT(g7918)
--	I27579 = NOT(g28184)
--	I29371 = NOT(g30325)
--	g12923 = NOT(I15542)
--	g31608 = NOT(g29653)
--	g18527 = NOT(I19345)
--	g20497 = NOT(g18065)
--	g32604 = NOT(g31154)
--	g34062 = NOT(g33711)
--	I28588 = NOT(g29368)
--	g32755 = NOT(g31672)
--	I30959 = NOT(g32021)
--	g10198 = NOT(I13672)
--	g12300 = NOT(I15144)
--	g11911 = NOT(g10022)
--	g16812 = NOT(g13555)
--	g21412 = NOT(g15758)
--	g32770 = NOT(g31710)
--	g34933 = NOT(g34916)
--	g14198 = NOT(g12180)
--	g32563 = NOT(g31554)
--	I32089 = NOT(g33665)
--	I33134 = NOT(g34906)
--	g13246 = NOT(g10939)
--	g20700 = NOT(g17873)
--	g20659 = NOT(g17873)
--	g34851 = NOT(I33075)
--	g20625 = NOT(g15348)
--	g10393 = NOT(g6991)
--	g24126 = NOT(g19935)
--	g24625 = NOT(g23135)
--	g14330 = NOT(I16486)
--	g24987 = NOT(g23630)
--	g8954 = NOT(g1079)
--	g7543 = NOT(I12033)
--	g31799 = NOT(g29385)
--	g23896 = NOT(g19210)
--	g25564 = NOT(g22312)
--	g8363 = NOT(g239)
--	g18894 = NOT(g16000)
--	g31813 = NOT(g29385)
--	g21228 = NOT(g17531)
--	g33799 = NOT(g33299)
--	g10365 = NOT(g6867)
--	g22224 = NOT(g19277)
--	g33813 = NOT(I31659)
--	g8032 = NOT(I12355)
--	g19517 = NOT(g16777)
--	g23228 = NOT(g21070)
--	I18373 = NOT(g13011)
--	g29906 = NOT(g28793)
--	g29348 = NOT(g28194)
--	g16795 = NOT(I18009)
--	g10960 = NOT(g9007)
--	I17675 = NOT(g13394)
--	g23011 = NOT(g20330)
--	g31798 = NOT(g29385)
--	g32767 = NOT(g30735)
--	g32794 = NOT(g30937)
--	I14623 = NOT(g8925)
--	g11147 = NOT(g8417)
--	g11754 = NOT(g8229)
--	I17154 = NOT(g13605)
--	I23680 = NOT(g23219)
--	g25183 = NOT(g22763)
--	g32899 = NOT(g31021)
--	g7534 = NOT(g1367)
--	g31805 = NOT(g29385)
--	g17224 = NOT(I18248)
--	g16514 = NOT(g14139)
--	g12885 = NOT(g10382)
--	g22495 = NOT(g19801)
--	g17308 = NOT(g14876)
--	g23582 = NOT(I22729)
--	g32633 = NOT(g31154)
--	g32898 = NOT(g30825)
--	I32659 = NOT(g34391)
--	g15048 = NOT(I16969)
--	g9620 = NOT(g6187)
--	g9462 = NOT(g6215)
--	I23336 = NOT(g22721)
--	I19756 = NOT(g17812)
--	g19362 = NOT(g16072)
--	g7927 = NOT(g4064)
--	g34574 = NOT(I32648)
--	g32719 = NOT(g31672)
--	I12041 = NOT(g2741)
--	g20060 = NOT(g16540)
--	g34047 = NOT(g33637)
--	g18979 = NOT(g16136)
--	g19523 = NOT(g16100)
--	g24060 = NOT(g21256)
--	g8912 = NOT(g4180)
--	I16120 = NOT(g11868)
--	g33934 = NOT(I31814)
--	g10708 = NOT(g7836)
--	g20197 = NOT(g16987)
--	g6928 = NOT(I11716)
--	I12746 = NOT(g4087)
--	g21379 = NOT(g17873)
--	g34311 = NOT(g34097)
--	I12493 = NOT(g5002)
--	g22976 = NOT(I22149)
--	g22985 = NOT(g20330)
--	g32718 = NOT(g30825)
--	g32521 = NOT(g31376)
--	g10087 = NOT(I13597)
--	g23925 = NOT(g21514)
--	g8357 = NOT(I12538)
--	g18978 = NOT(g16000)
--	g7946 = NOT(I12314)
--	g7660 = NOT(I12144)
--	g29653 = NOT(I27927)
--	I22729 = NOT(g21308)
--	g26820 = NOT(I25534)
--	g21050 = NOT(g17873)
--	g20527 = NOT(g18008)
--	I13597 = NOT(g4417)
--	g11367 = NOT(I14381)
--	g28918 = NOT(g27832)
--	g32832 = NOT(g30735)
--	I20321 = NOT(g16920)
--	g23378 = NOT(g21070)
--	g13394 = NOT(I15915)
--	I31491 = NOT(g33283)
--	g33761 = NOT(I31616)
--	g24527 = NOT(g22670)
--	g7903 = NOT(g969)
--	g30072 = NOT(I28301)
--	g17687 = NOT(g15042)
--	I31604 = NOT(g33176)
--	g28079 = NOT(I26578)
--	g10043 = NOT(g1632)
--	I13280 = NOT(g6140)
--	g7513 = NOT(g6315)
--	g26731 = NOT(g25470)
--	g34592 = NOT(I32684)
--	I11688 = NOT(g70)
--	I16698 = NOT(g12077)
--	g29333 = NOT(g28167)
--	g16473 = NOT(g13977)
--	I31770 = NOT(g33197)
--	g32861 = NOT(g31376)
--	g9842 = NOT(g3274)
--	g23944 = NOT(g19147)
--	g32573 = NOT(g30825)
--	g18094 = NOT(I18888)
--	g31013 = NOT(g29679)
--	I14589 = NOT(g8818)
--	g25213 = NOT(g23293)
--	g19437 = NOT(g16349)
--	g20503 = NOT(g15373)
--	g9298 = NOT(g5080)
--	g28598 = NOT(g27717)
--	I18909 = NOT(g16873)
--	g9392 = NOT(g5869)
--	g32926 = NOT(g31376)
--	I32855 = NOT(g34540)
--	g7178 = NOT(g4392)
--	g7436 = NOT(g5276)
--	I14836 = NOT(g9688)
--	g8626 = NOT(g4040)
--	g21681 = NOT(I21242)
--	g29963 = NOT(g28931)
--	g16724 = NOT(g14079)
--	g22842 = NOT(g19875)
--	g23681 = NOT(g21012)
--	I18117 = NOT(g13302)
--	g32612 = NOT(g30614)
--	g16325 = NOT(g13223)
--	g18877 = NOT(g15224)
--	I23309 = NOT(g21677)
--	g25452 = NOT(g22228)
--	g15371 = NOT(I17114)
--	g25047 = NOT(g23733)
--	g32099 = NOT(g31009)
--	g10375 = NOT(g6941)
--	I21288 = NOT(g18216)
--	g34820 = NOT(I33034)
--	g16920 = NOT(I18086)
--	g20714 = NOT(g15277)
--	g20450 = NOT(g15277)
--	g23429 = NOT(g20453)
--	g32701 = NOT(g31376)
--	g12076 = NOT(g9280)
--	g7335 = NOT(g2287)
--	g7831 = NOT(I12227)
--	I14119 = NOT(g7824)
--	g32777 = NOT(g31710)
--	g32534 = NOT(g30673)
--	g12721 = NOT(g10061)
--	g34152 = NOT(I32109)
--	g20707 = NOT(g18008)
--	g21428 = NOT(g15758)
--	I22622 = NOT(g21209)
--	g20910 = NOT(g15171)
--	g34846 = NOT(I33064)
--	g23793 = NOT(g19074)
--	g12054 = NOT(g7690)
--	g17392 = NOT(g14924)
--	g19600 = NOT(g16164)
--	g10337 = NOT(g5016)
--	g24819 = NOT(I23998)
--	g19781 = NOT(g16489)
--	g17489 = NOT(g12955)
--	I24334 = NOT(g22976)
--	g20496 = NOT(g17929)
--	g7805 = NOT(g4366)
--	g7916 = NOT(I12300)
--	g25051 = NOT(I24215)
--	g25072 = NOT(g23630)
--	g24818 = NOT(g23191)
--	g32462 = NOT(g30673)
--	I14749 = NOT(g10031)
--	g24979 = NOT(g22369)
--	g21690 = NOT(g16540)
--	g22830 = NOT(g20283)
--	g19952 = NOT(g15915)
--	g24055 = NOT(g19968)
--	g7749 = NOT(g996)
--	g19351 = NOT(g17367)
--	I12523 = NOT(g3794)
--	g23549 = NOT(g18833)
--	g27773 = NOT(I26378)
--	g20070 = NOT(g16173)
--	g20978 = NOT(g15595)
--	g24111 = NOT(g19890)
--	g28656 = NOT(g27742)
--	g9708 = NOT(g2741)
--	g24070 = NOT(g20014)
--	g24978 = NOT(g22342)
--	g34691 = NOT(I32843)
--	g29312 = NOT(g28877)
--	g20590 = NOT(g15426)
--	g22544 = NOT(g19589)
--	g22865 = NOT(g20330)
--	g23548 = NOT(g18833)
--	g8778 = NOT(I12758)
--	g29115 = NOT(g27779)
--	g7947 = NOT(g1500)
--	I20216 = NOT(g15862)
--	g24986 = NOT(g23590)
--	I14305 = NOT(g8805)
--	g9252 = NOT(g4304)
--	I26880 = NOT(g27527)
--	g23504 = NOT(g21468)
--	g13902 = NOT(g11389)
--	g13301 = NOT(g10862)
--	g31771 = NOT(I29337)
--	g19264 = NOT(I19802)
--	g18917 = NOT(g16077)
--	g19790 = NOT(g16971)
--	g20384 = NOT(g18008)
--	g12180 = NOT(g9477)
--	g9958 = NOT(g6148)
--	g29921 = NOT(g28864)
--	g13120 = NOT(g10632)
--	I18293 = NOT(g1079)
--	g24384 = NOT(g22885)
--	g25820 = NOT(g25051)
--	I26512 = NOT(g26817)
--	I17653 = NOT(g14276)
--	g20067 = NOT(g17328)
--	g32766 = NOT(g31376)
--	g6955 = NOT(I11726)
--	g29745 = NOT(g28500)
--	g24067 = NOT(g21256)
--	g24094 = NOT(g21143)
--	g11562 = NOT(g7648)
--	g17713 = NOT(g12947)
--	I18265 = NOT(g13350)
--	g34929 = NOT(I33179)
--	g27930 = NOT(I26451)
--	I12437 = NOT(g4999)
--	g27993 = NOT(I26503)
--	g8075 = NOT(g3742)
--	g32871 = NOT(g30937)
--	g30020 = NOT(g29097)
--	g30928 = NOT(I28908)
--	g22189 = NOT(I21769)
--	g8475 = NOT(I12608)
--	g26105 = NOT(I25146)
--	g9829 = NOT(g2250)
--	g12839 = NOT(g10350)
--	g6814 = NOT(g632)
--	g12930 = NOT(g12347)
--	g7873 = NOT(g1266)
--	g26743 = NOT(g25476)
--	g26827 = NOT(g24819)
--	g34583 = NOT(I32665)
--	g7632 = NOT(I12117)
--	g34928 = NOT(I33176)
--	g7095 = NOT(g6545)
--	I17636 = NOT(g14252)
--	g21057 = NOT(g15426)
--	g23002 = NOT(I22177)
--	g10079 = NOT(g1950)
--	g11290 = NOT(I14326)
--	g24150 = NOT(g19268)
--	g23057 = NOT(g20453)
--	I28594 = NOT(g29379)
--	g9911 = NOT(g2384)
--	g7495 = NOT(g4375)
--	g14545 = NOT(g12768)
--	g7437 = NOT(g5666)
--	g17610 = NOT(g15008)
--	I27253 = NOT(g27996)
--	I30995 = NOT(g32449)
--	g12838 = NOT(g10353)
--	g23128 = NOT(g20283)
--	I20569 = NOT(g16486)
--	I17852 = NOT(g3625)
--	g10078 = NOT(g1854)
--	g21245 = NOT(I20982)
--	g24019 = NOT(g19968)
--	g17189 = NOT(g14708)
--	g23245 = NOT(g20785)
--	I13287 = NOT(g110)
--	g26769 = NOT(g25400)
--	g8526 = NOT(g1526)
--	g19208 = NOT(g17367)
--	g20695 = NOT(I20781)
--	I20747 = NOT(g17141)
--	I31701 = NOT(g33164)
--	g21299 = NOT(g16600)
--	g30113 = NOT(g29154)
--	g9733 = NOT(g5736)
--	g10086 = NOT(g2193)
--	g23323 = NOT(g20283)
--	g23299 = NOT(I22400)
--	g9974 = NOT(g2518)
--	I32067 = NOT(g33661)
--	g17188 = NOT(I18224)
--	I11721 = NOT(g4145)
--	g17124 = NOT(g14051)
--	g17678 = NOT(I18653)
--	g34787 = NOT(I32991)
--	g26803 = NOT(g25389)
--	g12487 = NOT(g9340)
--	g20526 = NOT(g15171)
--	I22576 = NOT(g21282)
--	I28185 = NOT(g28803)
--	I18835 = NOT(g6365)
--	I13054 = NOT(g6744)
--	g24526 = NOT(g22942)
--	g19542 = NOT(g16349)
--	g30302 = NOT(g28924)
--	g7752 = NOT(g1542)
--	I16181 = NOT(g3672)
--	g18102 = NOT(I18912)
--	g8439 = NOT(g3129)
--	g9073 = NOT(g150)
--	g32629 = NOT(g31376)
--	g34302 = NOT(I32305)
--	I26989 = NOT(g27277)
--	I32150 = NOT(g33923)
--	g30105 = NOT(I28336)
--	g6836 = NOT(g1322)
--	g7917 = NOT(g1157)
--	I14630 = NOT(g7717)
--	g27279 = NOT(g26330)
--	g32472 = NOT(g30825)
--	g10159 = NOT(g4477)
--	g34827 = NOT(I33041)
--	g10532 = NOT(g10233)
--	g32628 = NOT(g31542)
--	g17093 = NOT(I18165)
--	g6918 = NOT(g3639)
--	g32911 = NOT(g31376)
--	g14125 = NOT(I16345)
--	g15344 = NOT(g14851)
--	g10158 = NOT(g2461)
--	g11403 = NOT(g7595)
--	g11547 = NOT(I14505)
--	g13895 = NOT(I16193)
--	g20917 = NOT(g15224)
--	I33140 = NOT(g34884)
--	I28883 = NOT(g30105)
--	g23232 = NOT(I22331)
--	g24866 = NOT(I24038)
--	g19905 = NOT(g15885)
--	I12790 = NOT(g4340)
--	I17609 = NOT(g13510)
--	g34769 = NOT(I32953)
--	I11655 = NOT(g1246)
--	g18876 = NOT(g15373)
--	g18885 = NOT(g15979)
--	g10353 = NOT(g6803)
--	g25046 = NOT(g23729)
--	g6993 = NOT(g4859)
--	g10295 = NOT(I13723)
--	g8919 = NOT(I12896)
--	g21697 = NOT(I21258)
--	g29013 = NOT(I27368)
--	I29981 = NOT(g31591)
--	g34768 = NOT(I32950)
--	g12039 = NOT(I14899)
--	g13715 = NOT(g10573)
--	I22745 = NOT(g19458)
--	g29214 = NOT(I27558)
--	g27038 = NOT(g25932)
--	g9206 = NOT(g5164)
--	g32591 = NOT(g30614)
--	I15572 = NOT(g10499)
--	g23995 = NOT(g19277)
--	g32776 = NOT(g31672)
--	g32785 = NOT(g31710)
--	I30989 = NOT(g32441)
--	g19565 = NOT(g16000)
--	g24077 = NOT(g20720)
--	g20706 = NOT(g18008)
--	I11734 = NOT(g4473)
--	g23880 = NOT(g19210)
--	g12038 = NOT(I14896)
--	g20597 = NOT(g17847)
--	I21042 = NOT(g15824)
--	g32754 = NOT(g30825)
--	I14570 = NOT(g7932)
--	g33435 = NOT(I30959)
--	g25282 = NOT(g22763)
--	I21189 = NOT(g17475)
--	g14336 = NOT(I16498)
--	g27187 = NOT(I25882)
--	g7296 = NOT(g5313)
--	g23512 = NOT(g20248)
--	g8616 = NOT(g2803)
--	g28752 = NOT(I27232)
--	g20923 = NOT(g15277)
--	g27975 = NOT(g26694)
--	g32859 = NOT(g30614)
--	g32825 = NOT(g30735)
--	g32950 = NOT(g31672)
--	g28954 = NOT(g27830)
--	g26710 = NOT(g25349)
--	g18660 = NOT(I19484)
--	g20624 = NOT(g18065)
--	g22455 = NOT(g19801)
--	g12975 = NOT(g12752)
--	g7532 = NOT(g1157)
--	I13694 = NOT(g117)
--	I16024 = NOT(g11171)
--	g32858 = NOT(g31327)
--	g33744 = NOT(I31604)
--	g7553 = NOT(g1274)
--	g8404 = NOT(g5005)
--	g15506 = NOT(I17131)
--	g31849 = NOT(g29385)
--	g8647 = NOT(g3416)
--	g14631 = NOT(g12239)
--	g10364 = NOT(g6869)
--	g19409 = NOT(g16431)
--	I14567 = NOT(g9708)
--	g12143 = NOT(I14999)
--	g20102 = NOT(g17533)
--	g16767 = NOT(I17989)
--	g20157 = NOT(g16886)
--	g25640 = NOT(I24781)
--	g12937 = NOT(g12419)
--	g28669 = NOT(g27705)
--	g26081 = NOT(g24619)
--	g8764 = NOT(g4826)
--	g22201 = NOT(g19277)
--	g24102 = NOT(g21143)
--	g23445 = NOT(I22564)
--	g31848 = NOT(g29385)
--	g18916 = NOT(g16053)
--	g24157 = NOT(I23315)
--	g32844 = NOT(g30937)
--	g9898 = NOT(g6444)
--	
--	g33848 = AND(g33261, g20384)
--	g28260 = AND(g27703, g26518)
--	g17617 = AND(g7885, g13326)
--	g18550 = AND(g2819, g15277)
--	g25768 = AND(g2912, g24560)
--	g25803 = AND(g24798, g21024)
--	g31141 = AND(g12224, g30038)
--	I26960 = AND(g24995, g26424, g22698)
--	g22075 = AND(g6247, g19210)
--	g18314 = AND(g1585, g16931)
--	g33652 = AND(g33393, g18889)
--	g18287 = AND(g1442, g16449)
--	g27410 = AND(g26549, g17527)
--	g16633 = AND(g5196, g14921)
--	g30248 = AND(g28743, g23938)
--	g34482 = AND(g34405, g18917)
--	g23498 = AND(g20234, g12998)
--	g28489 = AND(g27010, g12417)
--	g26356 = AND(g15581, g25523)
--	g18307 = AND(g1559, g16931)
--	g29771 = AND(g28322, g23242)
--	g30003 = AND(g28149, g9021)
--	g34710 = AND(g34553, g20903)
--	g16191 = AND(g5475, g14262)
--	g22623 = AND(g19337, g19470)
--	g21989 = AND(g5587, g19074)
--	g30204 = AND(g28670, g23868)
--	g13671 = AND(g4498, g10532)
--	g26826 = AND(g24907, g15747)
--	g27666 = AND(g26865, g23521)
--	I31246 = AND(g31672, g31839, g32810, g32811)
--	g18721 = AND(g15138, g16077)
--	g22037 = AND(g5941, g19147)
--	g25881 = AND(g3821, g24685)
--	g26380 = AND(g19572, g25547)
--	g33263 = AND(g32393, g25481)
--	g18596 = AND(g2941, g16349)
--	g32420 = AND(g31127, g19533)
--	g28488 = AND(g27969, g17713)
--	g27363 = AND(g10231, g26812)
--	g23056 = AND(g16052, g19860)
--	g27217 = AND(g26236, g8418, g2610)
--	g29683 = AND(g1821, g29046)
--	g18243 = AND(g1189, g16431)
--	g33332 = AND(g32217, g20608)
--	I17692 = AND(g14988, g11450, g6756)
--	g21988 = AND(g5583, g19074)
--	g26090 = AND(g1624, g25081)
--	g21924 = AND(g5057, g21468)
--	g28558 = AND(g7301, g27046)
--	g18431 = AND(g2185, g18008)
--	g26233 = AND(g2279, g25309)
--	I31071 = AND(g31170, g31808, g32557, g32558)
--	g26182 = AND(g9978, g25317)
--	g26651 = AND(g22707, g24425)
--	g12015 = AND(g1002, g7567)
--	g34081 = AND(g33706, g19552)
--	g27486 = AND(g26519, g17645)
--	g31962 = AND(g8033, g31013)
--	g24763 = AND(g17569, g22457)
--	g33406 = AND(g32355, g21399)
--	g18269 = AND(g15069, g16031)
--	g33361 = AND(g32257, g20911)
--	g15903 = AND(g13796, g13223)
--	g18773 = AND(g5694, g15615)
--	I31147 = AND(g32668, g32669, g32670, g32671)
--	g18341 = AND(g1648, g17873)
--	g29515 = AND(g28888, g22342)
--	g29882 = AND(g2361, g29151)
--	g18268 = AND(g1280, g16000)
--	g29991 = AND(g29179, g12922)
--	g21753 = AND(g3179, g20785)
--	g31500 = AND(g29802, g23449)
--	g18156 = AND(g572, g17533)
--	g18655 = AND(g15106, g14454)
--	g33500 = AND(g32744, I31196, I31197)
--	g24660 = AND(g22648, g19737)
--	g33833 = AND(g33093, g25852)
--	g32203 = AND(g4249, g31327)
--	g18180 = AND(g767, g17328)
--	g26513 = AND(g19501, g24365)
--	g17418 = AND(g9618, g14407)
--	I27409 = AND(g25556, g26424, g22698)
--	g34999 = AND(g34998, g23085)
--	g18670 = AND(g4621, g15758)
--	g34380 = AND(g34158, g20571)
--	g25482 = AND(g5752, g23816, I24597)
--	g32044 = AND(g31483, g20085)
--	I24684 = AND(g20014, g24033, g24034, g24035)
--	g16612 = AND(g5603, g14927)
--	g21736 = AND(g3065, g20330)
--	g11546 = AND(g7289, g4375)
--	g21887 = AND(g15101, g19801)
--	g30233 = AND(g28720, g23913)
--	g18734 = AND(g4966, g16826)
--	I31151 = AND(g30825, g31822, g32673, g32674)
--	g16324 = AND(g13657, g182)
--	I31172 = AND(g32703, g32704, g32705, g32706)
--	g18335 = AND(g1687, g17873)
--	g16701 = AND(g5547, g14845)
--	g22589 = AND(g19267, g19451)
--	g32281 = AND(g31257, g20500)
--	g34182 = AND(g33691, g24384)
--	g28255 = AND(g8515, g27983)
--	g16534 = AND(g5575, g14665)
--	g28679 = AND(g27572, g20638)
--	g11024 = AND(g5436, g9070)
--	g16098 = AND(g5148, g14238)
--	I13937 = AND(g7340, g7293, g7261)
--	g18993 = AND(g11224, g16172)
--	g24550 = AND(g3684, g23308)
--	g32301 = AND(g31276, g20547)
--	g14643 = AND(g11998, g12023)
--	g24314 = AND(g4515, g22228)
--	g22588 = AND(g79, g20078)
--	g21843 = AND(g3869, g21070)
--	g32120 = AND(g31639, g29941)
--	g24287 = AND(g4401, g22550)
--	g28124 = AND(g27368, g22842)
--	g15794 = AND(g3239, g14008)
--	g18667 = AND(g4601, g17367)
--	g18694 = AND(g4722, g16053)
--	g12179 = AND(g9745, g10027)
--	g24307 = AND(g4486, g22228)
--	g29584 = AND(g1706, g29018)
--	g27178 = AND(g25997, g16652)
--	g21764 = AND(g3227, g20785)
--	g11497 = AND(g6398, g7192)
--	g18131 = AND(g482, g16971)
--	g29206 = AND(g24124, I27528, I27529)
--	g13497 = AND(g2724, g12155)
--	g28686 = AND(g27574, g20650)
--	g32146 = AND(g31624, g29978)
--	g28939 = AND(g17321, g25184, g26424, g27421)
--	g24721 = AND(g17488, g22369)
--	g22119 = AND(g6581, g19277)
--	g21869 = AND(g4087, g19801)
--	g27186 = AND(g26195, g8316, g2342)
--	g31273 = AND(g30143, g27779)
--	g34513 = AND(g9003, g34346)
--	g21960 = AND(g5421, g21514)
--	g27676 = AND(g26377, g20627)
--	g27685 = AND(g13032, g25895)
--	g15633 = AND(g3841, g13584)
--	g33106 = AND(g32408, g18990)
--	g18487 = AND(g2441, g15426)
--	g27373 = AND(g26488, g17477)
--	g29759 = AND(g28308, g23226)
--	g22118 = AND(g6605, g19277)
--	g32290 = AND(g31267, g20525)
--	g11126 = AND(g6035, g10185)
--	g12186 = AND(g1178, g7519)
--	g28267 = AND(g7328, g2227, g27421)
--	g17401 = AND(g1083, g13143)
--	g21868 = AND(g4076, g19801)
--	g18619 = AND(g3466, g17062)
--	g18502 = AND(g2567, g15509)
--	g22022 = AND(g5873, g19147)
--	g34961 = AND(g34944, g23019)
--	g12953 = AND(g411, g11048)
--	g18557 = AND(g2771, g15277)
--	g33812 = AND(g23088, g33187, g9104)
--	g18210 = AND(g936, g15938)
--	g29758 = AND(g28306, g23222)
--	g17119 = AND(g5272, g14800)
--	g33463 = AND(g32477, I31011, I31012)
--	I31227 = AND(g32784, g32785, g32786, g32787)
--	g18618 = AND(g3457, g17062)
--	g18443 = AND(g2265, g18008)
--	g24773 = AND(g22832, g19872)
--	g21709 = AND(g283, g20283)
--	g18279 = AND(g1361, g16136)
--	g30026 = AND(g28476, g25064)
--	g33371 = AND(g32280, g21155)
--	g30212 = AND(g28687, g23879)
--	g16766 = AND(g6649, g12915)
--	g26387 = AND(g24813, g20231)
--	g27334 = AND(g12539, g26769)
--	g34212 = AND(g33761, g22689)
--	g28219 = AND(g9316, g27573)
--	g21708 = AND(g15049, g20283)
--	g18278 = AND(g1345, g16136)
--	I16111 = AND(g8691, g11409, g11381)
--	g26148 = AND(g25357, g11724, g11709, g11686)
--	g23708 = AND(g19050, g9104)
--	g16871 = AND(g6597, g14908)
--	g29345 = AND(g4749, g28376)
--	g22053 = AND(g6116, g21611)
--	g23471 = AND(g20148, g20523)
--	g26097 = AND(g5821, g25092)
--	g18469 = AND(g2399, g15224)
--	g24670 = AND(g5138, g23590)
--	g33795 = AND(g33138, g20782)
--	g28218 = AND(g27768, g26645)
--	g29940 = AND(g1740, g28758)
--	g26104 = AND(g2250, g25101)
--	g18286 = AND(g1404, g16164)
--	g22900 = AND(g17137, g19697)
--	g27762 = AND(g22472, g25226, g26424, g26218)
--	g15861 = AND(g3957, g14170)
--	g8690 = AND(g2941, g2936)
--	g27964 = AND(g25956, g22492)
--	g18468 = AND(g2393, g15224)
--	g25331 = AND(g5366, g22194, I24508)
--	g18306 = AND(g15074, g16931)
--	g12762 = AND(g4358, g8977)
--	g22036 = AND(g5937, g19147)
--	g25449 = AND(g6946, g22496)
--	g13060 = AND(g8587, g11110)
--	g31514 = AND(g20041, g29956)
--	g32403 = AND(g31117, g15842)
--	g27216 = AND(g26055, g16725)
--	g33514 = AND(g32844, I31266, I31267)
--	g22101 = AND(g6474, g18833)
--	g24930 = AND(g4826, g23948)
--	g29652 = AND(g2667, g29157)
--	g29804 = AND(g1592, g29014)
--	g17809 = AND(g7873, g13125)
--	I31281 = AND(g30735, g31845, g32861, g32862)
--	g28160 = AND(g26309, g27463)
--	g15612 = AND(g3143, g13530)
--	g25448 = AND(g11202, g22680)
--	g18815 = AND(g6523, g15483)
--	g30149 = AND(g28605, g21248)
--	g25961 = AND(g25199, g20682)
--	I27381 = AND(g25549, g26424, g22698)
--	g33507 = AND(g32795, I31231, I31232)
--	I31301 = AND(g31327, g31849, g32889, g32890)
--	g20131 = AND(g15170, g14309)
--	g15701 = AND(g3821, g13584)
--	g10705 = AND(g6850, g10219, g2689)
--	g18601 = AND(g3106, g16987)
--	g13411 = AND(g4955, g11834)
--	g18187 = AND(g794, g17328)
--	g18677 = AND(g4639, g15758)
--	g14610 = AND(g1484, g10935)
--	g28455 = AND(g27289, g20103)
--	g33421 = AND(g32374, g21455)
--	g21810 = AND(g3578, g20924)
--	g17177 = AND(g6657, g14984)
--	g21774 = AND(g3361, g20391)
--	g29332 = AND(g29107, g22170)
--	g23657 = AND(g19401, g11941)
--	g28617 = AND(g27533, g20552)
--	g34097 = AND(g33772, g9104, g18957)
--	g21955 = AND(g5385, g21514)
--	g23774 = AND(g14867, g21252)
--	g22064 = AND(g15162, g19210)
--	I24600 = AND(g6077, g6082, g9946)
--	I31146 = AND(g30735, g31821, g32666, g32667)
--	g25026 = AND(g22929, g10503)
--	g34104 = AND(g33916, g23639)
--	g27117 = AND(g26055, g16528)
--	g21879 = AND(g4132, g19801)
--	g34811 = AND(g14165, g34766)
--	g21970 = AND(g5401, g21514)
--	g18143 = AND(g586, g17533)
--	g24502 = AND(g23428, g13223)
--	g28201 = AND(g27499, g16720)
--	g19536 = AND(g518, g16768)
--	g19948 = AND(g17515, g16320)
--	g29962 = AND(g23616, g28959)
--	g21878 = AND(g4129, g19801)
--	I16695 = AND(g10207, g12523, g12463)
--	g32127 = AND(g31624, g29950)
--	g31541 = AND(g22536, g29348)
--	g24618 = AND(g22625, g19672)
--	g26229 = AND(g1724, g25275)
--	g33473 = AND(g32549, I31061, I31062)
--	g18169 = AND(g676, g17433)
--	g21886 = AND(g4153, g19801)
--	g27568 = AND(g26576, g17791)
--	g18791 = AND(g6044, g15634)
--	g31789 = AND(g30201, g24013)
--	g28467 = AND(g26993, g12295)
--	g28494 = AND(g27973, g17741)
--	g33789 = AND(g33159, g23022)
--	g21792 = AND(g3396, g20391)
--	g16591 = AND(g5256, g14879)
--	g22009 = AND(g5782, g21562)
--	g22665 = AND(g17174, g20905)
--	g18168 = AND(g681, g17433)
--	g18410 = AND(g2079, g15373)
--	g21967 = AND(g5456, g21514)
--	g21994 = AND(g5607, g19074)
--	g31788 = AND(g21352, g29385)
--	g33724 = AND(g14145, g33258)
--	g32376 = AND(g2689, g31710)
--	g19564 = AND(g17175, g13976)
--	g33359 = AND(g32252, g20853)
--	g25149 = AND(g14030, g23546)
--	g17693 = AND(g1306, g13291)
--	g22008 = AND(g5774, g21562)
--	g32103 = AND(g31609, g29905)
--	g24286 = AND(g4405, g22550)
--	g18479 = AND(g2449, g15426)
--	g18666 = AND(g4593, g17367)
--	g33829 = AND(g33240, g20164)
--	g18363 = AND(g1840, g17955)
--	g32095 = AND(g7619, g30825)
--	g18217 = AND(g15063, g16100)
--	g33434 = AND(g32239, g29702)
--	g24306 = AND(g4483, g22228)
--	g33358 = AND(g32249, g20778)
--	g25148 = AND(g16867, g23545)
--	g11496 = AND(g4382, g7495)
--	g15871 = AND(g3203, g13951)
--	g18478 = AND(g2445, g15426)
--	g30133 = AND(g28591, g21179)
--	g33828 = AND(g33090, g24411)
--	g28352 = AND(g10014, g27705)
--	g11111 = AND(g5297, g7004, g5283, g9780)
--	g14875 = AND(g1495, g10939)
--	g34133 = AND(g33845, g23958)
--	g21919 = AND(g15144, g21468)
--	g30229 = AND(g28716, g23904)
--	g25104 = AND(g16800, g23504)
--	g11978 = AND(g2629, g7462)
--	g26310 = AND(g2102, g25389)
--	g23919 = AND(g4122, g19546)
--	g32181 = AND(g31020, g19912)
--	g33121 = AND(g8748, g32212)
--	g18486 = AND(g2485, g15426)
--	g27230 = AND(g25906, g19558)
--	g27293 = AND(g9972, g26655)
--	g29613 = AND(g28208, g19763)
--	g28266 = AND(g23748, g27714)
--	g19062 = AND(g446, g16180)
--	g33344 = AND(g32228, g20670)
--	g14218 = AND(g875, g10632)
--	g21918 = AND(g5097, g21468)
--	g30228 = AND(g28715, g23903)
--	g26379 = AND(g19904, g25546)
--	g18556 = AND(g2823, g15277)
--	g25971 = AND(g1917, g24992)
--	g24187 = AND(g305, g22722)
--	g34228 = AND(g33750, g22942)
--	g30011 = AND(g29183, g12930)
--	g27265 = AND(g26785, g26759)
--	I31226 = AND(g29385, g32781, g32782, g32783)
--	g16844 = AND(g7212, g13000)
--	g18580 = AND(g2907, g16349)
--	g26050 = AND(g9630, g25047)
--	g27416 = AND(g8046, g26314, g9187, g504)
--	g26378 = AND(g19576, g25544)
--	g13384 = AND(g4944, g11804)
--	g29605 = AND(g2445, g28973)
--	g18223 = AND(g1030, g16100)
--	g23599 = AND(g19050, g9104)
--	g27992 = AND(g26800, g23964)
--	g22074 = AND(g6239, g19210)
--	g27391 = AND(g26549, g17505)
--	g24143 = AND(g17694, g21659)
--	g25368 = AND(g6946, g22408)
--	g27510 = AND(g26576, g17687)
--	g34582 = AND(g7764, g34313)
--	g32190 = AND(g142, g31233)
--	g26096 = AND(g9733, g25268)
--	g29951 = AND(g1874, g28786)
--	g18110 = AND(g441, g17015)
--	g34310 = AND(g14003, g34162)
--	g25850 = AND(g3502, g24636)
--	g15911 = AND(g3111, g13530)
--	g28588 = AND(g27489, g20499)
--	g28524 = AND(g6821, g27084)
--	I31127 = AND(g32638, g32639, g32640, g32641)
--	g18321 = AND(g1620, g17873)
--	g24884 = AND(g3401, g23555, I24051)
--	g30925 = AND(g29908, g23309)
--	g21817 = AND(g3606, g20924)
--	g11019 = AND(g5092, g9036)
--	g18179 = AND(g763, g17328)
--	g13019 = AND(g194, g11737)
--	g18531 = AND(g2719, g15277)
--	g30112 = AND(g28566, g20919)
--	g28477 = AND(g27966, g17676)
--	g33760 = AND(g33143, g20328)
--	g24410 = AND(g3817, g23139)
--	g32089 = AND(g27261, g31021)
--	g25229 = AND(g7636, g22654)
--	g30050 = AND(g22545, g28126)
--	g29795 = AND(g28344, g23257)
--	g34112 = AND(g22957, g9104, g33778)
--	g11018 = AND(g7655, g7643, g7627)
--	g18178 = AND(g758, g17328)
--	g18740 = AND(g4572, g17384)
--	g26857 = AND(g25062, g25049)
--	g34050 = AND(g33772, g22942)
--	g21977 = AND(g5535, g19074)
--	g22092 = AND(g6419, g18833)
--	g23532 = AND(g19400, g11852)
--	g23901 = AND(g19606, g7963)
--	g34378 = AND(g13095, g34053)
--	g16025 = AND(g446, g14063)
--	g33506 = AND(g32788, I31226, I31227)
--	I24530 = AND(g9501, g9733, g5747)
--	g32088 = AND(g27241, g31070)
--	g24666 = AND(g11753, g22975)
--	g22518 = AND(g12982, g19398)
--	g21783 = AND(g3419, g20391)
--	I31297 = AND(g32884, g32885, g32886, g32887)
--	g24217 = AND(g18200, g22594)
--	g18186 = AND(g753, g17328)
--	g15785 = AND(g3558, g14107)
--	g18676 = AND(g4358, g15758)
--	g18685 = AND(g4688, g15885)
--	g34386 = AND(g10800, g34060)
--	g18373 = AND(g1890, g15171)
--	g29514 = AND(g1608, g28780)
--	g24015 = AND(g19540, g10951)
--	g30096 = AND(g28546, g20770)
--	g22637 = AND(g19363, g19489)
--	g17176 = AND(g8616, g13008)
--	g34742 = AND(g9000, g34698)
--	g28616 = AND(g27532, g20551)
--	g34096 = AND(g22957, g9104, g33772)
--	g18654 = AND(g4146, g16249)
--	g16203 = AND(g5821, g14297)
--	g28313 = AND(g27231, g19766)
--	g27116 = AND(g26026, g16527)
--	I27509 = AND(g24084, g24085, g24086, g24087)
--	g21823 = AND(g3731, g20453)
--	g27615 = AND(g26789, g26770)
--	g18800 = AND(g6187, g15348)
--	g15859 = AND(g3610, g13923)
--	I31181 = AND(g29385, g32716, g32717, g32718)
--	g18417 = AND(g2116, g15373)
--	g24556 = AND(g4035, g23341)
--	g28285 = AND(g9657, g27717)
--	g34681 = AND(g34491, g19438)
--	I27508 = AND(g19935, g24082, g24083, g28033)
--	g15858 = AND(g3542, g14045)
--	g27041 = AND(g8519, g26330)
--	g32126 = AND(g31601, g29948)
--	g18334 = AND(g1696, g17873)
--	g27275 = AND(g25945, g19745)
--	g19756 = AND(g9899, g17154)
--	g33927 = AND(g33094, g21412)
--	g28254 = AND(g7268, g1668, g27395)
--	g27430 = AND(g26488, g17579)
--	g34857 = AND(g16540, g34813)
--	g10822 = AND(g4264, g8514)
--	g24223 = AND(g239, g22594)
--	g27493 = AND(g246, g26837)
--	g16957 = AND(g13064, g10418)
--	g25959 = AND(g1648, g24963)
--	g30730 = AND(g26346, g29778)
--	g25925 = AND(g24990, g23234)
--	g28466 = AND(g27960, g17637)
--	g25112 = AND(g10428, g23510)
--	g21966 = AND(g5406, g21514)
--	g18762 = AND(g5475, g17929)
--	g25050 = AND(g13056, g22312)
--	g20084 = AND(g11591, g16609)
--	g32339 = AND(g31474, g20672)
--	g31240 = AND(g14793, g30206)
--	g19350 = AND(g15968, g13505)
--	g34765 = AND(g34692, g20057)
--	g27340 = AND(g10199, g26784)
--	g27035 = AND(g26348, g1500)
--	g18423 = AND(g12851, g18008)
--	g29789 = AND(g28270, g10233)
--	g32338 = AND(g31466, g20668)
--	g33491 = AND(g32679, I31151, I31152)
--	g33903 = AND(g33447, g19146)
--	g24922 = AND(g4831, g23931)
--	g26129 = AND(g2384, g25121)
--	g18216 = AND(g967, g15979)
--	g24321 = AND(g4558, g22228)
--	g16699 = AND(g7134, g12933)
--	g27684 = AND(g26386, g20657)
--	g28642 = AND(g27555, g20598)
--	g18587 = AND(g2980, g16349)
--	g25096 = AND(g23778, g20560)
--	g29788 = AND(g28335, g23250)
--	g26128 = AND(g2319, g25120)
--	g14589 = AND(g10586, g10569)
--	g29535 = AND(g2303, g28871)
--	I31211 = AND(g31021, g31833, g32759, g32760)
--	g27517 = AND(g26400, g17707)
--	g10588 = AND(g7004, g5297)
--	g18909 = AND(g16226, g13570)
--	g32197 = AND(g31144, g20088)
--	g18543 = AND(g2779, g15277)
--	g26323 = AND(g10262, g25273)
--	g24186 = AND(g18102, g22722)
--	g14588 = AND(g11957, g11974)
--	g24676 = AND(g2748, g23782)
--	I16721 = AND(g10224, g12589, g12525)
--	g18117 = AND(g464, g17015)
--	g16427 = AND(g5216, g14876)
--	g25802 = AND(g8106, g24586)
--	g22083 = AND(g6287, g19210)
--	g32411 = AND(g31119, g13469)
--	g23023 = AND(g650, g20248)
--	g19691 = AND(g9614, g17085)
--	g24654 = AND(g11735, g22922)
--	g28630 = AND(g27544, g20575)
--	g29344 = AND(g29168, g18932)
--	g18569 = AND(g94, g16349)
--	g30002 = AND(g28481, g23487)
--	g27130 = AND(g26026, g16585)
--	g30057 = AND(g29144, g9462)
--	g22622 = AND(g19336, g19469)
--	g18568 = AND(g37, g16349)
--	g18747 = AND(g5138, g17847)
--	g25765 = AND(g24989, g24973)
--	g27362 = AND(g26080, g20036)
--	g31990 = AND(g31772, g18945)
--	g33899 = AND(g32132, g33335)
--	g18242 = AND(g962, g16431)
--	g10616 = AND(g7998, g174)
--	g27523 = AND(g26549, g17718)
--	g30245 = AND(g28733, g23935)
--	I31126 = AND(g30673, g31818, g32636, g32637)
--	g26232 = AND(g2193, g25396)
--	g33898 = AND(g33419, g15655)
--	g21816 = AND(g3602, g20924)
--	g18123 = AND(g479, g16886)
--	g18814 = AND(g6519, g15483)
--	g33719 = AND(g33141, g19433)
--	g24762 = AND(g655, g23573)
--	g10704 = AND(g2145, g10200, g2130)
--	g34533 = AND(g34318, g19731)
--	g18751 = AND(g5156, g17847)
--	g18807 = AND(g6386, g15656)
--	g21976 = AND(g5527, g19074)
--	g21985 = AND(g5571, g19074)
--	g15902 = AND(g441, g13975)
--	g18772 = AND(g5689, g15615)
--	g28555 = AND(g27429, g20373)
--	g33718 = AND(g33147, g19432)
--	g34298 = AND(g8679, g34132)
--	g28454 = AND(g26976, g12233)
--	g33521 = AND(g32895, I31301, I31302)
--	g18974 = AND(g174, g16127)
--	g26261 = AND(g24688, g10678, g8778, g8757)
--	g32315 = AND(g31306, g23517)
--	g24423 = AND(g4950, g22897)
--	g21752 = AND(g3171, g20785)
--	g27727 = AND(g22432, g25211, g26424, g26195)
--	I31296 = AND(g30937, g31848, g32882, g32883)
--	g18639 = AND(g3831, g17096)
--	g28570 = AND(g27456, g20434)
--	g28712 = AND(g27590, g20708)
--	g21954 = AND(g5381, g21514)
--	g27222 = AND(g26055, g13932)
--	g29760 = AND(g28309, g23227)
--	g33832 = AND(g33088, g27991)
--	g18230 = AND(g1111, g16326)
--	g29029 = AND(g14506, g25227, g26424, g27494)
--	g17139 = AND(g8635, g12967)
--	g18293 = AND(g1484, g16449)
--	g17653 = AND(g11547, g11592, g6789, I18620)
--	g15738 = AND(g1111, g13260)
--	g18638 = AND(g3827, g17096)
--	g27437 = AND(g26576, g17589)
--	g33440 = AND(g32250, g29719)
--	g32055 = AND(g10999, g30825)
--	g17138 = AND(g255, g13239)
--	g18265 = AND(g1270, g16000)
--	g25129 = AND(g17682, g23527)
--	g15699 = AND(g1437, g13861)
--	g30232 = AND(g28719, g23912)
--	g32111 = AND(g31616, g29922)
--	g18416 = AND(g2112, g15373)
--	g25057 = AND(g23275, g20511)
--	g32070 = AND(g10967, g30825)
--	g33861 = AND(g33271, g20502)
--	g28239 = AND(g27135, g19659)
--	g25128 = AND(g17418, g23525)
--	g17636 = AND(g10829, g13463)
--	g11916 = AND(g2227, g7328)
--	g33247 = AND(g32130, g19980)
--	g28567 = AND(g6832, g27101)
--	I31197 = AND(g32740, g32741, g32742, g32743)
--	g27347 = AND(g26400, g17390)
--	g18992 = AND(g8341, g16171)
--	g18391 = AND(g1982, g15171)
--	g24908 = AND(g3752, g23239, I24075)
--	g28238 = AND(g27133, g19658)
--	g21842 = AND(g3863, g21070)
--	g18510 = AND(g2625, g15509)
--	g30261 = AND(g28772, g23961)
--	g23392 = AND(g7247, g21430)
--	g24569 = AND(g5115, g23382)
--	g25323 = AND(g6888, g22359)
--	g31324 = AND(g30171, g27937)
--	g33099 = AND(g32395, g18944)
--	g13287 = AND(g1221, g11472)
--	g27600 = AND(g26755, g26725)
--	g10733 = AND(g3639, g6905, g3625, g8542)
--	g18579 = AND(g2984, g16349)
--	g31777 = AND(g21343, g29385)
--	g33701 = AND(g33162, g16305)
--	g24747 = AND(g17510, g22417)
--	g32067 = AND(g4727, g30614)
--	g21559 = AND(g16236, g10897)
--	g31272 = AND(g30117, g27742)
--	I16618 = AND(g10124, g12341, g12293)
--	g15632 = AND(g3494, g13555)
--	g28185 = AND(g27026, g19435)
--	g10874 = AND(g7791, g6219, g6227)
--	g18578 = AND(g2873, g16349)
--	g25775 = AND(g2922, g24568)
--	g23424 = AND(g7345, g21556)
--	g27351 = AND(g10218, g26804)
--	g27372 = AND(g26488, g17476)
--	g19768 = AND(g2803, g15833)
--	g14874 = AND(g1099, g10909)
--	g16671 = AND(g6275, g14817)
--	g21558 = AND(g15904, g13729)
--	g27821 = AND(g7680, g25892)
--	g32150 = AND(g31624, g29995)
--	g28154 = AND(g8492, g27306)
--	g18586 = AND(g2886, g16349)
--	g29649 = AND(g2241, g28678)
--	g33462 = AND(g32470, I31006, I31007)
--	g21830 = AND(g3774, g20453)
--	g26611 = AND(g24935, g20580)
--	g20751 = AND(g16260, g4836)
--	g10665 = AND(g209, g8292)
--	g28637 = AND(g22399, g27011)
--	g18442 = AND(g2259, g18008)
--	g32019 = AND(g30579, g22358)
--	g24772 = AND(g16287, g23061)
--	g29648 = AND(g2112, g29121)
--	g27264 = AND(g25941, g19714)
--	g22115 = AND(g6573, g19277)
--	g27137 = AND(g26026, g16606)
--	g21865 = AND(g3965, g21070)
--	g31140 = AND(g2102, g30037)
--	g32196 = AND(g27587, g31376)
--	g13942 = AND(g5897, g12512)
--	g24639 = AND(g6181, g23699)
--	g32018 = AND(g4146, g30937)
--	g26271 = AND(g1992, g25341)
--	g29604 = AND(g2315, g28966)
--	g30316 = AND(g29199, g7097, g6682)
--	g21713 = AND(g298, g20283)
--	g34499 = AND(g31288, g34339)
--	g24230 = AND(g901, g22594)
--	g13156 = AND(g10816, g10812, g10805)
--	g18116 = AND(g168, g17015)
--	g24293 = AND(g4438, g22550)
--	g18615 = AND(g3347, g17200)
--	g22052 = AND(g6113, g21611)
--	g10476 = AND(g7244, g7259, I13862)
--	g24638 = AND(g22763, g19690)
--	g29770 = AND(g28320, g23238)
--	g16190 = AND(g14626, g11810)
--	g29563 = AND(g1616, g28853)
--	I31202 = AND(g32747, g32748, g32749, g32750)
--	g34498 = AND(g13888, g34336)
--	g18720 = AND(g15137, g16795)
--	g26753 = AND(g16024, g24452)
--	I31257 = AND(g32826, g32827, g32828, g32829)
--	g25880 = AND(g8443, g24814)
--	g14555 = AND(g12521, g12356, g12307, I16671)
--	g24416 = AND(g4939, g22870)
--	g16520 = AND(g5909, g14965)
--	g21705 = AND(g209, g20283)
--	g30056 = AND(g29165, g12659)
--	g18275 = AND(g15070, g16136)
--	g26145 = AND(g11962, g25131)
--	I31111 = AND(g31070, g31815, g32615, g32616)
--	g18430 = AND(g2204, g18008)
--	g18746 = AND(g5134, g17847)
--	g27209 = AND(g26213, g8365, g2051)
--	g32402 = AND(g4888, g30990)
--	g18493 = AND(g2514, g15426)
--	g33871 = AND(g33281, g20546)
--	g30080 = AND(g28121, g20674)
--	g28215 = AND(g9264, g27565)
--	g26650 = AND(g10796, g24424)
--	g34080 = AND(g22957, g9104, g33750)
--	g16211 = AND(g5445, g14215)
--	g27208 = AND(g9037, g26598)
--	g18465 = AND(g2384, g15224)
--	g29767 = AND(g28317, g23236)
--	g29794 = AND(g28342, g23256)
--	g21188 = AND(g7666, g15705)
--	g33360 = AND(g32253, g20869)
--	g18237 = AND(g1146, g16326)
--	g29845 = AND(g28375, g23291)
--	g23188 = AND(g13994, g20025)
--	I16143 = AND(g8751, g11491, g11445)
--	g28439 = AND(g27273, g10233)
--	g18340 = AND(g1720, g17873)
--	g29899 = AND(g28428, g23375)
--	g29990 = AND(g29007, g9239)
--	g21939 = AND(g5224, g18997)
--	g25831 = AND(g3151, g24623)
--	g15784 = AND(g3235, g13977)
--	g18806 = AND(g6381, g15656)
--	g18684 = AND(g4681, g15885)
--	g26393 = AND(g19467, g25558)
--	g14567 = AND(g10568, g10552)
--	g24835 = AND(g8720, g23233)
--	g29633 = AND(g1978, g29085)
--	I31067 = AND(g32552, g32553, g32554, g32555)
--	g24014 = AND(g7933, g19063)
--	g15103 = AND(g4180, g14454)
--	g34753 = AND(g34676, g19586)
--	g21938 = AND(g5216, g18997)
--	g18142 = AND(g577, g17533)
--	g34342 = AND(g34103, g19998)
--	g30145 = AND(g28603, g21247)
--	g30031 = AND(g29071, g10540)
--	g27614 = AND(g26785, g26759)
--	g32256 = AND(g31249, g20382)
--	g18517 = AND(g2652, g15509)
--	g27436 = AND(g26576, g17588)
--	g30199 = AND(g28664, g23861)
--	g29718 = AND(g28512, g11136)
--	g29521 = AND(g1744, g28824)
--	g16700 = AND(g5208, g14838)
--	g31220 = AND(g30273, g25202)
--	g33472 = AND(g32542, I31056, I31057)
--	g16126 = AND(g5495, g14262)
--	g28284 = AND(g11398, g27994)
--	g10675 = AND(g3436, g8500)
--	g25989 = AND(g25258, g21012)
--	g27073 = AND(g7121, g3873, g3881, g26281)
--	g30198 = AND(g28662, g23860)
--	g32300 = AND(g31274, g20544)
--	g14185 = AND(g8686, g11744)
--	g25056 = AND(g12779, g23456)
--	g28304 = AND(g27226, g19753)
--	g33911 = AND(g33137, g10725)
--	g34198 = AND(g33688, g24491)
--	g26161 = AND(g2518, g25139)
--	g34529 = AND(g34306, g19634)
--	g21875 = AND(g4116, g19801)
--	g25988 = AND(g9510, g25016)
--	I31196 = AND(g30825, g31830, g32738, g32739)
--	g25924 = AND(g24976, g16846)
--	g27346 = AND(g26400, g17389)
--	g34528 = AND(g34305, g19617)
--	g17692 = AND(g1124, g13307)
--	g18130 = AND(g528, g16971)
--	g34696 = AND(g34531, g20004)
--	g18193 = AND(g837, g17821)
--	g22013 = AND(g5802, g21562)
--	g32157 = AND(g31646, g30021)
--	g34393 = AND(g34189, g21304)
--	g26259 = AND(g24430, g25232)
--	I24508 = AND(g9434, g9672, g5401)
--	g18362 = AND(g1834, g17955)
--	g23218 = AND(g20200, g16530)
--	g29861 = AND(g28390, g23313)
--	g29573 = AND(g1752, g28892)
--	g33071 = AND(g31591, g32404)
--	g21837 = AND(g3719, g20453)
--	g34764 = AND(g34691, g20009)
--	g22329 = AND(g11940, g20329)
--	g10883 = AND(g3355, g9061)
--	g18165 = AND(g650, g17433)
--	g23837 = AND(g21160, g10804)
--	g18523 = AND(g2675, g15509)
--	g26087 = AND(g5475, g25072)
--	g27034 = AND(g26328, g8609)
--	g13306 = AND(g441, g11048)
--	g31776 = AND(g21329, g29385)
--	g34365 = AND(g34149, g20451)
--	g26258 = AND(g12875, g25231)
--	g19651 = AND(g1111, g16119)
--	g33785 = AND(g33100, g20550)
--	g29926 = AND(g1604, g28736)
--	g34869 = AND(g34816, g19869)
--	g28139 = AND(g27337, g26054)
--	g22005 = AND(g5759, g21562)
--	g31147 = AND(g12286, g30054)
--	g28653 = AND(g7544, g27014)
--	g13038 = AND(g8509, g11034)
--	g27292 = AND(g1714, g26654)
--	g29612 = AND(g27875, g28633)
--	g24465 = AND(g3827, g23139)
--	g12641 = AND(g10295, g3171, g3179)
--	g22538 = AND(g14035, g20248)
--	g27153 = AND(g26055, g16629)
--	g33355 = AND(g32243, g20769)
--	g29324 = AND(g29078, g18883)
--	g34868 = AND(g34813, g19866)
--	g7396 = AND(g392, g441)
--	g25031 = AND(g20675, g23432)
--	g30161 = AND(g28614, g21275)
--	g18475 = AND(g12853, g15426)
--	g33859 = AND(g33426, g10531)
--	g26244 = AND(g24688, g8812, g10658, g8757)
--	g29534 = AND(g28965, g22457)
--	g33370 = AND(g32279, g21139)
--	g24983 = AND(g23217, g20238)
--	g27409 = AND(g26519, g17524)
--	g16855 = AND(g4392, g13107)
--	g18727 = AND(g4931, g16077)
--	g28415 = AND(g27250, g19963)
--	g24684 = AND(g11769, g22989)
--	g28333 = AND(g27239, g19787)
--	g33858 = AND(g33268, g20448)
--	g34709 = AND(g34549, g17242)
--	g18222 = AND(g1024, g16100)
--	g10501 = AND(g1233, g9007)
--	g16870 = AND(g6625, g14905)
--	g27136 = AND(g26026, g16605)
--	g27408 = AND(g26519, g17523)
--	g27635 = AND(g23032, g26281, g26424, g24996)
--	g21915 = AND(g5080, g21468)
--	g30225 = AND(g28705, g23897)
--	g31151 = AND(g10037, g30065)
--	g18437 = AND(g2241, g18008)
--	g24142 = AND(g17700, g21657)
--	I31001 = AND(g29385, g32456, g32457, g32458)
--	g31996 = AND(g31779, g18979)
--	g34225 = AND(g33744, g22942)
--	I31077 = AND(g32566, g32567, g32568, g32569)
--	g26602 = AND(g7487, g24453)
--	g30258 = AND(g28751, g23953)
--	g11937 = AND(g1936, g7362)
--	g15860 = AND(g3889, g14160)
--	g34087 = AND(g33766, g9104, g18957)
--	g23201 = AND(g14027, g20040)
--	g33844 = AND(g33257, g20327)
--	g33367 = AND(g32271, g21053)
--	I31256 = AND(g31021, g31841, g32824, g32825)
--	g18703 = AND(g4776, g16782)
--	g22100 = AND(g6466, g18833)
--	g18347 = AND(g1756, g17955)
--	g19717 = AND(g6527, g17122)
--	g14438 = AND(g1087, g10726)
--	g30043 = AND(g29106, g9392)
--	g18253 = AND(g1211, g16897)
--	g25132 = AND(g10497, g23528)
--	g30244 = AND(g28732, g23930)
--	g26171 = AND(g25357, g6856, g11709, g11686)
--	g15700 = AND(g3089, g13483)
--	I24051 = AND(g3380, g3385, g8492)
--	g18600 = AND(g3111, g16987)
--	g20193 = AND(g15578, g17264)
--	g18781 = AND(g5831, g18065)
--	g28585 = AND(g27063, g10530)
--	g24193 = AND(g336, g22722)
--	g28484 = AND(g27187, g10290, g21163, I26972)
--	g33420 = AND(g32373, g21454)
--	g30069 = AND(g29175, g12708)
--	g29766 = AND(g28316, g23235)
--	g18236 = AND(g15065, g16326)
--	g21782 = AND(g3416, g20391)
--	g17771 = AND(g13288, g13190)
--	g20165 = AND(g5156, g17733)
--	g34069 = AND(g8774, g33797)
--	g21984 = AND(g5563, g19074)
--	I31102 = AND(g32603, g32604, g32605, g32606)
--	g26994 = AND(g23032, g26226, g26424, g25557)
--	g27474 = AND(g8038, g26314, g518, g504)
--	g28554 = AND(g27426, g20372)
--	I31157 = AND(g32682, g32683, g32684, g32685)
--	g18351 = AND(g1760, g17955)
--	g18372 = AND(g1886, g15171)
--	g24523 = AND(g22318, g19468)
--	g32314 = AND(g31304, g23516)
--	g29871 = AND(g28400, g23332)
--	g33446 = AND(g32385, g21607)
--	g27711 = AND(g22369, g25193, g26424, g26166)
--	g16707 = AND(g6641, g15033)
--	g21419 = AND(g16681, g13595)
--	g32287 = AND(g2823, g30578)
--	g34774 = AND(g34695, g20180)
--	g18175 = AND(g744, g17328)
--	g18821 = AND(g15168, g15680)
--	g34955 = AND(g34931, g34320)
--	g27327 = AND(g2116, g26732)
--	g34375 = AND(g13077, g34049)
--	g16202 = AND(g86, g14197)
--	g28312 = AND(g27828, g26608)
--	g28200 = AND(g27652, g11383)
--	g32307 = AND(g31291, g23500)
--	g14566 = AND(g10566, g10551)
--	g32085 = AND(g27253, g31021)
--	I31066 = AND(g31070, g31807, g32550, g32551)
--	g29360 = AND(g27364, g28294)
--	g21822 = AND(g3727, g20453)
--	g22515 = AND(g12981, g19395)
--	I31231 = AND(g31376, g31836, g32789, g32790)
--	g22991 = AND(g645, g20248)
--	g27537 = AND(g26549, g17742)
--	g28115 = AND(g27354, g22759)
--	g31540 = AND(g29904, g23548)
--	g25087 = AND(g17307, g23489)
--	g32054 = AND(g10890, g30735)
--	g24475 = AND(g3831, g23139)
--	g7685 = AND(g4382, g4375)
--	g18264 = AND(g1263, g16000)
--	g18790 = AND(g6040, g15634)
--	g18137 = AND(g538, g17249)
--	I27513 = AND(g19984, g24089, g24090, g28034)
--	g18516 = AND(g2638, g15509)
--	g34337 = AND(g34095, g19881)
--	g24727 = AND(g13300, g23016)
--	g34171 = AND(g33925, g24360)
--	g16590 = AND(g5236, g14683)
--	g24222 = AND(g262, g22594)
--	g16986 = AND(g246, g13142)
--	g27303 = AND(g11996, g26681)
--	g11223 = AND(g8281, g8505)
--	g25043 = AND(g20733, g23447)
--	g32269 = AND(g31253, g20443)
--	g21853 = AND(g3917, g21070)
--	g28799 = AND(g21434, g26424, g25348, g27445)
--	g26079 = AND(g6199, g25060)
--	g34967 = AND(g34951, g23189)
--	g28813 = AND(g4104, g27038)
--	g29629 = AND(g28211, g19779)
--	g32341 = AND(g31472, g23610)
--	g31281 = AND(g30106, g27742)
--	g15870 = AND(g3231, g13948)
--	g26078 = AND(g5128, g25055)
--	g32156 = AND(g31639, g30018)
--	g25069 = AND(g23296, g20535)
--	g24703 = AND(g17592, g22369)
--	g31301 = AND(g30170, g27907)
--	g18209 = AND(g921, g15938)
--	g29628 = AND(g27924, g28648)
--	g33902 = AND(g33085, g13202)
--	g21836 = AND(g3805, g20453)
--	g31120 = AND(g1700, g29976)
--	g32180 = AND(g2791, g31638)
--	g23836 = AND(g4129, g19495)
--	g26086 = AND(g9672, g25255)
--	g28674 = AND(g27569, g20629)
--	g13321 = AND(g847, g11048)
--	g25068 = AND(g17574, g23477)
--	g25955 = AND(g24720, g19580)
--	g30919 = AND(g29898, g23286)
--	g18208 = AND(g930, g15938)
--	g16801 = AND(g5120, g14238)
--	g16735 = AND(g6235, g15027)
--	g23401 = AND(g7262, g21460)
--	g25879 = AND(g11135, g24683)
--	g24600 = AND(g22591, g19652)
--	g25970 = AND(g1792, g24991)
--	g31146 = AND(g12285, g30053)
--	g30010 = AND(g29035, g9274)
--	g30918 = AND(g8681, g29707)
--	g32335 = AND(g6199, g31566)
--	g11178 = AND(g6682, g7097, g6668, g10061)
--	g11740 = AND(g8769, g703)
--	g18542 = AND(g2787, g15277)
--	I18803 = AND(g13156, g11450, g6756)
--	g18453 = AND(g2315, g15224)
--	g29591 = AND(g28552, g11346)
--	g29785 = AND(g28332, g23248)
--	g31290 = AND(g29734, g23335)
--	g22114 = AND(g6565, g19277)
--	g26159 = AND(g2370, g25137)
--	g26125 = AND(g1894, g25117)
--	g21864 = AND(g3961, g21070)
--	g34079 = AND(g33703, g19532)
--	g22082 = AND(g6283, g19210)
--	g27390 = AND(g26549, g17504)
--	g18726 = AND(g4927, g16077)
--	g26977 = AND(g23032, g26261, g26424, g25550)
--	g30599 = AND(g18911, g29863)
--	g22107 = AND(g6411, g18833)
--	g30078 = AND(g28526, g20667)
--	g21749 = AND(g3155, g20785)
--	g26158 = AND(g2255, g25432)
--	g17725 = AND(g11547, g11592, g6789, I18716)
--	g26783 = AND(g25037, g21048)
--	I31287 = AND(g32870, g32871, g32872, g32873)
--	g18614 = AND(g3343, g17200)
--	g28692 = AND(g27578, g20661)
--	g28761 = AND(g21434, g26424, g25299, g27416)
--	g34078 = AND(g33699, g19531)
--	g18436 = AND(g2227, g18008)
--	g25967 = AND(g9373, g24986)
--	g30598 = AND(g18898, g29862)
--	g14585 = AND(g1141, g10905)
--	g29859 = AND(g28388, g23307)
--	I31307 = AND(g32898, g32899, g32900, g32901)
--	I31076 = AND(g30614, g31809, g32564, g32565)
--	g30086 = AND(g28536, g20704)
--	g21748 = AND(g15089, g20785)
--	g15707 = AND(g4082, g13506)
--	g15819 = AND(g3251, g14101)
--	g18607 = AND(g3139, g16987)
--	g34086 = AND(g20114, g33766, g9104)
--	g18320 = AND(g1616, g17873)
--	g24790 = AND(g7074, g23681)
--	g21276 = AND(g10157, g17625)
--	g21285 = AND(g7857, g16027)
--	g26295 = AND(g13070, g25266)
--	g29858 = AND(g28387, g23306)
--	g21704 = AND(g164, g20283)
--	g18274 = AND(g1311, g16031)
--	g22849 = AND(g1227, g19653)
--	g33366 = AND(g32268, g21010)
--	g27522 = AND(g26549, g17717)
--	g26823 = AND(g24401, g13106)
--	g15818 = AND(g3941, g14082)
--	g18530 = AND(g2715, g15277)
--	g25459 = AND(g6058, g23844, I24582)
--	g18593 = AND(g2999, g16349)
--	g18346 = AND(g1752, g17955)
--	g19716 = AND(g12100, g17121)
--	g21809 = AND(g3574, g20924)
--	g23254 = AND(g20056, g20110)
--	g28214 = AND(g27731, g26625)
--	g15111 = AND(g4281, g14454)
--	g22848 = AND(g19449, g19649)
--	g18122 = AND(g15052, g17015)
--	g23900 = AND(g1129, g19408)
--	g34322 = AND(g14188, g34174)
--	g14608 = AND(g12638, g12476, g12429, I16721)
--	g15978 = AND(g246, g14032)
--	g18565 = AND(g2852, g16349)
--	g26336 = AND(g10307, g25480)
--	g30125 = AND(g28581, g21056)
--	g18464 = AND(g2370, g15224)
--	g21808 = AND(g3570, g20924)
--	g29844 = AND(g28374, g23290)
--	g34532 = AND(g34314, g19710)
--	g15590 = AND(g3139, g13530)
--	g29367 = AND(g8575, g28325)
--	g28539 = AND(g27187, g12762)
--	g10921 = AND(g1548, g8685)
--	g27483 = AND(g26488, g17642)
--	g30158 = AND(g28613, g21274)
--	g33403 = AND(g32352, g21396)
--	g24422 = AND(g4771, g22896)
--	I31341 = AND(g31710, g31856, g32947, g32948)
--	g32278 = AND(g2811, g30572)
--	g27553 = AND(g26293, g23353)
--	g18641 = AND(g3841, g17096)
--	g18797 = AND(g6173, g15348)
--	g25079 = AND(g21011, g23483)
--	I31156 = AND(g31070, g31823, g32680, g32681)
--	g18292 = AND(g1472, g16449)
--	g16706 = AND(g6621, g14868)
--	g31226 = AND(g30282, g25218)
--	g32286 = AND(g31658, g29312)
--	g34561 = AND(g34368, g17410)
--	g16597 = AND(g6263, g15021)
--	g18153 = AND(g626, g17533)
--	g27326 = AND(g12048, g26731)
--	g25078 = AND(g23298, g20538)
--	g31481 = AND(g29768, g23417)
--	g32039 = AND(g31476, g20070)
--	g33715 = AND(g33135, g19416)
--	g32306 = AND(g31289, g23499)
--	g34295 = AND(g34057, g19370)
--	g33481 = AND(g32607, I31101, I31102)
--	g22135 = AND(g6657, g19277)
--	g27536 = AND(g26519, g17738)
--	g18409 = AND(g2084, g15373)
--	g27040 = AND(g7812, g6565, g6573, g26226)
--	g25086 = AND(g13941, g23488)
--	g21733 = AND(g3034, g20330)
--	g10674 = AND(g6841, g10200, g2130)
--	g18136 = AND(g550, g17249)
--	g18408 = AND(g2070, g15373)
--	g18635 = AND(g3808, g17096)
--	g24726 = AND(g15965, g23015)
--	g27252 = AND(g26733, g26703)
--	g24913 = AND(g4821, g23908)
--	g21874 = AND(g4112, g19801)
--	g25817 = AND(g24807, g21163)
--	g32187 = AND(g30672, g25287)
--	g26289 = AND(g2551, g25400)
--	g24436 = AND(g3125, g23067)
--	g25159 = AND(g4907, g22908)
--	g10732 = AND(g6850, g2697, g2689)
--	g22049 = AND(g6082, g21611)
--	g25125 = AND(g20187, g23520)
--	g27564 = AND(g26305, g23378)
--	g25901 = AND(g24853, g16290)
--	g26023 = AND(g9528, g25036)
--	I31131 = AND(g31542, g31819, g32643, g32644)
--	g34966 = AND(g34950, g23170)
--	g31490 = AND(g29786, g23429)
--	g10934 = AND(g9197, g7918)
--	g24607 = AND(g5817, g23666)
--	g25977 = AND(g25236, g20875)
--	g26288 = AND(g2259, g25309)
--	g33490 = AND(g32672, I31146, I31147)
--	g19681 = AND(g5835, g17014)
--	g24320 = AND(g6973, g22228)
--	g28235 = AND(g9467, g27592)
--	g26571 = AND(g10472, g24386)
--	g23166 = AND(g13959, g19979)
--	g23009 = AND(g20196, g14219)
--	g22048 = AND(g6052, g21611)
--	g26308 = AND(g6961, g25289)
--	g29203 = AND(g24095, I27513, I27514)
--	g18164 = AND(g699, g17433)
--	g28683 = AND(g27876, g20649)
--	g32143 = AND(g31646, g29967)
--	g31784 = AND(g30176, g24003)
--	g34364 = AND(g34048, g24366)
--	g33784 = AND(g33107, g20531)
--	g31376 = AND(g24952, g29814)
--	g31297 = AND(g30144, g27837)
--	g27183 = AND(g26055, g16658)
--	g33376 = AND(g32294, g21268)
--	g27673 = AND(g25769, g23541)
--	g22004 = AND(g5742, g21562)
--	g23008 = AND(g1570, g19783)
--	g33889 = AND(g33303, g20641)
--	g11123 = AND(g5644, g7028, g5630, g9864)
--	g24464 = AND(g3480, g23112)
--	I24027 = AND(g3029, g3034, g8426)
--	g16885 = AND(g6605, g14950)
--	g32169 = AND(g31014, g23046)
--	g18575 = AND(g2878, g16349)
--	g18474 = AND(g2287, g15224)
--	g29902 = AND(g28430, g23377)
--	g30289 = AND(g28884, g24000)
--	g29377 = AND(g28132, g19387)
--	g13807 = AND(g4504, g10606)
--	g18711 = AND(g15136, g15915)
--	g32168 = AND(g30597, g25185)
--	g32410 = AND(g4933, g30997)
--	g28991 = AND(g14438, g25209, g26424, g27469)
--	g13974 = AND(g6243, g12578)
--	g18327 = AND(g1636, g17873)
--	g24797 = AND(g22872, g19960)
--	g30023 = AND(g28508, g20570)
--	g21712 = AND(g294, g20283)
--	I24482 = AND(g9364, g9607, g5057)
--	g18109 = AND(g437, g17015)
--	g27508 = AND(g26549, g17684)
--	g16763 = AND(g6239, g14937)
--	g27634 = AND(g26805, g26793)
--	g34309 = AND(g13947, g34147)
--	g21914 = AND(g5077, g21468)
--	g24292 = AND(g4443, g22550)
--	g30224 = AND(g28704, g23896)
--	g18537 = AND(g6856, g15277)
--	I24710 = AND(g24071, g24072, g24073, g24074)
--	g34224 = AND(g33736, g22670)
--	g30308 = AND(g29178, g7004, g5297)
--	g22106 = AND(g6497, g18833)
--	I24552 = AND(g9733, g9316, g5747)
--	g29645 = AND(g1714, g29018)
--	I24003 = AND(g8097, g8334, g3045)
--	g17613 = AND(g11547, g11592, g11640, I18568)
--	g34571 = AND(g27225, g34299)
--	g18108 = AND(g433, g17015)
--	g14207 = AND(g8639, g11793)
--	g21907 = AND(g5033, g21468)
--	I31286 = AND(g30825, g31846, g32868, g32869)
--	I13862 = AND(g7232, g7219, g7258)
--	g15077 = AND(g2138, g12955)
--	g24409 = AND(g3484, g23112)
--	g25966 = AND(g9364, g24985)
--	I31306 = AND(g30614, g31850, g32896, g32897)
--	g13265 = AND(g9018, g11493)
--	g18283 = AND(g1384, g16136)
--	g15706 = AND(g13296, g13484)
--	g18606 = AND(g3133, g16987)
--	g18492 = AND(g2523, g15426)
--	g18303 = AND(g1536, g16489)
--	g24408 = AND(g23989, g18946)
--	g24635 = AND(g19874, g22883)
--	g34495 = AND(g34274, g19365)
--	g22033 = AND(g5925, g19147)
--	g27213 = AND(g26026, g16721)
--	g18750 = AND(g15145, g17847)
--	g31520 = AND(g29879, g23507)
--	I31187 = AND(g32726, g32727, g32728, g32729)
--	g33520 = AND(g32888, I31296, I31297)
--	g18982 = AND(g3835, g16159)
--	g18381 = AND(g1882, g15171)
--	g34687 = AND(g14181, g34543)
--	g21941 = AND(g5232, g18997)
--	g26842 = AND(g2894, g24522)
--	I27429 = AND(g25562, g26424, g22698)
--	g27452 = AND(g26400, g17600)
--	g21382 = AND(g10086, g17625)
--	g29632 = AND(g28899, g22417)
--	g31211 = AND(g10156, g30102)
--	g26195 = AND(g25357, g6856, g11709, g7558)
--	g34752 = AND(g34675, g19544)
--	g23675 = AND(g19050, g9104)
--	g18174 = AND(g739, g17328)
--	g27311 = AND(g12431, g26693)
--	g18796 = AND(g6167, g15348)
--	g28725 = AND(g27596, g20779)
--	g32084 = AND(g10948, g30825)
--	g32110 = AND(g31639, g29921)
--	g16596 = AND(g5941, g14892)
--	g28114 = AND(g25869, g27051)
--	g25571 = AND(I24694, I24695)
--	g33860 = AND(g33270, g20501)
--	g32321 = AND(g27613, g31376)
--	g16243 = AND(g6483, g14275)
--	g29661 = AND(g1687, g29015)
--	g29547 = AND(g1748, g28857)
--	g29895 = AND(g2495, g29170)
--	g28107 = AND(g27970, g18874)
--	g10683 = AND(g7289, g4438)
--	g32179 = AND(g31748, g27907)
--	g21935 = AND(g5196, g18997)
--	g18390 = AND(g1978, g15171)
--	g31497 = AND(g20041, g29930)
--	g33497 = AND(g32723, I31181, I31182)
--	g20109 = AND(g17954, g17616)
--	g24327 = AND(g4549, g22228)
--	g21883 = AND(g4141, g19801)
--	g32178 = AND(g31747, g27886)
--	g15876 = AND(g13512, g13223)
--	g24537 = AND(g22626, g10851)
--	g11116 = AND(g9960, g6466)
--	g20108 = AND(g15508, g11048)
--	g34842 = AND(g34762, g20168)
--	g18192 = AND(g817, g17821)
--	g22012 = AND(g5752, g21562)
--	g26544 = AND(g7446, g24357)
--	I27504 = AND(g24077, g24078, g24079, g24080)
--	I18620 = AND(g13156, g11450, g11498)
--	g25816 = AND(g8164, g24604)
--	g33700 = AND(g33148, g11012)
--	g33126 = AND(g9044, g32201)
--	g31987 = AND(g31767, g22198)
--	g29551 = AND(g2173, g28867)
--	g29572 = AND(g1620, g28885)
--	g26713 = AND(g25447, g20714)
--	I31217 = AND(g32768, g32769, g32770, g32771)
--	g34489 = AND(g34421, g19068)
--	g24283 = AND(g4411, g22550)
--	g18522 = AND(g2671, g15509)
--	g27350 = AND(g10217, g26803)
--	g18663 = AND(g4311, g17367)
--	g24606 = AND(g5489, g23630)
--	g25976 = AND(g9443, g25000)
--	g24303 = AND(g4369, g22228)
--	g16670 = AND(g5953, g14999)
--	g27820 = AND(g7670, g25932)
--	g34525 = AND(g34297, g19528)
--	g28141 = AND(g10831, g11797, g11261, g27163)
--	g34488 = AND(g34417, g18988)
--	g28652 = AND(g27282, g10288)
--	g13493 = AND(g9880, g11866)
--	g25374 = AND(g5366, g23789, I24527)
--	g31943 = AND(g4717, g30614)
--	I24505 = AND(g9607, g9229, g5057)
--	g21729 = AND(g3021, g20330)
--	g26610 = AND(g14198, g24405)
--	g33339 = AND(g32221, g20634)
--	g33943 = AND(g33384, g21609)
--	g31296 = AND(g30119, g27779)
--	g34558 = AND(g34353, g20578)
--	g16734 = AND(g5961, g14735)
--	g23577 = AND(g19444, g13033)
--	g18483 = AND(g2453, g15426)
--	g24750 = AND(g17662, g22472)
--	g32334 = AND(g31375, g23568)
--	g21728 = AND(g3010, g20330)
--	g33338 = AND(g32220, g20633)
--	g28263 = AND(g23747, g27711)
--	g16930 = AND(g239, g13132)
--	g23439 = AND(g13771, g20452)
--	g11035 = AND(g5441, g9800)
--	g18553 = AND(g2827, g15277)
--	g13035 = AND(g8497, g11033)
--	g26270 = AND(g1700, g25275)
--	g31969 = AND(g31189, g22139)
--	g29784 = AND(g28331, g23247)
--	g26124 = AND(g1811, g25116)
--	g22920 = AND(g19764, g19719)
--	g16667 = AND(g5268, g14659)
--	g20174 = AND(g5503, g17754)
--	g29376 = AND(g14002, g28504)
--	g27413 = AND(g26576, g17530)
--	g34865 = AND(g16540, g34836)
--	g16965 = AND(g269, g13140)
--	g18949 = AND(g10183, g17625)
--	g31968 = AND(g31757, g22168)
--	g18326 = AND(g1664, g17873)
--	g24796 = AND(g7097, g23714)
--	g11142 = AND(g6381, g10207)
--	g27691 = AND(g25778, g23609)
--	g17724 = AND(g11547, g11592, g11640, I18713)
--	g29354 = AND(g4961, g28421)
--	I27533 = AND(g21143, g24125, g24126, g24127)
--	g18536 = AND(g2748, g15277)
--	g23349 = AND(g13662, g20182)
--	g22121 = AND(g6593, g19277)
--	g29888 = AND(g28418, g23352)
--	g33855 = AND(g33265, g20441)
--	g14206 = AND(g8655, g11790)
--	g21906 = AND(g5022, g21468)
--	g18702 = AND(g15133, g16856)
--	g21348 = AND(g10121, g17625)
--	g18757 = AND(g5352, g15595)
--	g31527 = AND(g7553, g29343)
--	g23083 = AND(g16076, g19878)
--	g23348 = AND(g15570, g21393)
--	g15076 = AND(g2130, g12955)
--	g33870 = AND(g33280, g20545)
--	g33411 = AND(g32361, g21410)
--	g33527 = AND(g32939, I31331, I31332)
--	g26294 = AND(g4245, g25230)
--	I31321 = AND(g31376, g31852, g32919, g32920)
--	g16619 = AND(g6629, g14947)
--	g30042 = AND(g29142, g12601)
--	g18252 = AND(g990, g16897)
--	g18621 = AND(g3476, g17062)
--	g25559 = AND(g13004, g22649)
--	g30255 = AND(g28748, g23946)
--	g25488 = AND(g6404, g23865, I24603)
--	g28833 = AND(g21434, g26424, g25388, g27469)
--	g16618 = AND(g6609, g15039)
--	g34679 = AND(g14093, g34539)
--	g18564 = AND(g2844, g16349)
--	g30188 = AND(g28644, g23841)
--	g24192 = AND(g311, g22722)
--	g30124 = AND(g28580, g21055)
--	g16279 = AND(g4512, g14424)
--	g34678 = AND(g34490, g19431)
--	g27020 = AND(g4601, g25852)
--	g31503 = AND(g20041, g29945)
--	I18716 = AND(g13156, g11450, g6756)
--	I31186 = AND(g31376, g31828, g32724, g32725)
--	g33503 = AND(g32765, I31211, I31212)
--	g24663 = AND(g16621, g22974)
--	g33867 = AND(g33277, g20529)
--	g17682 = AND(g9742, g14637)
--	g34686 = AND(g34494, g19494)
--	g13523 = AND(g7046, g12246)
--	g18183 = AND(g781, g17328)
--	g18673 = AND(g4643, g15758)
--	g25865 = AND(g25545, g18991)
--	g26218 = AND(g25357, g6856, g7586, g11686)
--	g18397 = AND(g2004, g15373)
--	g30030 = AND(g29198, g12347)
--	g30267 = AND(g28776, g23967)
--	g34093 = AND(g20114, g33755, g9104)
--	g33450 = AND(g32266, g29737)
--	g22760 = AND(g9360, g20237)
--	g22134 = AND(g6653, g19277)
--	g27113 = AND(g25997, g16522)
--	g32242 = AND(g31245, g20324)
--	g18509 = AND(g2587, g15509)
--	g22029 = AND(g5901, g19147)
--	g31707 = AND(g30081, g23886)
--	g34065 = AND(g33813, g23148)
--	g33819 = AND(g23088, g33176, g9104)
--	g33707 = AND(g33174, g13346)
--	g18933 = AND(g16237, g13597)
--	g33910 = AND(g33134, g7836)
--	g24553 = AND(g22983, g19539)
--	g26160 = AND(g2453, g25138)
--	g28273 = AND(g27927, g23729)
--	g7696 = AND(g2955, g2950)
--	g18508 = AND(g2606, g15509)
--	g22028 = AND(g5893, g19147)
--	g27302 = AND(g1848, g26680)
--	g18634 = AND(g3813, g17096)
--	g21333 = AND(g1300, g15740)
--	g23415 = AND(g20077, g20320)
--	g27357 = AND(g26400, g17414)
--	g25042 = AND(g23262, g20496)
--	g31496 = AND(g2338, g30312)
--	g33818 = AND(g33236, g20113)
--	g24949 = AND(g23796, g20751)
--	g33496 = AND(g32714, I31176, I31177)
--	g19461 = AND(g11708, g16846)
--	g27105 = AND(g26026, g16511)
--	g24326 = AND(g4552, g22228)
--	g30219 = AND(g28698, g23887)
--	g17134 = AND(g5619, g14851)
--	g21852 = AND(g3909, g21070)
--	g15839 = AND(g3929, g13990)
--	g34875 = AND(g34836, g20073)
--	g28812 = AND(g26972, g13037)
--	g33111 = AND(g24005, g32421)
--	g34219 = AND(g33736, g22942)
--	g31070 = AND(g29814, g25985)
--	g19145 = AND(g8450, g16200)
--	g24536 = AND(g19516, g22635)
--	g29860 = AND(g28389, g23312)
--	g17506 = AND(g9744, g14505)
--	g25124 = AND(g4917, g22908)
--	g15694 = AND(g457, g13437)
--	g15838 = AND(g3602, g14133)
--	g21963 = AND(g5436, g21514)
--	g24702 = AND(g17464, g22342)
--	g34218 = AND(g33744, g22670)
--	g24757 = AND(g7004, g23563)
--	g31986 = AND(g31766, g22197)
--	g19736 = AND(g12136, g17136)
--	g24904 = AND(g11761, g23279)
--	g28234 = AND(g27877, g26686)
--	g32293 = AND(g2827, g30593)
--	I31216 = AND(g30937, g31834, g32766, g32767)
--	g25939 = AND(g24583, g19490)
--	g26277 = AND(g2547, g25400)
--	g18213 = AND(g952, g15979)
--	g32265 = AND(g2799, g30567)
--	g25030 = AND(g23251, g20432)
--	g25938 = AND(g8997, g24953)
--	g25093 = AND(g12831, g23493)
--	g31067 = AND(g29484, g22868)
--	g24564 = AND(g23198, g21163)
--	g29625 = AND(g28514, g14226)
--	g29987 = AND(g29197, g26424, g22763)
--	g19393 = AND(g691, g16325)
--	g16884 = AND(g6159, g14321)
--	g18574 = AND(g2882, g16349)
--	g23484 = AND(g20160, g20541)
--	g18452 = AND(g2311, g15224)
--	g18205 = AND(g904, g15938)
--	g31150 = AND(g1682, g30063)
--	g23554 = AND(g20390, g13024)
--	I31117 = AND(g32624, g32625, g32626, g32627)
--	g18311 = AND(g1554, g16931)
--	g33801 = AND(g33437, g25327)
--	g24673 = AND(g22659, g19748)
--	g33735 = AND(g33118, g19553)
--	g33877 = AND(g33287, g20563)
--	I24582 = AND(g9809, g9397, g6093)
--	g30915 = AND(g29886, g24778)
--	g29943 = AND(g2165, g28765)
--	g34470 = AND(g7834, g34325)
--	g16666 = AND(g5200, g14794)
--	g25875 = AND(g8390, g24809)
--	g31019 = AND(g29481, g22856)
--	I18765 = AND(g13156, g11450, g11498)
--	g29644 = AND(g28216, g19794)
--	g29338 = AND(g29145, g22181)
--	g30277 = AND(g28817, g23987)
--	g13063 = AND(g8567, g10808)
--	g31018 = AND(g29480, g22855)
--	g32014 = AND(g8715, g30673)
--	g29969 = AND(g28121, g20509)
--	g30075 = AND(g28525, g20662)
--	g26155 = AND(g1945, g25134)
--	g14221 = AND(g8686, g11823)
--	g21921 = AND(g5109, g21468)
--	g26822 = AND(g24841, g13116)
--	I31242 = AND(g32805, g32806, g32807, g32808)
--	g16486 = AND(g6772, g11592, g6789, I17692)
--	g18592 = AND(g2994, g16349)
--	g23921 = AND(g19379, g4146)
--	g18756 = AND(g5348, g15595)
--	g34075 = AND(g33692, g19517)
--	g31526 = AND(g22521, g29342)
--	g24634 = AND(g22634, g19685)
--	g30595 = AND(g18911, g29847)
--	g33526 = AND(g32932, I31326, I31327)
--	g24872 = AND(g23088, g9104)
--	g29968 = AND(g2433, g28843)
--	g21745 = AND(g3017, g20330)
--	g18780 = AND(g5827, g18065)
--	g12027 = AND(g9499, g9729)
--	g14613 = AND(g10602, g10585)
--	g27249 = AND(g25929, g19678)
--	g21799 = AND(g3530, g20924)
--	g29855 = AND(g2287, g29093)
--	g17770 = AND(g7863, g13189)
--	g21813 = AND(g3590, g20924)
--	g23799 = AND(g14911, g21279)
--	g27482 = AND(g26488, g17641)
--	g15815 = AND(g3594, g14075)
--	g28541 = AND(g27403, g20274)
--	g10947 = AND(g9200, g1430)
--	g18350 = AND(g1779, g17955)
--	I24603 = AND(g9892, g9467, g6439)
--	g33402 = AND(g32351, g21395)
--	g29870 = AND(g2421, g29130)
--	g29527 = AND(g28945, g22432)
--	g27710 = AND(g26422, g20904)
--	g21798 = AND(g3522, g20924)
--	g34782 = AND(g34711, g33888)
--	I27529 = AND(g28038, g24121, g24122, g24123)
--	g18820 = AND(g15166, g15563)
--	g26853 = AND(g94, g24533)
--	g28789 = AND(g21434, g26424, g25340, g27440)
--	g21973 = AND(g5511, g19074)
--	g32116 = AND(g31658, g29929)
--	g27204 = AND(g26026, g16689)
--	g33866 = AND(g33276, g20528)
--	g22899 = AND(g19486, g19695)
--	g21805 = AND(g3550, g20924)
--	g22990 = AND(g19555, g19760)
--	I27528 = AND(g20998, g24118, g24119, g24120)
--	g18152 = AND(g613, g17533)
--	g25915 = AND(g24926, g9602)
--	g32041 = AND(g13913, g31262)
--	g18396 = AND(g2008, g15373)
--	g22633 = AND(g19359, g19479)
--	g17767 = AND(g6772, g11592, g6789, I18765)
--	g18731 = AND(g15140, g16861)
--	g30266 = AND(g28775, g23966)
--	g28535 = AND(g11981, g27088)
--	g15937 = AND(g11950, g14387)
--	g25201 = AND(g12346, g23665)
--	g22191 = AND(g8119, g19875)
--	g16179 = AND(g6187, g14321)
--	g29867 = AND(g1996, g29117)
--	g29894 = AND(g2070, g29169)
--	g19069 = AND(g8397, g16186)
--	g21732 = AND(g3004, g20330)
--	g16531 = AND(g5232, g14656)
--	g13542 = AND(g10053, g11927)
--	g21934 = AND(g5220, g18997)
--	g18413 = AND(g2089, g15373)
--	g24912 = AND(g23687, g20682)
--	g26119 = AND(g11944, g25109)
--	g24311 = AND(g4498, g22228)
--	g16178 = AND(g5845, g14297)
--	g18691 = AND(g4727, g16053)
--	g15884 = AND(g3901, g14113)
--	g33689 = AND(g33144, g11006)
--	g32340 = AND(g31468, g23585)
--	g29581 = AND(g28462, g11796)
--	g32035 = AND(g4176, g30937)
--	g31280 = AND(g29717, g23305)
--	g17191 = AND(g1384, g13242)
--	g17719 = AND(g9818, g14675)
--	g21761 = AND(g3215, g20785)
--	g29315 = AND(g29188, g7051, g5990)
--	g27999 = AND(g23032, g26200, g26424, g25529)
--	g26864 = AND(g2907, g24548)
--	g26022 = AND(g25271, g20751)
--	g13436 = AND(g9721, g11811)
--	g18405 = AND(g2040, g15373)
--	g31300 = AND(g30148, g27858)
--	g30167 = AND(g28622, g23793)
--	g30194 = AND(g28651, g23849)
--	g30589 = AND(g18898, g29811)
--	I24690 = AND(g24043, g24044, g24045, g24046)
--	I24549 = AND(g5385, g5390, g9792)
--	g26749 = AND(g24494, g23578)
--	g27090 = AND(g25997, g16423)
--	g29202 = AND(g24088, I27508, I27509)
--	g25782 = AND(g2936, g24571)
--	g32142 = AND(g31616, g29965)
--	g13320 = AND(g417, g11048)
--	g26313 = AND(g12645, g25326)
--	g28291 = AND(g7411, g2070, g27469)
--	g29979 = AND(g23655, g28991)
--	g34588 = AND(g26082, g34323)
--	g22861 = AND(g19792, g19670)
--	g27651 = AND(g22448, g25781)
--	g34524 = AND(g9083, g34359)
--	g33102 = AND(g32399, g18978)
--	I31007 = AND(g32466, g32467, g32468, g32469)
--	g26276 = AND(g2461, g25476)
--	g26285 = AND(g1834, g25300)
--	g34401 = AND(g34199, g21383)
--	g34477 = AND(g26344, g34328)
--	g22045 = AND(g6069, g21611)
--	g18583 = AND(g2936, g16349)
--	g29590 = AND(g2625, g28615)
--	g34119 = AND(g20516, g9104, g33755)
--	g26254 = AND(g2413, g25349)
--	g31066 = AND(g29483, g22865)
--	g31231 = AND(g30290, g25239)
--	g29986 = AND(g28468, g23473)
--	g22099 = AND(g6462, g18833)
--	g27932 = AND(g25944, g19369)
--	g27331 = AND(g10177, g26754)
--	g30118 = AND(g28574, g21050)
--	g24820 = AND(g13944, g23978)
--	g26808 = AND(g25521, g21185)
--	g16762 = AND(g5901, g14930)
--	g20152 = AND(g11545, g16727)
--	g22534 = AND(g8766, g21389)
--	g29384 = AND(g26424, g22763, g28179)
--	g22098 = AND(g6459, g18833)
--	g32193 = AND(g30732, g25410)
--	I31116 = AND(g31154, g31816, g32622, g32623)
--	g24846 = AND(g3361, g23555, I24018)
--	g26101 = AND(g1760, g25098)
--	g33876 = AND(g33286, g20562)
--	g33885 = AND(g33296, g20609)
--	g26177 = AND(g2079, g25154)
--	g18113 = AND(g405, g17015)
--	g18787 = AND(g15158, g15634)
--	g32165 = AND(g31669, g27742)
--	g24731 = AND(g6519, g23733)
--	I31041 = AND(g31566, g31803, g32513, g32514)
--	g18282 = AND(g1379, g16136)
--	g34748 = AND(g34672, g19529)
--	g27505 = AND(g26519, g17681)
--	g27404 = AND(g26400, g17518)
--	g31763 = AND(g30127, g23965)
--	g18302 = AND(g1514, g16489)
--	g33511 = AND(g32823, I31251, I31252)
--	g15084 = AND(g2710, g12983)
--	g18357 = AND(g1816, g17955)
--	g19545 = AND(g3147, g16769)
--	g29877 = AND(g28405, g23340)
--	g15110 = AND(g4245, g14454)
--	g18105 = AND(g417, g17015)
--	g10724 = AND(g3689, g8728)
--	g22032 = AND(g5921, g19147)
--	g30254 = AND(g28747, g23944)
--	g18743 = AND(g5115, g17847)
--	g27212 = AND(g25997, g16717)
--	g10829 = AND(g7289, g4375)
--	I31237 = AND(g32798, g32799, g32800, g32801)
--	g21771 = AND(g3255, g20785)
--	g10828 = AND(g6888, g7640)
--	g18640 = AND(g3835, g17096)
--	g18769 = AND(g15151, g18062)
--	g22061 = AND(g6065, g21611)
--	g30101 = AND(g28551, g20780)
--	g30177 = AND(g28631, g23814)
--	g29526 = AND(g28938, g22384)
--	g17140 = AND(g8616, g12968)
--	g26630 = AND(g7592, g24419)
--	g34560 = AND(g34366, g17366)
--	g18768 = AND(g5503, g17929)
--	g18803 = AND(g15161, g15480)
--	g31480 = AND(g1644, g30296)
--	I31142 = AND(g32661, g32662, g32663, g32664)
--	g33480 = AND(g32600, I31096, I31097)
--	g24929 = AND(g23751, g20875)
--	g22871 = AND(g9523, g20871)
--	g26166 = AND(g25357, g11724, g11709, g7558)
--	g27723 = AND(g26512, g21049)
--	g15654 = AND(g3845, g13584)
--	g31314 = AND(g30183, g27937)
--	g28240 = AND(g27356, g17239)
--	g27149 = AND(g25997, g16623)
--	g30064 = AND(g28517, g20630)
--	g17766 = AND(g6772, g11592, g11640, I18762)
--	g27433 = AND(g26519, g17583)
--	g27387 = AND(g26488, g17499)
--	g15936 = AND(g475, g13999)
--	g25285 = AND(g22152, g13061)
--	g29866 = AND(g1906, g29116)
--	g27148 = AND(g25997, g16622)
--	g21882 = AND(g4057, g19801)
--	g21991 = AND(g5595, g19074)
--	g26485 = AND(g24968, g10502)
--	g23991 = AND(g19209, g21428)
--	g27097 = AND(g25867, g22526)
--	g33721 = AND(g33163, g19440)
--	g19656 = AND(g2807, g15844)
--	g27104 = AND(g25997, g16510)
--	g16751 = AND(g13155, g13065)
--	g16807 = AND(g6585, g14978)
--	g27646 = AND(g13094, g25773)
--	g25900 = AND(g24390, g19368)
--	g34874 = AND(g34833, g20060)
--	g23407 = AND(g9295, g20273)
--	g33243 = AND(g32124, g19947)
--	g28563 = AND(g11981, g27100)
--	g25466 = AND(g23574, g21346)
--	g19680 = AND(g12028, g17013)
--	g33431 = AND(g32364, g32377)
--	g16639 = AND(g6291, g14974)
--	g26712 = AND(g24508, g24463)
--	I17741 = AND(g14988, g11450, g11498)
--	g18662 = AND(g15126, g17367)
--	g32175 = AND(g31709, g27858)
--	g30166 = AND(g28621, g23792)
--	g30009 = AND(g29034, g10518)
--	g24302 = AND(g15124, g22228)
--	g16638 = AND(g6271, g14773)
--	g33269 = AND(g31970, g15582)
--	g34665 = AND(g34583, g19067)
--	g22472 = AND(g7753, g9285, g21289)
--	g18890 = AND(g10158, g17625)
--	g13492 = AND(g9856, g11865)
--	g27369 = AND(g25894, g25324)
--	g24743 = AND(g22708, g19789)
--	g30008 = AND(g29191, g12297)
--	g18249 = AND(g1216, g16897)
--	g33942 = AND(g33383, g21608)
--	g33341 = AND(g32223, g20640)
--	g18482 = AND(g2472, g15426)
--	g14506 = AND(g1430, g10755)
--	g29688 = AND(g2509, g28713)
--	I31006 = AND(g31376, g31796, g32464, g32465)
--	g29624 = AND(g28491, g8070)
--	g14028 = AND(g8673, g11797)
--	g18248 = AND(g15067, g16897)
--	g16841 = AND(g5913, g14858)
--	g18710 = AND(g15135, g17302)
--	g34476 = AND(g34399, g18891)
--	g34485 = AND(g34411, g18952)
--	g18552 = AND(g2815, g15277)
--	g24640 = AND(g6509, g23733)
--	g24769 = AND(g19619, g23058)
--	g19631 = AND(g1484, g16093)
--	g18204 = AND(g914, g15938)
--	I31222 = AND(g32775, g32776, g32777, g32778)
--	g27412 = AND(g26576, g17529)
--	g34555 = AND(g34349, g20512)
--	g18779 = AND(g5821, g18065)
--	g22071 = AND(g6251, g19210)
--	g24803 = AND(g22901, g20005)
--	g33734 = AND(g7806, g33136, I31593)
--	g30914 = AND(g29873, g20887)
--	g21759 = AND(g3199, g20785)
--	g15117 = AND(g4300, g14454)
--	g23725 = AND(g14772, g21138)
--	g18778 = AND(g5817, g18065)
--	g25874 = AND(g11118, g24665)
--	g27229 = AND(g26055, g16774)
--	g31993 = AND(g31774, g22214)
--	g21758 = AND(g3191, g20785)
--	g26176 = AND(g1964, g25467)
--	g26092 = AND(g9766, g25083)
--	g18786 = AND(g15156, g15345)
--	g27228 = AND(g26055, g16773)
--	g24881 = AND(g3050, g23211, I24048)
--	I31347 = AND(g32956, g32957, g32958, g32959)
--	g22859 = AND(g9456, g20734)
--	g26154 = AND(g1830, g25426)
--	g30239 = AND(g28728, g23923)
--	g17785 = AND(g13341, g10762)
--	g25166 = AND(g17506, g23571)
--	g31131 = AND(g2393, g30020)
--	g18647 = AND(g4040, g17271)
--	g34074 = AND(g33685, g19498)
--	g30594 = AND(g18898, g29846)
--	g18356 = AND(g1802, g17955)
--	g29876 = AND(g28404, g23339)
--	g29885 = AND(g28416, g23350)
--	g21744 = AND(g3103, g20330)
--	g30238 = AND(g28727, g23922)
--	g34567 = AND(g34377, g17491)
--	I31600 = AND(g31009, g8400, g7809)
--	g28440 = AND(g27274, g20059)
--	g18826 = AND(g7097, g15680)
--	g18380 = AND(g1926, g15171)
--	g19571 = AND(g3498, g16812)
--	g33487 = AND(g32649, I31131, I31132)
--	g22172 = AND(g8064, g19857)
--	g29854 = AND(g2197, g29092)
--	g21849 = AND(g3889, g21070)
--	g21940 = AND(g5228, g18997)
--	I31236 = AND(g30735, g31837, g32796, g32797)
--	g15814 = AND(g3574, g13920)
--	g31502 = AND(g2472, g29311)
--	g28573 = AND(g7349, g27059)
--	g25485 = AND(g6098, g22220, I24600)
--	g33502 = AND(g32758, I31206, I31207)
--	g29511 = AND(g1736, g28783)
--	g31210 = AND(g2509, g30100)
--	I31351 = AND(g30937, g31858, g32961, g32962)
--	g18233 = AND(g1094, g16326)
--	g28247 = AND(g27147, g19675)
--	g21848 = AND(g3913, g21070)
--	g15807 = AND(g3570, g13898)
--	g18182 = AND(g776, g17328)
--	g27310 = AND(g26574, g23059)
--	g18651 = AND(g15102, g16249)
--	g18672 = AND(g15127, g15758)
--	g34382 = AND(g34167, g20618)
--	g30185 = AND(g28640, g23838)
--	g34519 = AND(g34293, g19504)
--	g17151 = AND(g8659, g12996)
--	g21804 = AND(g3542, g20924)
--	g34185 = AND(g33702, g24389)
--	g27627 = AND(g13266, g25790)
--	g25570 = AND(I24689, I24690)
--	g27959 = AND(g25948, g19374)
--	g28612 = AND(g27524, g20539)
--	g34092 = AND(g33750, g9104, g18957)
--	g30154 = AND(g28611, g23769)
--	g28324 = AND(g9875, g27687)
--	g24482 = AND(g6875, g23055)
--	g31278 = AND(g29716, g23302)
--	g34518 = AND(g34292, g19503)
--	g32274 = AND(g31256, g20447)
--	g27050 = AND(g25789, g22338)
--	g27958 = AND(g25950, g22449)
--	g25907 = AND(g24799, g22519)
--	g24710 = AND(g22679, g19771)
--	g27378 = AND(g26089, g20052)
--	I31137 = AND(g32654, g32655, g32656, g32657)
--	g18331 = AND(g1682, g17873)
--	I27364 = AND(g25541, g26424, g22698)
--	g24552 = AND(g22487, g19538)
--	g33469 = AND(g32519, I31041, I31042)
--	g28251 = AND(g27826, g23662)
--	g30935 = AND(g8808, g29745)
--	g28272 = AND(g27721, g26548)
--	g31286 = AND(g30159, g27858)
--	g32122 = AND(g31646, g29944)
--	g18513 = AND(g2575, g15509)
--	g21332 = AND(g996, g15739)
--	g18449 = AND(g12852, g15224)
--	I26972 = AND(g25011, g26424, g22698)
--	g27386 = AND(g26488, g17498)
--	g19752 = AND(g2771, g15864)
--	g33468 = AND(g32512, I31036, I31037)
--	g15841 = AND(g4273, g13868)
--	g25567 = AND(I24674, I24675)
--	g27096 = AND(g26026, g16475)
--	g18448 = AND(g2153, g18008)
--	g29550 = AND(g28990, g22457)
--	g32034 = AND(g14124, g31239)
--	g25238 = AND(g12466, g23732)
--	g16806 = AND(g6247, g14971)
--	g29314 = AND(g29005, g22144)
--	g22059 = AND(g6148, g21611)
--	g21962 = AND(g5428, g21514)
--	g18505 = AND(g2583, g15509)
--	g21361 = AND(g7869, g16066)
--	g22025 = AND(g5905, g19147)
--	g18404 = AND(g2066, g15373)
--	g24786 = AND(g661, g23654)
--	g33815 = AND(g33449, g12911)
--	g32292 = AND(g31269, g20530)
--	g10898 = AND(g3706, g9100)
--	g18717 = AND(g4849, g15915)
--	g22058 = AND(g6098, g21611)
--	g31187 = AND(g10118, g30090)
--	g32153 = AND(g31646, g29999)
--	g24647 = AND(g19903, g22907)
--	g33677 = AND(g33443, g31937)
--	g31975 = AND(g31761, g22177)
--	g13252 = AND(g11561, g11511, g11469, g699)
--	g18212 = AND(g947, g15979)
--	g29596 = AND(g27823, g28620)
--	g24945 = AND(g23183, g20197)
--	g10719 = AND(g6841, g2138, g2130)
--	g16517 = AND(g5248, g14797)
--	g21833 = AND(g15096, g20453)
--	g30215 = AND(g28690, g23881)
--	g32409 = AND(g4754, g30996)
--	g14719 = AND(g4392, g10830)
--	g34215 = AND(g33778, g22670)
--	g30577 = AND(g26267, g29679)
--	g34577 = AND(g24577, g34307)
--	g25518 = AND(g6444, g23865, I24625)
--	g27428 = AND(g26400, g17576)
--	g13564 = AND(g4480, g12820)
--	g22044 = AND(g6058, g21611)
--	g26304 = AND(g2697, g25246)
--	g31143 = AND(g29506, g22999)
--	I24709 = AND(g21256, g24068, g24069, g24070)
--	I31021 = AND(g31070, g31799, g32485, g32486)
--	g24998 = AND(g17412, g23408)
--	g12730 = AND(g9024, g4349)
--	g27765 = AND(g4146, g25886)
--	g24651 = AND(g2741, g23472)
--	g24672 = AND(g19534, g22981)
--	g14832 = AND(g1489, g10939)
--	g29773 = AND(g28203, g10233)
--	g27690 = AND(g25784, g23607)
--	g16193 = AND(g6533, g14348)
--	g27549 = AND(g26576, g14785)
--	g31169 = AND(g10083, g30079)
--	g11397 = AND(g5360, g7139)
--	g18723 = AND(g4922, g16077)
--	g25883 = AND(g13728, g24699)
--	g28360 = AND(g27401, g19861)
--	g22120 = AND(g6585, g19277)
--	g33884 = AND(g33295, g20590)
--	g15116 = AND(g4297, g14454)
--	g18149 = AND(g608, g17533)
--	g27548 = AND(g26576, g17763)
--	g31168 = AND(g2241, g30077)
--	g32164 = AND(g30733, g25171)
--	g18433 = AND(g2197, g18008)
--	g33410 = AND(g32360, g21409)
--	g18387 = AND(g1955, g15171)
--	g24331 = AND(g6977, g22228)
--	g30083 = AND(g28533, g20698)
--	g13509 = AND(g9951, g11889)
--	g27504 = AND(g26519, g17680)
--	g18620 = AND(g3470, g17062)
--	g18148 = AND(g562, g17533)
--	g21947 = AND(g5256, g18997)
--	g30284 = AND(g28852, g23994)
--	g34083 = AND(g33714, g19573)
--	g34348 = AND(g34125, g20128)
--	I31593 = AND(g31003, g8350, g7788)
--	g33479 = AND(g32593, I31091, I31092)
--	g34284 = AND(g34046, g19351)
--	g21605 = AND(g13005, g15695)
--	I31346 = AND(g31021, g31857, g32954, g32955)
--	g33363 = AND(g32262, g20918)
--	g13508 = AND(g9927, g11888)
--	g18104 = AND(g392, g17015)
--	g18811 = AND(g6500, g15483)
--	g18646 = AND(g4031, g17271)
--	I31122 = AND(g32631, g32632, g32633, g32634)
--	g14612 = AND(g11971, g11993)
--	g31478 = AND(g29764, g23410)
--	g8234 = AND(g4515, g4521)
--	g31015 = AND(g29476, g22758)
--	g18343 = AND(g12847, g17955)
--	g24897 = AND(g3401, g23223, I24064)
--	g29839 = AND(g1728, g29045)
--	g30566 = AND(g26247, g29507)
--	g33478 = AND(g32584, I31086, I31087)
--	g24961 = AND(g23193, g20209)
--	g21812 = AND(g3586, g20924)
--	g17146 = AND(g5965, g14895)
--	g34566 = AND(g34376, g17489)
--	g28451 = AND(g27283, g20090)
--	g16222 = AND(g6513, g14348)
--	g31486 = AND(g29777, g23422)
--	g32327 = AND(g31319, g23544)
--	g29667 = AND(g2671, g29157)
--	g29838 = AND(g1636, g29044)
--	g27129 = AND(g26026, g16584)
--	g33486 = AND(g32642, I31126, I31127)
--	g32109 = AND(g31609, g29920)
--	g21951 = AND(g5272, g18997)
--	g26852 = AND(g24975, g24958)
--	g21972 = AND(g15152, g19074)
--	g27057 = AND(g7791, g6219, g6227, g26261)
--	g19610 = AND(g1141, g16069)
--	g18369 = AND(g12848, g15171)
--	g24717 = AND(g22684, g19777)
--	g27128 = AND(g25997, g16583)
--	g28246 = AND(g8572, g27976)
--	I31292 = AND(g32877, g32878, g32879, g32880)
--	g32108 = AND(g31631, g29913)
--	g30139 = AND(g28596, g21184)
--	g18368 = AND(g1728, g17955)
--	g34139 = AND(g33827, g23314)
--	g16703 = AND(g5889, g15002)
--	g22632 = AND(g19356, g19476)
--	g31223 = AND(g20028, g29689)
--	g21795 = AND(g3506, g20924)
--	g32283 = AND(g31259, g20506)
--	g27323 = AND(g26268, g23086)
--	g30138 = AND(g28595, g21182)
--	g27299 = AND(g26546, g23028)
--	g29619 = AND(g2269, g29060)
--	g32303 = AND(g27550, g31376)
--	g34138 = AND(g33929, g23828)
--	g11047 = AND(g6474, g9212)
--	g18412 = AND(g2098, g15373)
--	I31136 = AND(g29385, g32651, g32652, g32653)
--	g11205 = AND(g8217, g8439)
--	g13047 = AND(g8534, g11042)
--	g27298 = AND(g26573, g23026)
--	g29618 = AND(g28870, g22384)
--	g19383 = AND(g16893, g13223)
--	g34415 = AND(g34207, g21458)
--	g18133 = AND(g15055, g17249)
--	g23514 = AND(g20149, g11829)
--	g26484 = AND(g24946, g8841)
--	g33110 = AND(g32404, g32415)
--	g13912 = AND(g5551, g12450)
--	g34333 = AND(g9984, g34192)
--	g24723 = AND(g17490, g22384)
--	g31321 = AND(g30146, g27886)
--	g18229 = AND(g1099, g16326)
--	g33922 = AND(g33448, g7202)
--	g14061 = AND(g8715, g11834)
--	g33531 = AND(g32967, I31351, I31352)
--	g18228 = AND(g1061, g16129)
--	g24387 = AND(g3457, g22761)
--	g26312 = AND(g2704, g25264)
--	g34963 = AND(g34946, g23041)
--	g26200 = AND(g24688, g10678, g10658, g10627)
--	g32174 = AND(g31708, g27837)
--	g21163 = AND(g16321, g4878)
--	g21012 = AND(g16304, g4688)
--	g28151 = AND(g8426, g27295)
--	g18716 = AND(g4878, g15915)
--	g31186 = AND(g2375, g30088)
--	g33186 = AND(g32037, g22830)
--	g24646 = AND(g22640, g19711)
--	g33676 = AND(g33125, g7970)
--	g33373 = AND(g32288, g21205)
--	g16516 = AND(g5228, g14627)
--	g27697 = AND(g25785, g23649)
--	g18582 = AND(g2922, g16349)
--	g27995 = AND(g26809, g23985)
--	g31654 = AND(g29325, g13062)
--	g30576 = AND(g18898, g29800)
--	g22127 = AND(g6625, g19277)
--	g34585 = AND(g24705, g34316)
--	g34484 = AND(g34407, g18939)
--	g18310 = AND(g1333, g16931)
--	g29601 = AND(g1890, g28955)
--	g31936 = AND(g31213, g24005)
--	g33417 = AND(g32371, g21424)
--	I31327 = AND(g32928, g32929, g32930, g32931)
--	g21789 = AND(g3451, g20391)
--	g26799 = AND(g25247, g21068)
--	g29975 = AND(g28986, g10420)
--	g34554 = AND(g34347, g20495)
--	g18627 = AND(g15093, g17093)
--	g15863 = AND(g13762, g13223)
--	g18379 = AND(g1906, g15171)
--	g30200 = AND(g28665, g23862)
--	g21788 = AND(g3401, g20391)
--	g33334 = AND(g32219, g20613)
--	g18112 = AND(g182, g17015)
--	g16422 = AND(g8216, g13627)
--	g23724 = AND(g14767, g21123)
--	g25852 = AND(g4593, g24411)
--	g18378 = AND(g1932, g15171)
--	g22103 = AND(g15164, g18833)
--	g34115 = AND(g20516, g9104, g33750)
--	g21829 = AND(g3770, g20453)
--	g29937 = AND(g13044, g29196)
--	g14220 = AND(g8612, g11820)
--	g21920 = AND(g5062, g21468)
--	g23920 = AND(g4135, g19549)
--	g22095 = AND(g6428, g18833)
--	g16208 = AND(g3965, g14085)
--	g25963 = AND(g1657, g24978)
--	g28318 = AND(g27233, g19770)
--	g18386 = AND(g1964, g15171)
--	g30921 = AND(g29900, g24789)
--	g28227 = AND(g9397, g27583)
--	g21828 = AND(g3767, g20453)
--	g15703 = AND(g452, g13437)
--	g17784 = AND(g1152, g13215)
--	g23828 = AND(g9104, g19128)
--	g18603 = AND(g3119, g16987)
--	g21946 = AND(g5252, g18997)
--	g18742 = AND(g5120, g17847)
--	g27445 = AND(g8038, g26314, g9187, g504)
--	g33423 = AND(g32225, g29657)
--	g29884 = AND(g2555, g29153)
--	g23121 = AND(g19128, g9104)
--	g24229 = AND(g896, g22594)
--	g34745 = AND(g34669, g19482)
--	g27316 = AND(g2407, g26710)
--	g24228 = AND(g862, g22594)
--	g18681 = AND(g4653, g15885)
--	I31091 = AND(g29385, g32586, g32587, g32588)
--	g24011 = AND(g7939, g19524)
--	g32326 = AND(g31317, g23539)
--	g29666 = AND(g28980, g22498)
--	g17181 = AND(g1945, g13014)
--	g16614 = AND(g5945, g14933)
--	g17671 = AND(g7685, g13485)
--	g29363 = AND(g8458, g28444)
--	g23682 = AND(g16970, g20874)
--	g18802 = AND(g6195, g15348)
--	g18429 = AND(g2193, g18008)
--	g32040 = AND(g14122, g31243)
--	g24716 = AND(g15935, g23004)
--	I24680 = AND(g24029, g24030, g24031, g24032)
--	g33909 = AND(g33131, g10708)
--	g34184 = AND(g33698, g24388)
--	g18730 = AND(g4950, g16861)
--	g15821 = AND(g3598, g14110)
--	g27988 = AND(g26781, g23941)
--	g18793 = AND(g6159, g15348)
--	g18428 = AND(g2169, g18008)
--	g24582 = AND(g5808, g23402)
--	g33908 = AND(g33092, g18935)
--	g28281 = AND(g7362, g1936, g27440)
--	g16593 = AND(g5599, g14885)
--	g12924 = AND(g1570, g10980)
--	g27432 = AND(g26519, g17582)
--	g13020 = AND(g401, g11048)
--	g18765 = AND(g5489, g17929)
--	g28301 = AND(g27224, g19750)
--	g24310 = AND(g4495, g22228)
--	g16122 = AND(g9491, g14291)
--	g18690 = AND(g15130, g16053)
--	g28739 = AND(g21434, g26424, g25274, g27395)
--	g18549 = AND(g2799, g15277)
--	g11046 = AND(g9889, g6120)
--	g25921 = AND(g24936, g9664)
--	g13046 = AND(g6870, g11270)
--	g26207 = AND(g2638, g25170)
--	g24627 = AND(g22763, g19679)
--	g29580 = AND(g28519, g14186)
--	g21760 = AND(g3207, g20785)
--	g20112 = AND(g13540, g16661)
--	g31242 = AND(g29373, g25409)
--	g22089 = AND(g6311, g19210)
--	g27461 = AND(g26576, g17611)
--	g33242 = AND(g32123, g19931)
--	g18548 = AND(g2807, g15277)
--	g15873 = AND(g3550, g14072)
--	g28645 = AND(g27556, g20599)
--	I31192 = AND(g32733, g32734, g32735, g32736)
--	g27342 = AND(g12592, g26792)
--	g24378 = AND(g3106, g22718)
--	g16641 = AND(g6613, g14782)
--	g27145 = AND(g14121, g26382)
--	g22088 = AND(g6307, g19210)
--	g18504 = AND(g2579, g15509)
--	g22024 = AND(g5897, g19147)
--	g31123 = AND(g1834, g29994)
--	g32183 = AND(g2795, g31653)
--	g19266 = AND(g246, g16214)
--	g33814 = AND(g33098, g28144)
--	g28290 = AND(g23780, g27759)
--	g32397 = AND(g31068, g15830)
--	g13282 = AND(g3546, g11480)
--	g27650 = AND(g26519, g15479)
--	g29110 = AND(g27187, g12687, g20751, I27429)
--	g25973 = AND(g2342, g24994)
--	g18317 = AND(g12846, g17873)
--	g33807 = AND(g33112, g25452)
--	g31974 = AND(g31760, g22176)
--	g29321 = AND(g29033, g22148)
--	g33639 = AND(g33386, g18829)
--	g26241 = AND(g24688, g10678, g8778, g10627)
--	g34214 = AND(g33772, g22689)
--	g29531 = AND(g1664, g28559)
--	g31230 = AND(g30285, g20751)
--	g18129 = AND(g518, g16971)
--	g30207 = AND(g28680, g23874)
--	g16635 = AND(g5607, g14959)
--	g27696 = AND(g25800, g23647)
--	g34329 = AND(g14511, g34181)
--	g27330 = AND(g2541, g26744)
--	g27393 = AND(g26099, g20066)
--	g28427 = AND(g27258, g20008)
--	g24681 = AND(g16653, g22988)
--	g29178 = AND(g27163, g12687)
--	g29740 = AND(g2648, g29154)
--	g30005 = AND(g28230, g24394)
--	g22126 = AND(g6621, g19277)
--	g18128 = AND(g504, g16971)
--	g21927 = AND(g5164, g18997)
--	g26100 = AND(g1677, g25097)
--	g19588 = AND(g3849, g16853)
--	g33416 = AND(g32370, g21423)
--	g29685 = AND(g2084, g28711)
--	I31326 = AND(g30735, g31853, g32926, g32927)
--	g18245 = AND(g1193, g16431)
--	g27132 = AND(g26055, g16589)
--	g34538 = AND(g34330, g20054)
--	g18626 = AND(g3498, g17062)
--	g15913 = AND(g3933, g14021)
--	g24730 = AND(g6177, g23699)
--	g31992 = AND(g31773, g22213)
--	g18323 = AND(g1632, g17873)
--	g33841 = AND(g33254, g20268)
--	g18299 = AND(g1526, g16489)
--	g18533 = AND(g2729, g15277)
--	g28547 = AND(g6821, g27091)
--	g33510 = AND(g32816, I31246, I31247)
--	g24765 = AND(g17699, g22498)
--	g18298 = AND(g15073, g16489)
--	g27161 = AND(g26166, g8241, g1783)
--	g30241 = AND(g28729, g23926)
--	I31252 = AND(g32819, g32820, g32821, g32822)
--	g31579 = AND(g19128, g29814)
--	g18775 = AND(g7028, g15615)
--	g24549 = AND(g23162, g20887)
--	g28226 = AND(g27825, g26667)
--	g21755 = AND(g3203, g20785)
--	g29334 = AND(g29148, g18908)
--	g16474 = AND(g8280, g13666)
--	g23755 = AND(g14821, g21204)
--	g27259 = AND(g26755, g26725)
--	g19749 = AND(g732, g16646)
--	g32047 = AND(g27248, g31070)
--	g33835 = AND(g4340, g33413)
--	g9968 = AND(g1339, g1500)
--	g21770 = AND(g3251, g20785)
--	g32205 = AND(g30922, g28463)
--	g21981 = AND(g5543, g19074)
--	g22060 = AND(g6151, g21611)
--	g10902 = AND(g7858, g1129)
--	g18737 = AND(g4975, g16826)
--	g27087 = AND(g13872, g26284)
--	g28572 = AND(g27829, g15669)
--	g12259 = AND(g9480, g640)
--	g24504 = AND(g22226, g19410)
--	g32311 = AND(g31295, g20582)
--	g25207 = AND(g22513, g10621)
--	g29762 = AND(g28298, g10233)
--	g18232 = AND(g1124, g16326)
--	g34771 = AND(g34693, g20147)
--	g29964 = AND(g2008, g28830)
--	g16537 = AND(g5937, g14855)
--	g11027 = AND(g5097, g9724)
--	g30235 = AND(g28723, g23915)
--	I18713 = AND(g13156, g6767, g6756)
--	g25328 = AND(g5022, g23764, I24505)
--	g11890 = AND(g7499, g9155)
--	g24317 = AND(g4534, g22228)
--	g15797 = AND(g3909, g14139)
--	g18697 = AND(g4749, g16777)
--	g27043 = AND(g26335, g8632)
--	g32051 = AND(g31506, g10831)
--	g16283 = AND(g11547, g11592, g6789, I17606)
--	g29587 = AND(g2181, g28935)
--	I31062 = AND(g32545, g32546, g32547, g32548)
--	g18261 = AND(g1256, g16000)
--	g21767 = AND(g3239, g20785)
--	g21794 = AND(g15094, g20924)
--	g21845 = AND(g3881, g21070)
--	g12043 = AND(g1345, g7601)
--	g16303 = AND(g4527, g12921)
--	g10290 = AND(g4358, g4349)
--	g24002 = AND(g19613, g10971)
--	g21990 = AND(g5591, g19074)
--	g11003 = AND(g7880, g1300)
--	g18512 = AND(g2619, g15509)
--	g23990 = AND(g19610, g10951)
--	I27524 = AND(g28037, g24114, g24115, g24116)
--	g33720 = AND(g33161, g19439)
--	g19560 = AND(g15832, g1157, g10893)
--	g29909 = AND(g28435, g23388)
--	g27602 = AND(g23032, g26244, g26424, g24966)
--	g31275 = AND(g30147, g27800)
--	g34515 = AND(g34288, g19491)
--	g34414 = AND(g34206, g21457)
--	g28889 = AND(g17292, g25169, g26424, g27395)
--	g31746 = AND(g30093, g23905)
--	g27375 = AND(g26519, g17479)
--	g26206 = AND(g2523, g25495)
--	g31493 = AND(g29791, g23434)
--	g32350 = AND(g2697, g31710)
--	g21719 = AND(g358, g21037)
--	g33493 = AND(g32693, I31161, I31162)
--	g24323 = AND(g4546, g22228)
--	g24299 = AND(g4456, g22550)
--	g13778 = AND(g4540, g10597)
--	g13081 = AND(g8626, g11122)
--	g29569 = AND(g29028, g22498)
--	g21718 = AND(g370, g21037)
--	g33465 = AND(g32491, I31021, I31022)
--	g31237 = AND(g29366, g25325)
--	g10632 = AND(g7475, g7441, g890)
--	g24298 = AND(g4392, g22550)
--	g33237 = AND(g32394, g25198)
--	g32152 = AND(g31631, g29998)
--	g18445 = AND(g2273, g18008)
--	g24775 = AND(g17594, g22498)
--	g29568 = AND(g2571, g28950)
--	g29747 = AND(g28286, g23196)
--	g32396 = AND(g4698, g30983)
--	g33340 = AND(g32222, g20639)
--	g21832 = AND(g3787, g20453)
--	g18499 = AND(g2476, g15426)
--	g18316 = AND(g1564, g16931)
--	g33684 = AND(g33139, g13565)
--	g16840 = AND(g5467, g14262)
--	g31142 = AND(g2527, g30039)
--	g22055 = AND(g6128, g21611)
--	g18498 = AND(g2547, g15426)
--	g32413 = AND(g31121, g19518)
--	g19693 = AND(g6181, g17087)
--	g22111 = AND(g6549, g19277)
--	I31047 = AND(g32524, g32525, g32526, g32527)
--	g21861 = AND(g3949, g21070)
--	g34584 = AND(g24653, g34315)
--	g22070 = AND(g6243, g19210)
--	g13998 = AND(g6589, g12629)
--	g31517 = AND(g29849, g23482)
--	g26345 = AND(g13051, g25505)
--	g28426 = AND(g27257, g20006)
--	g33517 = AND(g32867, I31281, I31282)
--	g29751 = AND(g28297, g23216)
--	g29807 = AND(g28359, g23272)
--	I31311 = AND(g30673, g31851, g32903, g32904)
--	g29772 = AND(g28323, g23243)
--	g22590 = AND(g19274, g19452)
--	g16192 = AND(g6191, g14321)
--	g26849 = AND(g2994, g24527)
--	g29974 = AND(g29173, g12914)
--	g15711 = AND(g460, g13437)
--	g18611 = AND(g15090, g17200)
--	g27459 = AND(g26549, g17609)
--	g21926 = AND(g15147, g18997)
--	g18722 = AND(g4917, g16077)
--	g26399 = AND(g15572, g25566)
--	g25414 = AND(g5406, g22194, I24549)
--	g25991 = AND(g2060, g25023)
--	g23389 = AND(g9072, g19757)
--	g29639 = AND(g28510, g11618)
--	g15109 = AND(g4269, g14454)
--	g26848 = AND(g2950, g24526)
--	I16646 = AND(g10160, g12413, g12343)
--	g26398 = AND(g24946, g10474)
--	g22384 = AND(g9354, g9285, g20784)
--	g18432 = AND(g2223, g18008)
--	I24705 = AND(g24064, g24065, g24066, g24067)
--	g29638 = AND(g2583, g29025)
--	I31051 = AND(g31376, g31804, g32529, g32530)
--	g21701 = AND(g153, g20283)
--	I31072 = AND(g32559, g32560, g32561, g32562)
--	g18271 = AND(g1296, g16031)
--	g30082 = AND(g29181, g12752)
--	g34114 = AND(g33920, g23742)
--	g15108 = AND(g4264, g14454)
--	g21777 = AND(g3380, g20391)
--	g34758 = AND(g34683, g19657)
--	g26652 = AND(g10799, g24426)
--	g31130 = AND(g12191, g30019)
--	g22067 = AND(g6215, g19210)
--	g22094 = AND(g6398, g18833)
--	g34082 = AND(g33709, g19554)
--	g30107 = AND(g28560, g20909)
--	g21251 = AND(g13969, g17470)
--	I24679 = AND(g19968, g24026, g24027, g24028)
--	g33362 = AND(g32259, g20914)
--	g11449 = AND(g6052, g7175)
--	g27545 = AND(g26519, g17756)
--	g16483 = AND(g5224, g14915)
--	g18753 = AND(g15148, g15595)
--	g18461 = AND(g2307, g15224)
--	g31523 = AND(g7528, g29333)
--	g32020 = AND(g4157, g30937)
--	g18342 = AND(g1592, g17873)
--	g33523 = AND(g32909, I31311, I31312)
--	g29841 = AND(g28371, g23283)
--	g19914 = AND(g2815, g15853)
--	g29992 = AND(g29012, g10490)
--	g27599 = AND(g26337, g20033)
--	g34744 = AND(g34668, g19481)
--	g18145 = AND(g582, g17533)
--	g29510 = AND(g28856, g22342)
--	g32046 = AND(g10925, g30735)
--	g18199 = AND(g832, g17821)
--	g22019 = AND(g5857, g19147)
--	g27598 = AND(g25899, g10475)
--	g18650 = AND(g6928, g17271)
--	g18736 = AND(g4991, g16826)
--	g27086 = AND(g25836, g22495)
--	g31475 = AND(g29756, g23406)
--	g29579 = AND(g28457, g7964)
--	g17150 = AND(g8579, g12995)
--	I24030 = AND(g8390, g8016, g3396)
--	g33475 = AND(g32563, I31071, I31072)
--	g16536 = AND(g5917, g14996)
--	g18198 = AND(g15059, g17821)
--	g22018 = AND(g15157, g19147)
--	g18529 = AND(g2712, g15277)
--	g21997 = AND(g5619, g19074)
--	g32113 = AND(g31601, g29925)
--	g34398 = AND(g7684, g34070)
--	I31152 = AND(g32675, g32676, g32677, g32678)
--	g33727 = AND(g33115, g19499)
--	g24499 = AND(g22217, g19394)
--	g29578 = AND(g2491, g28606)
--	g33863 = AND(g33273, g20505)
--	g19594 = AND(g11913, g17268)
--	g29835 = AND(g28326, g24866)
--	g34141 = AND(g33932, g23828)
--	g16702 = AND(g5615, g14691)
--	g24316 = AND(g4527, g22228)
--	g31222 = AND(g2643, g30113)
--	g32282 = AND(g31258, g20503)
--	g27817 = AND(g22498, g25245, g26424, g26236)
--	g15796 = AND(g3586, g14015)
--	g18696 = AND(g4741, g16053)
--	g18330 = AND(g1668, g17873)
--	g32302 = AND(g31279, g23485)
--	g18393 = AND(g1917, g15171)
--	g24498 = AND(g14036, g23850)
--	g29586 = AND(g1886, g28927)
--	g16621 = AND(g8278, g13821)
--	g12817 = AND(g1351, g7601)
--	g21766 = AND(g3235, g20785)
--	g26833 = AND(g2852, g24509)
--	g26049 = AND(g9621, g25046)
--	g30263 = AND(g28773, g23962)
--	g32105 = AND(g4922, g30673)
--	g28658 = AND(g27563, g20611)
--	g18764 = AND(g5485, g17929)
--	g20056 = AND(g16291, g9007, g8954, g8903)
--	g18365 = AND(g1848, g17955)
--	g27158 = AND(g26609, g16645)
--	g21871 = AND(g4108, g19801)
--	g25107 = AND(g17643, g23508)
--	g22457 = AND(g7753, g7717, g21288)
--	g15840 = AND(g3949, g14142)
--	g18132 = AND(g513, g16971)
--	g26048 = AND(g5853, g25044)
--	g28339 = AND(g9946, g27693)
--	g30135 = AND(g28592, g21180)
--	g24722 = AND(g17618, g22417)
--	g34135 = AND(g33926, g23802)
--	I18782 = AND(g13156, g11450, g6756)
--	g7948 = AND(g1548, g1430)
--	g29615 = AND(g1844, g29049)
--	g16673 = AND(g6617, g14822)
--	g18161 = AND(g691, g17433)
--	g34962 = AND(g34945, g23020)
--	g19637 = AND(g5142, g16958)
--	g26613 = AND(g1361, g24518)
--	g18709 = AND(g59, g17302)
--	g22001 = AND(g5731, g21562)
--	g22077 = AND(g6263, g19210)
--	g25848 = AND(g25539, g18977)
--	g14190 = AND(g859, g10632)
--	g27336 = AND(g2675, g26777)
--	g30049 = AND(g13114, g28167)
--	g18259 = AND(g15068, g16000)
--	g29746 = AND(g28279, g20037)
--	g34500 = AND(g34276, g30568)
--	g18225 = AND(g1041, g16100)
--	g33351 = AND(g32236, g20707)
--	g33372 = AND(g32285, g21183)
--	g18708 = AND(g4818, g16782)
--	g28197 = AND(g27647, g11344)
--	g25804 = AND(g8069, g24587)
--	g18471 = AND(g2407, g15224)
--	g33821 = AND(g33238, g20153)
--	g26273 = AND(g2122, g25389)
--	g30048 = AND(g29193, g12945)
--	g22689 = AND(g18918, g9104)
--	g18258 = AND(g1221, g16897)
--	g16634 = AND(g5264, g14953)
--	g20887 = AND(g16282, g4864)
--	g23451 = AND(g13805, g20510)
--	g24199 = AND(g355, g22722)
--	g24650 = AND(g22641, g19718)
--	g23220 = AND(g19417, g20067)
--	g24887 = AND(g3712, g23239, I24054)
--	g30004 = AND(g28521, g25837)
--	I31046 = AND(g29385, g32521, g32522, g32523)
--	g22624 = AND(g19344, g19471)
--	g21911 = AND(g5046, g21468)
--	g30221 = AND(g28700, g23893)
--	g31790 = AND(g21299, g29385)
--	g33264 = AND(g31965, g21306)
--	g31516 = AND(g29848, g23476)
--	g24198 = AND(g351, g22722)
--	g33790 = AND(g33108, g20643)
--	g33516 = AND(g32860, I31276, I31277)
--	g29806 = AND(g28358, g23271)
--	g29684 = AND(g1982, g29085)
--	g18244 = AND(g1171, g16431)
--	g26234 = AND(g2657, g25514)
--	g22102 = AND(g6479, g18833)
--	g24843 = AND(g3010, g23211, I24015)
--	g33873 = AND(g33291, g20549)
--	g24330 = AND(g18661, g22228)
--	g22157 = AND(g14608, g18892)
--	g24393 = AND(g3808, g22844)
--	I24075 = AND(g3736, g3742, g8553)
--	I31282 = AND(g32863, g32864, g32865, g32866)
--	g25962 = AND(g9258, g24971)
--	g16213 = AND(g6772, g6782, g11640, I17552)
--	g24764 = AND(g17570, g22472)
--	g29517 = AND(g1870, g28827)
--	I31302 = AND(g32891, g32892, g32893, g32894)
--	I31357 = AND(g32970, g32971, g32972, g32973)
--	g21776 = AND(g3376, g20391)
--	g21785 = AND(g3431, g20391)
--	I27519 = AND(g28036, g24107, g24108, g24109)
--	g18602 = AND(g3115, g16987)
--	g18810 = AND(g6505, g15483)
--	g15757 = AND(g3207, g14066)
--	g18657 = AND(g4308, g17128)
--	g22066 = AND(g6209, g19210)
--	g18774 = AND(g5698, g15615)
--	g7918 = AND(g1205, g1087)
--	g18375 = AND(g1902, g15171)
--	g31209 = AND(g2084, g30097)
--	g33422 = AND(g32375, g21456)
--	g34106 = AND(g33917, g23675)
--	g32248 = AND(g31616, g30299)
--	g21754 = AND(g3195, g20785)
--	I27518 = AND(g20720, g24104, g24105, g24106)
--	g10625 = AND(g3431, g7926)
--	g27309 = AND(g26603, g23057)
--	g23754 = AND(g14816, g21189)
--	g28714 = AND(g27591, g20711)
--	g16047 = AND(g13322, g1500, g10699)
--	g25833 = AND(g8228, g24626)
--	g14126 = AND(g881, g10632)
--	g16205 = AND(g11547, g6782, g11640, I17542)
--	g27288 = AND(g26515, g23013)
--	g28315 = AND(g27232, g19769)
--	g33834 = AND(g33095, g29172)
--	g31208 = AND(g30262, g25188)
--	g32204 = AND(g4245, g31327)
--	g21859 = AND(g3941, g21070)
--	g21825 = AND(g3736, g20453)
--	g21950 = AND(g5268, g18997)
--	g26514 = AND(g7400, g25564)
--	g22876 = AND(g20136, g9104)
--	g18337 = AND(g1706, g17873)
--	g28202 = AND(g27659, g11413)
--	g30033 = AND(g29189, g12937)
--	g28257 = AND(g27179, g19686)
--	g21858 = AND(g3937, g21070)
--	g29362 = AND(g27379, g28307)
--	g18171 = AND(g728, g17433)
--	g30234 = AND(g28721, g23914)
--	g34371 = AND(g7450, g34044)
--	g24709 = AND(g16690, g23000)
--	g31542 = AND(g19050, g29814)
--	g31021 = AND(g26025, g29814)
--	g29523 = AND(g28930, g22417)
--	g23151 = AND(g18994, g7162)
--	g28111 = AND(g27343, g22716)
--	g14296 = AND(g2638, g11897)
--	g21996 = AND(g5615, g19074)
--	g24225 = AND(g246, g22594)
--	g15673 = AND(g182, g13437)
--	g18792 = AND(g7051, g15634)
--	g15847 = AND(g3191, g14005)
--	g23996 = AND(g19596, g10951)
--	g24708 = AND(g16474, g22998)
--	g14644 = AND(g10610, g10605)
--	g33913 = AND(g23088, g33204, g9104)
--	g16592 = AND(g5579, g14688)
--	g21844 = AND(g3873, g21070)
--	g21394 = AND(g13335, g15799)
--	g32356 = AND(g2704, g31710)
--	g29475 = AND(g14033, g28500)
--	g18459 = AND(g2331, g15224)
--	g18425 = AND(g2161, g18008)
--	g33905 = AND(g33089, g15574)
--	g33073 = AND(g32386, g18828)
--	g12687 = AND(g9024, g8977)
--	g25106 = AND(g17391, g23506)
--	g26541 = AND(g319, g24375)
--	g34514 = AND(g34286, g19480)
--	g15851 = AND(g3953, g14157)
--	g15872 = AND(g9095, g14234)
--	g18458 = AND(g2357, g15224)
--	g19139 = AND(g452, g16195)
--	g27374 = AND(g26519, g17478)
--	g33530 = AND(g32960, I31346, I31347)
--	g21420 = AND(g16093, g13596)
--	g34507 = AND(g34280, g19454)
--	g31122 = AND(g12144, g29993)
--	g32182 = AND(g31753, g27937)
--	g20069 = AND(g16312, g9051, g9011, g8955)
--	g33122 = AND(g8859, g32192)
--	g8530 = AND(g2902, g2907)
--	I31027 = AND(g32494, g32495, g32496, g32497)
--	I24524 = AND(g5041, g5046, g9716)
--	g33464 = AND(g32484, I31016, I31017)
--	I16129 = AND(g8728, g11443, g11411)
--	g20602 = AND(g10803, g15580)
--	g28150 = AND(g10862, g11834, g11283, g27187)
--	g16846 = AND(g14034, g12591, g11185)
--	g18545 = AND(g2783, g15277)
--	g25951 = AND(g24500, g19565)
--	g26325 = AND(g12644, g25370)
--	g24602 = AND(g16507, g22854)
--	g25972 = AND(g2217, g24993)
--	g18444 = AND(g2269, g18008)
--	g25033 = AND(g17500, g23433)
--	g25371 = AND(g5062, g22173, I24524)
--	g20375 = AND(g671, g16846)
--	g24657 = AND(g22644, g19730)
--	g24774 = AND(g718, g23614)
--	g16731 = AND(g7153, g12941)
--	g26829 = AND(g2844, g24505)
--	g27669 = AND(g26840, g13278)
--	g17480 = AND(g9683, g14433)
--	g19333 = AND(g464, g16223)
--	g29347 = AND(g29176, g22201)
--	g18599 = AND(g2955, g16349)
--	g22307 = AND(g20027, g21163)
--	g22076 = AND(g6255, g19210)
--	g22085 = AND(g6295, g19210)
--	g26358 = AND(g19522, g25528)
--	I27349 = AND(g25534, g26424, g22698)
--	g23025 = AND(g16021, g19798)
--	g27260 = AND(g26766, g26737)
--	g32331 = AND(g31322, g20637)
--	g31292 = AND(g29735, g23338)
--	g26828 = AND(g24919, g15756)
--	g27668 = AND(g1367, g25917)
--	g23540 = AND(g16866, g20622)
--	g18598 = AND(g3003, g16349)
--	g22054 = AND(g6120, g21611)
--	g28695 = AND(g27580, g20666)
--	g31153 = AND(g12336, g30068)
--	g27392 = AND(g26576, g17507)
--	g29600 = AND(g1840, g29049)
--	g26121 = AND(g6167, g25111)
--	g20171 = AND(g16479, g10476)
--	g34541 = AND(g34331, g20087)
--	g17307 = AND(g9498, g14343)
--	g15574 = AND(g4311, g13202)
--	g33409 = AND(g32359, g21408)
--	I24616 = AND(g6082, g6088, g9946)
--	g29952 = AND(g23576, g28939)
--	g27559 = AND(g26576, g17777)
--	g29351 = AND(g4771, g28406)
--	g27525 = AND(g26576, g17720)
--	g27488 = AND(g26549, g17648)
--	g18817 = AND(g6533, g15483)
--	g15912 = AND(g3562, g14018)
--	g14581 = AND(g12587, g12428, g12357, I16695)
--	g18322 = AND(g1608, g17873)
--	g33408 = AND(g32358, g21407)
--	I31081 = AND(g30673, g31810, g32571, g32572)
--	g24967 = AND(g23197, g20213)
--	g10707 = AND(g3787, g8561)
--	g18159 = AND(g671, g17433)
--	g27558 = AND(g26576, g17776)
--	g25507 = AND(g6098, g23844, I24616)
--	g22942 = AND(g9104, g20219)
--	g18125 = AND(g15053, g16886)
--	g18532 = AND(g2724, g15277)
--	g26291 = AND(g2681, g25439)
--	g30920 = AND(g29889, g21024)
--	I24704 = AND(g21193, g24061, g24062, g24063)
--	g19585 = AND(g17180, g14004)
--	g14202 = AND(g869, g10632)
--	g16929 = AND(g6505, g14348)
--	g18158 = AND(g667, g17433)
--	g14257 = AND(g8612, g11878)
--	g21957 = AND(g5390, g21514)
--	g18783 = AND(g5841, g18065)
--	g23957 = AND(g4138, g19589)
--	g29516 = AND(g28895, g22369)
--	g14496 = AND(g12411, g12244, g12197, I16618)
--	g22670 = AND(g20114, g9104)
--	g21739 = AND(g3080, g20330)
--	I31356 = AND(g31327, g31859, g32968, g32969)
--	g25163 = AND(g20217, g23566)
--	g18561 = AND(g2841, g15277)
--	g18656 = AND(g15120, g17128)
--	g30121 = AND(g28577, g21052)
--	g25012 = AND(g20644, g23419)
--	g18353 = AND(g1772, g17955)
--	g18295 = AND(g1489, g16449)
--	g21738 = AND(g3072, g20330)
--	g10590 = AND(g7246, g7392, I13937)
--	g17156 = AND(g305, g13385)
--	g17655 = AND(g7897, g13342)
--	g18680 = AND(g15128, g15885)
--	g18144 = AND(g590, g17533)
--	g18823 = AND(g6727, g15680)
--	g34344 = AND(g34107, g20038)
--	g21699 = AND(g142, g20283)
--	g28706 = AND(g27584, g20681)
--	g28597 = AND(g27515, g20508)
--	I31182 = AND(g32719, g32720, g32721, g32722)
--	g18336 = AND(g1700, g17873)
--	g24545 = AND(g3333, g23285)
--	g33474 = AND(g32556, I31066, I31067)
--	g28256 = AND(g11398, g27984)
--	g15820 = AND(g3578, g13955)
--	g28689 = AND(g27575, g20651)
--	g32149 = AND(g31658, g29983)
--	g27042 = AND(g25774, g19343)
--	g33711 = AND(g33176, g10727, g22332)
--	g30173 = AND(g28118, g13082)
--	g34291 = AND(g34055, g19366)
--	g31327 = AND(g19200, g29814)
--	g27255 = AND(g25936, g19689)
--	g28280 = AND(g23761, g27724)
--	g22131 = AND(g6641, g19277)
--	g29834 = AND(g28368, g23278)
--	g33327 = AND(g32208, g20561)
--	g34173 = AND(g33679, g24368)
--	I24064 = AND(g3385, g3391, g8492)
--	g29208 = AND(g24138, I27538, I27539)
--	g25788 = AND(g8010, g24579)
--	g32148 = AND(g31631, g29981)
--	g28624 = AND(g22357, g27009)
--	g28300 = AND(g27771, g26605)
--	g27270 = AND(g26805, g26793)
--	g32097 = AND(g25960, g31021)
--	I31331 = AND(g30825, g31854, g32933, g32934)
--	g27678 = AND(g947, g25830)
--	g18631 = AND(g3694, g17226)
--	g32104 = AND(g31616, g29906)
--	g7520 = AND(g2704, g2697, g2689)
--	g18364 = AND(g1844, g17955)
--	g32343 = AND(g31473, g20710)
--	g31283 = AND(g30156, g27837)
--	g27460 = AND(g26549, g17610)
--	g27686 = AND(g1291, g25849)
--	g25946 = AND(g24496, g19537)
--	g31492 = AND(g29790, g23431)
--	g24817 = AND(g22929, g7235)
--	g30029 = AND(g29164, g12936)
--	g33492 = AND(g32686, I31156, I31157)
--	g19674 = AND(g2819, g15867)
--	g24322 = AND(g4423, g22228)
--	g12939 = AND(g405, g11048)
--	g27030 = AND(g26343, g7947)
--	g20977 = AND(g10123, g17301)
--	g13299 = AND(g437, g11048)
--	g24532 = AND(g22331, g19478)
--	g32369 = AND(g2130, g31672)
--	g27267 = AND(g26026, g17124)
--	g27294 = AND(g9975, g26656)
--	g29614 = AND(g28860, g22369)
--	g30028 = AND(g29069, g9311)
--	g28231 = AND(g27187, g22763, g27074)
--	g24977 = AND(g23209, g20232)
--	g34506 = AND(g8833, g34354)
--	g16803 = AND(g5933, g14810)
--	g31750 = AND(g30103, g23925)
--	g29607 = AND(g28509, g14208)
--	g18289 = AND(g1448, g16449)
--	I31026 = AND(g31194, g31800, g32492, g32493)
--	g29320 = AND(g29068, g22147)
--	g33381 = AND(g11842, g32318)
--	I31212 = AND(g32761, g32762, g32763, g32764)
--	g29073 = AND(g27163, g10290, g21012, I27409)
--	g12065 = AND(g9557, g9805)
--	g18309 = AND(g1339, g16931)
--	g29530 = AND(g1612, g28820)
--	g24656 = AND(g11736, g22926)
--	g29593 = AND(g28470, g7985)
--	g33091 = AND(g32392, g18897)
--	g18288 = AND(g1454, g16449)
--	g18224 = AND(g1036, g16100)
--	g21715 = AND(g160, g20283)
--	g22039 = AND(g5949, g19147)
--	g29346 = AND(g4894, g28381)
--	g25173 = AND(g12234, g23589)
--	g24295 = AND(g4434, g22550)
--	g18571 = AND(g2856, g16349)
--	g18308 = AND(g6832, g16931)
--	g24680 = AND(g16422, g22986)
--	g27219 = AND(g26026, g16742)
--	g32412 = AND(g4765, g30998)
--	g24144 = AND(g17727, g21660)
--	g33796 = AND(g33117, g25267)
--	g19692 = AND(g12066, g17086)
--	I24555 = AND(g9559, g9809, g6093)
--	g29565 = AND(g1932, g28590)
--	g26604 = AND(g13248, g25051)
--	g17469 = AND(g4076, g13217)
--	g13737 = AND(g4501, g10571)
--	g22038 = AND(g5945, g19147)
--	g23551 = AND(g10793, g18948)
--	g23572 = AND(g20230, g20656)
--	g10917 = AND(g9174, g1087)
--	g12219 = AND(g1189, g7532)
--	g27218 = AND(g25997, g16740)
--	g30927 = AND(g29910, g24795)
--	g18495 = AND(g2533, g15426)
--	g33840 = AND(g33253, g20267)
--	g29641 = AND(g28520, g14237)
--	g29797 = AND(g28347, g23259)
--	g16662 = AND(g4552, g14753)
--	g13697 = AND(g11166, g8608)
--	g28660 = AND(g27824, g20623)
--	g18816 = AND(g6527, g15483)
--	g32011 = AND(g8287, g31134)
--	g27160 = AND(g14163, g26340)
--	g10706 = AND(g3338, g8691)
--	g15113 = AND(g4291, g14454)
--	g19207 = AND(g7803, g15992)
--	g18687 = AND(g4664, g15885)
--	g28456 = AND(g27290, g20104)
--	I31097 = AND(g32596, g32597, g32598, g32599)
--	g17601 = AND(g9616, g14572)
--	g22143 = AND(g19568, g10971)
--	g21784 = AND(g3423, g20391)
--	g22937 = AND(g753, g20540)
--	g26845 = AND(g24391, g21426)
--	g14256 = AND(g2079, g11872)
--	g21956 = AND(g5360, g21514)
--	g18752 = AND(g15146, g17926)
--	g27455 = AND(g26488, g17603)
--	g26395 = AND(g22547, g25561)
--	g30604 = AND(g18911, g29878)
--	g33522 = AND(g32902, I31306, I31307)
--	g18374 = AND(g1878, g15171)
--	g29635 = AND(g28910, g22432)
--	g21889 = AND(g4169, g19801)
--	g23103 = AND(g10143, g20765)
--	g27617 = AND(g23032, g26264, g26424, g24982)
--	g15105 = AND(g4235, g14454)
--	g21980 = AND(g5567, g19074)
--	g10624 = AND(g8387, g3072)
--	g28550 = AND(g12009, g27092)
--	g18643 = AND(g3849, g17096)
--	g7469 = AND(g4382, g4438)
--	g32310 = AND(g27577, g31376)
--	g16204 = AND(g6537, g14348)
--	g28314 = AND(g27552, g14205)
--	g21888 = AND(g4165, g19801)
--	g21824 = AND(g3706, g20453)
--	g26633 = AND(g24964, g20616)
--	g34563 = AND(g34372, g17465)
--	I17542 = AND(g13156, g6767, g6756)
--	g27201 = AND(g25997, g16685)
--	g27277 = AND(g26359, g14191)
--	I24675 = AND(g24022, g24023, g24024, g24025)
--	g33483 = AND(g32621, I31111, I31112)
--	g26719 = AND(g10709, g24438)
--	g24289 = AND(g4427, g22550)
--	g18669 = AND(g4608, g17367)
--	g32112 = AND(g31646, g29923)
--	g25927 = AND(g25004, g20375)
--	g32050 = AND(g11003, g30825)
--	g24309 = AND(g4480, g22228)
--	g33862 = AND(g33272, g20504)
--	g18260 = AND(g1252, g16000)
--	g28243 = AND(g27879, g23423)
--	g24288 = AND(g4417, g22550)
--	g27595 = AND(g26733, g26703)
--	g24224 = AND(g269, g22594)
--	g18668 = AND(g4322, g17367)
--	g27467 = AND(g269, g26832)
--	g27494 = AND(g8038, g26314, g518, g9077)
--	g31949 = AND(g1287, g30825)
--	g18392 = AND(g1988, g15171)
--	g29891 = AND(g28420, g23356)
--	g24308 = AND(g4489, g22228)
--	g21931 = AND(g5188, g18997)
--	g18195 = AND(g847, g17821)
--	g22015 = AND(g5719, g21562)
--	g18489 = AND(g2509, g15426)
--	g34395 = AND(g34193, g21336)
--	g31948 = AND(g30670, g18884)
--	g32096 = AND(g31601, g29893)
--	g28269 = AND(g27205, g19712)
--	g29575 = AND(g2066, g28604)
--	g15881 = AND(g3582, g13983)
--	g18559 = AND(g12856, g15277)
--	g25491 = AND(g23615, g21355)
--	g18525 = AND(g2610, g15509)
--	g18488 = AND(g2495, g15426)
--	g18424 = AND(g2165, g18008)
--	g28341 = AND(g27240, g19790)
--	g29711 = AND(g2541, g29134)
--	g33904 = AND(g33321, g21059)
--	g24495 = AND(g6928, g23127)
--	g28268 = AND(g8572, g27990)
--	g31252 = AND(g29643, g20101)
--	g29327 = AND(g29070, g22156)
--	g26861 = AND(g25021, g25003)
--	g33252 = AND(g32155, g20064)
--	g13080 = AND(g6923, g11357)
--	g18558 = AND(g2803, g15277)
--	g28655 = AND(g27561, g20603)
--	g30191 = AND(g28647, g23843)
--	g16233 = AND(g6137, g14251)
--	g29537 = AND(g28976, g22472)
--	g34191 = AND(g33713, g24404)
--	g16672 = AND(g6295, g15008)
--	g27822 = AND(g4157, g25893)
--	I27539 = AND(g28040, g24135, g24136, g24137)
--	g26389 = AND(g19949, g25553)
--	g18893 = AND(g16215, g16030)
--	g25981 = AND(g2051, g25007)
--	g24687 = AND(g5827, g23666)
--	I31011 = AND(g30735, g31797, g32471, g32472)
--	g27266 = AND(g26789, g26770)
--	g26612 = AND(g901, g24407)
--	I27538 = AND(g21209, g24132, g24133, g24134)
--	g26388 = AND(g19595, g25552)
--	g18544 = AND(g2791, g15277)
--	g26324 = AND(g2661, g25439)
--	g32428 = AND(g31133, g16261)
--	g29606 = AND(g28480, g8011)
--	g21024 = AND(g16306, g4871)
--	g18713 = AND(g4836, g15915)
--	g13461 = AND(g2719, g11819)
--	g22084 = AND(g6291, g19210)
--	g31183 = AND(g30249, g25174)
--	g26251 = AND(g1988, g25341)
--	g22110 = AND(g15167, g19277)
--	g24643 = AND(g22636, g19696)
--	g26272 = AND(g2036, g25470)
--	g33847 = AND(g33260, g20383)
--	g21860 = AND(g3945, g21070)
--	g16513 = AND(g8345, g13708)
--	g28694 = AND(g27579, g20664)
--	g29750 = AND(g28296, g23215)
--	g29982 = AND(g23656, g28998)
--	g29381 = AND(g28135, g19399)
--	g18610 = AND(g15088, g17059)
--	g34861 = AND(g16540, g34827)
--	g30247 = AND(g28735, g23937)
--	g18705 = AND(g4801, g16782)
--	g13887 = AND(g5204, g12402)
--	g25990 = AND(g9461, g25017)
--	g23497 = AND(g20169, g20569)
--	g33509 = AND(g32809, I31241, I31242)
--	g24669 = AND(g22653, g19742)
--	g31933 = AND(g939, g30735)
--	g30926 = AND(g29903, g21163)
--	g30045 = AND(g29200, g12419)
--	g18255 = AND(g1087, g16897)
--	g18189 = AND(g812, g17821)
--	g27588 = AND(g26690, g26673)
--	g15779 = AND(g13909, g11214)
--	g18679 = AND(g4633, g15758)
--	g31508 = AND(g29813, g23459)
--	g34389 = AND(g34170, g20715)
--	g17321 = AND(g1418, g13105)
--	I31112 = AND(g32617, g32618, g32619, g32620)
--	g34045 = AND(g33766, g22942)
--	g30612 = AND(g26338, g29597)
--	g33508 = AND(g32802, I31236, I31237)
--	g24668 = AND(g11754, g22979)
--	g21700 = AND(g150, g20283)
--	g30099 = AND(g28549, g20776)
--	g33872 = AND(g33282, g20548)
--	g18270 = AND(g1291, g16031)
--	g29796 = AND(g28345, g23258)
--	g17179 = AND(g1041, g13211)
--	g24392 = AND(g3115, g23067)
--	g22685 = AND(g11891, g20192)
--	g18188 = AND(g807, g17328)
--	g18124 = AND(g102, g16886)
--	g21987 = AND(g5579, g19074)
--	g18678 = AND(g66, g15758)
--	g34388 = AND(g10802, g34062)
--	g16026 = AND(g854, g14065)
--	g28557 = AND(g27772, g15647)
--	g34324 = AND(g14064, g34161)
--	g15081 = AND(g2689, g12983)
--	g13393 = AND(g703, g11048)
--	g16212 = AND(g6167, g14321)
--	g24195 = AND(g74, g22722)
--	g28210 = AND(g9229, g27554)
--	g32317 = AND(g5507, g31542)
--	g27119 = AND(g25877, g22542)
--	g30098 = AND(g28548, g20774)
--	g34701 = AND(g34536, g20179)
--	g10721 = AND(g3288, g6875, g3274, g8481)
--	g20559 = AND(g336, g15831)
--	g30251 = AND(g28745, g23940)
--	g34534 = AND(g34321, g19743)
--	g23658 = AND(g14687, g20852)
--	g30272 = AND(g28814, g23982)
--	g34098 = AND(g33744, g9104, g18957)
--	g19206 = AND(g460, g16206)
--	g15786 = AND(g13940, g11233)
--	g18460 = AND(g2351, g15224)
--	g18686 = AND(g4659, g15885)
--	g24559 = AND(g22993, g19567)
--	g18383 = AND(g1950, g15171)
--	g29840 = AND(g2153, g29056)
--	g24488 = AND(g6905, g23082)
--	I31096 = AND(g31376, g31812, g32594, g32595)
--	g24016 = AND(g14528, g21610)
--	g27118 = AND(g26055, g16529)
--	g22417 = AND(g7753, g9285, g21186)
--	g11960 = AND(g2495, g7424)
--	g32129 = AND(g31658, g29955)
--	g21943 = AND(g5240, g18997)
--	g25832 = AND(g8219, g24625)
--	g21296 = AND(g7879, g16072)
--	g24558 = AND(g22516, g19566)
--	g18267 = AND(g1266, g16000)
--	g18294 = AND(g15072, g16449)
--	g27616 = AND(g26349, g20449)
--	g26871 = AND(g25038, g25020)
--	g17654 = AND(g962, g13284)
--	g32128 = AND(g31631, g29953)
--	I17575 = AND(g13156, g11450, g6756)
--	g27313 = AND(g1982, g26701)
--	g29192 = AND(g27163, g10290)
--	g30032 = AND(g29072, g9326)
--	g21969 = AND(g5373, g21514)
--	g26360 = AND(g10589, g25533)
--	g25573 = AND(I24704, I24705)
--	g30140 = AND(g28600, g23749)
--	g27276 = AND(g9750, g26607)
--	g27285 = AND(g9912, g26632)
--	g29522 = AND(g28923, g22369)
--	g32323 = AND(g31311, g20610)
--	g24865 = AND(g11323, g23253)
--	g29663 = AND(g1950, g28693)
--	g34140 = AND(g33931, g23802)
--	g22762 = AND(g9305, g20645)
--	g15651 = AND(g429, g13414)
--	g21968 = AND(g5459, g21514)
--	g10655 = AND(g8440, g3423)
--	g15672 = AND(g433, g13458)
--	g27305 = AND(g10041, g26683)
--	g25926 = AND(g25005, g24839)
--	g24713 = AND(g5831, g23666)
--	g25045 = AND(g17525, g23448)
--	g18219 = AND(g969, g16100)
--	g27254 = AND(g25935, g19688)
--	g30061 = AND(g1036, g28188)
--	g33311 = AND(g31942, g12925)
--	g21855 = AND(g3925, g21070)
--	g34061 = AND(g33800, g23076)
--	g14180 = AND(g872, g10632)
--	g23855 = AND(g4112, g19455)
--	g22216 = AND(g13660, g20000)
--	g18218 = AND(g1008, g16100)
--	g21870 = AND(g4093, g19801)
--	I17606 = AND(g14988, g11450, g6756)
--	g28601 = AND(g27506, g20514)
--	g28677 = AND(g27571, g20635)
--	g27036 = AND(g26329, g11038)
--	g29553 = AND(g2437, g28911)
--	g26629 = AND(g14173, g24418)
--	g27177 = AND(g25997, g16651)
--	g27560 = AND(g26299, g20191)
--	g34871 = AND(g34823, g19908)
--	g24189 = AND(g324, g22722)
--	g31756 = AND(g30114, g23942)
--	g24679 = AND(g13289, g22985)
--	g11244 = AND(g8346, g8566)
--	g29949 = AND(g23575, g28924)
--	g32232 = AND(g31241, g20266)
--	g20188 = AND(g5849, g17772)
--	g18160 = AND(g645, g17433)
--	g29326 = AND(g29105, g22155)
--	g10838 = AND(g7738, g5527, g5535)
--	g28143 = AND(g27344, g26083)
--	g31780 = AND(g30163, g23999)
--	g25462 = AND(g6404, g22300, I24585)
--	g24188 = AND(g316, g22722)
--	g22117 = AND(g6597, g19277)
--	g29536 = AND(g28969, g22432)
--	g22000 = AND(g5727, g21562)
--	g21867 = AND(g4082, g19801)
--	g18455 = AND(g2327, g15224)
--	g24686 = AND(g5485, g23630)
--	g24939 = AND(g23771, g21012)
--	g29757 = AND(g28305, g23221)
--	I31317 = AND(g32914, g32915, g32916, g32917)
--	g33350 = AND(g32235, g20702)
--	g32261 = AND(g31251, g20386)
--	g18617 = AND(g3462, g17062)
--	g18470 = AND(g2403, g15224)
--	g20093 = AND(g15372, g14584)
--	g33820 = AND(g33075, g26830)
--	g29621 = AND(g2449, g28994)
--	I24576 = AND(g5390, g5396, g9792)
--	I24585 = AND(g9621, g9892, g6439)
--	g10619 = AND(g3080, g7907)
--	g21714 = AND(g278, g20283)
--	g23581 = AND(g20183, g11900)
--	g24294 = AND(g4452, g22550)
--	g31152 = AND(g10039, g30067)
--	g25061 = AND(g17586, g23461)
--	I31002 = AND(g32459, g32460, g32461, g32462)
--	g18201 = AND(g15061, g15938)
--	g33846 = AND(g33259, g20380)
--	I31057 = AND(g32538, g32539, g32540, g32541)
--	g21707 = AND(g191, g20283)
--	g21819 = AND(g3614, g20924)
--	g29564 = AND(g1882, g28896)
--	g18277 = AND(g1312, g16136)
--	g14210 = AND(g4392, g10590)
--	g21910 = AND(g5016, g21468)
--	g26147 = AND(g6513, g25133)
--	g30220 = AND(g28699, g23888)
--	g28666 = AND(g27567, g20625)
--	g33731 = AND(g33116, g19520)
--	g28217 = AND(g27733, g23391)
--	g22123 = AND(g6609, g19277)
--	g21818 = AND(g3610, g20924)
--	g17747 = AND(g6772, g11592, g11640, I18740)
--	g21979 = AND(g5559, g19074)
--	g16896 = AND(g262, g13120)
--	g27665 = AND(g26872, g23519)
--	g30246 = AND(g28734, g23936)
--	g25871 = AND(g8334, g24804)
--	g20875 = AND(g16281, g4681)
--	g18595 = AND(g2927, g16349)
--	g28478 = AND(g27007, g12345)
--	g18467 = AND(g2380, g15224)
--	g18494 = AND(g2527, g15426)
--	g19500 = AND(g504, g16712)
--	g24219 = AND(g225, g22594)
--	g26858 = AND(g2970, g24540)
--	g21978 = AND(g5551, g19074)
--	g11967 = AND(g311, g7802)
--	g18623 = AND(g3484, g17062)
--	g20218 = AND(g6541, g17815)
--	g30071 = AND(g29184, g12975)
--	g17123 = AND(g225, g13209)
--	g24218 = AND(g872, g22594)
--	g21986 = AND(g5575, g19074)
--	g34071 = AND(g8854, g33799)
--	g18782 = AND(g5835, g18065)
--	g27485 = AND(g26519, g17644)
--	g28556 = AND(g27431, g20374)
--	g29509 = AND(g1600, g28755)
--	g32316 = AND(g31307, g23522)
--	g33405 = AND(g32354, g21398)
--	g21741 = AND(g15086, g20330)
--	g26844 = AND(g25261, g21418)
--	g18419 = AND(g2051, g15373)
--	g27454 = AND(g26488, g17602)
--	g26394 = AND(g22530, g25560)
--	g18352 = AND(g1798, g17955)
--	g29634 = AND(g2108, g29121)
--	g29851 = AND(g1668, g29079)
--	g29872 = AND(g28401, g23333)
--	g28223 = AND(g27338, g17194)
--	g15104 = AND(g6955, g14454)
--	g34754 = AND(g34677, g19602)
--	g18155 = AND(g15056, g17533)
--	g21067 = AND(g10085, g17625)
--	g18418 = AND(g2122, g15373)
--	g18822 = AND(g6723, g15680)
--	g30825 = AND(g29814, g22332)
--	g19613 = AND(g1437, g16713)
--	g32056 = AND(g27271, g31021)
--	g18266 = AND(g1274, g16000)
--	g11010 = AND(g4698, g8933)
--	g34859 = AND(g16540, g34820)
--	g18170 = AND(g661, g17433)
--	I31232 = AND(g32791, g32792, g32793, g32794)
--	g10677 = AND(g4141, g7611)
--	g22992 = AND(g1227, g19765)
--	g34370 = AND(g34067, g10554)
--	I24674 = AND(g19919, g24019, g24020, g24021)
--	g21801 = AND(g3554, g20924)
--	g28110 = AND(g27974, g18886)
--	g21735 = AND(g3057, g20330)
--	g21877 = AND(g6888, g19801)
--	g23801 = AND(g1448, g19362)
--	g34858 = AND(g16540, g34816)
--	g30151 = AND(g28607, g21249)
--	g30172 = AND(g28625, g21286)
--	g24915 = AND(g23087, g20158)
--	I31261 = AND(g30937, g31842, g32831, g32832)
--	g27594 = AND(g26721, g26694)
--	g28531 = AND(g27722, g15608)
--	g17391 = AND(g9556, g14378)
--	g22835 = AND(g15803, g19633)
--	g28178 = AND(g27019, g19397)
--	g18167 = AND(g718, g17433)
--	g18194 = AND(g843, g17821)
--	g18589 = AND(g2902, g16349)
--	g22014 = AND(g5805, g21562)
--	g34367 = AND(g7404, g34042)
--	g31787 = AND(g21281, g29385)
--	g34394 = AND(g34190, g21305)
--	g25071 = AND(g12804, g23478)
--	g33113 = AND(g31964, g22339)
--	g33787 = AND(g33103, g20595)
--	g32342 = AND(g6545, g31579)
--	g29574 = AND(g2016, g28931)
--	g31282 = AND(g30130, g27779)
--	g22007 = AND(g5770, g21562)
--	g15850 = AND(g3606, g14151)
--	g29205 = AND(g24117, I27523, I27524)
--	g18588 = AND(g2970, g16349)
--	g18524 = AND(g2681, g15509)
--	g28676 = AND(g27570, g20632)
--	g32145 = AND(g31609, g29977)
--	g14791 = AND(g1146, g10909)
--	g32031 = AND(g31372, g13464)
--	g24467 = AND(g13761, g23047)
--	g27519 = AND(g26488, g17710)
--	g33357 = AND(g32247, g20775)
--	g27185 = AND(g26190, g8302, g1917)
--	g25147 = AND(g20202, g23542)
--	g32199 = AND(g30916, g25506)
--	g18401 = AND(g2036, g15373)
--	g28654 = AND(g1030, g27108)
--	g33105 = AND(g26298, g32138)
--	g14168 = AND(g887, g10632)
--	g18477 = AND(g2429, g15426)
--	g26203 = AND(g1632, g25337)
--	g33743 = AND(g33119, g19574)
--	g16802 = AND(g5567, g14807)
--	g18119 = AND(g475, g17015)
--	g27518 = AND(g26488, g17709)
--	g27154 = AND(g26055, g16630)
--	g34319 = AND(g9535, g34156)
--	g32198 = AND(g4253, g31327)
--	g22116 = AND(g6589, g19277)
--	g16730 = AND(g5212, g14723)
--	g24984 = AND(g22929, g12818)
--	g18118 = AND(g471, g17015)
--	g21866 = AND(g4072, g19801)
--	g21917 = AND(g5092, g21468)
--	g30227 = AND(g28708, g23899)
--	g31769 = AND(g30141, g23986)
--	g23917 = AND(g1472, g19428)
--	g33640 = AND(g33387, g18831)
--	g26281 = AND(g24688, g8812, g8778, g8757)
--	g32330 = AND(g31320, g20631)
--	g29592 = AND(g28469, g11832)
--	g30059 = AND(g28106, g12467)
--	g22720 = AND(g9253, g20619)
--	I31316 = AND(g29385, g32911, g32912, g32913)
--	g30025 = AND(g28492, g23502)
--	g25151 = AND(g17719, g23549)
--	g16765 = AND(g6581, g15045)
--	g15716 = AND(g468, g13437)
--	g18749 = AND(g5148, g17847)
--	g22041 = AND(g5957, g19147)
--	g26301 = AND(g2145, g25244)
--	g13656 = AND(g278, g11144)
--	g18616 = AND(g6875, g17200)
--	g18313 = AND(g1430, g16931)
--	g33803 = AND(g33231, g20071)
--	g24822 = AND(g3010, g23534, I24003)
--	g26120 = AND(g9809, g25293)
--	g30058 = AND(g29180, g12950)
--	g16690 = AND(g8399, g13867)
--	g11144 = AND(g239, g8136, g246, I14198)
--	g18748 = AND(g5142, g17847)
--	g8643 = AND(g2927, g2922)
--	g25367 = AND(g6946, g22407)
--	I31056 = AND(g30735, g31805, g32536, g32537)
--	g21706 = AND(g222, g20283)
--	g18276 = AND(g1351, g16136)
--	g18285 = AND(g1395, g16164)
--	g29350 = AND(g4939, g28395)
--	g26146 = AND(g9892, g25334)
--	g30203 = AND(g28668, g23864)
--	g18704 = AND(g4793, g16782)
--	g34203 = AND(g33726, g24537)
--	g18305 = AND(g1521, g16489)
--	g33881 = AND(g33292, g20586)
--	g30044 = AND(g29174, g12944)
--	g18254 = AND(g1236, g16897)
--	g18809 = AND(g7074, g15656)
--	g21923 = AND(g5029, g21468)
--	g22340 = AND(g19605, g13522)
--	g32161 = AND(g3151, g31154)
--	g22035 = AND(g5933, g19147)
--	g28587 = AND(g27487, g20498)
--	g26290 = AND(g2595, g25498)
--	g18466 = AND(g2389, g15224)
--	g23280 = AND(g19417, g20146)
--	g27215 = AND(g26055, g16724)
--	g27501 = AND(g26400, g17673)
--	g15112 = AND(g4284, g14454)
--	I31271 = AND(g29385, g32846, g32847, g32848)
--	g30281 = AND(g28850, g23992)
--	g18808 = AND(g6390, g15656)
--	g25420 = AND(g6058, g22220, I24555)
--	g24194 = AND(g106, g22722)
--	g24589 = AND(g5471, g23630)
--	g34281 = AND(g34043, g19276)
--	g29731 = AND(g2089, g29118)
--	g22142 = AND(g7957, g19140)
--	g27439 = AND(g232, g26831)
--	g34301 = AND(g34064, g19415)
--	g18177 = AND(g749, g17328)
--	g18560 = AND(g2837, g15277)
--	g30120 = AND(g28576, g21051)
--	g28543 = AND(g27735, g15628)
--	g24588 = AND(g5142, g23590)
--	g32087 = AND(g1291, g30825)
--	g34120 = AND(g33930, g25158)
--	I31342 = AND(g32949, g32950, g32951, g32952)
--	g32258 = AND(g31624, g30303)
--	g28117 = AND(g8075, g27245)
--	g18642 = AND(g15097, g17096)
--	g25059 = AND(g20870, g23460)
--	g33890 = AND(g33310, g20659)
--	g19788 = AND(g9983, g17216)
--	I31031 = AND(g30614, g31801, g32499, g32500)
--	g16128 = AND(g14333, g14166)
--	g34146 = AND(g33788, g20091)
--	g34738 = AND(g34660, g33442)
--	g33249 = AND(g32144, g20026)
--	g34562 = AND(g34369, g17411)
--	g28569 = AND(g27453, g20433)
--	g21066 = AND(g10043, g17625)
--	g25058 = AND(g23276, g20513)
--	g16245 = AND(g14278, g14708)
--	g32043 = AND(g31482, g16173)
--	g33482 = AND(g32614, I31106, I31107)
--	g32244 = AND(g31609, g30297)
--	g31710 = AND(g29814, g19128)
--	g33248 = AND(g32131, g19996)
--	g10676 = AND(g8506, g3774)
--	I27514 = AND(g24091, g24092, g24093, g24094)
--	g18733 = AND(g15141, g16877)
--	g27083 = AND(g25819, g22456)
--	g27348 = AND(g26488, g17392)
--	g33710 = AND(g14037, g33246)
--	g22130 = AND(g6637, g19277)
--	g27284 = AND(g9908, g26631)
--	g24864 = AND(g11201, g22305)
--	g22193 = AND(g19880, g20682)
--	g28242 = AND(g27769, g23626)
--	g21876 = AND(g4119, g19801)
--	g21885 = AND(g4122, g19801)
--	g26547 = AND(g13283, g25027)
--	g10654 = AND(g3085, g8434)
--	g11023 = AND(g9669, g5084)
--	g15857 = AND(g3199, g14038)
--	g23885 = AND(g4132, g19513)
--	g27304 = AND(g2273, g26682)
--	g24749 = AND(g17511, g22432)
--	g32069 = AND(g10878, g30735)
--	g12284 = AND(g1532, g7557)
--	g14654 = AND(g7178, g10476)
--	g24313 = AND(g4504, g22228)
--	g22165 = AND(g15594, g18903)
--	g18630 = AND(g3689, g17226)
--	g21854 = AND(g3921, g21070)
--	g15793 = AND(g3219, g13873)
--	g18693 = AND(g4717, g16053)
--	g23854 = AND(g4093, g19506)
--	g31778 = AND(g21369, g29385)
--	g24748 = AND(g17656, g22457)
--	g26226 = AND(g24688, g8812, g10658, g10627)
--	g32068 = AND(g31515, g10862)
--	g33081 = AND(g32388, g18875)
--	g17193 = AND(g2504, g13023)
--	g21763 = AND(g3223, g20785)
--	g18166 = AND(g655, g17433)
--	g24285 = AND(g4388, g22550)
--	g25902 = AND(g24398, g19373)
--	g18665 = AND(g4584, g17367)
--	I31132 = AND(g32645, g32646, g32647, g32648)
--	g31786 = AND(g30189, g24010)
--	g25957 = AND(g17190, g24960)
--	g24704 = AND(g17593, g22384)
--	g25377 = AND(g5712, g22210, I24530)
--	g33786 = AND(g33130, g20572)
--	g24305 = AND(g4477, g22228)
--	g16737 = AND(g6645, g15042)
--	g26572 = AND(g7443, g24439)
--	g22006 = AND(g5767, g21562)
--	g28639 = AND(g27767, g20597)
--	g24900 = AND(g3752, g23582, I24067)
--	g33647 = AND(g33390, g18878)
--	g32337 = AND(g31465, g20663)
--	g27139 = AND(g26055, g16608)
--	g28293 = AND(g7424, g2495, g27474)
--	g33356 = AND(g32245, g20772)
--	g22863 = AND(g9547, g20388)
--	g27653 = AND(g26549, g15562)
--	g28638 = AND(g27551, g20583)
--	g32171 = AND(g31706, g27800)
--	I31161 = AND(g30614, g31824, g32687, g32688)
--	g18476 = AND(g2433, g15426)
--	g18485 = AND(g2465, g15426)
--	g29787 = AND(g28334, g23249)
--	g26127 = AND(g2236, g25119)
--	g27138 = AND(g26055, g16607)
--	g28265 = AND(g11367, g27989)
--	g34661 = AND(g34575, g18907)
--	g18555 = AND(g2834, g15277)
--	g18454 = AND(g2303, g15224)
--	g25290 = AND(g5022, g22173, I24482)
--	g14216 = AND(g7631, g10608)
--	g21916 = AND(g5084, g21468)
--	g30226 = AND(g28707, g23898)
--	g18570 = AND(g2848, g16349)
--	g18712 = AND(g4843, g15915)
--	g33233 = AND(g32094, g23005)
--	g31182 = AND(g30240, g20682)
--	g31672 = AND(g29814, g19050)
--	g27333 = AND(g10180, g26765)
--	g24642 = AND(g8290, g22898)
--	g34226 = AND(g33914, g21467)
--	g14587 = AND(g10584, g10567)
--	g29743 = AND(g28206, g10233)
--	I31087 = AND(g32580, g32581, g32582, g32583)
--	g34715 = AND(g34570, g33375)
--	g34481 = AND(g34404, g18916)
--	g23314 = AND(g9104, g19200)
--	g32425 = AND(g31668, g21604)
--	g26103 = AND(g2185, g25100)
--	g34572 = AND(g34387, g33326)
--	g10543 = AND(g8238, g437)
--	g26095 = AND(g11923, g25090)
--	g27963 = AND(g25952, g16047)
--	g23076 = AND(g19128, g9104)
--	g29640 = AND(g28498, g8125)
--	g25366 = AND(g7733, g22406)
--	g29769 = AND(g28319, g23237)
--	g18239 = AND(g1135, g16326)
--	g21721 = AND(g385, g21037)
--	g33331 = AND(g32216, g20607)
--	g27664 = AND(g1024, g25911)
--	g18567 = AND(g2894, g16349)
--	g18594 = AND(g12858, g16349)
--	g31513 = AND(g2606, g29318)
--	g32010 = AND(g31785, g22303)
--	g33513 = AND(g32837, I31261, I31262)
--	g29803 = AND(g28414, g26836)
--	g18238 = AND(g1152, g16326)
--	g26181 = AND(g2652, g25157)
--	g26671 = AND(g316, g24429)
--	g28586 = AND(g27484, g20497)
--	g24630 = AND(g23255, g14149)
--	g31961 = AND(g31751, g22154)
--	g33897 = AND(g33315, g20777)
--	g17781 = AND(g6772, g11592, g6789, I18785)
--	g31505 = AND(g30195, g24379)
--	g28442 = AND(g27278, g20072)
--	g33505 = AND(g32779, I31221, I31222)
--	g18382 = AND(g1936, g15171)
--	g24009 = AND(g19671, g10971)
--	g33404 = AND(g32353, g21397)
--	g29881 = AND(g2040, g29150)
--	g21773 = AND(g3263, g20785)
--	g18519 = AND(g2648, g15509)
--	g11016 = AND(g4888, g8984)
--	g21942 = AND(g5236, g18997)
--	g13525 = AND(g10019, g11911)
--	g18176 = AND(g732, g17328)
--	g18185 = AND(g790, g17328)
--	g22063 = AND(g6109, g21611)
--	g18675 = AND(g4349, g15758)
--	g34385 = AND(g34168, g20642)
--	g33717 = AND(g14092, g33306)
--	g24008 = AND(g7909, g19502)
--	g32086 = AND(g7597, g30735)
--	g30095 = AND(g28545, g20768)
--	g31212 = AND(g20028, g29669)
--	g28116 = AND(g27366, g26183)
--	g18518 = AND(g2657, g15509)
--	g18154 = AND(g622, g17533)
--	g27312 = AND(g12019, g26700)
--	g24892 = AND(g11559, g23264)
--	g26190 = AND(g25357, g11724, g7586, g11686)
--	g24485 = AND(g10710, g22319)
--	g24476 = AND(g18879, g22330)
--	I31337 = AND(g32942, g32943, g32944, g32945)
--	g16611 = AND(g5583, g14727)
--	g27115 = AND(g26026, g16526)
--	g11893 = AND(g1668, g7268)
--	g13830 = AND(g11543, g11424, g11395, I16143)
--	g22873 = AND(g19854, g19683)
--	g25551 = AND(g23822, g21511)
--	g18637 = AND(g3821, g17096)
--	g25572 = AND(I24699, I24700)
--	I31171 = AND(g31528, g31826, g32701, g32702)
--	g30181 = AND(g28636, g23821)
--	g30671 = AND(g29319, g22317)
--	g18935 = AND(g4322, g15574)
--	g32322 = AND(g31308, g20605)
--	g24555 = AND(g23184, g21024)
--	g29662 = AND(g1848, g29049)
--	g9217 = AND(g632, g626)
--	g21734 = AND(g3040, g20330)
--	g32159 = AND(g31658, g30040)
--	g24712 = AND(g19592, g23001)
--	g29890 = AND(g28419, g23355)
--	g24914 = AND(g8721, g23301)
--	g21839 = AND(g3763, g20453)
--	g21930 = AND(g5180, g18997)
--	g25127 = AND(g13997, g23524)
--	g21993 = AND(g5603, g19074)
--	g32158 = AND(g31658, g30022)
--	g22209 = AND(g19907, g20751)
--	g15856 = AND(g9056, g14223)
--	g15995 = AND(g13314, g1157, g10666)
--	g33723 = AND(g14091, g33299)
--	g28237 = AND(g9492, g27597)
--	g21838 = AND(g3747, g20453)
--	g22834 = AND(g102, g19630)
--	g15880 = AND(g3211, g13980)
--	g31149 = AND(g29508, g23021)
--	g21965 = AND(g15149, g21514)
--	g26088 = AND(g6545, g25080)
--	g26024 = AND(g2619, g25039)
--	g22208 = AND(g19906, g20739)
--	g29710 = AND(g2380, g29094)
--	g28035 = AND(g24103, I26530, I26531)
--	g29552 = AND(g2223, g28579)
--	g33433 = AND(g32238, g29694)
--	g23131 = AND(g13919, g19930)
--	g32295 = AND(g27931, g31376)
--	g10841 = AND(g8509, g8567)
--	g29204 = AND(g24110, I27518, I27519)
--	g31148 = AND(g2661, g30055)
--	g30190 = AND(g28646, g23842)
--	g13042 = AND(g433, g11048)
--	g16199 = AND(g3614, g14051)
--	g18215 = AND(g943, g15979)
--	g25103 = AND(g4927, g22908)
--	g27184 = AND(g26628, g13756)
--	g16736 = AND(g6303, g15036)
--	g18501 = AND(g12854, g15509)
--	g18729 = AND(g15139, g16821)
--	g22021 = AND(g5869, g19147)
--	g27674 = AND(g26873, g23543)
--	g25980 = AND(g1926, g25006)
--	g18577 = AND(g2988, g16349)
--	g33104 = AND(g26296, g32137)
--	g25095 = AND(g23319, g20556)
--	g33811 = AND(g33439, g17573)
--	g33646 = AND(g33389, g18876)
--	g19767 = AND(g16810, g14203)
--	g32336 = AND(g31596, g11842)
--	g34520 = AND(g34294, g19505)
--	g23619 = AND(g19453, g13045)
--	g33343 = AND(g32227, g20665)
--	g21557 = AND(g12980, g15674)
--	g18728 = AND(g4939, g16821)
--	g18439 = AND(g2250, g18008)
--	g30089 = AND(g28538, g20709)
--	g24941 = AND(g23171, g20190)
--	g26126 = AND(g1959, g25118)
--	g30211 = AND(g28685, g23878)
--	g11939 = AND(g2361, g7380)
--	g23618 = AND(g19388, g11917)
--	g25181 = AND(g23405, g20696)
--	g34089 = AND(g22957, g9104, g33744)
--	g16843 = AND(g6251, g14864)
--	g18438 = AND(g2236, g18008)
--	g34211 = AND(g33891, g21349)
--	g26250 = AND(g1902, g25429)
--	g13383 = AND(g4765, g11797)
--	g24675 = AND(g17568, g22342)
--	g29647 = AND(g28934, g22457)
--	g30024 = AND(g28497, g23501)
--	g33369 = AND(g32277, g21060)
--	I24048 = AND(g3034, g3040, g8426)
--	g17726 = AND(g1467, g13315)
--	g16764 = AND(g6307, g14776)
--	g34088 = AND(g33736, g9104, g18957)
--	g13030 = AND(g429, g11048)
--	g22073 = AND(g6235, g19210)
--	g18349 = AND(g1768, g17955)
--	g14586 = AND(g11953, g11970)
--	g13294 = AND(g1564, g11513)
--	I31086 = AND(g31554, g31811, g32578, g32579)
--	g29380 = AND(g28134, g19396)
--	g33368 = AND(g32275, g21057)
--	g34860 = AND(g16540, g34823)
--	g16869 = AND(g6259, g14902)
--	g27692 = AND(g26392, g20697)
--	g28130 = AND(g27353, g23063)
--	g28193 = AND(g8851, g27629)
--	g26339 = AND(g225, g24836)
--	g25931 = AND(g24574, g19477)
--	g18906 = AND(g13568, g16264)
--	g18348 = AND(g1744, g17955)
--	g24637 = AND(g16586, g22884)
--	g19521 = AND(g513, g16739)
--	g22122 = AND(g6601, g19277)
--	g12692 = AND(g10323, g3522, g3530)
--	g12761 = AND(g969, g7567)
--	g18284 = AND(g15071, g16164)
--	g16868 = AND(g5813, g14297)
--	g34497 = AND(g34275, g33072)
--	g28165 = AND(g27018, g22455)
--	g28523 = AND(g27704, g15585)
--	g18304 = AND(g1542, g16489)
--	g29182 = AND(g27163, g12730)
--	g29651 = AND(g2537, g29134)
--	g33412 = AND(g32362, g21411)
--	I31322 = AND(g32921, g32922, g32923, g32924)
--	g16161 = AND(g5841, g14297)
--	g15611 = AND(g471, g13437)
--	g15722 = AND(g464, g13437)
--	g18622 = AND(g3480, g17062)
--	g22034 = AND(g5929, g19147)
--	g15080 = AND(g12855, g12983)
--	g18566 = AND(g2860, g16349)
--	g30126 = AND(g28582, g21058)
--	g14615 = AND(g10604, g10587)
--	g27214 = AND(g26026, g13901)
--	g34700 = AND(g34535, g20129)
--	g31229 = AND(g30288, g23949)
--	g10720 = AND(g2704, g10219, g2689)
--	g21815 = AND(g3598, g20924)
--	g30250 = AND(g28744, g23939)
--	g27329 = AND(g12052, g26743)
--	g32309 = AND(g5160, g31528)
--	g27207 = AND(g26055, g16692)
--	g33896 = AND(g33314, g20771)
--	g31228 = AND(g20028, g29713)
--	g27539 = AND(g26576, g17745)
--	g29331 = AND(g29143, g22169)
--	g32224 = AND(g4300, g31327)
--	g34658 = AND(g34574, g18896)
--	g23187 = AND(g13989, g20010)
--	g26855 = AND(g2960, g24535)
--	g21975 = AND(g5523, g19074)
--	g27328 = AND(g12482, g26736)
--	g25089 = AND(g23317, g20553)
--	g32308 = AND(g31293, g23503)
--	g20215 = AND(g16479, g10476)
--	g29513 = AND(g28448, g14095)
--	g18139 = AND(g542, g17249)
--	g27538 = AND(g26549, g14744)
--	g18653 = AND(g4176, g16249)
--	g24501 = AND(g14000, g23182)
--	g24729 = AND(g22719, g23018)
--	g25088 = AND(g17601, g23491)
--	g17292 = AND(g1075, g13093)
--	g11160 = AND(g6336, g7074, g6322, g10003)
--	g17153 = AND(g6311, g14943)
--	I24033 = AND(g8219, g8443, g3747)
--	g18138 = AND(g546, g17249)
--	I26531 = AND(g24099, g24100, g24101, g24102)
--	g21937 = AND(g5208, g18997)
--	I17552 = AND(g13156, g11450, g11498)
--	g34338 = AND(g34099, g19905)
--	g24728 = AND(g16513, g23017)
--	g16244 = AND(g11547, g11592, g6789, I17585)
--	I31336 = AND(g31672, g31855, g32940, g32941)
--	g14035 = AND(g699, g11048)
--	g15650 = AND(g8362, g13413)
--	g34969 = AND(g34960, g19570)
--	g10684 = AND(g7998, g411)
--	g28703 = AND(g27925, g20680)
--	g18636 = AND(g3817, g17096)
--	g18415 = AND(g2108, g15373)
--	g31310 = AND(g30157, g27886)
--	g18333 = AND(g1691, g17873)
--	g30060 = AND(g29146, g10581)
--	g21791 = AND(g3368, g20391)
--	g28253 = AND(g23719, g27700)
--	g21884 = AND(g4104, g19801)
--	g11915 = AND(g1802, g7315)
--	g34968 = AND(g34952, g23203)
--	g23884 = AND(g4119, g19510)
--	g30197 = AND(g28661, g23859)
--	g31959 = AND(g4907, g30673)
--	g33379 = AND(g30984, g32364)
--	g19462 = AND(g7850, g14182, g14177, g16646)
--	g25126 = AND(g16839, g23523)
--	g25987 = AND(g9501, g25015)
--	I31017 = AND(g32480, g32481, g32482, g32483)
--	g13277 = AND(g3195, g11432)
--	g28236 = AND(g8515, g27971)
--	g34870 = AND(g34820, g19882)
--	g34527 = AND(g34303, g19603)
--	g24284 = AND(g4375, g22550)
--	g18664 = AND(g4332, g17367)
--	g27235 = AND(g25910, g19579)
--	g24304 = AND(g12875, g22228)
--	g26819 = AND(g106, g24490)
--	g27683 = AND(g25770, g23567)
--	g24622 = AND(g19856, g22866)
--	g33742 = AND(g7828, g33142, I31600)
--	g26257 = AND(g4253, g25197)
--	g31944 = AND(g31745, g22146)
--	g11037 = AND(g6128, g9184)
--	g18576 = AND(g2868, g16349)
--	g18585 = AND(g2960, g16349)
--	g14193 = AND(g7178, g10590)
--	g18484 = AND(g2491, g15426)
--	g22109 = AND(g6455, g18833)
--	g32260 = AND(g31250, g20385)
--	g28264 = AND(g7315, g1802, g27416)
--	g34503 = AND(g34278, g19437)
--	g34867 = AND(g34826, g20145)
--	g25969 = AND(g9310, g24987)
--	g18554 = AND(g2831, g15277)
--	g29620 = AND(g2399, g29097)
--	g33681 = AND(g33129, g7991)
--	g22108 = AND(g6439, g18833)
--	g18609 = AND(g3147, g16987)
--	g27414 = AND(g255, g26827)
--	g32195 = AND(g30734, g25451)
--	g24139 = AND(g17619, g21653)
--	g25968 = AND(g25215, g20739)
--	g18312 = AND(g1579, g16931)
--	g33802 = AND(g33097, g14545)
--	g33429 = AND(g32231, g29676)
--	g33857 = AND(g33267, g20445)
--	g29646 = AND(g1816, g28675)
--	g30315 = AND(g29182, g7028, g5644)
--	g34581 = AND(g22864, g34312)
--	g18608 = AND(g15087, g16987)
--	g27407 = AND(g26488, g17522)
--	g18115 = AND(g460, g17015)
--	I27534 = AND(g28039, g24128, g24129, g24130)
--	g33730 = AND(g7202, g4621, g33127, g4633)
--	g32016 = AND(g8522, g31138)
--	g33428 = AND(g32230, g29672)
--	g34707 = AND(g34544, g20579)
--	g30202 = AND(g28667, g23863)
--	g25870 = AND(g24840, g16182)
--	g30257 = AND(g28750, g23952)
--	g25411 = AND(g5062, g23764, I24546)
--	g26094 = AND(g24936, g9664)
--	g31765 = AND(g30128, g23968)
--	g24415 = AND(g4760, g22869)
--	g7763 = AND(g2965, g2960)
--	g24333 = AND(g4512, g22228)
--	g29369 = AND(g28209, g22341)
--	g14222 = AND(g8655, g11826)
--	g21922 = AND(g5112, g21468)
--	g22982 = AND(g19535, g19747)
--	g30111 = AND(g28565, g20917)
--	g18745 = AND(g5128, g17847)
--	g33690 = AND(g33146, g16280)
--	g30070 = AND(g29167, g9529)
--	g34111 = AND(g33733, g22936)
--	g18799 = AND(g6181, g15348)
--	g22091 = AND(g6415, g18833)
--	g23531 = AND(g10760, g18930)
--	g13853 = AND(g4549, g10620)
--	g18813 = AND(g6513, g15483)
--	g30590 = AND(g18911, g29812)
--	g21740 = AND(g3085, g20330)
--	g16599 = AND(g6601, g15030)
--	g26019 = AND(g5507, g25032)
--	g25503 = AND(g6888, g22529)
--	g18798 = AND(g6177, g15348)
--	g28542 = AND(g27405, g20275)
--	g31504 = AND(g29370, g10553)
--	g28453 = AND(g27582, g10233)
--	g27206 = AND(g26055, g16691)
--	g33504 = AND(g32772, I31216, I31217)
--	g24664 = AND(g22652, g19741)
--	g29850 = AND(g28340, g24893)
--	g19911 = AND(g14707, g17748)
--	g34741 = AND(g8899, g34697)
--	g16598 = AND(g6283, g14899)
--	g15810 = AND(g3937, g14055)
--	g13524 = AND(g9995, g11910)
--	g17091 = AND(g8659, g12940)
--	g18184 = AND(g785, g17328)
--	g21953 = AND(g5377, g21514)
--	g18805 = AND(g6377, g15656)
--	g18674 = AND(g4340, g15758)
--	g23373 = AND(g13699, g20195)
--	g30094 = AND(g28544, g20767)
--	g27759 = AND(g22457, g25224, g26424, g26213)
--	g25581 = AND(g19338, g24150)
--	g25450 = AND(g6888, g22497)
--	g32042 = AND(g27244, g31070)
--	g21800 = AND(g3546, g20924)
--	g24484 = AND(g16288, g23208)
--	g29896 = AND(g2599, g29171)
--	g27114 = AND(g25997, g16523)
--	g32255 = AND(g31248, g20381)
--	g31129 = AND(g1968, g30017)
--	g32189 = AND(g30824, g25369)
--	g21936 = AND(g5200, g18997)
--	g18732 = AND(g4961, g16877)
--	g27435 = AND(g26549, g17585)
--	g18934 = AND(g3133, g16096)
--	g30735 = AND(g29814, g22319)
--	g24554 = AND(g22490, g19541)
--	g27107 = AND(g26055, g16514)
--	g32270 = AND(g31254, g20444)
--	g16125 = AND(g5152, g14238)
--	g16532 = AND(g5252, g14841)
--	g25818 = AND(g8124, g24605)
--	g28530 = AND(g27383, g20240)
--	g31128 = AND(g12187, g30016)
--	g32188 = AND(g27586, g31376)
--	g25979 = AND(g24517, g19650)
--	g28346 = AND(g27243, g19800)
--	g7251 = AND(g452, g392)
--	g24312 = AND(g4501, g22228)
--	g18692 = AND(g4732, g16053)
--	g18761 = AND(g5471, g17929)
--	g33245 = AND(g32125, g19961)
--	g24608 = AND(g6500, g23425)
--	g25978 = AND(g9391, g25001)
--	g13313 = AND(g475, g11048)
--	g15967 = AND(g3913, g14058)
--	g30196 = AND(g28659, g23858)
--	g31323 = AND(g30150, g27907)
--	g29582 = AND(g27766, g28608)
--	g31299 = AND(g30123, g27800)
--	g17192 = AND(g1677, g13022)
--	g34196 = AND(g33682, g24485)
--	g21762 = AND(g3219, g20785)
--	g21964 = AND(g5441, g21514)
--	g25986 = AND(g5160, g25013)
--	g32030 = AND(g4172, g30937)
--	g24921 = AND(g23721, g20739)
--	I31016 = AND(g30825, g31798, g32478, g32479)
--	g31298 = AND(g30169, g27886)
--	g34526 = AND(g34300, g19569)
--	g18400 = AND(g2012, g15373)
--	g10873 = AND(g3004, g9015)
--	g26077 = AND(g9607, g25233)
--	g24745 = AND(g650, g23550)
--	g29627 = AND(g28493, g11884)
--	g18214 = AND(g939, g15979)
--	g28292 = AND(g23781, g27762)
--	g29959 = AND(g28953, g12823)
--	g22862 = AND(g1570, g19673)
--	g28153 = AND(g26424, g22763, g27031)
--	g18329 = AND(g1612, g17873)
--	g25067 = AND(g4722, g22885)
--	g25094 = AND(g23318, g20554)
--	g18207 = AND(g925, g15938)
--	g26689 = AND(g15754, g24431)
--	g29378 = AND(g28137, g22493)
--	g13808 = AND(g4543, g10607)
--	g18539 = AND(g2763, g15277)
--	g11036 = AND(g9806, g5774)
--	g26280 = AND(g13051, g25248)
--	g18328 = AND(g1657, g17873)
--	g27263 = AND(g25940, g19713)
--	g21909 = AND(g5041, g21468)
--	g31232 = AND(g30294, g23972)
--	g25150 = AND(g17480, g23547)
--	g22040 = AND(g5953, g19147)
--	g25801 = AND(g8097, g24585)
--	g26300 = AND(g1968, g25341)
--	g34866 = AND(g34819, g20106)
--	g28136 = AND(g27382, g23135)
--	g18538 = AND(g2759, g15277)
--	g15079 = AND(g2151, g12955)
--	g27332 = AND(g12538, g26758)
--	g29603 = AND(g2265, g29060)
--	g24674 = AND(g446, g23496)
--	g29742 = AND(g28288, g10233)
--	g21908 = AND(g5037, g21468)
--	g15078 = AND(g10361, g12955)
--	g33697 = AND(g33160, g13330)
--	g30001 = AND(g28490, g23486)
--	g31995 = AND(g28274, g30569)
--	g33856 = AND(g33266, g20442)
--	g26102 = AND(g1825, g25099)
--	g12135 = AND(g9684, g9959)
--	g31261 = AND(g14754, g30259)
--	g26157 = AND(g2093, g25136)
--	g27406 = AND(g26488, g17521)
--	g34077 = AND(g22957, g9104, g33736)
--	g27962 = AND(g25954, g19597)
--	g27361 = AND(g26519, g17419)
--	g33880 = AND(g33290, g20568)
--	I31042 = AND(g32515, g32516, g32517, g32518)
--	g18241 = AND(g1183, g16431)
--	g34706 = AND(g34496, g10570)
--	g21747 = AND(g3061, g20330)
--	g32160 = AND(g31001, g22995)
--	g30256 = AND(g28749, g23947)
--	g25526 = AND(g23720, g21400)
--	g28164 = AND(g8651, g27528)
--	g26231 = AND(g1854, g25300)
--	g33512 = AND(g32830, I31256, I31257)
--	g14913 = AND(g1442, g10939)
--	g27500 = AND(g26400, g17672)
--	g29857 = AND(g28386, g23304)
--	g15817 = AND(g3921, g13929)
--	g14614 = AND(g11975, g11997)
--	g24761 = AND(g22751, g19852)
--	g19540 = AND(g1124, g15904)
--	g21814 = AND(g3594, g20924)
--	g18771 = AND(g5685, g15615)
--	g16023 = AND(g3813, g13584)
--	g16224 = AND(g14583, g14232)
--	g11166 = AND(g8363, g269, g8296, I14225)
--	g18235 = AND(g1141, g16326)
--	g21751 = AND(g3167, g20785)
--	g21807 = AND(g3566, g20924)
--	g21772 = AND(g3259, g20785)
--	g26854 = AND(g2868, g24534)
--	g15783 = AND(g3215, g14098)
--	g21974 = AND(g5517, g19074)
--	g22062 = AND(g6093, g21611)
--	g18683 = AND(g4674, g15885)
--	g25866 = AND(g3853, g24648)
--	g24400 = AND(g3466, g23112)
--	g27221 = AND(g26055, g16747)
--	g33831 = AND(g23088, g33149, g9104)
--	g28327 = AND(g27365, g19785)
--	g29549 = AND(g2012, g28900)
--	g34102 = AND(g33912, g23599)
--	g26511 = AND(g19265, g24364)
--	g34157 = AND(g33794, g20159)
--	g23639 = AND(g19050, g9104)
--	I31267 = AND(g32840, g32841, g32842, g32843)
--	g10565 = AND(g8182, g424)
--	g28537 = AND(g6832, g27089)
--	g31499 = AND(g29801, g23446)
--	g33499 = AND(g32737, I31191, I31192)
--	g14565 = AND(g11934, g11952)
--	g29548 = AND(g1798, g28575)
--	g23293 = AND(g9104, g19200)
--	g24329 = AND(g4462, g22228)
--	g30066 = AND(g28518, g20636)
--	g22851 = AND(g496, g19654)
--	g28108 = AND(g7975, g27237)
--	g30231 = AND(g28718, g23907)
--	g15823 = AND(g3945, g14116)
--	g34066 = AND(g33730, g19352)
--	g10034 = AND(g1521, g1500)
--	g25077 = AND(g23297, g20536)
--	g33498 = AND(g32730, I31186, I31187)
--	g23265 = AND(g20069, g20132)
--	g24328 = AND(g4567, g22228)
--	g28283 = AND(g7380, g2361, g27445)
--	g18515 = AND(g2643, g15509)
--	g23416 = AND(g20082, g20321)
--	g18414 = AND(g2102, g15373)
--	g31989 = AND(g31770, g22200)
--	g14641 = AND(g11994, g12020)
--	g28303 = AND(g7462, g2629, g27494)
--	g27106 = AND(g26026, g16512)
--	g21841 = AND(g3857, g21070)
--	g21992 = AND(g5599, g19074)
--	g34876 = AND(g34844, g20534)
--	g18407 = AND(g2016, g15373)
--	g25923 = AND(g24443, g19443)
--	g31988 = AND(g31768, g22199)
--	g33722 = AND(g33175, g19445)
--	g33924 = AND(g33335, g33346)
--	g32419 = AND(g4955, g31000)
--	g15966 = AND(g3462, g13555)
--	g28982 = AND(g27163, g12687, g20682, I27349)
--	g31271 = AND(g29706, g23300)
--	g12812 = AND(g518, g9158)
--	g34763 = AND(g34689, g19915)
--	g15631 = AND(g168, g13437)
--	g27033 = AND(g25767, g19273)
--	g27371 = AND(g26400, g17473)
--	g32418 = AND(g31126, g16239)
--	g26287 = AND(g2138, g25225)
--	g27234 = AND(g26055, g16814)
--	g25102 = AND(g4727, g22885)
--	g21835 = AND(g3802, g20453)
--	g32170 = AND(g31671, g27779)
--	g13567 = AND(g10102, g11948)
--	g22047 = AND(g6077, g21611)
--	g26307 = AND(g13070, g25288)
--	g26085 = AND(g11906, g25070)
--	g29626 = AND(g28584, g11415)
--	g33461 = AND(g32463, I31001, I31002)
--	g16669 = AND(g5611, g14993)
--	g33342 = AND(g32226, g20660)
--	g29323 = AND(g28539, g6905, g3639)
--	g23007 = AND(g681, g20248)
--	g31145 = AND(g9970, g30052)
--	g18441 = AND(g2246, g18008)
--	g18584 = AND(g2950, g16349)
--	g24771 = AND(g7028, g23605)
--	g18206 = AND(g918, g15938)
--	g29533 = AND(g28958, g22417)
--	g12795 = AND(g1312, g7601)
--	g16668 = AND(g5543, g14962)
--	g16842 = AND(g6279, g14861)
--	g17574 = AND(g9554, g14546)
--	g33887 = AND(g33298, g20615)
--	g18759 = AND(g5467, g17929)
--	g22051 = AND(g6105, g21611)
--	g22072 = AND(g6259, g19210)
--	g18725 = AND(g4912, g16077)
--	g32167 = AND(g3853, g31194)
--	g32194 = AND(g30601, g28436)
--	g25876 = AND(g3470, g24667)
--	g33529 = AND(g32953, I31341, I31342)
--	I31201 = AND(g31672, g31831, g32745, g32746)
--	g27507 = AND(g26549, g17683)
--	I31277 = AND(g32856, g32857, g32858, g32859)
--	g18114 = AND(g452, g17015)
--	g28192 = AND(g8891, g27415)
--	g18758 = AND(g7004, g15595)
--	g31528 = AND(g19050, g29814)
--	g26341 = AND(g24746, g20105)
--	g18435 = AND(g2173, g18008)
--	g33528 = AND(g32946, I31336, I31337)
--	g34287 = AND(g11370, g34124)
--	g19661 = AND(g5489, g16969)
--	g33843 = AND(g33256, g20325)
--	g21720 = AND(g376, g21037)
--	g33330 = AND(g32211, g20588)
--	g26156 = AND(g2028, g25135)
--	g18107 = AND(g429, g17015)
--	g27421 = AND(g8038, g26314, g9187, g9077)
--	g34085 = AND(g33761, g9104, g18957)
--	g28663 = AND(g27566, g20624)
--	g32401 = AND(g31116, g13432)
--	g34076 = AND(g33694, g19519)
--	g30596 = AND(g30279, g18947)
--	g26180 = AND(g2587, g25156)
--	g26670 = AND(g13385, g24428)
--	g21746 = AND(g3045, g20330)
--	g33365 = AND(g32267, g20994)
--	g32119 = AND(g31609, g29939)
--	g30243 = AND(g28731, g23929)
--	g31132 = AND(g29504, g22987)
--	g18744 = AND(g5124, g17847)
--	g34054 = AND(g33778, g22942)
--	g31960 = AND(g31749, g22153)
--	g33869 = AND(g33279, g20543)
--	g14537 = AND(g10550, g10529)
--	g18345 = AND(g1736, g17955)
--	g19715 = AND(g9679, g17120)
--	I31037 = AND(g32508, g32509, g32510, g32511)
--	g29856 = AND(g28385, g23303)
--	g17780 = AND(g6772, g11592, g11640, I18782)
--	g21465 = AND(g16155, g13663)
--	g18399 = AND(g2024, g15373)
--	g29880 = AND(g1936, g29149)
--	g33868 = AND(g33278, g20542)
--	g26839 = AND(g2988, g24516)
--	g27541 = AND(g26278, g23334)
--	g30269 = AND(g28778, g23970)
--	g22846 = AND(g9386, g20676)
--	g21983 = AND(g5555, g19074)
--	g28553 = AND(g27187, g10290)
--	g25456 = AND(g5752, g22210, I24579)
--	g18398 = AND(g2020, g15373)
--	g29512 = AND(g2161, g28793)
--	g32313 = AND(g31303, g23515)
--	I31352 = AND(g32963, g32964, g32965, g32966)
--	g21806 = AND(g3558, g20924)
--	g26838 = AND(g2860, g24515)
--	g18141 = AND(g568, g17533)
--	g30268 = AND(g28777, g23969)
--	g18652 = AND(g4172, g16249)
--	g18804 = AND(g15163, g15656)
--	g34341 = AND(g34101, g19952)
--	g25916 = AND(g24432, g19434)
--	g16610 = AND(g5260, g14918)
--	g16705 = AND(g6299, g15024)
--	g17152 = AND(g8635, g12997)
--	g31225 = AND(g30276, g21012)
--	g32276 = AND(g31646, g30313)
--	g27724 = AND(g22417, g25208, g26424, g26190)
--	g34655 = AND(g34573, g18885)
--	I31266 = AND(g31327, g31843, g32838, g32839)
--	g27359 = AND(g26488, g17416)
--	g30180 = AND(g28635, g23820)
--	g27325 = AND(g12478, g26724)
--	g30670 = AND(g11330, g29359)
--	g31471 = AND(g29754, g23399)
--	g32305 = AND(g31287, g20567)
--	g32053 = AND(g14176, g31509)
--	g33471 = AND(g32535, I31051, I31052)
--	g34180 = AND(g33716, g24373)
--	g33087 = AND(g32391, g18888)
--	g18263 = AND(g1249, g16000)
--	g32254 = AND(g31247, g20379)
--	g27535 = AND(g26519, g17737)
--	g26487 = AND(g15702, g24359)
--	g27434 = AND(g26549, g17584)
--	g27358 = AND(g26400, g17415)
--	g25076 = AND(g12805, g23479)
--	g25085 = AND(g4912, g22908)
--	g18332 = AND(g1677, g17873)
--	g19784 = AND(g2775, g15877)
--	g28252 = AND(g27159, g19682)
--	g12920 = AND(g1227, g10960)
--	g18135 = AND(g136, g17249)
--	g34335 = AND(g8461, g34197)
--	g25054 = AND(g12778, g23452)
--	g24725 = AND(g19587, g23012)
--	g30930 = AND(g29915, g23342)
--	g32036 = AND(g31469, g13486)
--	g27121 = AND(g136, g26326)
--	g29316 = AND(g28528, g6875, g3288)
--	g19354 = AND(g471, g16235)
--	g33244 = AND(g32190, g23152)
--	g32177 = AND(g30608, g25214)
--	g18406 = AND(g2060, g15373)
--	g13349 = AND(g4933, g11780)
--	I31167 = AND(g32696, g32697, g32698, g32699)
--	I18785 = AND(g13156, g6767, g11498)
--	g26279 = AND(g4249, g25213)
--	g18361 = AND(g1821, g17955)
--	g24758 = AND(g6523, g23733)
--	g23130 = AND(g728, g20248)
--	g34667 = AND(g34471, g33424)
--	g34694 = AND(g34530, g19885)
--	g17405 = AND(g1422, g13137)
--	g11083 = AND(g8836, g802)
--	g34965 = AND(g34949, g23084)
--	g30131 = AND(g28589, g21178)
--	g31069 = AND(g29793, g14150)
--	g19671 = AND(g1454, g16155)
--	g29989 = AND(g29006, g10489)
--	g18500 = AND(g2421, g15426)
--	g22020 = AND(g5863, g19147)
--	g27682 = AND(g25777, g23565)
--	g23165 = AND(g13954, g19964)
--	g28183 = AND(g27024, g19421)
--	g28673 = AND(g1373, g27122)
--	g33810 = AND(g33427, g12768)
--	g27291 = AND(g11969, g26653)
--	g29611 = AND(g28540, g14209)
--	g33657 = AND(g30991, g33443)
--	g26286 = AND(g2126, g25389)
--	g29988 = AND(g29187, g12235)
--	g29924 = AND(g13031, g29190)
--	g34487 = AND(g34416, g18983)
--	g13566 = AND(g7092, g12358)
--	g22046 = AND(g6073, g21611)
--	g26306 = AND(g13087, g25286)
--	g24849 = AND(g4165, g22227)
--	g33879 = AND(g33289, g20566)
--	g24940 = AND(g5011, g23971)
--	g24399 = AND(g3133, g23067)
--	g34502 = AND(g26363, g34343)
--	g30210 = AND(g28684, g23877)
--	g34557 = AND(g34352, g20555)
--	g23006 = AND(g19575, g19776)
--	g23475 = AND(g19070, g8971)
--	g33878 = AND(g33288, g20565)
--	I31022 = AND(g32487, g32488, g32489, g32490)
--	g18221 = AND(g1018, g16100)
--	g22113 = AND(g6561, g19277)
--	g21863 = AND(g3957, g21070)
--	g26815 = AND(g4108, g24528)
--	g24141 = AND(g17657, g21656)
--	g34279 = AND(g34231, g19208)
--	g11139 = AND(g5990, g7051, g5976, g9935)
--	g33886 = AND(g33297, g20614)
--	g27134 = AND(g25997, g16602)
--	g30278 = AND(g28818, g23988)
--	g27029 = AND(g26327, g11031)
--	g18613 = AND(g3338, g17200)
--	g31792 = AND(g30214, g24017)
--	g32166 = AND(g31007, g23029)
--	g32009 = AND(g31782, g22224)
--	g25993 = AND(g2610, g25025)
--	g31967 = AND(g31755, g22167)
--	g31994 = AND(g31775, g22215)
--	g22105 = AND(g6494, g18833)
--	I31276 = AND(g31376, g31844, g32854, g32855)
--	g27028 = AND(g26342, g1157)
--	g29199 = AND(g27187, g12687)
--	g32008 = AND(g31781, g22223)
--	g25965 = AND(g2208, g24980)
--	g29650 = AND(g28949, g22472)
--	g29736 = AND(g28522, g10233)
--	g16160 = AND(g5499, g14262)
--	g29887 = AND(g28417, g23351)
--	g21703 = AND(g146, g20283)
--	g18273 = AND(g1287, g16031)
--	g24332 = AND(g4459, g22228)
--	g18106 = AND(g411, g17015)
--	g20135 = AND(g16258, g16695)
--	g18605 = AND(g3129, g16987)
--	g13415 = AND(g837, g11048)
--	g21347 = AND(g1339, g15750)
--	g13333 = AND(g4743, g11755)
--	g33425 = AND(g32380, g21466)
--	g28213 = AND(g27720, g23380)
--	g15679 = AND(g3470, g13555)
--	g18812 = AND(g6509, g15483)
--	g10948 = AND(g7880, g1478)
--	g18463 = AND(g2375, g15224)
--	g33919 = AND(g33438, g10795)
--	g24406 = AND(g13623, g22860)
--	g29528 = AND(g2429, g28874)
--	I31036 = AND(g30673, g31802, g32506, g32507)
--	g24962 = AND(g23194, g20210)
--	g29843 = AND(g28373, g23289)
--	g21781 = AND(g3408, g20391)
--	g29330 = AND(g29114, g18894)
--	g16617 = AND(g6287, g14940)
--	g25502 = AND(g6946, g22527)
--	g15678 = AND(g1094, g13846)
--	I31101 = AND(g30735, g31813, g32601, g32602)
--	I31177 = AND(g32710, g32711, g32712, g32713)
--	g18951 = AND(g3484, g16124)
--	g30187 = AND(g28643, g23840)
--	g18371 = AND(g1870, g15171)
--	g8721 = AND(g385, g376, g365)
--	g28205 = AND(g27516, g16746)
--	g18234 = AND(g1129, g16326)
--	g34187 = AND(g33708, g24397)
--	g17769 = AND(g1146, g13188)
--	g21952 = AND(g5366, g21514)
--	g28311 = AND(g9792, g27679)
--	g23372 = AND(g16448, g20194)
--	g29869 = AND(g2331, g29129)
--	g21821 = AND(g3723, g20453)
--	g17768 = AND(g13325, g10741)
--	I26530 = AND(g26365, g24096, g24097, g24098)
--	g18795 = AND(g6163, g15348)
--	g30937 = AND(g22626, g29814)
--	g29868 = AND(g2227, g29128)
--	g27649 = AND(g10820, g25820)
--	g34143 = AND(g33934, g23828)
--	g16595 = AND(g5921, g14697)
--	g21790 = AND(g3454, g20391)
--	g24004 = AND(g37, g21225)
--	g33086 = AND(g32390, g18887)
--	g27648 = AND(g25882, g8974)
--	g24221 = AND(g232, g22594)
--	g27491 = AND(g26576, g17652)
--	g26486 = AND(g4423, g24358)
--	g18514 = AND(g2629, g15509)
--	g29709 = AND(g2116, g29121)
--	g34169 = AND(g33804, g31227)
--	g21873 = AND(g6946, g19801)
--	g18507 = AND(g2595, g15509)
--	g22027 = AND(g5889, g19147)
--	g23873 = AND(g21222, g10815)
--	g15875 = AND(g3961, g13963)
--	g30168 = AND(g28623, g23794)
--	g29708 = AND(g1955, g29082)
--	g33817 = AND(g33235, g20102)
--	g11115 = AND(g6133, g9954)
--	g33322 = AND(g32202, g20450)
--	g34410 = AND(g34204, g21427)
--	g27981 = AND(g26751, g23924)
--	g25815 = AND(g8155, g24603)
--	g31125 = AND(g29502, g22973)
--	g32176 = AND(g2779, g31623)
--	I31166 = AND(g30673, g31825, g32694, g32695)
--	g26223 = AND(g24688, g10678, g10658, g8757)
--	g31977 = AND(g31764, g22179)
--	g33532 = AND(g32974, I31356, I31357)
--	g33901 = AND(g33317, g20920)
--	g34479 = AND(g34403, g18905)
--	g34666 = AND(g34587, g19144)
--	g25187 = AND(g12296, g23629)
--	g18163 = AND(g79, g17433)
--	g15837 = AND(g3255, g14127)
--	g32154 = AND(g31277, g14184)
--	g34363 = AND(g34148, g20389)
--	g25975 = AND(g9434, g24999)
--	g34217 = AND(g33736, g22876)
--	g22710 = AND(g19358, g19600)
--	g30015 = AND(g29040, g10519)
--	g21834 = AND(g3752, g20453)
--	g22003 = AND(g5736, g21562)
--	g34478 = AND(g34402, g18904)
--	g28152 = AND(g26297, g27279)
--	g26084 = AND(g24926, g9602)
--	g28846 = AND(g21434, g26424, g25399, g27474)
--	g24812 = AND(g19662, g22192)
--	g19855 = AND(g2787, g15962)
--	g33353 = AND(g32240, g20732)
--	g25143 = AND(g4922, g22908)
--	g34486 = AND(g34412, g18953)
--	g18541 = AND(g2767, g15277)
--	g27395 = AND(g8046, g26314, g9187, g9077)
--	g33680 = AND(g33128, g4688)
--	g18473 = AND(g2342, g15224)
--	g27262 = AND(g25997, g17092)
--	g26179 = AND(g2504, g25155)
--	g12794 = AND(g1008, g7567)
--	I17529 = AND(g13156, g11450, g6756)
--	g34556 = AND(g34350, g20537)
--	g18789 = AND(g6035, g15634)
--	g21453 = AND(g16713, g13625)
--	g22081 = AND(g6279, g19210)
--	g29602 = AND(g2020, g28962)
--	g29810 = AND(g28259, g11317)
--	g29774 = AND(g28287, g10233)
--	g34580 = AND(g29539, g34311)
--	g26178 = AND(g2389, g25473)
--	g16194 = AND(g11547, g6782, g11640, I17529)
--	g27633 = AND(g13076, g25766)
--	g21913 = AND(g5069, g21468)
--	g29375 = AND(g13946, g28370)
--	g30223 = AND(g28702, g23895)
--	g13805 = AND(g11489, g11394, g11356, I16129)
--	g18788 = AND(g6031, g15634)
--	g18724 = AND(g4907, g16077)
--	g25884 = AND(g11153, g24711)
--	g18359 = AND(g1825, g17955)
--	g34223 = AND(g33744, g22876)
--	g18325 = AND(g1624, g17873)
--	g26186 = AND(g24580, g23031)
--	g23436 = AND(g676, g20375)
--	g18535 = AND(g2741, g15277)
--	g18434 = AND(g2217, g18008)
--	g18358 = AND(g1811, g17955)
--	g31966 = AND(g31754, g22166)
--	g30084 = AND(g28534, g20700)
--	g27521 = AND(g26519, g14700)
--	g29337 = AND(g29166, g22180)
--	g17786 = AND(g1489, g13216)
--	g30110 = AND(g28564, g20916)
--	g25479 = AND(g22646, g9917)
--	g34084 = AND(g9214, g33851)
--	g15075 = AND(g12850, g12955)
--	g31017 = AND(g29479, g22841)
--	g34110 = AND(g33732, g22935)
--	g25217 = AND(g12418, g23698)
--	g33364 = AND(g32264, g20921)
--	g18121 = AND(g424, g17015)
--	g22090 = AND(g6404, g18833)
--	g30179 = AND(g28634, g23819)
--	g24507 = AND(g22304, g19429)
--	g18344 = AND(g1740, g17955)
--	g19581 = AND(g15843, g1500, g10918)
--	g34179 = AND(g33686, g24372)
--	g27440 = AND(g8046, g26314, g518, g504)
--	g21464 = AND(g16181, g10872)
--	g28020 = AND(g23032, g26241, g26424, g25542)
--	g28583 = AND(g12009, g27112)
--	g30178 = AND(g28632, g23815)
--	g9479 = AND(g305, g324)
--	g24421 = AND(g3835, g23139)
--	g34178 = AND(g33712, g24361)
--	g34740 = AND(g34664, g19414)
--	g16616 = AND(g6267, g14741)
--	g10756 = AND(g3990, g6928, g3976, g8595)
--	g18682 = AND(g4646, g15885)
--	I31176 = AND(g31579, g31827, g32708, g32709)
--	g30186 = AND(g28641, g23839)
--	g27247 = AND(g2759, g26745)
--	I31092 = AND(g32589, g32590, g32591, g32592)
--	g18291 = AND(g1437, g16449)
--	g24012 = AND(g14496, g21561)
--	g17182 = AND(g8579, g13016)
--	g21797 = AND(g3518, g20924)
--	g34186 = AND(g33705, g24396)
--	g34685 = AND(g14164, g34550)
--	g25580 = AND(g19268, g24149)
--	g18173 = AND(g736, g17328)
--	g27389 = AND(g26519, g17503)
--	g34953 = AND(g34935, g19957)
--	g27045 = AND(g10295, g3171, g3179, g26244)
--	g31309 = AND(g30132, g27837)
--	I24699 = AND(g21127, g24054, g24055, g24056)
--	g32083 = AND(g947, g30735)
--	g32348 = AND(g2145, g31672)
--	g23292 = AND(g19879, g16726)
--	g25223 = AND(g22523, g10652)
--	g16704 = AND(g5957, g15018)
--	g27612 = AND(g25887, g8844)
--	g31224 = AND(g30280, g23932)
--	g32284 = AND(g31260, g20507)
--	g28113 = AND(g8016, g27242)
--	g26423 = AND(g19488, g24356)
--	g27099 = AND(g14094, g26352)
--	g15822 = AND(g3925, g13960)
--	g27388 = AND(g26519, g17502)
--	g27324 = AND(g10150, g26720)
--	g24541 = AND(g22626, g10851)
--	g32304 = AND(g31284, g20564)
--	g30936 = AND(g8830, g29916)
--	g28282 = AND(g23762, g27727)
--	g12099 = AND(g9619, g9888)
--	g27534 = AND(g26488, g17735)
--	g27098 = AND(g25868, g22528)
--	g28302 = AND(g23809, g27817)
--	g25084 = AND(g4737, g22885)
--	g27251 = AND(g26721, g26694)
--	g27272 = AND(g26055, g17144)
--	g25110 = AND(g10427, g23509)
--	g16808 = AND(g6653, g14825)
--	g19384 = AND(g667, g16310)
--	g18760 = AND(g5462, g17929)
--	g18134 = AND(g534, g17249)
--	g25922 = AND(g24959, g20065)
--	g34334 = AND(g34090, g19865)
--	g24788 = AND(g11384, g23111)
--	g31495 = AND(g1913, g30309)
--	g24724 = AND(g17624, g22432)
--	g29599 = AND(g1710, g29018)
--	g33495 = AND(g32707, I31171, I31172)
--	g22717 = AND(g9291, g20212)
--	g16177 = AND(g5128, g14238)
--	g24325 = AND(g4543, g22228)
--	g25179 = AND(g16928, g23611)
--	g26543 = AND(g12910, g24377)
--	I27503 = AND(g19890, g24075, g24076, g28032)
--	g18506 = AND(g2571, g15509)
--	g22026 = AND(g5913, g19147)
--	g27462 = AND(g26576, g17612)
--	g33816 = AND(g33234, g20096)
--	g29598 = AND(g28823, g22342)
--	g16642 = AND(g6633, g14981)
--	g25178 = AND(g20241, g23608)
--	g15589 = AND(g411, g13334)
--	g32139 = AND(g31601, g29960)
--	g27032 = AND(g7704, g5180, g5188, g26200)
--	g34964 = AND(g34947, g23060)
--	g33687 = AND(g33132, g4878)
--	g31976 = AND(g31762, g22178)
--	g31985 = AND(g4722, g30614)
--	g19735 = AND(g9740, g17135)
--	g27140 = AND(g25885, g22593)
--	g30216 = AND(g28691, g23882)
--	g27997 = AND(g26813, g23995)
--	g28768 = AND(g21434, g26424, g25308, g27421)
--	g15836 = AND(g3187, g14104)
--	g31752 = AND(g30104, g23928)
--	g34216 = AND(g33778, g22689)
--	g31374 = AND(g29748, g23390)
--	g29322 = AND(g29192, g7074, g6336)
--	g33374 = AND(g32289, g21221)
--	g16733 = AND(g5893, g14889)
--	I18671 = AND(g13156, g11450, g6756)
--	g29532 = AND(g1878, g28861)
--	g29901 = AND(g28429, g23376)
--	g32333 = AND(g31326, g23559)
--	g15119 = AND(g4249, g14454)
--	g20682 = AND(g16238, g4646)
--	g13771 = AND(g11441, g11355, g11302, I16111)
--	g25417 = AND(g5712, g23816, I24552)
--	g23474 = AND(g13830, g20533)
--	g24682 = AND(g22662, g19754)
--	g22149 = AND(g14581, g18880)
--	g29783 = AND(g28329, g23246)
--	g21711 = AND(g291, g20283)
--	g26123 = AND(g1696, g25382)
--	g15118 = AND(g4253, g14454)
--	g34909 = AND(g34856, g20130)
--	g24291 = AND(g18660, g22550)
--	g30000 = AND(g23685, g29029)
--	g29656 = AND(g28515, g11666)
--	g34117 = AND(g33742, g19755)
--	g15749 = AND(g1454, g13273)
--	g18649 = AND(g4049, g17271)
--	g22097 = AND(g6451, g18833)
--	g27360 = AND(g26488, g17417)
--	g33842 = AND(g33255, g20322)
--	g18240 = AND(g15066, g16431)
--	g22104 = AND(g6444, g18833)
--	g17149 = AND(g232, g13255)
--	g33392 = AND(g32344, g21362)
--	g18648 = AND(g4045, g17271)
--	g18491 = AND(g2518, g15426)
--	g31489 = AND(g2204, g30305)
--	g26230 = AND(g1768, g25385)
--	g25964 = AND(g1783, g24979)
--	g33489 = AND(g32665, I31141, I31142)
--	g21606 = AND(g15959, g13763)
--	g27162 = AND(g26171, g8259, g2208)
--	g34568 = AND(g34379, g17512)
--	g34747 = AND(g34671, g19527)
--	g23606 = AND(g16927, g20679)
--	g29336 = AND(g4704, g28363)
--	g15704 = AND(g3440, g13504)
--	g30242 = AND(g28730, g23927)
--	g18604 = AND(g3125, g16987)
--	g21303 = AND(g10120, g17625)
--	g16485 = AND(g5563, g14924)
--	g18755 = AND(g5343, g15595)
--	g31525 = AND(g29892, g23526)
--	g31488 = AND(g1779, g30302)
--	g31016 = AND(g29478, g22840)
--	g33525 = AND(g32925, I31321, I31322)
--	g33488 = AND(g32658, I31136, I31137)
--	g28249 = AND(g27152, g19677)
--	g15809 = AND(g3917, g14154)
--	g18770 = AND(g15153, g15615)
--	g22369 = AND(g9354, g7717, g20783)
--	g18563 = AND(g2890, g16349)
--	g18981 = AND(g11206, g16158)
--	g21750 = AND(g3161, g20785)
--	g28248 = AND(g27150, g19676)
--	g29966 = AND(g23617, g28970)
--	g28710 = AND(g27589, g20703)
--	g15808 = AND(g3590, g14048)
--	g21982 = AND(g5547, g19074)
--	g27451 = AND(g26400, g17599)
--	g26391 = AND(g19593, g25555)
--	I26948 = AND(g24981, g26424, g22698)
--	g23381 = AND(g7239, g21413)
--	g27220 = AND(g26026, g16743)
--	g33830 = AND(g33382, g20166)
--	g29631 = AND(g1682, g28656)
--	g32312 = AND(g31302, g20591)
--	g32200 = AND(g27468, g31376)
--	g33893 = AND(g33313, g20706)
--	g28204 = AND(g26098, g27654)
--	g27628 = AND(g26400, g18061)
--	g34751 = AND(g34674, g19543)
--	g29364 = AND(g27400, g28321)
--	g10827 = AND(g8914, g4258)
--	g25909 = AND(g8745, g24875)
--	g32115 = AND(g31631, g29928)
--	g25543 = AND(g23795, g21461)
--	g12220 = AND(g1521, g7535)
--	g27246 = AND(g26690, g26673)
--	g33865 = AND(g33275, g20526)
--	g21796 = AND(g3512, g20924)
--	g30230 = AND(g28717, g23906)
--	g25908 = AND(g24782, g22520)
--	g18767 = AND(g15150, g17929)
--	g18794 = AND(g6154, g15348)
--	g34230 = AND(g33761, g22942)
--	g18395 = AND(g12849, g15373)
--	g32052 = AND(g31507, g13885)
--	g18262 = AND(g1259, g16000)
--	g22133 = AND(g6649, g19277)
--	g25569 = AND(I24684, I24685)
--	g21840 = AND(g15099, g21070)
--	g25568 = AND(I24679, I24680)
--	g18633 = AND(g6905, g17226)
--	g17133 = AND(g10683, g13222)
--	g34841 = AND(g34761, g20080)
--	g18191 = AND(g827, g17821)
--	g18719 = AND(g4894, g16795)
--	g22011 = AND(g15154, g21562)
--	g15874 = AND(g3893, g14079)
--	g24649 = AND(g6527, g23733)
--	g29571 = AND(g28452, g11762)
--	g11114 = AND(g5689, g10160)
--	g31270 = AND(g29692, g23282)
--	g16519 = AND(g5591, g14804)
--	g16176 = AND(g14596, g11779)
--	g16185 = AND(g3263, g14011)
--	g25123 = AND(g4732, g22885)
--	g18718 = AND(g4854, g15915)
--	g15693 = AND(g269, g13474)
--	g18521 = AND(g2667, g15509)
--	g31188 = AND(g20028, g29653)
--	g25814 = AND(g24760, g13323)
--	g27370 = AND(g26400, g17472)
--	g31124 = AND(g2259, g29997)
--	g32184 = AND(g30611, g25249)
--	g28998 = AND(g17424, g25212, g26424, g27474)
--	g33124 = AND(g8945, g32296)
--	g33678 = AND(g33149, g10710, g22319)
--	g24491 = AND(g10727, g22332)
--	g24903 = AND(g128, g23889)
--	g28233 = AND(g27827, g23411)
--	g16518 = AND(g5571, g14956)
--	g28182 = AND(g8770, g27349)
--	g25772 = AND(g24944, g24934)
--	g28672 = AND(g7577, g27017)
--	g24755 = AND(g16022, g23030)
--	g27151 = AND(g26026, g16626)
--	g34578 = AND(g24578, g34308)
--	g16637 = AND(g5949, g14968)
--	g22310 = AND(g19662, g20235)
--	g18440 = AND(g2255, g18008)
--	g13345 = AND(g4754, g11773)
--	g26275 = AND(g2417, g25349)
--	g30007 = AND(g29141, g12929)
--	I24546 = AND(g5046, g5052, g9716)
--	g34586 = AND(g11025, g34317)
--	g18573 = AND(g2898, g16349)
--	g29687 = AND(g2407, g29097)
--	g22112 = AND(g6555, g19277)
--	g18247 = AND(g1178, g16431)
--	g29985 = AND(g28127, g20532)
--	g10890 = AND(g7858, g1105)
--	g21862 = AND(g3953, g21070)
--	g22050 = AND(g6088, g21611)
--	g23553 = AND(g19413, g11875)
--	g18389 = AND(g1974, g15171)
--	g29752 = AND(g28516, g10233)
--	I31312 = AND(g32905, g32906, g32907, g32908)
--	g29954 = AND(g2299, g28796)
--	g21949 = AND(g5264, g18997)
--	g15712 = AND(g3791, g13521)
--	g18612 = AND(g3329, g17200)
--	g15914 = AND(g3905, g14024)
--	g25992 = AND(g2485, g25024)
--	g18388 = AND(g1968, g15171)
--	g19660 = AND(g12001, g16968)
--	g18324 = AND(g1644, g17873)
--	g24794 = AND(g11414, g23138)
--	g31219 = AND(g30265, g20875)
--	g34116 = AND(g33933, g25140)
--	g24395 = AND(g4704, g22845)
--	g25510 = AND(g6444, g22300, I24619)
--	g18701 = AND(g4771, g16856)
--	g26684 = AND(g25407, g20673)
--	g21948 = AND(g5260, g18997)
--	g22096 = AND(g6434, g18833)
--	g32400 = AND(g4743, g30989)
--	g18777 = AND(g5808, g18065)
--	g18534 = AND(g2735, g15277)
--	I14198 = AND(g225, g8237, g232, g8180)
--	g32013 = AND(g8673, g30614)
--	g30041 = AND(g28511, g23518)
--	I31052 = AND(g32531, g32532, g32533, g32534)
--	g18251 = AND(g996, g16897)
--	g21702 = AND(g157, g20283)
--	g31218 = AND(g30271, g23909)
--	g16729 = AND(g5240, g14720)
--	g18272 = AND(g1283, g16031)
--	g21757 = AND(g3187, g20785)
--	g25579 = AND(g19422, g24147)
--	g30275 = AND(g28816, g23984)
--	I24700 = AND(g24057, g24058, g24059, g24060)
--	g27227 = AND(g26026, g16771)
--	g33837 = AND(g33251, g20233)
--	I24625 = AND(g6428, g6434, g10014)
--	g32207 = AND(g31221, g23323)
--	g26517 = AND(g15708, g24367)
--	g34746 = AND(g34670, g19526)
--	g34493 = AND(g34273, g19360)
--	g25578 = AND(g19402, g24146)
--	g15567 = AND(g392, g13312)
--	g27025 = AND(g26334, g7917)
--	g24191 = AND(g319, g22722)
--	g24719 = AND(g681, g23530)
--	g18462 = AND(g2361, g15224)
--	g25014 = AND(g17474, g23420)
--	g32328 = AND(g5853, g31554)
--	g29668 = AND(g28527, g14255)
--	g29842 = AND(g28372, g23284)
--	g27540 = AND(g26576, g17746)
--	g23564 = AND(g16882, g20648)
--	g27058 = AND(g10323, g3522, g3530, g26264)
--	g30035 = AND(g22539, g28120)
--	g18140 = AND(g559, g17533)
--	g34340 = AND(g34100, g19950)
--	g27203 = AND(g26026, g16688)
--	g19596 = AND(g1094, g16681)
--	g26130 = AND(g24890, g19772)
--	g29525 = AND(g2169, g28837)
--	g21847 = AND(g3905, g21070)
--	g34684 = AND(g14178, g34545)
--	g10999 = AND(g7880, g1472)
--	g13833 = AND(g4546, g10613)
--	I18819 = AND(g13156, g11450, g11498)
--	g26362 = AND(g19557, g25538)
--	g27044 = AND(g7766, g5873, g5881, g26241)
--	g31470 = AND(g29753, g23398)
--	g23397 = AND(g11154, g20239)
--	g33470 = AND(g32528, I31046, I31047)
--	g33915 = AND(g33140, g7846)
--	g32241 = AND(g31244, g20323)
--	g26165 = AND(g11980, g25153)
--	g17793 = AND(g6772, g11592, g6789, I18803)
--	g10998 = AND(g8567, g8509, g8451, g7650)
--	g18766 = AND(g5495, g17929)
--	g13048 = AND(g8558, g11043)
--	g23062 = AND(g718, g20248)
--	g27281 = AND(g9830, g26615)
--	g24861 = AND(g3712, g23582, I24033)
--	g24573 = AND(g17198, g23716)
--	g34517 = AND(g34290, g19493)
--	g28148 = AND(g27355, g26093)
--	g14233 = AND(g8639, g11855)
--	g21933 = AND(g5212, g18997)
--	g27301 = AND(g11992, g26679)
--	I14225 = AND(g8457, g255, g8406, g262)
--	g27957 = AND(g25947, g15995)
--	g7804 = AND(g2975, g2970)
--	g25041 = AND(g23261, g20494)
--	g13221 = AND(g6946, g11425)
--	g27120 = AND(g25878, g22543)
--	g17690 = AND(g11547, g11592, g11640, I18671)
--	g29865 = AND(g1802, g29115)
--	g21851 = AND(g3901, g21070)
--	g21872 = AND(g4098, g19801)
--	g23872 = AND(g19389, g4157)
--	g15883 = AND(g9180, g14258)
--	g18360 = AND(g1830, g17955)
--	g31467 = AND(g30162, g27937)
--	g31494 = AND(g29792, g23435)
--	g28343 = AND(g27380, g19799)
--	I24527 = AND(g9672, g9264, g5401)
--	g19655 = AND(g2729, g16966)
--	g33467 = AND(g32505, I31031, I31032)
--	g33494 = AND(g32700, I31166, I31167)
--	g24324 = AND(g4540, g22228)
--	g27146 = AND(g26148, g8187, g1648)
--	g27645 = AND(g26488, g15344)
--	g26863 = AND(g24974, g24957)
--	g18447 = AND(g2208, g18008)
--	g30193 = AND(g28650, g23848)
--	g24777 = AND(g11345, g23066)
--	g27699 = AND(g26396, g20766)
--	g16653 = AND(g8343, g13850)
--	g18162 = AND(g686, g17433)
--	g25983 = AND(g2476, g25009)
--	g29610 = AND(g28483, g8026)
--	g30165 = AND(g28619, g23788)
--	g22129 = AND(g6633, g19277)
--	g34523 = AND(g9162, g34351)
--	g22002 = AND(g5706, g21562)
--	g22057 = AND(g15159, g21611)
--	g17317 = AND(g1079, g13124)
--	g22128 = AND(g6629, g19277)
--	g33352 = AND(g32237, g20712)
--	I31207 = AND(g32754, g32755, g32756, g32757)
--	g16636 = AND(g5929, g14768)
--	g18629 = AND(g3680, g17226)
--	g25142 = AND(g4717, g22885)
--	g18451 = AND(g2295, g15224)
--	g26347 = AND(g262, g24850)
--	g18472 = AND(g2413, g15224)
--	g32414 = AND(g4944, g30999)
--	g29188 = AND(g27163, g12762)
--	g33418 = AND(g32372, g21425)
--	g33822 = AND(g33385, g20157)
--	g18220 = AND(g1002, g16100)
--	g26253 = AND(g2327, g25435)
--	g30006 = AND(g29032, g9259)
--	g31266 = AND(g30129, g27742)
--	g31170 = AND(g19128, g29814)
--	g21452 = AND(g16119, g13624)
--	g18628 = AND(g15095, g17226)
--	g27427 = AND(g26400, g17575)
--	g34475 = AND(g27450, g34327)
--	g17057 = AND(g446, g13173)
--	g24140 = AND(g17663, g21654)
--	g22299 = AND(g19999, g21024)
--	g29686 = AND(g2246, g29057)
--	g24997 = AND(g22929, g10419)
--	g18246 = AND(g1199, g16431)
--	g21912 = AND(g5052, g21468)
--	g29383 = AND(g28138, g19412)
--	g30222 = AND(g28701, g23894)
--	g34863 = AND(g16540, g34833)
--	g28133 = AND(g27367, g23108)
--	g22298 = AND(g19997, g21012)
--	g26236 = AND(g25357, g6856, g7586, g7558)
--	g28229 = AND(g27345, g17213)
--	g19487 = AND(g499, g16680)
--	g29938 = AND(g23552, g28889)
--	g26351 = AND(g239, g24869)
--	g28228 = AND(g27126, g19636)
--	g25130 = AND(g23358, g20600)
--	g26821 = AND(g24821, g13103)
--	g27661 = AND(g26576, g15568)
--	I31241 = AND(g30825, g31838, g32803, g32804)
--	g27547 = AND(g26549, g17759)
--	g18591 = AND(g2965, g16349)
--	g31194 = AND(g19128, g29814)
--	g31167 = AND(g10080, g30076)
--	g18776 = AND(g5813, g18065)
--	g18785 = AND(g5849, g18065)
--	g15083 = AND(g10362, g12983)
--	g21756 = AND(g3211, g20785)
--	g18147 = AND(g599, g17533)
--	g25165 = AND(g14062, g23570)
--	g30253 = AND(g28746, g23943)
--	g16484 = AND(g5244, g14755)
--	g18754 = AND(g5339, g15595)
--	g31524 = AND(g29897, g20593)
--	g33524 = AND(g32918, I31316, I31317)
--	g18355 = AND(g1748, g17955)
--	g26264 = AND(g24688, g8812, g8778, g10627)
--	g33836 = AND(g33096, g27020)
--	g21780 = AND(g3391, g20391)
--	g29875 = AND(g28403, g23337)
--	g32206 = AND(g30609, g25524)
--	g26516 = AND(g24968, g8876)
--	g13507 = AND(g7023, g12198)
--	g27481 = AND(g26400, g14630)
--	g30600 = AND(g30287, g18975)
--	g18825 = AND(g6736, g15680)
--	g18950 = AND(g11193, g16123)
--	g18370 = AND(g1874, g15171)
--	g31477 = AND(g29763, g23409)
--	g33401 = AND(g32349, g21381)
--	g33477 = AND(g32577, I31081, I31082)
--	g20162 = AND(g8737, g16750)
--	g30236 = AND(g28724, g23916)
--	g14148 = AND(g884, g10632)
--	g29837 = AND(g28369, g20144)
--	g14097 = AND(g878, g10632)
--	g21820 = AND(g3712, g20453)
--	g11163 = AND(g6727, g10224)
--	I24067 = AND(g3731, g3736, g8553)
--	g9906 = AND(g996, g1157)
--	g18151 = AND(g617, g17533)
--	g31118 = AND(g29490, g22906)
--	g18172 = AND(g15058, g17328)
--	g28627 = AND(g27543, g20574)
--	g32114 = AND(g31624, g29927)
--	g28959 = AND(g17401, g25194, g26424, g27440)
--	g30175 = AND(g28629, g23813)
--	g32082 = AND(g4917, g30673)
--	g33864 = AND(g33274, g20524)
--	g27127 = AND(g25997, g16582)
--	g21846 = AND(g3897, g21070)
--	g28112 = AND(g27352, g26162)
--	g32107 = AND(g31624, g29912)
--	g15653 = AND(g3119, g13530)
--	g24629 = AND(g6163, g23699)
--	g23396 = AND(g20051, g20229)
--	g18367 = AND(g1783, g17955)
--	g18394 = AND(g1862, g15171)
--	g31313 = AND(g30160, g27907)
--	g24451 = AND(g3476, g23112)
--	g21731 = AND(g3029, g20330)
--	g24220 = AND(g255, g22594)
--	g20628 = AND(g1046, g15789)
--	g27490 = AND(g26576, g17651)
--	g13541 = AND(g7069, g12308)
--	g30264 = AND(g28774, g23963)
--	g34063 = AND(g33806, g23121)
--	g13473 = AND(g9797, g11841)
--	g30137 = AND(g28594, g21181)
--	g19601 = AND(g16198, g11149)
--	g24628 = AND(g5835, g23666)
--	g32345 = AND(g2138, g31672)
--	g34137 = AND(g33928, g23802)
--	g31285 = AND(g30134, g27800)
--	g34516 = AND(g34289, g19492)
--	g27376 = AND(g26549, g17481)
--	g27385 = AND(g26400, g17497)
--	g33704 = AND(g33176, g10710, g22319)
--	g29617 = AND(g2024, g28987)
--	g31305 = AND(g29741, g23354)
--	I24695 = AND(g24050, g24051, g24052, g24053)
--	I24018 = AND(g8155, g8390, g3396)
--	g27103 = AND(g25997, g16509)
--	g33305 = AND(g31935, g17811)
--	g22831 = AND(g19441, g19629)
--	g23691 = AND(g14731, g20993)
--	g26542 = AND(g13102, g24376)
--	g34873 = AND(g34830, g20046)
--	g26021 = AND(g9568, g25035)
--	g18420 = AND(g1996, g15373)
--	g15852 = AND(g13820, g13223)
--	g27095 = AND(g25997, g16473)
--	g18319 = AND(g1600, g17873)
--	g33809 = AND(g33432, g30184)
--	g33900 = AND(g33316, g20913)
--	g33466 = AND(g32498, I31026, I31027)
--	g16184 = AND(g9285, g14183)
--	g16805 = AND(g7187, g12972)
--	g21405 = AND(g13377, g15811)
--	g16674 = AND(g6637, g15014)
--	g29201 = AND(g24081, I27503, I27504)
--	g32141 = AND(g31639, g29963)
--	g22316 = AND(g2837, g20270)
--	g18318 = AND(g1604, g17873)
--	g18446 = AND(g2279, g18008)
--	g33808 = AND(g33109, g22161)
--	g24785 = AND(g7051, g23645)
--	g18227 = AND(g1052, g16129)
--	g7777 = AND(g723, g822, g817)
--	g27181 = AND(g26026, g16655)
--	g30209 = AND(g28682, g23876)
--	g22498 = AND(g7753, g7717, g21334)
--	g33101 = AND(g32398, g18976)
--	g19791 = AND(g14253, g17189)
--	g24754 = AND(g19604, g23027)
--	g29595 = AND(g28475, g11833)
--	g29494 = AND(g9073, g28479)
--	g30208 = AND(g28681, g23875)
--	g16732 = AND(g5555, g14882)
--	g21929 = AND(g5176, g18997)
--	g32263 = AND(g31631, g30306)
--	g18540 = AND(g2775, g15277)
--	g10896 = AND(g1205, g8654)
--	g22056 = AND(g6133, g21611)
--	g26274 = AND(g2130, g25210)
--	g29623 = AND(g28496, g11563)
--	g32332 = AND(g31325, g23558)
--	I31206 = AND(g31710, g31832, g32752, g32753)
--	g21928 = AND(g5170, g18997)
--	g22080 = AND(g6275, g19210)
--	g25063 = AND(g13078, g22325)
--	g24858 = AND(g3361, g23223, I24030)
--	g29782 = AND(g28328, g23245)
--	g18203 = AND(g911, g15938)
--	g26122 = AND(g24557, g19762)
--	g16761 = AND(g7170, g12947)
--	g29984 = AND(g2567, g28877)
--	g34542 = AND(g34332, g20089)
--	g22432 = AND(g9354, g7717, g21187)
--	g12931 = AND(g392, g11048)
--	g29352 = AND(g4950, g28410)
--	g25873 = AND(g24854, g16197)
--	g30614 = AND(g20154, g29814)
--	I24597 = AND(g5736, g5742, g9875)
--	I31082 = AND(g32573, g32574, g32575, g32576)
--	g18281 = AND(g1373, g16136)
--	g27520 = AND(g26519, g17714)
--	g21787 = AND(g15091, g20391)
--	g15115 = AND(g2946, g14454)
--	I31107 = AND(g32610, g32611, g32612, g32613)
--	g22342 = AND(g9354, g9285, g21287)
--	g18301 = AND(g1532, g16489)
--	g30607 = AND(g30291, g18989)
--	g32049 = AND(g10902, g30735)
--	I24689 = AND(g20841, g24040, g24041, g24042)
--	g26292 = AND(g2689, g25228)
--	g33693 = AND(g33145, g13594)
--	g18377 = AND(g1894, g15171)
--	g19556 = AND(g11932, g16809)
--	g30073 = AND(g1379, g28194)
--	g22145 = AND(g14555, g18832)
--	g18120 = AND(g457, g17015)
--	g26153 = AND(g24565, g19780)
--	g18739 = AND(g5008, g16826)
--	g21302 = AND(g956, g15731)
--	g22031 = AND(g5917, g19147)
--	g27546 = AND(g26549, g17758)
--	g30274 = AND(g28815, g23983)
--	g31166 = AND(g1816, g30074)
--	g34073 = AND(g8948, g33823)
--	g10925 = AND(g7858, g956)
--	g16207 = AND(g9839, g14204)
--	g27211 = AND(g25997, g16716)
--	g32048 = AND(g31498, g13869)
--	g16539 = AND(g11547, g6782, g6789, I17741)
--	g21743 = AND(g3100, g20330)
--	g21827 = AND(g3759, g20453)
--	g11029 = AND(g5782, g9103)
--	g17753 = AND(g13281, g13175)
--	g18146 = AND(g595, g17533)
--	g18738 = AND(g15142, g16826)
--	g13029 = AND(g8359, g11030)
--	g15745 = AND(g686, g13223)
--	g18645 = AND(g15100, g17271)
--	g30122 = AND(g28578, g21054)
--	g24420 = AND(g23997, g18980)
--	g24319 = AND(g4561, g22228)
--	g29853 = AND(g1862, g29081)
--	g16538 = AND(g6255, g15005)
--	g17145 = AND(g7469, g13249)
--	g26635 = AND(g25321, g20617)
--	g11028 = AND(g9730, g5428)
--	g18699 = AND(g4760, g16816)
--	g34565 = AND(g34374, g17471)
--	g15813 = AND(g3247, g14069)
--	g31485 = AND(g29776, g23421)
--	g29589 = AND(g2575, g28977)
--	g33892 = AND(g33312, g20701)
--	g18290 = AND(g1467, g16449)
--	g17199 = AND(g2236, g13034)
--	g24318 = AND(g4555, g22228)
--	g33476 = AND(g32570, I31076, I31077)
--	g33485 = AND(g32635, I31121, I31122)
--	g21769 = AND(g3247, g20785)
--	g30034 = AND(g29077, g10541)
--	g22843 = AND(g9429, g20272)
--	g24227 = AND(g890, g22594)
--	g18698 = AND(g15131, g16777)
--	I31141 = AND(g31376, g31820, g32659, g32660)
--	g25453 = AND(g5406, g23789, I24576)
--	g29588 = AND(g2311, g28942)
--	g29524 = AND(g2004, g28864)
--	g29836 = AND(g28425, g26841)
--	g21768 = AND(g3243, g20785)
--	g21803 = AND(g3538, g20924)
--	g28245 = AND(g11367, g27975)
--	g15805 = AND(g3243, g14041)
--	g28626 = AND(g27542, g20573)
--	g30153 = AND(g28610, g23768)
--	g28299 = AND(g9716, g27670)
--	g27700 = AND(g22342, g25182, g26424, g26148)
--	g22132 = AND(g6645, g19277)
--	g29477 = AND(g14090, g28441)
--	g32273 = AND(g31255, g20446)
--	g32106 = AND(g31601, g29911)
--	g18427 = AND(g2181, g18008)
--	g14681 = AND(g4392, g10476)
--	g19740 = AND(g2783, g15907)
--	g20203 = AND(g6195, g17789)
--	g33907 = AND(g23088, g33219, g9104)
--	g18366 = AND(g1854, g17955)
--	I31332 = AND(g32935, g32936, g32937, g32938)
--	g21881 = AND(g4064, g19801)
--	g27658 = AND(g22491, g25786)
--	g18632 = AND(g3698, g17226)
--	g25905 = AND(g24879, g16311)
--	g17365 = AND(g7650, g13036)
--	g22161 = AND(g13202, g19071)
--	g33074 = AND(g32387, g18830)
--	g34136 = AND(g33850, g23293)
--	g33239 = AND(g32117, g19902)
--	g25530 = AND(g23750, g21414)
--	g27339 = AND(g26400, g17308)
--	g29749 = AND(g28295, g23214)
--	g29616 = AND(g1974, g29085)
--	g7511 = AND(g2145, g2138, g2130)
--	g26711 = AND(g25446, g20713)
--	g31238 = AND(g29583, g20053)
--	g32234 = AND(g31601, g30292)
--	g25122 = AND(g23374, g20592)
--	g18403 = AND(g2028, g15373)
--	g18547 = AND(g121, g15277)
--	g25565 = AND(g13013, g22660)
--	g24301 = AND(g6961, g22228)
--	g28232 = AND(g27732, g23586)
--	g20739 = AND(g16259, g4674)
--	g13491 = AND(g6999, g12160)
--	g22087 = AND(g6303, g19210)
--	g30164 = AND(g28618, g23787)
--	g31941 = AND(g1283, g30825)
--	g33941 = AND(g33380, g21560)
--	g18226 = AND(g15064, g16129)
--	g21890 = AND(g4125, g19801)
--	g13604 = AND(g4495, g10487)
--	g31519 = AND(g29864, g23490)
--	g18715 = AND(g4871, g15915)
--	g27968 = AND(g25958, g19614)
--	g28697 = AND(g27581, g20669)
--	g31185 = AND(g10114, g30087)
--	g18481 = AND(g2461, g15426)
--	g33519 = AND(g32881, I31291, I31292)
--	g29809 = AND(g28362, g23274)
--	g33675 = AND(g33164, g10727, g22332)
--	g24645 = AND(g22639, g19709)
--	g28261 = AND(g27878, g23695)
--	g26606 = AND(g1018, g24510)
--	g28880 = AND(g21434, g26424, g25438, g27494)
--	g18551 = AND(g2811, g15277)
--	g22043 = AND(g5965, g19147)
--	g26303 = AND(g2685, g25439)
--	g31518 = AND(g20041, g29970)
--	g31154 = AND(g19128, g29814)
--	g18572 = AND(g2864, g16349)
--	g33518 = AND(g32874, I31286, I31287)
--	g29808 = AND(g28361, g23273)
--	g21710 = AND(g287, g20283)
--	I31221 = AND(g31327, g31835, g32773, g32774)
--	g24290 = AND(g4430, g22550)
--	g29036 = AND(g27163, g12762, g20875, I27381)
--	g27411 = AND(g26549, g17528)
--	g34474 = AND(g20083, g34326)
--	g24698 = AND(g22664, g19761)
--	g21779 = AND(g3385, g20391)
--	g26750 = AND(g24514, g24474)
--	g12527 = AND(g8680, g667)
--	g23779 = AND(g1105, g19355)
--	g18127 = AND(g499, g16971)
--	g22069 = AND(g6227, g19210)
--	g25408 = AND(g22682, g9772)
--	g30109 = AND(g28562, g20912)
--	g26381 = AND(g4456, g25548)
--	g34109 = AND(g33918, g23708)
--	g29642 = AND(g27954, g28669)
--	g33883 = AND(g33294, g20589)
--	g21778 = AND(g3355, g20391)
--	g22068 = AND(g6219, g19210)
--	g26091 = AND(g1691, g25082)
--	g18490 = AND(g2504, g15426)
--	g30108 = AND(g28561, g20910)
--	g32163 = AND(g3502, g31170)
--	g32012 = AND(g8297, g31233)
--	g34108 = AND(g22957, g9104, g33766)
--	g24427 = AND(g4961, g22919)
--	g21786 = AND(g3436, g20391)
--	g27503 = AND(g26488, g14668)
--	I24054 = AND(g8443, g8075, g3747)
--	g30283 = AND(g28851, g23993)
--	I31106 = AND(g30825, g31814, g32608, g32609)
--	g18784 = AND(g15155, g18065)
--	g18376 = AND(g1913, g15171)
--	g18385 = AND(g1959, g15171)
--	g29733 = AND(g2675, g29157)
--	g18297 = AND(g1478, g16449)
--	g17810 = AND(g1495, g13246)
--	g18103 = AND(g401, g17015)
--	g10626 = AND(g4057, g7927)
--	g34492 = AND(g34272, g33430)
--	g13633 = AND(g4567, g10509)
--	g25164 = AND(g16883, g23569)
--	g21945 = AND(g5248, g18997)
--	g28499 = AND(g27982, g17762)
--	g18354 = AND(g1792, g17955)
--	g29874 = AND(g28402, g23336)
--	g27714 = AND(g22384, g25195, g26424, g26171)
--	g21826 = AND(g3742, g20453)
--	g21999 = AND(g5723, g21562)
--	g26390 = AND(g4423, g25554)
--	g31501 = AND(g2047, g29310)
--	g18824 = AND(g6732, g15680)
--	g27315 = AND(g12022, g26709)
--	g33501 = AND(g32751, I31201, I31202)
--	g29630 = AND(g28212, g19781)
--	g24403 = AND(g4894, g22858)
--	g29693 = AND(g28207, g10233)
--	g30982 = AND(g8895, g29933)
--	g34750 = AND(g34673, g19542)
--	g16759 = AND(g5587, g14761)
--	g18181 = AND(g772, g17328)
--	g21998 = AND(g5712, g21562)
--	g18671 = AND(g4628, g15758)
--	g34381 = AND(g34166, g20594)
--	g23998 = AND(g19631, g10971)
--	g33728 = AND(g22626, g10851, g33187)
--	g27202 = AND(g25997, g13876)
--	g19568 = AND(g1467, g15959)
--	g30091 = AND(g28127, g20716)
--	g32325 = AND(g31316, g23538)
--	g29665 = AND(g2375, g28696)
--	g16758 = AND(g5220, g14758)
--	g34091 = AND(g22957, g9104, g33761)
--	g24226 = AND(g446, g22594)
--	g13832 = AND(g8880, g10612)
--	g28722 = AND(g27955, g20738)
--	g28924 = AND(g17317, g25183, g26424, g27416)
--	g30174 = AND(g28628, g23812)
--	g29008 = AND(g27163, g12730, g20739, I27364)
--	g12979 = AND(g424, g11048)
--	g24551 = AND(g17148, g23331)
--	g24572 = AND(g5462, g23393)
--	g33349 = AND(g32233, g20699)
--	g25108 = AND(g23345, g20576)
--	g21932 = AND(g5204, g18997)
--	g32121 = AND(g31616, g29942)
--	g18426 = AND(g2177, g18008)
--	g33906 = AND(g33084, g22311)
--	g13247 = AND(g8964, g11316)
--	g29555 = AND(g29004, g22498)
--	g21513 = AND(g16196, g10882)
--	g18190 = AND(g822, g17821)
--	g22010 = AND(g5787, g21562)
--	g23513 = AND(g19430, g13007)
--	g34390 = AND(g34172, g21069)
--	g10856 = AND(g4269, g8967)
--	g11045 = AND(g5787, g9883)
--	g15882 = AND(g3554, g13986)
--	g27384 = AND(g26400, g17496)
--	g29570 = AND(g2763, g28598)
--	g29712 = AND(g2643, g28726)
--	I24694 = AND(g20982, g24047, g24048, g24049)
--	g33304 = AND(g32427, g31971)
--	g14261 = AND(g4507, g10738)
--	g18520 = AND(g2661, g15509)
--	g21961 = AND(g5424, g21514)
--	g22079 = AND(g6271, g19210)
--	g27094 = AND(g25997, g16472)
--	g30192 = AND(g28649, g23847)
--	g31566 = AND(g19050, g29814)
--	g13324 = AND(g854, g11326)
--	g29907 = AND(g2629, g29177)
--	g32291 = AND(g31268, g20527)
--	g16804 = AND(g5905, g14813)
--	g21404 = AND(g16069, g13569)
--	g28199 = AND(g27479, g16684)
--	g22078 = AND(g6267, g19210)
--	g23404 = AND(g20063, g20247)
--	g32173 = AND(g160, g31134)
--	g18546 = AND(g2795, g15277)
--	g25982 = AND(g2351, g25008)
--	I31012 = AND(g32473, g32474, g32475, g32476)
--	g18211 = AND(g15062, g15979)
--	g21717 = AND(g15051, g21037)
--	g28198 = AND(g26649, g27492)
--	g24297 = AND(g4455, g22550)
--	g22086 = AND(g6299, g19210)
--	g25091 = AND(g12830, g23492)
--	g20095 = AND(g8873, g16632)
--	I24619 = AND(g6423, g6428, g10014)
--	g29567 = AND(g2357, g28593)
--	g29594 = AND(g28529, g14192)
--	g12735 = AND(g7121, g3873, g3881)
--	g31139 = AND(g12221, g30036)
--	g28528 = AND(g27187, g12730)
--	g28330 = AND(g27238, g19786)
--	g26252 = AND(g2283, g25309)
--	g11032 = AND(g9354, g7717)
--	g34483 = AND(g34406, g18938)
--	g18497 = AND(g2541, g15426)
--	g32029 = AND(g31318, g16482)
--	g24671 = AND(g5481, g23630)
--	g14831 = AND(g1152, g10909)
--	g22125 = AND(g6617, g19277)
--	g29382 = AND(g26424, g22763, g28172)
--	g27526 = AND(g26576, g17721)
--	g34862 = AND(g16540, g34830)
--	g29519 = AND(g2295, g28840)
--	g32028 = AND(g30569, g29339)
--	g19578 = AND(g16183, g11130)
--	g33415 = AND(g32368, g21422)
--	g22158 = AND(g13698, g19609)
--	g14316 = AND(g2370, g11920)
--	g33333 = AND(g32218, g20612)
--	g18700 = AND(g15132, g16816)
--	g17817 = AND(g11547, g6782, g11640, I18819)
--	g18126 = AND(g15054, g16971)
--	g18659 = AND(g4366, g17183)
--	g18625 = AND(g15092, g17062)
--	g18987 = AND(g182, g16162)
--	g29518 = AND(g28906, g22384)
--	g18250 = AND(g6821, g16897)
--	g24931 = AND(g23153, g20178)
--	g15114 = AND(g4239, g14454)
--	g25192 = AND(g20276, g23648)
--	g26847 = AND(g2873, g24525)
--	g34948 = AND(g16540, g34935)
--	g18658 = AND(g15121, g17183)
--	g27457 = AND(g26519, g17606)
--	g26397 = AND(g19475, g25563)
--	g15082 = AND(g2697, g12983)
--	g23387 = AND(g16506, g20211)
--	g31963 = AND(g30731, g18895)
--	g29637 = AND(g2533, g29134)
--	g22680 = AND(g19530, g7781)
--	g34702 = AND(g34537, g20208)
--	g15107 = AND(g4258, g14454)
--	g23148 = AND(g19128, g9104)
--	g34757 = AND(g34682, g19635)
--	g17783 = AND(g7851, g13110)
--	g25522 = AND(g6888, g22544)
--	I31121 = AND(g30614, g31817, g32629, g32630)
--	g24190 = AND(g329, g22722)
--	g18339 = AND(g1714, g17873)
--	g18943 = AND(g269, g16099)
--	g29883 = AND(g2465, g29152)
--	g18296 = AND(g1495, g16449)
--	g21811 = AND(g3582, g20924)
--	g28225 = AND(g27770, g23400)
--	g23104 = AND(g661, g20248)
--	g23811 = AND(g4087, g19364)
--	g23646 = AND(g16959, g20737)
--	g18644 = AND(g15098, g17125)
--	g28471 = AND(g27187, g12762, g21024, I26960)
--	g16221 = AND(g5791, g14231)
--	g18338 = AND(g1710, g17873)
--	g30564 = AND(g21358, g29385)
--	g9967 = AND(g1178, g1157)
--	g28258 = AND(g27182, g19687)
--	g21971 = AND(g5417, g21514)
--	g34564 = AND(g34373, g17466)
--	g15849 = AND(g3538, g14136)
--	g31484 = AND(g29775, g23418)
--	g24546 = AND(g22447, g19523)
--	g33484 = AND(g32628, I31116, I31117)
--	g16613 = AND(g5925, g14732)
--	I31291 = AND(g31021, g31847, g32875, g32876)
--	g15848 = AND(g3259, g13892)
--	g19275 = AND(g7823, g16044)
--	g31554 = AND(g19050, g29814)
--	g30673 = AND(g20175, g29814)
--	g27256 = AND(g25937, g19698)
--	g19746 = AND(g9816, g17147)
--	g28244 = AND(g27926, g26715)
--	g34183 = AND(g33695, g24385)
--	g18197 = AND(g854, g17821)
--	g22017 = AND(g5763, g21562)
--	g15652 = AND(g174, g13437)
--	g15804 = AND(g3223, g13889)
--	g34397 = AND(g7673, g34068)
--	g25949 = AND(g24701, g19559)
--	g27280 = AND(g9825, g26614)
--	g31312 = AND(g30136, g27858)
--	g29577 = AND(g2441, g28946)
--	g30062 = AND(g13129, g28174)
--	g27300 = AND(g12370, g26672)
--	g10736 = AND(g4040, g8751)
--	g10887 = AND(g7812, g6565, g6573)
--	g31115 = AND(g29487, g22882)
--	g18411 = AND(g2093, g15373)
--	g25536 = AND(g23770, g21431)
--	g25040 = AND(g12738, g23443)
--	g26213 = AND(g25357, g11724, g7586, g7558)
--	g34509 = AND(g34283, g19473)
--	g21850 = AND(g3893, g21070)
--	g28602 = AND(g27509, g20515)
--	g23412 = AND(g7297, g21510)
--	g28657 = AND(g27562, g20606)
--	g25904 = AND(g14001, g24791)
--	g33921 = AND(g33187, g9104, g19200)
--	g19684 = AND(g2735, g17297)
--	g34508 = AND(g34282, g19472)
--	g10528 = AND(g1576, g9051)
--	g34872 = AND(g34827, g19954)
--	I18740 = AND(g13156, g11450, g11498)
--	g24700 = AND(g645, g23512)
--	g28970 = AND(g17405, g25196, g26424, g27445)
--	g24659 = AND(g5134, g23590)
--	g14528 = AND(g12459, g12306, g12245, I16646)
--	g26205 = AND(g2098, g25492)
--	g23229 = AND(g18994, g4521)
--	g16234 = AND(g6772, g6782, g11640, I17575)
--	g29349 = AND(g4760, g28391)
--	g22309 = AND(g1478, g19751)
--	g20658 = AND(g1389, g15800)
--	g18503 = AND(g2563, g15509)
--	g22023 = AND(g5881, g19147)
--	g26311 = AND(g2527, g25400)
--	g24658 = AND(g22645, g19732)
--	I24015 = AND(g8334, g7975, g3045)
--	g10869 = AND(g7766, g5873, g5881)
--	g22308 = AND(g1135, g19738)
--	g28171 = AND(g27016, g19385)
--	g33798 = AND(g33227, g20058)
--	g21716 = AND(g301, g20283)
--	g30213 = AND(g28688, g23880)
--	g24296 = AND(g4382, g22550)
--	g18581 = AND(g2912, g16349)
--	g18714 = AND(g4864, g15915)
--	g26051 = AND(g24896, g14169)
--	g18450 = AND(g2299, g15224)
--	g31184 = AND(g1950, g30085)
--	g34213 = AND(g33766, g22689)
--	g18315 = AND(g1548, g16931)
--	g33805 = AND(g33232, g20079)
--	g33674 = AND(g33164, g10710, g22319)
--	g24644 = AND(g11714, g22903)
--	g29622 = AND(g2579, g29001)
--	g29566 = AND(g2307, g28907)
--	g18707 = AND(g15134, g16782)
--	g18819 = AND(g6541, g15483)
--	g18910 = AND(g16227, g16075)
--	g18202 = AND(g907, g15938)
--	g30047 = AND(g29109, g9407)
--	g18257 = AND(g1205, g16897)
--	g26780 = AND(g4098, g24437)
--	g30205 = AND(g28671, g23869)
--	g32191 = AND(g27593, g31376)
--	g18818 = AND(g15165, g15483)
--	g18496 = AND(g2537, g15426)
--	g34205 = AND(g33729, g24541)
--	g31934 = AND(g31670, g18827)
--	g18111 = AND(g174, g17015)
--	g21959 = AND(g5413, g21514)
--	g21925 = AND(g5073, g21468)
--	g26350 = AND(g13087, g25517)
--	g25872 = AND(g3119, g24655)
--	g28919 = AND(g27663, g21295)
--	g14708 = AND(g74, g12369)
--	I18762 = AND(g13156, g6767, g11498)
--	g28458 = AND(g27187, g12730, g20887, I26948)
--	g24197 = AND(g347, g22722)
--	g24855 = AND(g3050, g23534, I24027)
--	g27660 = AND(g24688, g26424, g22763)
--	g16163 = AND(g14254, g14179)
--	g22752 = AND(g15792, g19612)
--	g15613 = AND(g3490, g13555)
--	g18590 = AND(g2917, g16349)
--	g21958 = AND(g5396, g21514)
--	g21378 = AND(g7887, g16090)
--	g23050 = AND(g655, g20248)
--	g28010 = AND(g23032, g26223, g26424, g25535)
--	g23958 = AND(g9104, g19200)
--	g24411 = AND(g4584, g22161)
--	g30051 = AND(g28513, g20604)
--	g26846 = AND(g37, g24524)
--	g18741 = AND(g15143, g17384)
--	g34072 = AND(g33839, g24872)
--	g23386 = AND(g20034, g20207)
--	g30592 = AND(g30270, g18929)
--	g18384 = AND(g1945, g15171)
--	g29636 = AND(g2403, g29097)
--	g21742 = AND(g3050, g20330)
--	g17752 = AND(g7841, g13174)
--	g27480 = AND(g26400, g17638)
--	g34756 = AND(g34680, g19618)
--	g23742 = AND(g19128, g9104)
--	g28599 = AND(g27027, g8922)
--	g21944 = AND(g5244, g18997)
--	g33400 = AND(g32347, g21380)
--	g29852 = AND(g1772, g29080)
--	g17643 = AND(g9681, g14599)
--	g15812 = AND(g3227, g13915)
--	g13319 = AND(g4076, g8812, g10658, g8757)
--	g27314 = AND(g12436, g26702)
--	g24503 = AND(g22225, g19409)
--	g27287 = AND(g26545, g23011)
--	g32045 = AND(g31491, g16187)
--	I24685 = AND(g24036, g24037, g24038, g24039)
--	g33329 = AND(g32210, g20585)
--	g31207 = AND(g30252, g20739)
--	g18150 = AND(g604, g17533)
--	g10657 = AND(g8451, g4064)
--	g18801 = AND(g15160, g15348)
--	g18735 = AND(g4983, g16826)
--	g25574 = AND(I24709, I24710)
--	g27085 = AND(g25835, g22494)
--	g32324 = AND(g31315, g23537)
--	g29664 = AND(g2273, g29060)
--	g33328 = AND(g32209, g20584)
--	g21802 = AND(g3562, g20924)
--	g22489 = AND(g12954, g19386)
--	g21857 = AND(g3933, g21070)
--	g23802 = AND(g9104, g19050)
--	g16535 = AND(g5595, g14848)
--	g20581 = AND(g10801, g15571)
--	g10970 = AND(g854, g9582)
--	g23857 = AND(g19626, g7908)
--	g13059 = AND(g6900, g11303)
--	g13025 = AND(g8431, g11026)
--	g30152 = AND(g28609, g23767)
--	g24581 = AND(g5124, g23590)
--	g24714 = AND(g6173, g23699)
--	g32098 = AND(g4732, g30614)
--	g24450 = AND(g3129, g23067)
--	g21730 = AND(g3025, g20330)
--	g24315 = AND(g4521, g22228)
--	g21793 = AND(g3412, g20391)
--	g32272 = AND(g31639, g30310)
--	g22525 = AND(g13006, g19411)
--	g28159 = AND(g8553, g27317)
--	I31262 = AND(g32833, g32834, g32835, g32836)
--	g10878 = AND(g7858, g1135)
--	g18196 = AND(g703, g17821)
--	g22016 = AND(g5747, g21562)
--	g28125 = AND(g27381, g26209)
--	g15795 = AND(g3566, g14130)
--	g18695 = AND(g4737, g16053)
--	g28532 = AND(g27394, g20265)
--	g34396 = AND(g34194, g21337)
--	I18568 = AND(g13156, g11450, g11498)
--	g24707 = AND(g13295, g22997)
--	g30731 = AND(g11374, g29361)
--	g29576 = AND(g2177, g28903)
--	g29585 = AND(g1756, g28920)
--	g21765 = AND(g3231, g20785)
--	g28158 = AND(g26424, g22763, g27037)
--	I27523 = AND(g20857, g24111, g24112, g24113)
--	g18526 = AND(g2555, g15509)
--	g27269 = AND(g25943, g19734)
--	g29554 = AND(g28997, g22472)
--	g23690 = AND(g14726, g20978)
--	g19372 = AND(g686, g16289)
--	g26020 = AND(g9559, g25034)
--	g33241 = AND(g32173, g23128)
--	g34413 = AND(g34094, g22670)
--	g17424 = AND(g1426, g13176)
--	g11044 = AND(g5343, g10124)
--	I31191 = AND(g30735, g31829, g32731, g32732)
--	g27341 = AND(g10203, g26788)
--	g10967 = AND(g7880, g1448)
--	g29609 = AND(g28482, g11861)
--	g27268 = AND(g25942, g19733)
--	g32032 = AND(g31373, g16515)
--	g25780 = AND(g25532, g25527)
--	g15507 = AND(g10970, g13305)
--	g32140 = AND(g31609, g29961)
--	g28144 = AND(g4608, g27020)
--	g18402 = AND(g2047, g15373)
--	g18457 = AND(g2319, g15224)
--	g24590 = AND(g6154, g23413)
--	g29608 = AND(g28568, g11385)
--	g27180 = AND(g26026, g16654)
--	g19516 = AND(g7824, g16097)
--	g20094 = AND(g8872, g16631)
--	g27335 = AND(g12087, g26776)
--	g33683 = AND(g33149, g10727, g22332)
--	g13738 = AND(g8880, g10572)
--	g25152 = AND(g23383, g20626)
--	g22042 = AND(g5961, g19147)
--	g26302 = AND(g2393, g25349)
--	g26357 = AND(g22547, g25525)
--	g29799 = AND(g28271, g10233)
--	g30583 = AND(g19666, g29355)
--	g16760 = AND(g5559, g14764)
--	g27667 = AND(g26361, g20601)
--	I31247 = AND(g32812, g32813, g32814, g32815)
--	g18706 = AND(g4785, g16782)
--	g18597 = AND(g2975, g16349)
--	g27965 = AND(g25834, g13117)
--	g13290 = AND(g3897, g11534)
--	g29798 = AND(g28348, g23260)
--	g22124 = AND(g6613, g19277)
--	g27131 = AND(g26055, g16588)
--	g30046 = AND(g29108, g10564)
--	g18256 = AND(g1242, g16897)
--	g29973 = AND(g28981, g9206)
--	g18689 = AND(g15129, g16752)
--	g31991 = AND(g4912, g30673)
--	g33515 = AND(g32853, I31271, I31272)
--	g33882 = AND(g33293, g20587)
--	g18280 = AND(g1367, g16136)
--	g29805 = AND(g28357, g23270)
--	g33414 = AND(g32367, g21421)
--	g22686 = AND(g19335, g19577)
--	g22939 = AND(g9708, g21062)
--	g18688 = AND(g4704, g16752)
--	g18624 = AND(g3490, g17062)
--	g32162 = AND(g31002, g23014)
--	g18300 = AND(g1306, g16489)
--	g24196 = AND(g333, g22722)
--	g33407 = AND(g32357, g21406)
--	g34113 = AND(g33734, g19744)
--	g27502 = AND(g26488, g17677)
--	I31251 = AND(g31710, g31840, g32817, g32818)
--	g11427 = AND(g5706, g7158)
--	g22030 = AND(g5909, g19147)
--	I31272 = AND(g32849, g32850, g32851, g32852)
--	g22938 = AND(g19782, g19739)
--	g27557 = AND(g26549, g17774)
--	g22093 = AND(g6423, g18833)
--	g23533 = AND(g19436, g13015)
--	g11366 = AND(g5016, g10338)
--	g27210 = AND(g26218, g8373, g2476)
--	g21298 = AND(g7697, g15825)
--	g29732 = AND(g2514, g29131)
--	g28289 = AND(g27734, g26575)
--	g21775 = AND(g3372, g20391)
--	I16671 = AND(g10185, g12461, g12415)
--	g13632 = AND(g10232, g12228)
--	g18157 = AND(g15057, g17433)
--	g23775 = AND(g14872, g21267)
--	g22065 = AND(g6203, g19210)
--	g34105 = AND(g33778, g9104, g18957)
--	g28224 = AND(g27163, g22763, g27064)
--	g34743 = AND(g8951, g34703)
--	I17585 = AND(g14988, g11450, g11498)
--	g28571 = AND(g27458, g20435)
--	g24402 = AND(g4749, g22857)
--	g29761 = AND(g28310, g23228)
--	I31032 = AND(g32501, g32502, g32503, g32504)
--	g18231 = AND(g1105, g16326)
--	g21737 = AND(g3068, g20330)
--	g32246 = AND(g31246, g20326)
--	g27469 = AND(g8046, g26314, g518, g9077)
--	g22219 = AND(g19953, g20887)
--	g25928 = AND(g25022, g23436)
--	g8583 = AND(g2917, g2912)
--	g27286 = AND(g6856, g26634)
--	g33441 = AND(g32251, g29722)
--	g31206 = AND(g30260, g23890)
--	g10656 = AND(g3782, g7952)
--	g27039 = AND(g7738, g5527, g5535, g26223)
--	g22218 = AND(g19951, g20875)
--	g28495 = AND(g27012, g12465)
--	g32071 = AND(g27236, g31070)
--	I31061 = AND(g30825, g31806, g32543, g32544)
--	g21856 = AND(g3929, g21070)
--	g10823 = AND(g7704, g5180, g5188)
--	g14295 = AND(g1811, g11894)
--	g21995 = AND(g5611, g19074)
--	g31759 = AND(g21291, g29385)
--	g23856 = AND(g4116, g19483)
--	g14680 = AND(g12024, g12053)
--	g33759 = AND(g33123, g22847)
--	g33725 = AND(g22626, g10851, g33176)
--	g24001 = AND(g19651, g10951)
--	g21880 = AND(g4135, g19801)
--	g29329 = AND(g7995, g28353)
--	g25113 = AND(g23346, g20577)
--	g18511 = AND(g2599, g15509)
--	g29207 = AND(g24131, I27533, I27534)
--	g25787 = AND(g24792, g20887)
--	g32147 = AND(g31616, g29980)
--	g18763 = AND(g5481, g17929)
--	g31758 = AND(g30115, g23945)
--	g33114 = AND(g22139, g31945)
--	g24706 = AND(g15910, g22996)
--	g26249 = AND(g1858, g25300)
--	g33758 = AND(g33133, g20269)
--	g22160 = AND(g8005, g19795)
--	g27601 = AND(g26766, g26737)
--	g33082 = AND(g32389, g18877)
--	g21512 = AND(g16225, g10881)
--	g29328 = AND(g28553, g6928, g3990)
--	g27677 = AND(g13021, g25888)
--	g25357 = AND(g23810, g23786)
--	g29538 = AND(g2563, g28914)
--	g11127 = AND(g6479, g10022)
--	g24923 = AND(g23129, g20167)
--	g25105 = AND(g13973, g23505)
--	g10966 = AND(g9226, g7948)
--	g31744 = AND(g30092, g23902)
--	g24688 = AND(g22681, g22663)
--	g26204 = AND(g1720, g25275)
--	g24624 = AND(g16524, g22867)
--	g24300 = AND(g15123, g22228)
--	I24579 = AND(g5731, g5736, g9875)
--	g26779 = AND(g24497, g23620)
--	g33345 = AND(g32229, g20671)
--	g32151 = AND(g31639, g29996)
--	g32172 = AND(g2767, g31608)
--	I31162 = AND(g32689, g32690, g32691, g32692)
--	g31940 = AND(g943, g30735)
--	g18456 = AND(g2338, g15224)
--	g33849 = AND(g33262, g20387)
--	g30027 = AND(g29104, g12550)
--	g33399 = AND(g32346, g21379)
--	g21831 = AND(g3782, g20453)
--	g26778 = AND(g25501, g20923)
--	g34662 = AND(g34576, g18931)
--	g16845 = AND(g6593, g15011)
--	g11956 = AND(g2070, g7411)
--	g18480 = AND(g2437, g15426)
--	
--	g32367 = OR(g29880, g31309)
--	g34890 = OR(g34863, g21674)
--	g28668 = OR(g27411, g16617)
--	g34249 = OR(g34110, g21702)
--	g13095 = OR(g11374, g1287)
--	g30482 = OR(g30230, g21978)
--	g24231 = OR(g22589, g18201)
--	g13888 = OR(g2941, g11691)
--	g26945 = OR(g26379, g24283)
--	g30552 = OR(g30283, g22123)
--	g34003 = OR(g33866, g18452)
--	g23989 = OR(g20581, g17179)
--	g29235 = OR(g28110, g18260)
--	g28525 = OR(g27284, g26176)
--	g34204 = OR(g33832, g33833)
--	I28566 = OR(g29201, g29202, g29203, g28035)
--	g14309 = OR(g10320, g11048)
--	I30330 = OR(g29385, g31376, g30735, g30825)
--	g24854 = OR(g21453, g24002)
--	g30081 = OR(g28454, g11366)
--	g32227 = OR(g31146, g29648)
--	g33962 = OR(g33822, g18123)
--	g19575 = OR(g15693, g13042)
--	g27556 = OR(g26097, g24687)
--	g25662 = OR(g24656, g21787)
--	g28544 = OR(g27300, g26229)
--	g30356 = OR(g30096, g18365)
--	g27580 = OR(g26159, g24749)
--	g34647 = OR(g34558, g18820)
--	g26932 = OR(g26684, g18549)
--	I31859 = OR(g33501, g33502, g33503, g33504)
--	g33049 = OR(g31966, g21929)
--	g30380 = OR(g30161, g18492)
--	g34826 = OR(g34742, g34685)
--	g16926 = OR(g14061, g11804, g11780)
--	I25736 = OR(g12, g22150, g20277)
--	I31858 = OR(g33497, g33498, g33499, g33500)
--	g33048 = OR(g31960, g21928)
--	g7684 = OR(g4072, g4176)
--	g25710 = OR(g25031, g21961)
--	g28610 = OR(g27347, g16484)
--	g26897 = OR(g26611, g18176)
--	g34090 = OR(g33676, g33680)
--	g26961 = OR(g26280, g24306)
--	g28705 = OR(g27460, g16672)
--	g28042 = OR(g24148, g26879)
--	g30672 = OR(g13737, g29752)
--	g34233 = OR(g32455, g33951)
--	g13211 = OR(g11294, g7567)
--	g33004 = OR(g32246, g18431)
--	g31221 = OR(g29494, g28204)
--	g23198 = OR(g20214, g20199, I22298)
--	I31844 = OR(g33474, g33475, g33476, g33477)
--	g27179 = OR(g25816, g24409)
--	g28188 = OR(g22535, g27108)
--	g33613 = OR(g33248, g18649)
--	g34331 = OR(g27121, g34072)
--	g30513 = OR(g30200, g22034)
--	g30449 = OR(g29845, g21858)
--	g33947 = OR(g32438, g33457)
--	g34449 = OR(g34279, g18662)
--	g25647 = OR(g24725, g21740)
--	g24243 = OR(g22992, g18254)
--	g33273 = OR(g32122, g29553)
--	g28030 = OR(g24018, g26874)
--	g33605 = OR(g33352, g18521)
--	g25945 = OR(g24427, g22307)
--	g28093 = OR(g27981, g21951)
--	g30448 = OR(g29809, g21857)
--	g34897 = OR(g34861, g21682)
--	g34448 = OR(g34365, g18553)
--	g30505 = OR(g30168, g22026)
--	g29114 = OR(g27646, g26602)
--	g30404 = OR(g29758, g21763)
--	g28065 = OR(g27299, g21792)
--	g27800 = OR(g17321, g26703)
--	g24269 = OR(g23131, g18613)
--	g34404 = OR(g34182, g25102)
--	g33951 = OR(g33469, I31838, I31839)
--	g33972 = OR(g33941, g18335)
--	g24341 = OR(g23564, g18771)
--	g33033 = OR(g32333, g21843)
--	g24268 = OR(g23025, g18612)
--	g25651 = OR(g24680, g21744)
--	g25672 = OR(g24647, g21829)
--	g33234 = OR(g32039, g32043)
--	g34026 = OR(g33715, g18682)
--	g32427 = OR(g8928, g30583)
--	g13296 = OR(g10626, g10657)
--	g23087 = OR(g19487, g15852)
--	g29849 = OR(g26049, g28273)
--	g13969 = OR(g11448, g8913)
--	g26343 = OR(g1514, g24609)
--	g19522 = OR(g17057, g14180)
--	g29848 = OR(g28260, g26077)
--	g24335 = OR(g22165, g18678)
--	g26971 = OR(g26325, g24333)
--	g34723 = OR(g34710, g18139)
--	g30433 = OR(g29899, g21817)
--	g34149 = OR(g33760, g19674)
--	g30387 = OR(g30151, g18524)
--	g24965 = OR(g22667, g23825)
--	g32226 = OR(g31145, g29645)
--	g29263 = OR(g28239, g18617)
--	g34620 = OR(g34529, g18582)
--	g34148 = OR(g33758, g19656)
--	g25717 = OR(g25106, g21968)
--	g27543 = OR(g26085, g24670)
--	g30104 = OR(g28478, g11427)
--	g33012 = OR(g32274, g18483)
--	g19949 = OR(g17671, g14681)
--	g30343 = OR(g29344, g18278)
--	g34646 = OR(g34557, g18803)
--	g24557 = OR(g22308, g19207)
--	g24210 = OR(g22900, g18125)
--	g27569 = OR(g26124, g24721)
--	g34971 = OR(g34869, g34962)
--	g33541 = OR(g33101, g18223)
--	g31473 = OR(g26180, g29666)
--	g28075 = OR(g27083, g21877)
--	g30369 = OR(g30066, g18439)
--	g24443 = OR(g23917, g21378)
--	g19904 = OR(g17636, g14654)
--	g23171 = OR(g19536, g15903)
--	g24279 = OR(g23218, g15105)
--	g26896 = OR(g26341, g18171)
--	g34369 = OR(g26279, g34136)
--	g28595 = OR(g27335, g26290)
--	g14030 = OR(g11037, g11046)
--	g30368 = OR(g30098, g18435)
--	g24278 = OR(g23201, g18648)
--	g25723 = OR(g25033, g22006)
--	g28623 = OR(g27361, g16520)
--	g34368 = OR(g26274, g34135)
--	g33788 = OR(g33122, g32041)
--	g31325 = OR(g29625, g29639)
--	g32385 = OR(g31480, g29938)
--	g31920 = OR(g31493, g22045)
--	g32980 = OR(g32254, g18198)
--	g30412 = OR(g29885, g21771)
--	g33535 = OR(g33233, g21711)
--	g24468 = OR(g10925, g22400)
--	g32354 = OR(g29854, g31285)
--	g34850 = OR(g34841, g18185)
--	g34412 = OR(g34187, g25143)
--	g28419 = OR(g27221, g15884)
--	g27974 = OR(g26544, g25063)
--	g33946 = OR(g32434, g33456)
--	g25646 = OR(g24706, g21739)
--	g28418 = OR(g27220, g15882)
--	g20187 = OR(g16202, g13491)
--	g26959 = OR(g26381, g24299)
--	g26925 = OR(g25939, g18301)
--	g34011 = OR(g33884, g18479)
--	g26958 = OR(g26395, g24297)
--	g29273 = OR(g28269, g18639)
--	g31291 = OR(g29581, g29593)
--	g17570 = OR(g14419, g14397, g11999, I18495)
--	g33291 = OR(g32154, g13477)
--	g26386 = OR(g24719, g23023)
--	g32426 = OR(g26105, g26131, g30613)
--	g28194 = OR(g22540, g27122)
--	g28589 = OR(g27331, g26285)
--	g26944 = OR(g26130, g18658)
--	g20169 = OR(g16184, g13460)
--	g27579 = OR(g26157, g24748)
--	g29234 = OR(g28415, g18239)
--	g30379 = OR(g30089, g18491)
--	g34627 = OR(g34534, g18644)
--	g27578 = OR(g26155, g24747)
--	g17594 = OR(g14450, g14420, g12025, I18543)
--	g28401 = OR(g27212, g15871)
--	g31760 = OR(g30007, g30027)
--	g34379 = OR(g26312, g34143)
--	g33029 = OR(g32332, g21798)
--	g32211 = OR(g31124, g29603)
--	g30378 = OR(g30125, g18487)
--	g21901 = OR(g21251, g15115)
--	g20217 = OR(g16221, g13523)
--	g33028 = OR(g32325, g21797)
--	g30386 = OR(g30139, g18523)
--	g24363 = OR(g7831, g22138)
--	g26793 = OR(g24478, g7520)
--	g28118 = OR(g27821, g26815)
--	g13526 = OR(g209, g10685, g301)
--	g24478 = OR(g11003, g22450)
--	g34603 = OR(g34561, g15075)
--	g25716 = OR(g25088, g21967)
--	g28749 = OR(g27523, g16764)
--	g26690 = OR(g10776, g24433)
--	g25582 = OR(g21662, g24152)
--	g28748 = OR(g27522, g16763)
--	g28704 = OR(g27459, g16671)
--	g24580 = OR(g22340, g13096)
--	g31927 = OR(g31500, g22091)
--	g30429 = OR(g29844, g21813)
--	g28305 = OR(g27103, g15793)
--	g28053 = OR(g27393, g18168)
--	g32987 = OR(g32311, g18323)
--	g32250 = OR(g30598, g29351)
--	g34802 = OR(g34757, g18589)
--	g25627 = OR(g24503, g18247)
--	g30428 = OR(g29807, g21812)
--	g34730 = OR(g34658, g18271)
--	g34793 = OR(g34744, g18570)
--	I26643 = OR(g27073, g27058, g27045, g27040)
--	g13077 = OR(g11330, g943)
--	I18492 = OR(g14538, g14513, g14446)
--	g28101 = OR(g27691, g22062)
--	g33240 = OR(g32052, g32068)
--	g13597 = OR(g9247, g11149)
--	g28560 = OR(g27311, g26249)
--	g31903 = OR(g31374, g21911)
--	g30549 = OR(g30215, g22120)
--	g25603 = OR(g24698, g18114)
--	g25742 = OR(g25093, g22057)
--	g31755 = OR(g29991, g30008)
--	g33604 = OR(g33345, g18520)
--	g30548 = OR(g30204, g22119)
--	g10589 = OR(g7223, g7201)
--	g29325 = OR(g28813, g27820)
--	g13300 = OR(g10656, g10676)
--	g31770 = OR(g30034, g30047)
--	g30504 = OR(g30253, g22025)
--	g28064 = OR(g27298, g21781)
--	g33563 = OR(g33361, g18383)
--	g33981 = OR(g33856, g18371)
--	g25681 = OR(g24710, g18636)
--	g28733 = OR(g27507, g16735)
--	g26299 = OR(g24551, g22665)
--	g30317 = OR(g29208, I28566, I28567)
--	g25730 = OR(g25107, g22013)
--	g22304 = OR(g21347, g17693)
--	g14119 = OR(g10776, g8703)
--	g31767 = OR(g30031, g30043)
--	g33794 = OR(g33126, g32053)
--	g34002 = OR(g33857, g18451)
--	g33262 = OR(g32112, g29528)
--	g31899 = OR(g31470, g21907)
--	g34057 = OR(g33911, g33915)
--	g28665 = OR(g27409, g16614)
--	g30128 = OR(g28495, g11497)
--	g33990 = OR(g33882, g18399)
--	g24334 = OR(g23991, g18676)
--	g25690 = OR(g24864, g21889)
--	g26737 = OR(g24460, g10720)
--	g29291 = OR(g28660, g18767)
--	g31898 = OR(g31707, g21906)
--	g34626 = OR(g34533, g18627)
--	g30533 = OR(g30203, g22079)
--	g22653 = OR(g18993, g15654)
--	g30298 = OR(g28245, g27251)
--	g23687 = OR(g21384, g21363, I22830)
--	g26880 = OR(g26610, g24186)
--	g24216 = OR(g23416, g18197)
--	g23374 = OR(g19767, g13514)
--	g32202 = OR(g31069, g13410)
--	g22636 = OR(g18943, g15611)
--	g26512 = OR(g24786, g23130)
--	g32257 = OR(g31184, g29708)
--	g13660 = OR(g8183, g12527)
--	g32979 = OR(g32181, g18177)
--	g29506 = OR(g28148, g25880)
--	g34232 = OR(g33451, g33944)
--	g32978 = OR(g32197, g18145)
--	g28074 = OR(g27119, g21876)
--	g33573 = OR(g33343, g18415)
--	g31247 = OR(g29513, g13324)
--	g28594 = OR(g27334, g26289)
--	g31926 = OR(g31765, g22090)
--	g32986 = OR(g31996, g18280)
--	g27253 = OR(g24661, g26052)
--	g33389 = OR(g32272, g29964)
--	g33045 = OR(g32206, g24328)
--	g22664 = OR(g19139, g15694)
--	g34856 = OR(g34811, g34743)
--	g25626 = OR(g24499, g18235)
--	g33612 = OR(g33247, g18633)
--	g34261 = OR(g34074, g18688)
--	g34880 = OR(g34867, g18153)
--	g8921 = OR(I12902, I12903)
--	g30512 = OR(g30191, g22033)
--	g33534 = OR(g33186, g21700)
--	g27236 = OR(g24620, g25974)
--	g32094 = OR(g30612, g29363)
--	g31251 = OR(g25973, g29527)
--	g22585 = OR(g20915, g21061)
--	g33251 = OR(g32096, g29509)
--	g24242 = OR(g22834, g18253)
--	g33272 = OR(g32121, g29551)
--	g28092 = OR(g27666, g21924)
--	I30124 = OR(g31070, g31154, g30614, g30673)
--	g28518 = OR(g27281, g26158)
--	g21893 = OR(g20094, g18655)
--	g29240 = OR(g28655, g18328)
--	g26080 = OR(g19393, g24502)
--	I12583 = OR(g1157, g1239, g990)
--	g25737 = OR(g25045, g22052)
--	g26924 = OR(g26153, g18291)
--	g30445 = OR(g29772, g21854)
--	g33032 = OR(g32326, g21842)
--	g34445 = OR(g34382, g18548)
--	g30499 = OR(g30261, g21995)
--	g33997 = OR(g33871, g18427)
--	g25697 = OR(g25086, g21916)
--	g25856 = OR(g25518, g25510, g25488, g25462)
--	g30498 = OR(g30251, g21994)
--	g25261 = OR(g23348, g20193)
--	g33061 = OR(g32334, g22050)
--	g24265 = OR(g22316, g18560)
--	g26342 = OR(g8407, g24591)
--	g31766 = OR(g30029, g30042)
--	g31871 = OR(g30596, g18279)
--	g30611 = OR(g13671, g29743)
--	g24841 = OR(g21420, g23998)
--	g34611 = OR(g34508, g18565)
--	g23255 = OR(g19655, g16122)
--	g34722 = OR(g34707, g18137)
--	g26887 = OR(g26542, g24193)
--	g28729 = OR(g27502, g16732)
--	g28577 = OR(g27326, g26272)
--	g24510 = OR(g22488, g7567)
--	g30432 = OR(g29888, g21816)
--	g28728 = OR(g27501, g16730)
--	g29262 = OR(g28327, g18608)
--	g27542 = OR(g16190, g26094)
--	g27453 = OR(g25976, g24606)
--	g23383 = OR(g19756, g16222)
--	g24578 = OR(g2882, g23825)
--	g30461 = OR(g30219, g21932)
--	g30342 = OR(g29330, g18261)
--	g34461 = OR(g34291, g18681)
--	g26365 = OR(g25504, g25141)
--	I18452 = OR(g14514, g14448, g14418)
--	g26960 = OR(g26258, g24304)
--	g34031 = OR(g33735, g18705)
--	g31472 = OR(g29642, g28352)
--	g28083 = OR(g27249, g18689)
--	g28348 = OR(g27139, g15823)
--	g34199 = OR(g33820, g33828)
--	g32280 = OR(g24790, g31225)
--	g9984 = OR(g4300, g4242)
--	g34887 = OR(g34865, g21670)
--	g31911 = OR(g31784, g21969)
--	g30529 = OR(g30212, g22075)
--	g33628 = OR(g33071, g32450)
--	g27274 = OR(g15779, g25915)
--	g31246 = OR(g25965, g29518)
--	g25611 = OR(g24931, g18128)
--	g19356 = OR(g17784, g14874)
--	g25722 = OR(g25530, g18768)
--	g28622 = OR(g27360, g16519)
--	g28566 = OR(g27316, g26254)
--	g30528 = OR(g30202, g22074)
--	g9483 = OR(g1008, g969)
--	g30393 = OR(g29986, g21748)
--	g27122 = OR(g22537, g25917)
--	g34843 = OR(g33924, g34782)
--	g34330 = OR(g34069, g33717)
--	g30365 = OR(g30158, g18412)
--	g24275 = OR(g23474, g18645)
--	g29247 = OR(g28694, g18410)
--	g31591 = OR(g29358, g29353)
--	g31785 = OR(g30071, g30082)
--	g33591 = OR(g33082, g18474)
--	g24430 = OR(g23151, g8234)
--	g24746 = OR(g22588, g19461)
--	g32231 = OR(g30590, g29346)
--	g25753 = OR(g25165, g22100)
--	g31754 = OR(g29989, g30006)
--	g28138 = OR(g27964, g27968)
--	g24237 = OR(g22515, g18242)
--	g33950 = OR(g32450, g33460)
--	g29777 = OR(g28227, g28234)
--	g24340 = OR(g24016, g18770)
--	g25650 = OR(g24663, g21743)
--	g25736 = OR(g25536, g18785)
--	g29251 = OR(g28679, g18464)
--	g29272 = OR(g28346, g18638)
--	g28636 = OR(g27376, g16538)
--	g19449 = OR(g15567, g12939)
--	g28852 = OR(g27559, g16871)
--	g34259 = OR(g34066, g18679)
--	g30471 = OR(g30175, g21942)
--	g33996 = OR(g33862, g18426)
--	g34708 = OR(g33381, g34572)
--	g26657 = OR(g24908, g24900, g24887, g24861)
--	g25696 = OR(g25012, g21915)
--	g26955 = OR(g26391, g24293)
--	g34258 = OR(g34211, g18675)
--	g24517 = OR(g22158, g18906)
--	g26879 = OR(g25580, g25581)
--	g26970 = OR(g26308, g24332)
--	g25764 = OR(g25551, g18819)
--	g28664 = OR(g27408, g16613)
--	g26878 = OR(g25578, g25579)
--	g16867 = OR(g13493, g11045)
--	g25960 = OR(g24566, g24678)
--	g34043 = OR(g33903, g33905)
--	g26886 = OR(g26651, g24192)
--	g25868 = OR(g25450, g23885)
--	g28576 = OR(g27325, g26271)
--	g31319 = OR(g29612, g28324)
--	g27575 = OR(g26147, g24731)
--	g26967 = OR(g26350, g24319)
--	g33318 = OR(g31969, g32434)
--	g34602 = OR(g34489, g18269)
--	g25709 = OR(g25014, g21960)
--	g30375 = OR(g30149, g18466)
--	g34657 = OR(g33114, g34497)
--	g28609 = OR(g27346, g16483)
--	g33227 = OR(g32029, g32031)
--	g9536 = OR(g1351, g1312)
--	g33059 = OR(g31987, g22021)
--	g33025 = OR(g32162, g21780)
--	g25708 = OR(g25526, g18751)
--	g34970 = OR(g34868, g34961)
--	I29986 = OR(g31070, g31194, g30614, g30673)
--	g23822 = OR(g20218, g16929)
--	g33540 = OR(g33099, g18207)
--	g27108 = OR(g22522, g25911)
--	g33058 = OR(g31976, g22020)
--	g30337 = OR(g29334, g18220)
--	g32243 = OR(g31166, g29683)
--	g26919 = OR(g25951, g18267)
--	g28052 = OR(g27710, g18167)
--	g27283 = OR(g25922, g25924)
--	g26918 = OR(g25931, g18243)
--	g28745 = OR(g27519, g16760)
--	g15968 = OR(g13038, g10677)
--	I31854 = OR(g33492, g33493, g33494, g33495)
--	g33044 = OR(g32199, g24327)
--	g34792 = OR(g34750, g18569)
--	g32268 = OR(g24785, g31219)
--	g23194 = OR(g19564, g19578)
--	g33281 = OR(g32142, g29576)
--	g31902 = OR(g31744, g21910)
--	g30459 = OR(g29314, g21926)
--	g30425 = OR(g29770, g21809)
--	g33957 = OR(g33523, I31868, I31869)
--	g24347 = OR(g23754, g18790)
--	g34459 = OR(g34415, g18673)
--	g25602 = OR(g24673, g18113)
--	g12982 = OR(g12220, g9968)
--	g25657 = OR(g24624, g21782)
--	g24253 = OR(g22525, g18300)
--	g25774 = OR(g25223, g12043)
--	g29246 = OR(g28710, g18406)
--	g30458 = OR(g30005, g24330)
--	g34458 = OR(g34396, g18671)
--	g33562 = OR(g33414, g18379)
--	g34010 = OR(g33872, g18478)
--	g24236 = OR(g22489, g18241)
--	g25878 = OR(g25503, g23920)
--	g28732 = OR(g27505, g16734)
--	g33699 = OR(g32409, g33433)
--	g32993 = OR(g32255, g18352)
--	g30545 = OR(g30268, g22116)
--	g30444 = OR(g29901, g21853)
--	g29776 = OR(g28225, g22846)
--	g24952 = OR(g21326, g21340, I24117)
--	g24351 = OR(g23774, g18807)
--	g33290 = OR(g32149, g29589)
--	g26901 = OR(g26362, g24218)
--	g34444 = OR(g34389, g18546)
--	g24821 = OR(g21404, g23990)
--	g29754 = OR(g28215, g28218)
--	g34599 = OR(g34542, g18149)
--	g32131 = OR(g24495, g30926)
--	g20063 = OR(g15978, g13313)
--	g34598 = OR(g34541, g18136)
--	g15910 = OR(g13025, g10654)
--	g24264 = OR(g22310, g18559)
--	g23276 = OR(g19681, g16161)
--	g27663 = OR(g26323, g24820)
--	g28400 = OR(g27211, g15870)
--	g32210 = OR(g31123, g29600)
--	g21900 = OR(g20977, g15114)
--	g16866 = OR(g13492, g11044)
--	g28329 = OR(g27128, g15813)
--	g30532 = OR(g30193, g22078)
--	g32279 = OR(g31220, g31224)
--	g34125 = OR(g33724, g33124)
--	g22652 = OR(g18992, g15653)
--	g13762 = OR(g499, g12527)
--	g34977 = OR(g34873, g34966)
--	g25010 = OR(g23267, g2932)
--	g31895 = OR(g31505, g24296)
--	g28328 = OR(g27127, g15812)
--	g33547 = OR(g33349, g18331)
--	g34158 = OR(g33784, g19740)
--	g24209 = OR(g23415, g18122)
--	g34783 = OR(g33110, g34667)
--	g28538 = OR(g27294, g26206)
--	g26966 = OR(g26345, g24318)
--	g25545 = OR(g23551, g20658)
--	g30561 = OR(g30284, g22132)
--	g7673 = OR(g4153, g4172)
--	g30353 = OR(g30095, g18355)
--	g24208 = OR(g23404, g18121)
--	g25599 = OR(g24914, g21721)
--	g34353 = OR(g26088, g34114)
--	g29319 = OR(g28812, g14453)
--	g25598 = OR(g24904, g21720)
--	g33551 = OR(g33446, g18342)
--	g33572 = OR(g33339, g18414)
--	g30336 = OR(g29324, g18203)
--	g29227 = OR(g28456, g18169)
--	g13543 = OR(g10543, g10565)
--	I31839 = OR(g33465, g33466, g33467, g33468)
--	I31838 = OR(g33461, g33462, g33463, g33464)
--	g28100 = OR(g27690, g22051)
--	g20905 = OR(g7216, g17264)
--	g34631 = OR(g34562, g15118)
--	g30364 = OR(g30086, g18411)
--	g34017 = OR(g33880, g18504)
--	g24274 = OR(g23187, g18631)
--	g13242 = OR(g11336, g7601)
--	g33956 = OR(g33514, I31863, I31864)
--	g24346 = OR(g23725, g18789)
--	g33297 = OR(g32157, g29621)
--	g25656 = OR(g24945, g18609)
--	g31889 = OR(g31118, g21822)
--	g33980 = OR(g33843, g18370)
--	g24565 = OR(g22309, g19275)
--	g21892 = OR(g19788, g15104)
--	g25680 = OR(g24794, g21839)
--	g16876 = OR(g14028, g11773, g11755)
--	g29281 = OR(g28541, g18743)
--	g31888 = OR(g31067, g21821)
--	g20034 = OR(g15902, g13299)
--	g29301 = OR(g28686, g18797)
--	g27509 = OR(g26023, g24640)
--	g34289 = OR(g26847, g34218)
--	g24641 = OR(g22151, g22159)
--	g34023 = OR(g33796, g24320)
--	g34288 = OR(g26846, g34217)
--	g32217 = OR(g31129, g29616)
--	g26954 = OR(g26380, g24292)
--	I18449 = OR(g14512, g14445, g14415)
--	g31931 = OR(g31494, g22095)
--	g29290 = OR(g28569, g18764)
--	g25631 = OR(g24554, g18275)
--	g30495 = OR(g30222, g21991)
--	g32223 = OR(g31142, g29637)
--	g29366 = OR(g13738, g28439)
--	g27574 = OR(g26145, g24730)
--	g34976 = OR(g34872, g34965)
--	g26392 = OR(g24745, g23050)
--	g27205 = OR(g25833, g24421)
--	g33546 = OR(g33402, g18327)
--	g30374 = OR(g30078, g18465)
--	g16076 = OR(g13081, g10736)
--	g34374 = OR(g26294, g34139)
--	I30728 = OR(g32345, g32350, g32056, g32018)
--	g33024 = OR(g32324, g21752)
--	g34643 = OR(g34554, g18752)
--	g28435 = OR(g27234, g15967)
--	g28082 = OR(g27369, g24315)
--	g26893 = OR(g26753, g24199)
--	g29226 = OR(g28455, g18159)
--	g28744 = OR(g27518, g16759)
--	g34260 = OR(g34113, g18680)
--	g28345 = OR(g27137, g15821)
--	g29481 = OR(g28117, g28125)
--	g30392 = OR(g30091, g18558)
--	g30489 = OR(g30250, g21985)
--	g33625 = OR(g33373, g18809)
--	g32373 = OR(g29894, g31321)
--	g33987 = OR(g33847, g18396)
--	g31250 = OR(g25972, g29526)
--	g25687 = OR(g24729, g21882)
--	g30559 = OR(g30269, g22130)
--	g30525 = OR(g30266, g22071)
--	g30488 = OR(g30197, g21984)
--	g30424 = OR(g29760, g21808)
--	g25752 = OR(g25079, g22099)
--	g34016 = OR(g33867, g18503)
--	g30558 = OR(g30258, g22129)
--	g27152 = OR(g24393, g25817)
--	g33296 = OR(g32156, g29617)
--	g25643 = OR(g24602, g21736)
--	g29490 = OR(g25832, g28136)
--	g16839 = OR(g13473, g11035)
--	g28332 = OR(g27130, g15815)
--	g30544 = OR(g30257, g22115)
--	g33969 = OR(g33864, g18321)
--	g25669 = OR(g24657, g18624)
--	g28135 = OR(g27959, g27963)
--	g29297 = OR(g28683, g18784)
--	g33060 = OR(g31992, g22022)
--	g33968 = OR(g33855, g18320)
--	g26939 = OR(g25907, g21884)
--	g25668 = OR(g24646, g18623)
--	g33197 = OR(g32342, I30745, I30746)
--	g28361 = OR(g27153, g15839)
--	g32216 = OR(g31128, g29615)
--	g27405 = OR(g24572, g25968)
--	g26938 = OR(g26186, g21883)
--	g31870 = OR(g30607, g18262)
--	I28147 = OR(g2946, g24561, g28220)
--	g24840 = OR(g21419, g23996)
--	g34610 = OR(g34507, g18564)
--	g24390 = OR(g23779, g21285)
--	g30189 = OR(g23401, g28543)
--	g28049 = OR(g27684, g18164)
--	g34255 = OR(g34120, g24302)
--	g34189 = OR(g33801, g33808)
--	g30270 = OR(g28624, g27664)
--	g28048 = OR(g27362, g18163)
--	g20522 = OR(g691, g16893)
--	g26875 = OR(g21652, g25575)
--	g32117 = OR(g24482, g30914)
--	I23163 = OR(g20982, g21127, g21193, g21256)
--	g31894 = OR(g30671, g21870)
--	g31867 = OR(g31238, g18175)
--	g30460 = OR(g30207, g21931)
--	g30383 = OR(g30138, g18513)
--	g34460 = OR(g34301, g18677)
--	g30093 = OR(g28467, g11397)
--	g34030 = OR(g33727, g18704)
--	g25713 = OR(g25147, g21964)
--	g28613 = OR(g27350, g26310)
--	g33581 = OR(g33333, g18443)
--	g33714 = OR(g32419, g33450)
--	g29520 = OR(g28291, g28281, g28264, g28254)
--	g34267 = OR(g34079, g18728)
--	g34294 = OR(g26855, g34225)
--	g31315 = OR(g29607, g29623)
--	g33315 = OR(g29665, g32175)
--	g31910 = OR(g31471, g21957)
--	g13006 = OR(g12284, g10034)
--	g25610 = OR(g24923, g18127)
--	g31257 = OR(g29531, g28253)
--	g25705 = OR(g25069, g18744)
--	g28605 = OR(g27341, g26302)
--	g33257 = OR(g32108, g29519)
--	g32123 = OR(g30915, g30919)
--	g33979 = OR(g33942, g18361)
--	g33055 = OR(g31986, g21976)
--	g16187 = OR(g8822, g13486)
--	g25679 = OR(g24728, g21836)
--	g33070 = OR(g32010, g22114)
--	g33978 = OR(g33892, g18356)
--	g25678 = OR(g24709, g21835)
--	g26915 = OR(g25900, g18230)
--	g33590 = OR(g33358, g18470)
--	g15965 = OR(g13035, g10675)
--	g28371 = OR(g27177, g15847)
--	I30745 = OR(g31777, g32321, g32069, g32084)
--	g32230 = OR(g30589, g29345)
--	g33986 = OR(g33639, g18387)
--	g24252 = OR(g22518, g18299)
--	g25686 = OR(g24712, g21881)
--	g33384 = OR(g32248, g29943)
--	g33067 = OR(g31989, g22111)
--	g12768 = OR(g7785, g7202)
--	g29250 = OR(g28695, g18460)
--	g32992 = OR(g32242, g18351)
--	g32391 = OR(g31502, g29982)
--	g30455 = OR(g30041, g21864)
--	g34455 = OR(g34284, g18668)
--	g11372 = OR(g490, g482, g8038)
--	g31877 = OR(g31278, g21732)
--	g30470 = OR(g30165, g21941)
--	g34617 = OR(g34526, g18579)
--	g22648 = OR(g18987, g15652)
--	I12611 = OR(g1500, g1582, g1333)
--	g29296 = OR(g28586, g18781)
--	g33019 = OR(g32339, g18536)
--	g30201 = OR(g23412, g28557)
--	g33018 = OR(g32312, g18525)
--	I30761 = OR(g32071, g32167, g32067, g32082)
--	g30467 = OR(g30185, g21938)
--	g30494 = OR(g30209, g21990)
--	g34467 = OR(g34341, g18717)
--	g34494 = OR(g26849, g34413)
--	g29197 = OR(g27187, g27163)
--	g34623 = OR(g34525, g18585)
--	g34037 = OR(g33803, g18734)
--	I30400 = OR(g31021, g30937, g31327, g30614)
--	g27248 = OR(g24880, g25953)
--	g30984 = OR(g29765, g29755)
--	g27552 = OR(g26092, g24676)
--	g31917 = OR(g31478, g22003)
--	g30419 = OR(g29759, g21803)
--	g31866 = OR(g31252, g18142)
--	g30352 = OR(g30094, g18340)
--	g27779 = OR(g17317, g26694)
--	g25617 = OR(g25466, g18189)
--	g24213 = OR(g23220, g18186)
--	g23184 = OR(g20198, g20185, I22280)
--	g28724 = OR(g27491, g16707)
--	g34352 = OR(g26079, g34109)
--	g28359 = OR(g27151, g15838)
--	g30418 = OR(g29751, g21802)
--	g32275 = OR(g31210, g29732)
--	g31001 = OR(g29360, g28151)
--	g28358 = OR(g27149, g15837)
--	g34266 = OR(g34076, g18719)
--	g33001 = OR(g32282, g18404)
--	g34170 = OR(g33790, g19855)
--	g24205 = OR(g23006, g18109)
--	g33706 = OR(g32412, g33440)
--	g33597 = OR(g33344, g18495)
--	g32237 = OR(g31153, g29667)
--	g31256 = OR(g25983, g29537)
--	g33256 = OR(g32107, g29517)
--	g25595 = OR(g24835, g21717)
--	g31923 = OR(g31763, g22048)
--	g32983 = OR(g31990, g18222)
--	g19879 = OR(g15841, g13265)
--	g28344 = OR(g27136, g15820)
--	g22832 = OR(g19354, g15722)
--	g33280 = OR(g32141, g29574)
--	g25623 = OR(g24552, g18219)
--	g20051 = OR(g15936, g13306)
--	g25037 = OR(g23103, g19911)
--	g33624 = OR(g33371, g18808)
--	g34167 = OR(g33786, g19768)
--	g34194 = OR(g33811, g33815)
--	g26616 = OR(g24881, g24855, g24843, g24822)
--	g19337 = OR(g17770, g17785)
--	g28682 = OR(g27430, g16635)
--	g29257 = OR(g28228, g18600)
--	I23755 = OR(g22904, g22927, g22980, g23444)
--	g30524 = OR(g30255, g22070)
--	g27233 = OR(g25876, g24451)
--	g16800 = OR(g13436, g11027)
--	g29496 = OR(g28567, g27615)
--	g27182 = OR(g25818, g24410)
--	g30401 = OR(g29782, g21760)
--	g30477 = OR(g30239, g21948)
--	g26305 = OR(g24556, g24564)
--	g24350 = OR(g23755, g18806)
--	g26809 = OR(g24930, g24939)
--	g33066 = OR(g32341, g22096)
--	g26900 = OR(g26819, g24217)
--	g33231 = OR(g32032, g32036)
--	g29741 = OR(g28205, g15883)
--	g32130 = OR(g30921, g30925)
--	g34022 = OR(g33873, g18538)
--	g28134 = OR(g27958, g27962)
--	g31876 = OR(g31125, g21731)
--	g31885 = OR(g31017, g21779)
--	g32362 = OR(g29870, g31301)
--	g34616 = OR(g34519, g18577)
--	g25589 = OR(g21690, g24159)
--	g29801 = OR(g25987, g28251)
--	g29735 = OR(g28202, g10898)
--	g25588 = OR(g21686, g24158)
--	g34305 = OR(g25775, g34050)
--	g25836 = OR(g25368, g23856)
--	g27026 = OR(g26828, g17726)
--	g34254 = OR(g34116, g24301)
--	g30466 = OR(g30174, g21937)
--	g34809 = OR(g33677, g34738)
--	g34900 = OR(g34860, g21686)
--	g26733 = OR(g10776, g24447)
--	g34466 = OR(g34337, g18716)
--	g34808 = OR(g34765, g18599)
--	g32222 = OR(g31141, g29636)
--	g23771 = OR(g21432, g21416, I22912)
--	g26874 = OR(I25612, I25613)
--	g34036 = OR(g33722, g18715)
--	g30560 = OR(g30278, g22131)
--	g34101 = OR(g33693, g33700)
--	g31916 = OR(g31756, g22002)
--	g34642 = OR(g34482, g18725)
--	g25749 = OR(g25094, g18800)
--	g25616 = OR(g25096, g18172)
--	g28649 = OR(g27390, g16597)
--	g33550 = OR(g33342, g18338)
--	g32347 = OR(g29839, g31273)
--	g33314 = OR(g29663, g32174)
--	g31287 = OR(g29578, g28292)
--	g15800 = OR(g10821, g13242)
--	g32253 = OR(g24771, g31207)
--	g25748 = OR(g25078, g18799)
--	g33287 = OR(g32146, g29586)
--	g34064 = OR(g33919, g33922)
--	g30733 = OR(g13807, g29773)
--	g31307 = OR(g29596, g28311)
--	g33076 = OR(g32336, g32446)
--	g34733 = OR(g34678, g18651)
--	g26892 = OR(g26719, g24198)
--	g25704 = OR(g25173, g21925)
--	g22447 = OR(g21464, g12761)
--	g33596 = OR(g33341, g18494)
--	g33054 = OR(g31975, g21975)
--	g32236 = OR(g31152, g29664)
--	g8790 = OR(I12782, I12783)
--	g32351 = OR(g29851, g31281)
--	g32372 = OR(g29884, g31314)
--	g34630 = OR(g34560, g15117)
--	g34693 = OR(g34513, g34310)
--	g24282 = OR(g23407, g18657)
--	g26914 = OR(g25949, g18227)
--	g29706 = OR(g28198, g27208)
--	g8461 = OR(g301, g534)
--	g31269 = OR(g26024, g29569)
--	g34166 = OR(g33785, g19752)
--	g34009 = OR(g33863, g18477)
--	g19336 = OR(g17769, g14831)
--	g26907 = OR(g26513, g24224)
--	g29256 = OR(g28597, g18533)
--	g31773 = OR(g30044, g30056)
--	I30399 = OR(g29385, g31376, g30735, g30825)
--	g31268 = OR(g29552, g28266)
--	g32264 = OR(g31187, g29711)
--	g34008 = OR(g33849, g18476)
--	g29280 = OR(g28530, g18742)
--	g33268 = OR(g32116, g29538)
--	g30476 = OR(g30229, g21947)
--	g30485 = OR(g30166, g21981)
--	g29300 = OR(g28666, g18796)
--	g31670 = OR(g29937, g28573)
--	g8904 = OR(g1779, g1798)
--	I31863 = OR(g33506, g33507, g33508, g33509)
--	g30555 = OR(g30227, g22126)
--	g30454 = OR(g29909, g21863)
--	g34454 = OR(g34414, g18667)
--	g25733 = OR(g25108, g18778)
--	g13091 = OR(g329, g319, g10796)
--	g22591 = OR(g18893, g18909)
--	g27133 = OR(g25788, g24392)
--	g28719 = OR(g27485, g16703)
--	g28191 = OR(g27217, g27210, g27186, g27162)
--	g31930 = OR(g31769, g22094)
--	g32209 = OR(g31122, g29599)
--	g33993 = OR(g33646, g18413)
--	g25630 = OR(g24532, g18263)
--	g28718 = OR(g27483, g16702)
--	g25693 = OR(g24627, g18707)
--	g29231 = OR(g28301, g18229)
--	g33694 = OR(g32402, g33429)
--	g32208 = OR(g31120, g29584)
--	g33965 = OR(g33805, g18179)
--	I12783 = OR(g4204, g4207, g4210, g4180)
--	g25665 = OR(g24708, g21790)
--	g34239 = OR(g32845, g33957)
--	g34238 = OR(g32780, g33956)
--	g23345 = OR(g19735, g16203)
--	g26883 = OR(g26670, g24189)
--	I23162 = OR(g19919, g19968, g20014, g20841)
--	g33619 = OR(g33359, g18758)
--	g33557 = OR(g33331, g18363)
--	g29763 = OR(g28217, g22762)
--	g30382 = OR(g30137, g18498)
--	g30519 = OR(g30264, g22040)
--	g33618 = OR(g33353, g18757)
--	g28389 = OR(g27206, g15860)
--	g30176 = OR(g23392, g28531)
--	g28045 = OR(g27378, g18141)
--	g30092 = OR(g28466, g16699)
--	g31279 = OR(g29571, g29579)
--	g24249 = OR(g22624, g18294)
--	g33279 = OR(g32140, g29573)
--	g25712 = OR(g25126, g21963)
--	g28099 = OR(g27992, g22043)
--	g30518 = OR(g30254, g22039)
--	I22280 = OR(g20271, g20150, g20134)
--	g28388 = OR(g27204, g15859)
--	g16430 = OR(g182, g13657)
--	g28701 = OR(g27455, g16669)
--	g24248 = OR(g22710, g18286)
--	g33278 = OR(g32139, g29572)
--	g12925 = OR(g8928, g10511)
--	g28777 = OR(g27539, g16807)
--	g28534 = OR(g27292, g26204)
--	g28098 = OR(g27683, g22016)
--	g32346 = OR(g29838, g31272)
--	g34637 = OR(g34478, g18694)
--	g24204 = OR(g22990, g18108)
--	g33286 = OR(g32145, g29585)
--	g31468 = OR(g29641, g29656)
--	g31306 = OR(g29595, g29610)
--	I31873 = OR(g33524, g33525, g33526, g33527)
--	g33039 = OR(g32187, g24312)
--	g29480 = OR(g28115, g22172)
--	g27742 = OR(g17292, g26673)
--	g22318 = OR(g21394, g17783)
--	g25594 = OR(g24772, g21708)
--	g33038 = OR(g32184, g24311)
--	g29287 = OR(g28555, g18760)
--	g29307 = OR(g28706, g18814)
--	g28140 = OR(I26643, I26644)
--	g26349 = OR(g24630, g13409)
--	g33601 = OR(g33422, g18508)
--	g25941 = OR(g24416, g22219)
--	g33187 = OR(g32014, I30740, I30741)
--	g33975 = OR(g33860, g18346)
--	g27429 = OR(g25969, g24589)
--	g26906 = OR(g26423, g24223)
--	g25675 = OR(g24769, g21832)
--	g29243 = OR(g28657, g18358)
--	g26348 = OR(g8466, g24609)
--	g30501 = OR(g29327, g22018)
--	g28061 = OR(g27287, g21735)
--	g34729 = OR(g34666, g18270)
--	g32408 = OR(g31541, g30073)
--	g30439 = OR(g29761, g21848)
--	g34728 = OR(g34661, g18214)
--	g34439 = OR(g34344, g18181)
--	g29269 = OR(g28249, g18634)
--	g25637 = OR(g24618, g18307)
--	g24233 = OR(g22590, g18236)
--	g25935 = OR(g24402, g22208)
--	g30438 = OR(g29890, g21847)
--	g19525 = OR(g7696, g16811)
--	g19488 = OR(g16965, g14148)
--	g34438 = OR(g34348, g18150)
--	g29268 = OR(g28343, g18625)
--	I25613 = OR(g25571, g25572, g25573, g25574)
--	g31884 = OR(g31290, g21778)
--	g33791 = OR(g33379, g32430)
--	g30349 = OR(g30051, g18333)
--	g34349 = OR(g26019, g34104)
--	g8417 = OR(g1056, g1116, I12583)
--	g30348 = OR(g30083, g18329)
--	g22645 = OR(g18982, g15633)
--	g34906 = OR(g34857, g21694)
--	g29734 = OR(g28201, g15872)
--	g30304 = OR(g28255, g27259)
--	g33015 = OR(g32343, g18507)
--	g34622 = OR(g34520, g18584)
--	g25729 = OR(g25091, g22012)
--	g26636 = OR(g24897, g24884, g24858, g24846)
--	g28629 = OR(g27371, g16532)
--	g25577 = OR(g24143, g24144)
--	g28220 = OR(g23495, I26741, I26742)
--	g25728 = OR(g25076, g22011)
--	g28628 = OR(g27370, g16531)
--	g33556 = OR(g33329, g18362)
--	g24212 = OR(g23280, g18155)
--	g26963 = OR(g26306, g24308)
--	g33580 = OR(g33330, g18442)
--	g29487 = OR(g25815, g28133)
--	g23795 = OR(g20203, g16884)
--	g28071 = OR(g27085, g21873)
--	g29502 = OR(g28139, g25871)
--	g27533 = OR(g26078, g24659)
--	I29351 = OR(g29328, g29323, g29316, g30316)
--	g28591 = OR(g27332, g26286)
--	g25906 = OR(g25559, g24014)
--	g28776 = OR(g27538, g13974)
--	g30415 = OR(g29843, g21799)
--	g30333 = OR(g29834, g21699)
--	g34636 = OR(g34476, g18693)
--	g22547 = OR(g16855, g20215)
--	g29279 = OR(g28442, g18741)
--	g31922 = OR(g31525, g22047)
--	g32982 = OR(g31948, g18208)
--	g33321 = OR(g29712, g32182)
--	g25622 = OR(g24546, g18217)
--	g29278 = OR(g28626, g18740)
--	g19267 = OR(g17752, g17768)
--	g22226 = OR(g21333, g17655)
--	g24433 = OR(g10878, g22400)
--	g20148 = OR(g16128, g13393)
--	g29286 = OR(g28542, g18759)
--	g27232 = OR(g25874, g24450)
--	g7404 = OR(g933, g939)
--	g29306 = OR(g28689, g18813)
--	g28172 = OR(g27469, g27440, g27416, g27395)
--	g33685 = OR(g32396, g33423)
--	g7764 = OR(g2999, g2932)
--	g33953 = OR(g33487, I31848, I31849)
--	g24343 = OR(g23724, g18773)
--	g26921 = OR(g25955, g18285)
--	g25653 = OR(g24664, g18602)
--	g32390 = OR(g31501, g29979)
--	g27261 = OR(g24544, g25996)
--	g30484 = OR(g30154, g21980)
--	g30554 = OR(g30216, g22125)
--	g22490 = OR(g21513, g12795)
--	g13820 = OR(g11184, g9187, g12527)
--	g26813 = OR(g24940, g24949)
--	g15727 = OR(g13383, g13345, g13333, g11010)
--	g25636 = OR(g24507, g18305)
--	g30609 = OR(g13633, g29742)
--	g34609 = OR(g34503, g18563)
--	g28420 = OR(g27222, g13290)
--	g30608 = OR(g13604, g29736)
--	g28319 = OR(g27115, g15807)
--	g30115 = OR(g28489, g11449)
--	g29143 = OR(g27650, g17146)
--	g34608 = OR(g34568, g15082)
--	g17490 = OR(g14364, g14337, g11958, I18421)
--	g26805 = OR(g10776, g24478)
--	g31762 = OR(g30011, g30030)
--	g23358 = OR(g19746, g16212)
--	I30760 = OR(g31778, g32295, g32046, g32050)
--	g31964 = OR(g31654, g14544)
--	g33964 = OR(g33817, g18146)
--	g25664 = OR(g24681, g21789)
--	g28059 = OR(g27042, g18276)
--	g29791 = OR(g28233, g22859)
--	g16021 = OR(g13047, g10706)
--	g26934 = OR(g26845, g18556)
--	g28058 = OR(g27235, g18268)
--	g29168 = OR(g27658, g26613)
--	g33587 = OR(g33363, g18463)
--	g24896 = OR(g22863, g19684)
--	g34799 = OR(g34751, g18578)
--	g25585 = OR(g21674, g24155)
--	g25576 = OR(g24141, g24142)
--	g29479 = OR(g28113, g28116)
--	g34798 = OR(g34754, g18575)
--	g31909 = OR(g31750, g21956)
--	g28044 = OR(g27256, g18130)
--	g33543 = OR(g33106, g18281)
--	g19595 = OR(g17149, g14218)
--	g29478 = OR(g28111, g22160)
--	g19467 = OR(g16896, g14097)
--	g25609 = OR(g24915, g18126)
--	g34805 = OR(g34748, g18594)
--	g31908 = OR(g31519, g21955)
--	g33000 = OR(g32270, g18403)
--	g29486 = OR(g28537, g27595)
--	g32252 = OR(g31183, g31206)
--	g25608 = OR(g24643, g18120)
--	g33569 = OR(g33415, g18402)
--	g30732 = OR(g13778, g29762)
--	g27271 = OR(g24547, g26053)
--	I18495 = OR(g14539, g14515, g14449)
--	g34732 = OR(g34686, g18593)
--	g26329 = OR(g8526, g24609)
--	g33568 = OR(g33409, g18395)
--	g25745 = OR(g25150, g22060)
--	g29223 = OR(g28341, g18131)
--	g26328 = OR(g1183, g24591)
--	g28562 = OR(g27313, g26251)
--	g14844 = OR(g10776, g8703)
--	g34761 = OR(g34679, g34506)
--	g28699 = OR(g27452, g16667)
--	g27031 = OR(g26213, g26190, g26166, g26148)
--	g33123 = OR(g31962, g30577)
--	I30755 = OR(g30564, g32303, g32049, g32055)
--	g28698 = OR(g27451, g16666)
--	g31751 = OR(g29975, g29990)
--	g31772 = OR(g30035, g28654)
--	g30400 = OR(g29766, g21759)
--	g33974 = OR(g33846, g18345)
--	g30214 = OR(g23424, g28572)
--	g34013 = OR(g33901, g18488)
--	g25805 = OR(g25453, g25414, g25374, g25331)
--	g25674 = OR(g24755, g21831)
--	g31293 = OR(g29582, g28299)
--	g33293 = OR(g32151, g29602)
--	g30539 = OR(g30267, g22085)
--	g34207 = OR(g33835, g33304)
--	g22659 = OR(g19062, g15673)
--	g22625 = OR(g18910, g18933)
--	g25732 = OR(g25201, g22017)
--	g34005 = OR(g33883, g18454)
--	g28632 = OR(g27373, g16535)
--	g33265 = OR(g32113, g29530)
--	g30538 = OR(g30256, g22084)
--	g29373 = OR(g13832, g28453)
--	I30262 = OR(g31672, g31710, g31021, g30937)
--	g33992 = OR(g33900, g18408)
--	g25761 = OR(g25152, g18812)
--	g28661 = OR(g27406, g16611)
--	g28403 = OR(g27214, g13282)
--	g22644 = OR(g18981, g15632)
--	I12782 = OR(g4188, g4194, g4197, g4200)
--	g33579 = OR(g33357, g18437)
--	g14044 = OR(g10776, g8703)
--	g28715 = OR(g27480, g16700)
--	I30718 = OR(g32348, g32356, g32097, g32020)
--	g33578 = OR(g33410, g18433)
--	g31014 = OR(g29367, g28160)
--	g27225 = OR(g2975, g26364)
--	g33014 = OR(g32305, g18499)
--	g23770 = OR(g20188, g16868)
--	g26882 = OR(g26650, g24188)
--	g28551 = OR(g27305, g26234)
--	g31007 = OR(g29364, g28159)
--	g27258 = OR(g25905, g15749)
--	g34100 = OR(g33690, g33697)
--	g33586 = OR(g33416, g18459)
--	g33007 = OR(g32331, g18455)
--	g25539 = OR(g23531, g20628)
--	g13662 = OR(g10896, g10917)
--	g34235 = OR(g32585, g33953)
--	g27244 = OR(g24652, g25995)
--	g28490 = OR(g27262, g16185)
--	g33116 = OR(g32403, g32411)
--	g33615 = OR(g33113, g21871)
--	g23262 = OR(g19661, g16126)
--	g21899 = OR(g20162, g15113)
--	g30515 = OR(g30223, g22036)
--	g30414 = OR(g30002, g21794)
--	g28385 = OR(g27201, g15857)
--	g33041 = OR(g32189, g24323)
--	g28297 = OR(g27096, g15785)
--	g21898 = OR(g20152, g15112)
--	g34882 = OR(g34876, g18659)
--	g28103 = OR(g27696, g22097)
--	g24245 = OR(g22849, g18256)
--	g33275 = OR(g32127, g29564)
--	g28095 = OR(g27674, g21970)
--	g30407 = OR(g29794, g21766)
--	g34407 = OR(g34185, g25124)
--	g27970 = OR(g26514, g25050)
--	g31465 = OR(g26156, g29647)
--	g26759 = OR(g24468, g7511)
--	g26725 = OR(g24457, g10719)
--	g28671 = OR(g27413, g16619)
--	g33983 = OR(g33877, g18373)
--	g22707 = OR(g20559, g17156)
--	g33035 = OR(g32019, g21872)
--	g27886 = OR(g14438, g26759)
--	g25683 = OR(g24669, g18641)
--	g29242 = OR(g28674, g18354)
--	g26082 = OR(g2898, g24561)
--	g11380 = OR(g8583, g8530)
--	g30441 = OR(g29787, g21850)
--	g34441 = OR(g34381, g18540)
--	g24232 = OR(g22686, g18228)
--	g34206 = OR(g33834, g33836)
--	g26940 = OR(g25908, g21886)
--	I25612 = OR(g25567, g25568, g25569, g25570)
--	g34725 = OR(g34700, g18183)
--	g24261 = OR(g22862, g18314)
--	g29230 = OR(g28107, g18202)
--	g27458 = OR(g24590, g25989)
--	g29293 = OR(g28570, g18777)
--	g30114 = OR(g28488, g16761)
--	g30435 = OR(g30025, g21840)
--	g29265 = OR(g28318, g18620)
--	g28546 = OR(g27302, g26231)
--	g28089 = OR(g27269, g18731)
--	g23251 = OR(g19637, g16098)
--	g28211 = OR(g27029, g27034)
--	g34107 = OR(g33710, g33121)
--	g19555 = OR(g15672, g13030)
--	g28088 = OR(g27264, g18729)
--	g30345 = OR(g29644, g18302)
--	g30399 = OR(g29757, g21758)
--	g34849 = OR(g34842, g18154)
--	g34399 = OR(g34178, g25067)
--	g25584 = OR(g21670, g24154)
--	g28497 = OR(g27267, g16199)
--	g33006 = OR(g32291, g18447)
--	g30398 = OR(g29749, g21757)
--	g26962 = OR(g26295, g24307)
--	g26361 = OR(g24674, g22991)
--	g23997 = OR(g20602, g17191)
--	g30141 = OR(g28499, g16844)
--	g34804 = OR(g34740, g18591)
--	g28700 = OR(g27454, g16668)
--	g25759 = OR(g25166, g22106)
--	g28659 = OR(g27404, g16610)
--	g25725 = OR(g25127, g22008)
--	g28625 = OR(g27363, g26324)
--	g14888 = OR(g10776, g8703)
--	g32357 = OR(g29865, g31296)
--	g27159 = OR(g25814, g12953)
--	g27532 = OR(g16176, g26084)
--	g25758 = OR(g25151, g22105)
--	g34263 = OR(g34078, g18699)
--	g34332 = OR(g34071, g33723)
--	g33703 = OR(g32410, g33434)
--	g28296 = OR(g27095, g15784)
--	g31253 = OR(g25980, g29533)
--	g27561 = OR(g26100, g24702)
--	g33253 = OR(g32103, g29511)
--	g25744 = OR(g25129, g22059)
--	g28644 = OR(g27387, g16593)
--	g30406 = OR(g29783, g21765)
--	g24432 = OR(g23900, g21361)
--	g30361 = OR(g30109, g18391)
--	g34406 = OR(g34184, g25123)
--	g24271 = OR(g23451, g18628)
--	g33600 = OR(g33418, g18501)
--	g25940 = OR(g24415, g22218)
--	g31781 = OR(g30058, g30069)
--	g23162 = OR(g20184, g20170, I22267)
--	g33236 = OR(g32044, g32045)
--	g30500 = OR(g29326, g21996)
--	g29275 = OR(g28165, g21868)
--	g28060 = OR(g27616, g18532)
--	g33952 = OR(g33478, I31843, I31844)
--	g24342 = OR(g23691, g18772)
--	g25652 = OR(g24777, g21747)
--	g26947 = OR(g26394, g24285)
--	g8905 = OR(g2204, g2223)
--	g29237 = OR(g28185, g18289)
--	g28527 = OR(g27286, g26182)
--	g33063 = OR(g31988, g22066)
--	g34004 = OR(g33879, g18453)
--	g26951 = OR(g26390, g24289)
--	g26972 = OR(g26780, g25229)
--	g31873 = OR(g31270, g21728)
--	g19501 = OR(g16986, g14168)
--	g34613 = OR(g34515, g18567)
--	g32249 = OR(g31169, g29687)
--	g30605 = OR(g29529, g29520)
--	g27289 = OR(g25925, g25927)
--	g34273 = OR(g27765, g34203)
--	g34605 = OR(g34566, g15077)
--	g18879 = OR(g17365, g14423)
--	g28581 = OR(g27329, g26276)
--	g27224 = OR(g25870, g15678)
--	g30463 = OR(g30140, g21934)
--	g27571 = OR(g26127, g24723)
--	g28707 = OR(g27461, g16673)
--	g34463 = OR(g34338, g18686)
--	g23825 = OR(g20705, g20781)
--	g30371 = OR(g30099, g18445)
--	g28818 = OR(g27549, g13998)
--	g34033 = OR(g33821, g18708)
--	g34234 = OR(g32520, g33952)
--	g28055 = OR(g27560, g18190)
--	g33542 = OR(g33102, g18265)
--	g33021 = OR(g32302, g21749)
--	g24259 = OR(g23008, g18312)
--	g28070 = OR(g27050, g21867)
--	g31913 = OR(g31485, g21999)
--	g18994 = OR(g16303, g13632)
--	g24471 = OR(g10999, g22450)
--	g34795 = OR(g34753, g18572)
--	g25613 = OR(g25181, g18140)
--	g24258 = OR(g22851, g18311)
--	g33614 = OR(g33249, g18650)
--	g17511 = OR(g14396, g14365, g11976, I18452)
--	g32999 = OR(g32337, g18401)
--	g33607 = OR(g33091, g18526)
--	g31905 = OR(g31746, g21952)
--	g31320 = OR(g26125, g29632)
--	g30514 = OR(g30211, g22035)
--	g32380 = OR(g29907, g31467)
--	g31274 = OR(g29565, g28280)
--	g25605 = OR(g24743, g18116)
--	g29222 = OR(g28252, g18105)
--	g24244 = OR(g23349, g18255)
--	g33274 = OR(g32126, g29563)
--	g30507 = OR(g30190, g22028)
--	g32998 = OR(g32300, g18393)
--	g28094 = OR(g27673, g21959)
--	g28067 = OR(g27309, g21827)
--	g33593 = OR(g33417, g18482)
--	g26789 = OR(g10776, g24471)
--	g32233 = OR(g31150, g29661)
--	g12954 = OR(g12186, g9906)
--	g23319 = OR(g19717, g16193)
--	g30421 = OR(g29784, g21805)
--	g33565 = OR(g33338, g18389)
--	g34421 = OR(g27686, g34198)
--	g26359 = OR(g24651, g22939)
--	g28735 = OR(g27510, g16737)
--	g23318 = OR(g19716, g16192)
--	g30163 = OR(g23381, g28523)
--	g33034 = OR(g32340, g21844)
--	g26920 = OR(g25865, g18283)
--	g34012 = OR(g33886, g18480)
--	g29253 = OR(g28697, g18490)
--	g24879 = OR(g21465, g24009)
--	g33292 = OR(g32150, g29601)
--	g26946 = OR(g26389, g24284)
--	g30541 = OR(g30281, g22087)
--	g30473 = OR(g30196, g21944)
--	g24337 = OR(g23540, g18754)
--	g27489 = OR(g24608, g26022)
--	g29236 = OR(g28313, g18287)
--	g28526 = OR(g27285, g26178)
--	g26344 = OR(g2927, g25010)
--	g27016 = OR(g26821, g14585)
--	g30359 = OR(g30075, g18385)
--	g34724 = OR(g34702, g18152)
--	g28402 = OR(g27213, g15873)
--	g30535 = OR(g30225, g22081)
--	g30434 = OR(g30024, g21818)
--	g19576 = OR(g17138, g14202)
--	g30358 = OR(g30108, g18381)
--	g34535 = OR(g34309, g34073)
--	g29264 = OR(g28248, g18618)
--	g29790 = OR(g25975, g28242)
--	g16928 = OR(g13525, g11127)
--	g27544 = OR(g26087, g24671)
--	g33164 = OR(g32203, I30727, I30728)
--	g17268 = OR(g9220, g14387)
--	g24919 = OR(g21606, g22143)
--	g30344 = OR(g29630, g18298)
--	g31891 = OR(g31305, g21824)
--	g28077 = OR(g27120, g21879)
--	g33891 = OR(g33264, g33269)
--	g31474 = OR(g29668, g13583)
--	g33575 = OR(g33086, g18420)
--	g24444 = OR(g10890, g22400)
--	g30291 = OR(g28672, g27685)
--	g25789 = OR(g25285, g14543)
--	g32387 = OR(g31489, g29952)
--	g25724 = OR(g25043, g22007)
--	g28688 = OR(g27435, g16639)
--	g33537 = OR(g33244, g21716)
--	g22487 = OR(g21512, g12794)
--	g28102 = OR(g27995, g22089)
--	g33283 = OR(g31995, g30318)
--	g27383 = OR(g24569, g25961)
--	g33606 = OR(g33369, g18522)
--	g31303 = OR(g29592, g29606)
--	g33303 = OR(g32159, g29638)
--	g34029 = OR(g33798, g18703)
--	g26927 = OR(g26711, g18539)
--	g30506 = OR(g30179, g22027)
--	g28066 = OR(g27553, g21819)
--	g21895 = OR(g20135, g15108)
--	g34028 = OR(g33720, g18684)
--	g32368 = OR(g29881, g31310)
--	g33982 = OR(g33865, g18372)
--	g25682 = OR(g24658, g18640)
--	g29274 = OR(g28360, g18642)
--	g24561 = OR(I23755, I23756)
--	g24353 = OR(g23682, g18822)
--	g26903 = OR(g26388, g24220)
--	g35000 = OR(g34953, g34999)
--	g11737 = OR(g8359, g8292)
--	g9012 = OR(g2047, g2066)
--	g26755 = OR(g10776, g24457)
--	g28511 = OR(g27272, g16208)
--	g32229 = OR(g31148, g29652)
--	g26770 = OR(g24471, g10732)
--	g24336 = OR(g24012, g18753)
--	g27837 = OR(g17401, g26725)
--	g33390 = OR(g32276, g29968)
--	g32228 = OR(g31147, g29651)
--	g25760 = OR(g25238, g22109)
--	g29292 = OR(g28556, g18776)
--	g34649 = OR(g33111, g34492)
--	g34240 = OR(g32910, g33958)
--	g30491 = OR(g30178, g21987)
--	g34903 = OR(g34859, g21690)
--	g23297 = OR(g19692, g16178)
--	g34604 = OR(g34563, g15076)
--	g26899 = OR(g26844, g18199)
--	g30563 = OR(g29347, g22134)
--	g26898 = OR(g26387, g18194)
--	g28085 = OR(g27263, g18700)
--	g28076 = OR(g27098, g21878)
--	g28721 = OR(g27488, g16705)
--	g28596 = OR(g27336, g26291)
--	g28054 = OR(g27723, g18170)
--	g33553 = OR(g33403, g18350)
--	g15803 = OR(g12924, g10528)
--	g22217 = OR(g21302, g17617)
--	g33949 = OR(g32446, g33459)
--	g31326 = OR(g29627, g29640)
--	g32386 = OR(g31488, g29949)
--	g30395 = OR(g29841, g21754)
--	g34794 = OR(g34746, g18571)
--	g25649 = OR(g24654, g21742)
--	I26644 = OR(g27057, g27044, g27039, g27032)
--	g27037 = OR(g26236, g26218, g26195, g26171)
--	g34262 = OR(g34075, g18697)
--	g33536 = OR(g33241, g21715)
--	g33040 = OR(g32164, g24313)
--	g33948 = OR(g32442, g33458)
--	g25648 = OR(g24644, g21741)
--	g28773 = OR(g27535, g16803)
--	g31757 = OR(g29992, g30010)
--	g31904 = OR(g31780, g21923)
--	g34633 = OR(g34481, g18690)
--	g25604 = OR(g24717, g18115)
--	g25755 = OR(g25192, g22102)
--	g33621 = OR(g33365, g18775)
--	g34719 = OR(g34701, g18133)
--	g28180 = OR(g20242, g27511)
--	g28670 = OR(g27412, g16618)
--	g26926 = OR(g26633, g18531)
--	g32429 = OR(g30318, g31794)
--	g30521 = OR(g29331, g22042)
--	g14511 = OR(g10685, g546)
--	g33564 = OR(g33332, g18388)
--	g26099 = OR(g24506, g22538)
--	g29283 = OR(g28627, g18746)
--	g28734 = OR(g27508, g16736)
--	g28335 = OR(g27132, g15818)
--	g29303 = OR(g28703, g18801)
--	g24374 = OR(g19345, g24004)
--	g30440 = OR(g29771, g21849)
--	g34440 = OR(g34364, g24226)
--	g25767 = OR(g25207, g12015)
--	g28667 = OR(g27410, g16616)
--	g33062 = OR(g31977, g22065)
--	g22531 = OR(g20773, g20922)
--	g27589 = OR(g26177, g24763)
--	g16448 = OR(g13287, g10934)
--	g30389 = OR(g29969, g18554)
--	g24260 = OR(g23373, g18313)
--	g27524 = OR(g26050, g24649)
--	g25633 = OR(g24420, g18282)
--	g31872 = OR(g31524, g18535)
--	g24842 = OR(g7804, g22669)
--	g30388 = OR(g30023, g18534)
--	g34612 = OR(g34514, g18566)
--	g25719 = OR(g25089, g18761)
--	g28619 = OR(g27358, g16517)
--	g34099 = OR(g33684, g33689)
--	g30534 = OR(g30213, g22080)
--	g19441 = OR(g15507, g12931)
--	g25718 = OR(g25187, g21971)
--	g28618 = OR(g27357, g16516)
--	g34251 = OR(g34157, g18147)
--	g28279 = OR(g27087, g25909)
--	g26766 = OR(g10776, g24460)
--	g30462 = OR(g30228, g21933)
--	g23296 = OR(g19691, g16177)
--	g34462 = OR(g34334, g18685)
--	g28286 = OR(g27090, g15757)
--	g32245 = OR(g31167, g29684)
--	g34032 = OR(g33816, g18706)
--	g28306 = OR(g27104, g15794)
--	g33574 = OR(g33362, g18416)
--	g33047 = OR(g31944, g21927)
--	I26741 = OR(g22881, g22905, g22928, g27402)
--	g31912 = OR(g31752, g21998)
--	g31311 = OR(g26103, g29618)
--	g23197 = OR(g19571, g15966)
--	g25612 = OR(g24941, g18132)
--	g28815 = OR(g27546, g16842)
--	g29483 = OR(g25801, g28130)
--	g16811 = OR(g8690, g13914)
--	g25701 = OR(g25054, g21920)
--	I30055 = OR(g31070, g31170, g30614, g30673)
--	g24705 = OR(g2890, g23267)
--	g33051 = OR(g32316, g21958)
--	g24255 = OR(g22835, g18308)
--	g33592 = OR(g33412, g18475)
--	g30360 = OR(g30145, g18386)
--	g24270 = OR(g23165, g18614)
--	g26911 = OR(g26612, g24230)
--	I30741 = OR(g32085, g32030, g32224, g32013)
--	g30447 = OR(g29798, g21856)
--	g21894 = OR(g20112, g15107)
--	g34447 = OR(g34363, g18552)
--	g32995 = OR(g32330, g18375)
--	g24460 = OR(g10967, g22450)
--	g29904 = OR(g28312, g26146)
--	g13657 = OR(g7251, g10616)
--	g29252 = OR(g28712, g18486)
--	g28884 = OR(g27568, g16885)
--	g26785 = OR(g10776, g24468)
--	g24267 = OR(g23439, g18611)
--	g30451 = OR(g29877, g21860)
--	g30472 = OR(g30186, g21943)
--	I30735 = OR(g32369, g32376, g32089, g32035)
--	g34629 = OR(g34495, g18654)
--	g17569 = OR(g14416, g14394, g11995, I18492)
--	g34451 = OR(g34393, g18664)
--	g34628 = OR(g34493, g18653)
--	g34911 = OR(g34909, g18188)
--	g26950 = OR(g26357, g24288)
--	g22751 = OR(g19333, g15716)
--	g27008 = OR(g26866, g21370, I25736)
--	g22639 = OR(g18950, g15612)
--	g27555 = OR(g26095, g24686)
--	g28580 = OR(g27328, g26275)
--	g29508 = OR(g28152, g27041)
--	g8476 = OR(g1399, g1459, I12611)
--	g20160 = OR(g16163, g13415)
--	g30355 = OR(g30131, g18360)
--	g27570 = OR(g26126, g24722)
--	g31929 = OR(g31540, g22093)
--	g32989 = OR(g32241, g18326)
--	g30370 = OR(g30135, g18440)
--	g25629 = OR(g24962, g18258)
--	g27907 = OR(g17424, g26770)
--	g16959 = OR(g13542, g11142)
--	g31020 = OR(g29375, g28164)
--	g31928 = OR(g31517, g22092)
--	g14187 = OR(g8871, g11771)
--	g32988 = OR(g32232, g18325)
--	g28084 = OR(g27254, g18698)
--	g33020 = OR(g32160, g21734)
--	g33583 = OR(g33074, g18448)
--	g25628 = OR(g24600, g18249)
--	g25911 = OR(g22514, g24510)
--	g27239 = OR(g25881, g24465)
--	g19605 = OR(g15707, g13063)
--	g33046 = OR(g32308, g21912)
--	g32271 = OR(g31209, g29731)
--	g34172 = OR(g33795, g19914)
--	g28179 = OR(g27494, g27474, g27445, g27421)
--	g27567 = OR(g26121, g24714)
--	g27238 = OR(g25879, g24464)
--	g17510 = OR(g14393, g14362, g11972, I18449)
--	g30394 = OR(g29805, g21753)
--	g30367 = OR(g30133, g18418)
--	g24201 = OR(g22848, g18104)
--	g24277 = OR(g23188, g18647)
--	g25591 = OR(g24642, g21705)
--	g33282 = OR(g32143, g29577)
--	g28186 = OR(g27209, g27185, g27161, g27146)
--	g28685 = OR(g27433, g16637)
--	g31302 = OR(g29590, g28302)
--	g28373 = OR(g27180, g15849)
--	g25754 = OR(g25179, g22101)
--	g30420 = OR(g29769, g21804)
--	g28417 = OR(g27219, g15881)
--	g24782 = OR(g23857, g23872)
--	g30446 = OR(g29788, g21855)
--	g34446 = OR(g34390, g18550)
--	g34318 = OR(g25850, g34063)
--	g28334 = OR(g27131, g15817)
--	g29756 = OR(g22717, g28223)
--	g24352 = OR(g22157, g18821)
--	g26902 = OR(g26378, g24219)
--	g26957 = OR(g26517, g24295)
--	g34025 = OR(g33927, g18672)
--	g31768 = OR(g30033, g30045)
--	g26377 = OR(g24700, g23007)
--	g30540 = OR(g30275, g22086)
--	g13295 = OR(g10625, g10655)
--	g15582 = OR(g8977, g12925)
--	g24266 = OR(g22329, g18561)
--	g32132 = OR(g31487, g31479)
--	g9535 = OR(g209, g538)
--	g31881 = OR(g31018, g21775)
--	g28216 = OR(g27036, g27043)
--	g24853 = OR(g21452, g24001)
--	g22684 = OR(g19206, g15703)
--	g32259 = OR(g31185, g29709)
--	g30377 = OR(g30124, g18472)
--	g32225 = OR(g30576, g29336)
--	g34957 = OR(g34948, g21662)
--	g34377 = OR(g26304, g34141)
--	g33027 = OR(g32314, g21796)
--	I22912 = OR(g21555, g21364, g21357)
--	g31890 = OR(g31143, g21823)
--	g24401 = OR(g23811, g21298)
--	g30562 = OR(g30289, g22133)
--	g31249 = OR(g25971, g29523)
--	g19359 = OR(g17786, g14875)
--	g34645 = OR(g34556, g18786)
--	g19535 = OR(g15651, g13020)
--	g31248 = OR(g25970, g29522)
--	g28747 = OR(g27521, g13942)
--	g34290 = OR(g26848, g34219)
--	g33552 = OR(g33400, g18343)
--	g13289 = OR(g10619, g10624)
--	g33003 = OR(g32323, g18429)
--	g33204 = OR(g32317, I30750, I30751)
--	g26895 = OR(g26783, g18148)
--	g31779 = OR(g30050, g28673)
--	I31843 = OR(g33470, g33471, g33472, g33473)
--	g10800 = OR(g7517, g952)
--	g19344 = OR(g17771, g14832)
--	g27566 = OR(g26119, g24713)
--	g28814 = OR(g27545, g16841)
--	g30427 = OR(g29796, g21811)
--	g20276 = OR(g16243, g13566)
--	g29583 = OR(g28182, g27099)
--	g32375 = OR(g29896, g31324)
--	g14936 = OR(g10776, g8703)
--	g30366 = OR(g30122, g18417)
--	I30054 = OR(g29385, g31376, g30735, g30825)
--	g24276 = OR(g23083, g18646)
--	g28751 = OR(g27526, g16766)
--	g28772 = OR(g27534, g16802)
--	g34366 = OR(g26257, g34133)
--	I31869 = OR(g33519, g33520, g33521, g33522)
--	g34632 = OR(g34565, g15119)
--	g25739 = OR(g25149, g22054)
--	g24254 = OR(g23265, g18306)
--	I31868 = OR(g33515, g33516, g33517, g33518)
--	g28230 = OR(g27669, g14261)
--	g33945 = OR(g32430, g33455)
--	g25738 = OR(g25059, g22053)
--	g25645 = OR(g24679, g21738)
--	g30547 = OR(g30194, g22118)
--	g30403 = OR(g29750, g21762)
--	g33999 = OR(g33893, g18436)
--	g33380 = OR(g32234, g29926)
--	g25699 = OR(g25125, g21918)
--	g34403 = OR(g34180, g25085)
--	g29282 = OR(g28617, g18745)
--	g28416 = OR(g27218, g15880)
--	g16261 = OR(g7898, g13469)
--	g32994 = OR(g32290, g18367)
--	g33998 = OR(g33878, g18428)
--	g29302 = OR(g28601, g18798)
--	g25698 = OR(g25104, g21917)
--	g29105 = OR(g27645, g17134)
--	g30481 = OR(g30221, g21977)
--	g7932 = OR(g4072, g4153)
--	g26956 = OR(g26487, g24294)
--	g30551 = OR(g30235, g22122)
--	I30734 = OR(g31790, g32191, g32086, g32095)
--	g26889 = OR(g26689, g24195)
--	g31932 = OR(g31792, g22107)
--	g26888 = OR(g26671, g24194)
--	g23721 = OR(g21401, g21385, I22852)
--	g25632 = OR(g24558, g18277)
--	g28578 = OR(g27327, g26273)
--	g30127 = OR(g28494, g16805)
--	g29768 = OR(g22760, g28229)
--	g34127 = OR(g33657, g32438)
--	g31897 = OR(g31237, g24322)
--	g30490 = OR(g30167, g21986)
--	g33961 = OR(g33789, g21712)
--	g25661 = OR(g24754, g21786)
--	g27484 = OR(g25988, g24628)
--	g30376 = OR(g30112, g18471)
--	g30385 = OR(g30172, g18518)
--	g26931 = OR(g26778, g18547)
--	g30103 = OR(g28477, g16731)
--	g34376 = OR(g26301, g34140)
--	g34297 = OR(g26858, g34228)
--	g34103 = OR(g33701, g33707)
--	g33026 = OR(g32307, g21795)
--	g30354 = OR(g30064, g18359)
--	g22516 = OR(g21559, g12817)
--	g34980 = OR(g34969, g18587)
--	g33212 = OR(g32328, I30755, I30756)
--	g25715 = OR(g25071, g21966)
--	g8679 = OR(g222, g199)
--	g34095 = OR(g33681, g33687)
--	g30824 = OR(g13833, g29789)
--	g28720 = OR(g27486, g16704)
--	g28041 = OR(g24145, g26878)
--	g17264 = OR(g7118, g14309)
--	g28430 = OR(g27229, g15914)
--	g32125 = OR(g30918, g29376)
--	g28746 = OR(g27520, g16762)
--	g32977 = OR(g32169, g21710)
--	g19604 = OR(g15704, g13059)
--	I30469 = OR(g31672, g31710, g31021, g30937)
--	g29249 = OR(g28658, g18438)
--	g26089 = OR(g24501, g22534)
--	g24907 = OR(g21558, g24015)
--	I30468 = OR(g29385, g31376, g30735, g30825)
--	g29482 = OR(g28524, g27588)
--	g34931 = OR(g2984, g34912)
--	g29248 = OR(g28677, g18434)
--	g33149 = OR(g32204, I30717, I30718)
--	g30426 = OR(g29785, g21810)
--	g32353 = OR(g29853, g31283)
--	g33387 = OR(g32263, g29954)
--	g24239 = OR(g22752, g18250)
--	g9055 = OR(g2606, g2625)
--	g28684 = OR(g27432, g16636)
--	g32144 = OR(g30927, g30930)
--	g33620 = OR(g33360, g18774)
--	g34190 = OR(g33802, g33810)
--	g24238 = OR(g23254, g18248)
--	g30520 = OR(g30272, g22041)
--	g28517 = OR(g27280, g26154)
--	g30546 = OR(g30277, g22117)
--	g33971 = OR(g33890, g18330)
--	g29786 = OR(g22843, g28240)
--	g25671 = OR(g24637, g21828)
--	g34024 = OR(g33807, g24331)
--	g13938 = OR(g11213, g11191)
--	g24518 = OR(g22517, g7601)
--	g22530 = OR(g16751, g20171)
--	g28362 = OR(g27154, g15840)
--	g30497 = OR(g30242, g21993)
--	g24935 = OR(g22937, g19749)
--	I12903 = OR(g4222, g4219, g4216, g4213)
--	g29233 = OR(g28171, g18234)
--	g26969 = OR(g26313, g24329)
--	I18421 = OR(g14447, g14417, g14395)
--	g32289 = OR(g24796, g31230)
--	g22641 = OR(g18974, g15631)
--	g34625 = OR(g34532, g18610)
--	g26968 = OR(g26307, g24321)
--	g17464 = OR(g14334, g14313, g11935, I18385)
--	g31896 = OR(g31242, g24305)
--	g34250 = OR(g34111, g21713)
--	g32288 = OR(g31226, g31229)
--	g28727 = OR(g27500, g16729)
--	g16258 = OR(g13247, g10856)
--	g33011 = OR(g32338, g18481)
--	g30339 = OR(g29629, g18244)
--	g24215 = OR(g23484, g18196)
--	g24577 = OR(g2856, g22531)
--	g30338 = OR(g29613, g18240)
--	g34644 = OR(g34555, g18769)
--	g33582 = OR(g33351, g18444)
--	g19534 = OR(g15650, g13019)
--	g27241 = OR(g24584, g25984)
--	g28347 = OR(g27138, g15822)
--	g29717 = OR(g28200, g10883)
--	g33310 = OR(g29631, g32165)
--	g26894 = OR(g25979, g18129)
--	g33627 = OR(g33376, g18826)
--	g31925 = OR(g31789, g22061)
--	g32976 = OR(g32207, g21704)
--	g32985 = OR(g31963, g18266)
--	g24349 = OR(g23646, g18805)
--	g16810 = OR(g13461, g11032)
--	g25700 = OR(g25040, g21919)
--	g28600 = OR(g27339, g16427)
--	g25659 = OR(g24707, g21784)
--	g25625 = OR(g24553, g18226)
--	g20083 = OR(g2902, g17058)
--	g30527 = OR(g30192, g22073)
--	g30411 = OR(g29872, g21770)
--	g33050 = OR(g31974, g21930)
--	g32374 = OR(g29895, g31323)
--	g33958 = OR(g33532, I31873, I31874)
--	g24348 = OR(g22149, g18804)
--	g34411 = OR(g34186, g25142)
--	g16970 = OR(g13567, g11163)
--	g25658 = OR(g24635, g21783)
--	g28372 = OR(g27178, g15848)
--	g23217 = OR(g19588, g16023)
--	g33386 = OR(g32258, g29951)
--	g26910 = OR(g26571, g24228)
--	g33603 = OR(g33372, g18515)
--	g25943 = OR(g24423, g22299)
--	I30740 = OR(g31776, g32188, g32083, g32087)
--	g13623 = OR(g482, g12527)
--	g25644 = OR(g24622, g21737)
--	g30503 = OR(g30243, g22024)
--	g28063 = OR(g27541, g21773)
--	g34894 = OR(g34862, g21678)
--	g29148 = OR(g27651, g26606)
--	g32392 = OR(g31513, g30000)
--	g27515 = OR(g26051, g13431)
--	g30450 = OR(g29861, g21859)
--	g24653 = OR(g2848, g22585)
--	g34450 = OR(g34281, g18663)
--	g13155 = OR(g11496, g11546)
--	g31793 = OR(g28031, g30317)
--	g34819 = OR(g34741, g34684)
--	g34257 = OR(g34226, g18674)
--	g28209 = OR(g27223, g27141)
--	g30496 = OR(g30231, g21992)
--	g8956 = OR(g1913, g1932)
--	g34979 = OR(g34875, g34968)
--	g34055 = OR(g33909, g33910)
--	g33549 = OR(g33328, g18337)
--	g28208 = OR(g27025, g27028)
--	g26877 = OR(g21658, g25577)
--	g34978 = OR(g34874, g34967)
--	g33548 = OR(g33327, g18336)
--	g27584 = OR(g26165, g24758)
--	g25867 = OR(g25449, g23884)
--	g25894 = OR(g24817, g23229)
--	g30384 = OR(g30101, g18517)
--	g31317 = OR(g29611, g29626)
--	g33317 = OR(g29688, g32179)
--	g29229 = OR(g28532, g18191)
--	g25714 = OR(g25056, g21965)
--	g28614 = OR(g27351, g26311)
--	g25707 = OR(g25041, g18749)
--	g25819 = OR(g25323, g23836)
--	g28607 = OR(g27342, g26303)
--	g29228 = OR(g28426, g18173)
--	g25910 = OR(g25565, g22142)
--	g28320 = OR(g27116, g15808)
--	g31002 = OR(g29362, g28154)
--	g28073 = OR(g27097, g21875)
--	g33002 = OR(g32304, g18419)
--	g33057 = OR(g31968, g22019)
--	g34801 = OR(g34756, g18588)
--	g34735 = OR(g34709, g15116)
--	g32124 = OR(g24488, g30920)
--	g29716 = OR(g28199, g15856)
--	g24200 = OR(g22831, g18103)
--	g31245 = OR(g25964, g29516)
--	g34019 = OR(g33889, g18506)
--	g26917 = OR(g26122, g18233)
--	g15792 = OR(g12920, g10501)
--	g26866 = OR(g20204, g20242, g24363)
--	g28565 = OR(g27315, g26253)
--	g33626 = OR(g33374, g18825)
--	g33323 = OR(g31936, g32442)
--	g34695 = OR(g34523, g34322)
--	g25590 = OR(g21694, g24160)
--	g34018 = OR(g33887, g18505)
--	g30526 = OR(g30181, g22072)
--	g32267 = OR(g31208, g31218)
--	g32294 = OR(g31231, g31232)
--	g33298 = OR(g32158, g29622)
--	g25741 = OR(g25178, g22056)
--	g28641 = OR(g27385, g16591)
--	g31775 = OR(g30048, g30059)
--	I30123 = OR(g29385, g31376, g30735, g30825)
--	g8957 = OR(g2338, g2357)
--	g24799 = OR(g23901, g23921)
--	g30402 = OR(g29871, g21761)
--	g24813 = OR(g22685, g19594)
--	I30751 = OR(g32042, g32161, g31943, g31959)
--	g30457 = OR(g29369, g21885)
--	g34402 = OR(g34179, g25084)
--	g34457 = OR(g34394, g18670)
--	g26923 = OR(g25923, g18290)
--	g32219 = OR(g31131, g29620)
--	g33232 = OR(g32034, g30936)
--	g25735 = OR(g25077, g18783)
--	g25877 = OR(g25502, g23919)
--	g28635 = OR(g27375, g16537)
--	g32218 = OR(g31130, g29619)
--	g27135 = OR(g24387, g25803)
--	g33995 = OR(g33848, g18425)
--	g34001 = OR(g33844, g18450)
--	g33261 = OR(g32111, g29525)
--	g25695 = OR(g24998, g21914)
--	g31880 = OR(g31280, g21774)
--	g30597 = OR(g13564, g29693)
--	g34256 = OR(g34173, g24303)
--	g29802 = OR(g28243, g22871)
--	g34280 = OR(g26833, g34213)
--	g29730 = OR(g28150, g28141)
--	g30300 = OR(g28246, g27252)
--	g29793 = OR(g28237, g27247)
--	g34624 = OR(g34509, g18592)
--	g34300 = OR(g26864, g34230)
--	g15125 = OR(g10363, g13605)
--	g26876 = OR(g21655, g25576)
--	g26885 = OR(g26541, g24191)
--	g23751 = OR(g21415, g21402, I22880)
--	g25917 = OR(g22524, g24518)
--	g32277 = OR(g31211, g29733)
--	g24214 = OR(g23471, g18195)
--	g31316 = OR(g29609, g29624)
--	g33316 = OR(g29685, g32178)
--	g22634 = OR(g18934, g15590)
--	g24207 = OR(g23396, g18119)
--	g22872 = OR(g19372, g19383)
--	I29985 = OR(g29385, g31376, g30735, g30825)
--	I22958 = OR(g21603, g21386, g21365)
--	g34231 = OR(g33898, g33902)
--	g29504 = OR(g28143, g25875)
--	g25706 = OR(g25030, g18748)
--	g25597 = OR(g24892, g21719)
--	g32037 = OR(g30566, g29329)
--	g33989 = OR(g33870, g18398)
--	g33056 = OR(g32327, g22004)
--	g13570 = OR(g9223, g11130)
--	g25689 = OR(g24849, g21888)
--	g13914 = OR(g8643, g11380)
--	g33611 = OR(g33243, g18632)
--	g31924 = OR(g31486, g22049)
--	g32984 = OR(g31934, g18264)
--	g33988 = OR(g33861, g18397)
--	g25688 = OR(g24812, g21887)
--	g28750 = OR(g27525, g16765)
--	g25624 = OR(g24408, g18224)
--	g26916 = OR(g25916, g18232)
--	g30511 = OR(g30180, g22032)
--	g20241 = OR(g16233, g13541)
--	g32352 = OR(g29852, g31282)
--	I30746 = OR(g32047, g31985, g31991, g32309)
--	g24241 = OR(g22920, g18252)
--	g33271 = OR(g32120, g29549)
--	g27972 = OR(g26131, g26105)
--	g32155 = OR(g30935, g29475)
--	g15017 = OR(g10776, g8703)
--	g28091 = OR(g27665, g21913)
--	g32266 = OR(g30604, g29354)
--	g29245 = OR(g28676, g18384)
--	g26721 = OR(g10776, g24444)
--	g29299 = OR(g28587, g18794)
--	g33031 = OR(g32315, g21841)
--	g30456 = OR(g29378, g21869)
--	g34456 = OR(g34395, g18669)
--	g29298 = OR(g28571, g18793)
--	g24235 = OR(g22632, g18238)
--	g13941 = OR(g11019, g11023)
--	g31887 = OR(g31292, g21820)
--	g28390 = OR(g27207, g15861)
--	g30480 = OR(g29321, g21972)
--	g30916 = OR(g13853, g29799)
--	g29775 = OR(g25966, g28232)
--	I26523 = OR(g20720, g20857, g20998, g21143)
--	g25885 = OR(g25522, g23957)
--	g30550 = OR(g30226, g22121)
--	g30314 = OR(g28268, g27266)
--	g23615 = OR(g20109, g20131)
--	g30287 = OR(g28653, g27677)
--	g34314 = OR(g25831, g34061)
--	g30307 = OR(g28256, g27260)
--	g33393 = OR(g32286, g29984)
--	g23720 = OR(g20165, g16801)
--	I12902 = OR(g4235, g4232, g4229, g4226)
--	g25763 = OR(g25113, g18817)
--	g29232 = OR(g28183, g18231)
--	g31764 = OR(g30015, g30032)
--	g23275 = OR(g19680, g16160)
--	g34721 = OR(g34696, g18135)
--	g31869 = OR(g30592, g18221)
--	I30193 = OR(g31070, g30614, g30673, g31528)
--	g30431 = OR(g29875, g21815)
--	g33960 = OR(g33759, g21701)
--	g25660 = OR(g24726, g21785)
--	g29261 = OR(g28247, g18605)
--	g31868 = OR(g30600, g18204)
--	g26335 = OR(g1526, g24609)
--	g19572 = OR(g17133, g14193)
--	g22152 = OR(g21188, g17469)
--	g26930 = OR(g26799, g18544)
--	g34269 = OR(g34083, g18732)
--	g30341 = OR(g29380, g18246)
--	g26694 = OR(g24444, g10704)
--	g26965 = OR(g26336, g24317)
--	g33709 = OR(g32414, g33441)
--	g34268 = OR(g34082, g18730)
--	g31259 = OR(g25992, g29554)
--	g32285 = OR(g31222, g29740)
--	g33259 = OR(g32109, g29521)
--	g28536 = OR(g27293, g26205)
--	I30727 = OR(g31759, g32196, g31933, g31941)
--	g31258 = OR(g25991, g29550)
--	g24206 = OR(g23386, g18110)
--	g13728 = OR(g6804, g12527)
--	g28702 = OR(g27457, g16670)
--	g30734 = OR(g13808, g29774)
--	I22298 = OR(g20371, g20161, g20151)
--	g30335 = OR(g29746, g18174)
--	g34734 = OR(g34681, g18652)
--	g25721 = OR(g25057, g18766)
--	g28621 = OR(g27359, g16518)
--	g25596 = OR(g24865, g21718)
--	I31853 = OR(g33488, g33489, g33490, g33491)
--	g33043 = OR(g32195, g24325)
--	g31244 = OR(g25963, g29515)
--	g20082 = OR(g16026, g13321)
--	g28564 = OR(g27314, g26252)
--	g23193 = OR(g19556, g15937)
--	I23756 = OR(g23457, g23480, g23494, g23511)
--	g26278 = OR(g24545, g24549)
--	g33069 = OR(g32009, g22113)
--	g33602 = OR(g33425, g18511)
--	g25942 = OR(g24422, g22298)
--	g31774 = OR(g30046, g30057)
--	g7834 = OR(g2886, g2946)
--	g30487 = OR(g30187, g21983)
--	g31375 = OR(g29628, g28339)
--	g33068 = OR(g31994, g22112)
--	g33955 = OR(g33505, I31858, I31859)
--	g24345 = OR(g23606, g18788)
--	g25655 = OR(g24645, g18607)
--	g31879 = OR(g31475, g21745)
--	g30502 = OR(g30232, g22023)
--	g28062 = OR(g27288, g21746)
--	g30557 = OR(g30247, g22128)
--	g33970 = OR(g33868, g18322)
--	g34619 = OR(g34528, g18581)
--	I22880 = OR(g21509, g21356, g21351)
--	g25670 = OR(g24967, g18626)
--	g29271 = OR(g28333, g18637)
--	g31878 = OR(g31015, g21733)
--	I31864 = OR(g33510, g33511, g33512, g33513)
--	g30443 = OR(g29808, g21852)
--	g34618 = OR(g34527, g18580)
--	g24398 = OR(g23801, g21296)
--	g30279 = OR(g28637, g27668)
--	g34443 = OR(g34385, g18545)
--	g25734 = OR(g25058, g18782)
--	g28634 = OR(g27374, g16536)
--	g28851 = OR(g27558, g16870)
--	g31886 = OR(g31481, g21791)
--	g29753 = OR(g28213, g22720)
--	g25839 = OR(g25507, g25485, g25459, g25420)
--	g34278 = OR(g26829, g34212)
--	g30469 = OR(g30153, g21940)
--	g33967 = OR(g33842, g18319)
--	g33994 = OR(g33841, g18424)
--	g27506 = OR(g26021, g24639)
--	g30286 = OR(g28191, g28186)
--	g25694 = OR(g24638, g18738)
--	g25667 = OR(g24682, g18619)
--	g24263 = OR(g23497, g18529)
--	g34286 = OR(g26842, g34216)
--	g30468 = OR(g30238, g21939)
--	g34468 = OR(g34342, g18718)
--	g34039 = OR(g33743, g18736)
--	g34306 = OR(g25782, g34054)
--	g29529 = OR(g28303, g28293, g28283, g28267)
--	g22640 = OR(g18951, g15613)
--	g34038 = OR(g33731, g18735)
--	g31919 = OR(g31758, g22044)
--	g32454 = OR(g30322, g31795)
--	g25619 = OR(g24961, g18193)
--	g15124 = OR(g13605, g4581)
--	g26884 = OR(g26511, g24190)
--	g28574 = OR(g27324, g26270)
--	g31918 = OR(g31786, g22015)
--	g28047 = OR(g27676, g18160)
--	g33010 = OR(g32301, g18473)
--	g34601 = OR(g34488, g18211)
--	g29764 = OR(g28219, g28226)
--	g25618 = OR(g25491, g18192)
--	g34975 = OR(g34871, g34964)
--	g24500 = OR(g24011, g21605)
--	g33545 = OR(g33399, g18324)
--	g9013 = OR(g2472, g2491)
--	g26363 = OR(g2965, g24965)
--	g33599 = OR(g33087, g18500)
--	g32239 = OR(g30595, g29350)
--	g28051 = OR(g27699, g18166)
--	g27240 = OR(g25883, g24467)
--	g28072 = OR(g27086, g21874)
--	g33598 = OR(g33364, g18496)
--	g32238 = OR(g30594, g29349)
--	I29352 = OR(g29322, g29315, g30315, g30308)
--	g28592 = OR(g27333, g26288)
--	I31874 = OR(g33528, g33529, g33530, g33531)
--	g34791 = OR(g34771, g18184)
--	g22662 = OR(g19069, g15679)
--	g34884 = OR(g34858, g21666)
--	g29259 = OR(g28304, g18603)
--	g29225 = OR(g28451, g18158)
--	g30410 = OR(g29857, g21769)
--	g31322 = OR(g26128, g29635)
--	g14062 = OR(g11047, g11116)
--	g34168 = OR(g33787, g19784)
--	g27563 = OR(g26104, g24704)
--	g29258 = OR(g28238, g18601)
--	g31901 = OR(g31516, g21909)
--	g33159 = OR(g32016, g30730)
--	g30479 = OR(g29320, g21950)
--	g33977 = OR(g33876, g18348)
--	g30363 = OR(g30121, g18407)
--	g25601 = OR(g24660, g18112)
--	g12981 = OR(g12219, g9967)
--	g24273 = OR(g23166, g18630)
--	g25677 = OR(g24684, g21834)
--	g31783 = OR(I29351, I29352)
--	g23209 = OR(g19585, g19601)
--	g30478 = OR(g30248, g21949)
--	g34015 = OR(g33858, g18502)
--	g29244 = OR(g28692, g18380)
--	g33561 = OR(g33408, g18376)
--	g30486 = OR(g30177, g21982)
--	g31295 = OR(g26090, g29598)
--	g26922 = OR(g25902, g18288)
--	g28731 = OR(g27504, g16733)
--	g33295 = OR(g32153, g29605)
--	g31144 = OR(g29477, g28193)
--	g25937 = OR(g24406, g22216)
--	g30556 = OR(g30236, g22127)
--	g24234 = OR(g22622, g18237)
--	g13973 = OR(g11024, g11028)
--	g29068 = OR(g27628, g17119)
--	g25791 = OR(g25411, g25371, g25328, g25290)
--	g28691 = OR(g27437, g16642)
--	g29879 = OR(g28289, g26096)
--	g26953 = OR(g26486, g24291)
--	g28405 = OR(g27216, g15875)
--	g33966 = OR(g33837, g18318)
--	g25666 = OR(g24788, g21793)
--	g33017 = OR(g32292, g18510)
--	g26800 = OR(g24922, g24929)
--	g34321 = OR(g25866, g34065)
--	g30531 = OR(g30274, g22077)
--	g23346 = OR(g19736, g16204)
--	g29792 = OR(g28235, g28244)
--	g12832 = OR(g10347, g10348)
--	g13761 = OR(g490, g12527)
--	g16022 = OR(g13048, g10707)
--	g26334 = OR(g1171, g24591)
--	g28046 = OR(g27667, g18157)
--	g32349 = OR(g29840, g31275)
--	g31289 = OR(g29580, g29591)
--	g30373 = OR(g30111, g18461)
--	g33289 = OR(g32148, g29588)
--	g22331 = OR(g21405, g17809)
--	g26964 = OR(g26259, g24316)
--	g34373 = OR(g26292, g34138)
--	g33023 = OR(g32313, g21751)
--	g31288 = OR(g2955, g29914)
--	g23153 = OR(g19521, g15876)
--	g33288 = OR(g32147, g29587)
--	g31308 = OR(g26101, g29614)
--	g33571 = OR(g33367, g18409)
--	g30417 = OR(g29874, g21801)
--	g34800 = OR(g34752, g18586)
--	g34417 = OR(g27678, g34196)
--	g28357 = OR(g27148, g15836)
--	g30334 = OR(g29837, g18143)
--	g28105 = OR(g27997, g22135)
--	g28743 = OR(g27517, g16758)
--	g29078 = OR(g27633, g26572)
--	g26909 = OR(g26543, g24227)
--	I18385 = OR(g14413, g14391, g14360)
--	g34762 = OR(g34687, g34524)
--	g25740 = OR(g25164, g22055)
--	g26908 = OR(g26358, g24225)
--	g28640 = OR(g27384, g16590)
--	g30423 = OR(g29887, g21807)
--	g33976 = OR(g33869, g18347)
--	g33985 = OR(g33896, g18382)
--	g24946 = OR(g22360, g22409, g8130)
--	g25676 = OR(g24668, g21833)
--	g25685 = OR(g24476, g21866)
--	I30750 = OR(g31788, g32310, g32054, g32070)
--	g33954 = OR(g33496, I31853, I31854)
--	g21891 = OR(g19948, g15103)
--	g24344 = OR(g22145, g18787)
--	g25654 = OR(g24634, g18606)
--	g25936 = OR(g24403, g22209)
--	g30543 = OR(g29338, g22110)
--	I26522 = OR(g19890, g19935, g19984, g26365)
--	g31260 = OR(g25993, g29555)
--	g34000 = OR(g33943, g18441)
--	g26751 = OR(g24903, g24912)
--	g33260 = OR(g32110, g29524)
--	g29295 = OR(g28663, g18780)
--	g31668 = OR(g29924, g28558)
--	g14583 = OR(g10685, g542)
--	g25762 = OR(g25095, g18816)
--	g28662 = OR(g27407, g16612)
--	g26293 = OR(g24550, g24555)
--	g33559 = OR(g33073, g18368)
--	I30192 = OR(g29385, g31376, g30735, g30825)
--	g33016 = OR(g32284, g18509)
--	g25587 = OR(g21682, g24157)
--	g33558 = OR(g33350, g18364)
--	g23750 = OR(g20174, g16840)
--	g31893 = OR(g31490, g21837)
--	g34807 = OR(g34764, g18596)
--	g34974 = OR(g34870, g34963)
--	g31865 = OR(g31149, g21709)
--	g33544 = OR(g33392, g18317)
--	g34639 = OR(g34486, g18722)
--	g12911 = OR(g10278, g12768)
--	g30293 = OR(g28236, g27246)
--	g23796 = OR(g21462, g21433, I22958)
--	g28778 = OR(g27540, g16808)
--	g16239 = OR(g7892, g13432)
--	g34293 = OR(g26854, g34224)
--	g34638 = OR(g34484, g18721)
--	g34265 = OR(g34117, g18711)
--	g30416 = OR(g29858, g21800)
--	g27591 = OR(g26181, g24765)
--	g34416 = OR(g34191, g25159)
--	g29289 = OR(g28642, g18763)
--	g25747 = OR(g25130, g18795)
--	g28647 = OR(g27389, g16596)
--	g33610 = OR(g33242, g18616)
--	g29309 = OR(g28722, g18818)
--	g30391 = OR(g30080, g18557)
--	g33042 = OR(g32193, g24324)
--	g27147 = OR(g25802, g24399)
--	g31255 = OR(g25982, g29536)
--	g29288 = OR(g28630, g18762)
--	g33255 = OR(g32106, g29514)
--	g29224 = OR(g28919, g18156)
--	g30510 = OR(g30263, g22031)
--	g29308 = OR(g28612, g18815)
--	g24240 = OR(g22861, g18251)
--	g33270 = OR(g32119, g29547)
--	g28090 = OR(g27275, g18733)
--	g30579 = OR(g30173, g14571)
--	g27858 = OR(g17405, g26737)
--	g25751 = OR(g25061, g22098)
--	g28651 = OR(g27392, g16599)
--	g29495 = OR(g28563, g27614)
--	g33383 = OR(g32244, g29940)
--	g25639 = OR(g25122, g18530)
--	g34014 = OR(g33647, g18493)
--	g33030 = OR(g32166, g21826)
--	g31267 = OR(g29548, g28263)
--	g25638 = OR(g24977, g18316)
--	g34007 = OR(g33640, g18467)
--	g16883 = OR(g13509, g11115)
--	g33267 = OR(g32115, g29535)
--	g33294 = OR(g32152, g29604)
--	g27394 = OR(g25957, g24573)
--	g28331 = OR(g27129, g15814)
--	g30442 = OR(g29797, g21851)
--	g33065 = OR(g32008, g22068)
--	g34442 = OR(g34380, g18542)
--	g28513 = OR(g27276, g26123)
--	g31875 = OR(g31066, g21730)
--	g29643 = OR(g28192, g27145)
--	g34615 = OR(g34516, g18576)
--	g33219 = OR(g32335, I30760, I30761)
--	g24262 = OR(g23387, g18315)
--	g28404 = OR(g27215, g15874)
--	g34720 = OR(g34694, g18134)
--	g34041 = OR(g33829, g18739)
--	g28717 = OR(g27482, g16701)
--	g30430 = OR(g29859, g21814)
--	g30493 = OR(g30198, g21989)
--	g28212 = OR(g27030, g27035)
--	g29260 = OR(g28315, g18604)
--	g25835 = OR(g25367, g23855)
--	g30465 = OR(g30164, g21936)
--	g34465 = OR(g34295, g18712)
--	g25586 = OR(g21678, g24156)
--	g34237 = OR(g32715, g33955)
--	g30340 = OR(g29377, g18245)
--	g29489 = OR(g28550, g27601)
--	g34035 = OR(g33721, g18714)
--	g29488 = OR(g28547, g27600)
--	g34806 = OR(g34763, g18595)
--	g23183 = OR(g19545, g15911)
--	g28723 = OR(g27490, g16706)
--	g33617 = OR(g33263, g24326)
--	g31915 = OR(g31520, g22001)
--	g25615 = OR(g24803, g18162)
--	g30517 = OR(g30244, g22038)
--	g28387 = OR(g27203, g15858)
--	g31277 = OR(g29570, g28285)
--	g25720 = OR(g25042, g18765)
--	g24247 = OR(g22623, g18259)
--	g33277 = OR(g32129, g29568)
--	g14182 = OR(g11741, g11721, g753)
--	g15935 = OR(g13029, g10665)
--	g28097 = OR(g27682, g22005)
--	g28104 = OR(g27697, g22108)
--	g25746 = OR(g25217, g22063)
--	g28646 = OR(g27388, g16595)
--	g33595 = OR(g33368, g18489)
--	g32235 = OR(g31151, g29662)
--	g27562 = OR(g26102, g24703)
--	g33623 = OR(g33370, g18792)
--	I30756 = OR(g32088, g32163, g32098, g32105)
--	g33037 = OR(g32177, g24310)
--	g30362 = OR(g30120, g18392)
--	g34193 = OR(g33809, g33814)
--	g24251 = OR(g22637, g18296)
--	g24272 = OR(g23056, g18629)
--	g31782 = OR(g30060, g30070)
--	g27290 = OR(g25926, g25928)
--	g28369 = OR(g27160, g25938)
--	g30523 = OR(g30245, g22069)
--	g33984 = OR(g33881, g18374)
--	g25684 = OR(g24983, g18643)
--	g29255 = OR(g28714, g18516)
--	g28368 = OR(g27158, g27184)
--	g26703 = OR(g24447, g10705)
--	g29270 = OR(g28258, g18635)
--	g32991 = OR(g32322, g18349)
--	g30475 = OR(g30220, g21946)
--	g34006 = OR(g33897, g18462)
--	g28850 = OR(g27557, g16869)
--	g33266 = OR(g32114, g29532)
--	g23574 = OR(g20093, g20108)
--	g13972 = OR(g11232, g11203)
--	g34727 = OR(g34655, g18213)
--	g26781 = OR(g24913, g24921)
--	g30437 = OR(g29876, g21846)
--	g26952 = OR(g26360, g24290)
--	g29294 = OR(g28645, g18779)
--	g29267 = OR(g28257, g18622)
--	g19619 = OR(g15712, g13080)
--	g8863 = OR(g1644, g1664)
--	g19557 = OR(g17123, g14190)
--	I22830 = OR(g21429, g21338, g21307)
--	g27403 = OR(g25962, g24581)
--	g33589 = OR(g33340, g18469)
--	g30347 = OR(g29383, g18304)
--	g28716 = OR(g27481, g13887)
--	g34347 = OR(g25986, g34102)
--	g33588 = OR(g33334, g18468)
--	g34253 = OR(g34171, g24300)
--	g27226 = OR(g25872, g24436)
--	g28582 = OR(g27330, g26277)
--	g34600 = OR(g34538, g18182)
--	g24447 = OR(g10948, g22450)
--	g14387 = OR(g9086, g11048)
--	g34781 = OR(g33431, g34715)
--	g27551 = OR(g26091, g24675)
--	g27572 = OR(g26129, g24724)
--	g33119 = OR(g32420, g32428)
--	g28310 = OR(g27107, g15797)
--	g34236 = OR(g32650, g33954)
--	g30351 = OR(g30084, g18339)
--	g30372 = OR(g30110, g18446)
--	g25727 = OR(g25163, g22010)
--	g33118 = OR(g32413, g32418)
--	g34372 = OR(g26287, g34137)
--	g31864 = OR(g31271, g21703)
--	g33022 = OR(g32306, g21750)
--	g26422 = OR(g24774, g23104)
--	g31749 = OR(g29974, g29988)
--	g16052 = OR(g13060, g10724)
--	g7450 = OR(g1277, g1283)
--	g28050 = OR(g27692, g18165)
--	g33616 = OR(g33237, g24314)
--	g33313 = OR(g29649, g32171)
--	g30516 = OR(g30233, g22037)
--	g34264 = OR(g34081, g18701)
--	g28386 = OR(g27202, g13277)
--	g34790 = OR(g34774, g18151)
--	g31276 = OR(g29567, g28282)
--	g25703 = OR(g25087, g21922)
--	g28603 = OR(g27340, g26300)
--	g24246 = OR(g23372, g18257)
--	g33276 = OR(g32128, g29566)
--	g28096 = OR(g27988, g21997)
--	g32399 = OR(g31527, g30062)
--	g33053 = OR(g31967, g21974)
--	g31254 = OR(g25981, g29534)
--	g27980 = OR(g26105, g26131)
--	g33254 = OR(g32104, g29512)
--	g31900 = OR(g31484, g21908)
--	g31466 = OR(g26160, g29650)
--	g32398 = OR(g31526, g30061)
--	I22267 = OR(g20236, g20133, g20111)
--	g25600 = OR(g24650, g18111)
--	g26913 = OR(g25848, g18225)
--	g28681 = OR(g27428, g16634)
--	g23405 = OR(g19791, g16245)
--	g29277 = OR(g28440, g18710)
--	g30422 = OR(g29795, g21806)
--	g33036 = OR(g32168, g24309)
--	g28429 = OR(g27228, g15913)
--	g33560 = OR(g33404, g18369)
--	g24355 = OR(g23799, g18824)
--	g28730 = OR(g27503, g13912)
--	g26905 = OR(g26397, g24222)
--	g25821 = OR(g25482, g25456, g25417, g25377)
--	g28428 = OR(g27227, g15912)
--	g30542 = OR(g29337, g22088)
--	g30453 = OR(g29902, g21862)
--	g33064 = OR(g31993, g22067)
--	g19363 = OR(g17810, g14913)
--	g28690 = OR(g27436, g16641)
--	g34021 = OR(g33652, g18519)
--	g34453 = OR(g34410, g18666)
--	g27426 = OR(g25967, g24588)
--	g28549 = OR(g27304, g26233)
--	g24151 = OR(g18088, g21661)
--	g33733 = OR(g33105, g32012)
--	g32361 = OR(g29869, g31300)
--	g34726 = OR(g34665, g18212)
--	g28548 = OR(g27303, g26232)
--	g31874 = OR(g31016, g21729)
--	g30436 = OR(g29860, g21845)
--	g19486 = OR(g15589, g12979)
--	g34614 = OR(g34518, g18568)
--	g29266 = OR(g28330, g18621)
--	g34607 = OR(g34567, g15081)
--	g30530 = OR(g30224, g22076)
--	g28317 = OR(g27114, g15805)
--	g33009 = OR(g32273, g18458)
--	g34274 = OR(g27822, g34205)
--	g30346 = OR(g29381, g18303)
--	g25834 = OR(g25366, g23854)
--	g27024 = OR(g26826, g17692)
--	I31849 = OR(g33483, g33484, g33485, g33486)
--	g33008 = OR(g32261, g18457)
--	g30464 = OR(g30152, g21935)
--	g32221 = OR(g31140, g29634)
--	g34464 = OR(g34340, g18687)
--	g31892 = OR(g31019, g21825)
--	I31848 = OR(g33479, g33480, g33481, g33482)
--	g28057 = OR(g27033, g18218)
--	g34034 = OR(g33719, g18713)
--	g33555 = OR(g33355, g18357)
--	g34641 = OR(g34479, g18724)
--	g34797 = OR(g34747, g18574)
--	g25726 = OR(g25148, g22009)
--	g33570 = OR(g33420, g18405)
--	g31914 = OR(g31499, g22000)
--	g34292 = OR(g26853, g34223)
--	g28323 = OR(g27118, g15810)
--	g33914 = OR(g33305, g33311)
--	g34153 = OR(g33899, g33451)
--	g27126 = OR(g24378, g25787)
--	g25614 = OR(g24797, g18161)
--	g28533 = OR(g27291, g26203)
--	g31907 = OR(g31492, g21954)
--	g30409 = OR(g29842, g21768)
--	g27250 = OR(g25901, g15738)
--	g26891 = OR(g26652, g24197)
--	g24203 = OR(g22982, g18107)
--	g25607 = OR(g24773, g18118)
--	g10802 = OR(g7533, g1296)
--	g15732 = OR(g13411, g13384, g13349, g11016)
--	g28775 = OR(g27537, g16806)
--	g30408 = OR(g29806, g21767)
--	g29864 = OR(g28272, g26086)
--	g34635 = OR(g34485, g18692)
--	g25593 = OR(g24716, g21707)
--	g33567 = OR(g33081, g18394)
--	g33594 = OR(g33421, g18485)
--	g32371 = OR(g29883, g31313)
--	g29313 = OR(g28284, g27270)
--	g24281 = OR(g23397, g18656)
--	g33238 = OR(g32048, g32051)
--	g26327 = OR(g8462, g24591)
--	g22225 = OR(g21332, g17654)
--	g29748 = OR(g28210, g28214)
--	g22708 = OR(g19266, g15711)
--	g29276 = OR(g28616, g18709)
--	g29285 = OR(g28639, g18750)
--	g29305 = OR(g28602, g18811)
--	g29254 = OR(g28725, g18512)
--	g33176 = OR(g32198, I30734, I30735)
--	g16882 = OR(g13508, g11114)
--	g30474 = OR(g30208, g21945)
--	g25635 = OR(g24504, g18293)
--	g31883 = OR(g31132, g21777)
--	g30537 = OR(g30246, g22083)
--	g19587 = OR(g15700, g13046)
--	I30331 = OR(g31672, g31710, g31021, g30937)
--	g34537 = OR(g34324, g34084)
--	g13794 = OR(g7396, g10684)
--	g34283 = OR(g26839, g34215)
--	g30492 = OR(g30188, g21988)
--	g34606 = OR(g34564, g15080)
--	g34303 = OR(g25768, g34045)
--	g28316 = OR(g27113, g15804)
--	g27581 = OR(g26161, g24750)
--	g27450 = OR(g2917, g26483)
--	I30717 = OR(g31787, g32200, g31940, g31949)
--	g33577 = OR(g33405, g18430)
--	g30381 = OR(g30126, g18497)
--	g25575 = OR(g24139, g24140)
--	g28056 = OR(g27230, g18210)
--	g32359 = OR(g29867, g31298)
--	g27257 = OR(g25904, g24498)
--	g29166 = OR(g27653, g17153)
--	g25711 = OR(g25105, g21962)
--	g28611 = OR(g27348, g16485)
--	g24715 = OR(g22189, g22207)
--	g32358 = OR(g29866, g31297)
--	g34796 = OR(g34745, g18573)
--	g29892 = OR(g28300, g26120)
--	g27590 = OR(g26179, g24764)
--	g29476 = OR(g28108, g28112)
--	g29485 = OR(g28535, g27594)
--	g31906 = OR(g31477, g21953)
--	g30390 = OR(g29985, g18555)
--	g32344 = OR(g29804, g31266)
--	g31284 = OR(g29575, g28290)
--	g25606 = OR(g24761, g18117)
--	g28342 = OR(g27134, g15819)
--	g31304 = OR(g29594, g29608)
--	g29914 = OR(g22531, g22585, I28147)
--	g21897 = OR(g20095, g15111)
--	g33622 = OR(g33366, g18791)
--	g33566 = OR(g33356, g18390)
--	g25750 = OR(g25543, g18802)
--	g26949 = OR(g26356, g24287)
--	g28650 = OR(g27391, g16598)
--	g30522 = OR(g29332, g22064)
--	g27150 = OR(g25804, g24400)
--	g34663 = OR(g32028, g34500)
--	g29239 = OR(g28427, g18297)
--	g26948 = OR(g26399, g24286)
--	g24354 = OR(g23775, g18823)
--	g27019 = OR(g26822, g14610)
--	g26904 = OR(g26393, g24221)
--	g29238 = OR(g28178, g18292)
--	g30483 = OR(g30241, g21979)
--	g30553 = OR(g30205, g22124)
--	g22901 = OR(g19384, g15745)
--	g28132 = OR(g27932, g27957)
--	g13997 = OR(g11029, g11036)
--	g29176 = OR(g27661, g17177)
--	g30536 = OR(g30234, g22082)
--	g26673 = OR(g24433, g10674)
--	g34040 = OR(g33818, g18737)
--	g33963 = OR(g33830, g18124)
--	g25663 = OR(g24666, g21788)
--	g34252 = OR(g34146, g18180)
--	g34621 = OR(g34517, g18583)
--	g28708 = OR(g27462, g16674)
--	g26933 = OR(g26808, g18551)
--	g28087 = OR(g27255, g18720)
--	g33576 = OR(g33401, g18423)
--	g33585 = OR(g33411, g18456)
--	g24211 = OR(g23572, g18138)
--	g28043 = OR(g27323, g21714)
--	g33554 = OR(g33407, g18353)
--	g32240 = OR(g24757, g31182)
--	g30397 = OR(g29747, g21756)
--	I26742 = OR(g23430, g23445, g23458, g23481)
--	g33609 = OR(g33239, g18615)
--	g29501 = OR(g28583, g27634)
--	g33312 = OR(g29646, g32170)
--	g30509 = OR(g30210, g22030)
--	g33608 = OR(g33322, g18537)
--	g28069 = OR(g27564, g21865)
--	g33115 = OR(g32397, g32401)
--	g25702 = OR(g25068, g21921)
--	g25757 = OR(g25132, g22104)
--	g28774 = OR(g27536, g16804)
--	g30508 = OR(g30199, g22029)
--	g31921 = OR(g31508, g22046)
--	g28068 = OR(g27310, g21838)
--	g32981 = OR(g32425, g18206)
--	g28375 = OR(g27183, g15851)
--	g33052 = OR(g31961, g21973)
--	g34634 = OR(g34483, g18691)
--	g25621 = OR(g24523, g18205)
--	g31745 = OR(g29959, g29973)
--	g21896 = OR(g20084, g15110)
--	g24250 = OR(g22633, g18295)
--	g26912 = OR(g25946, g18209)
--	g27231 = OR(g25873, g15699)
--	g29284 = OR(g28554, g18747)
--	g32395 = OR(g31523, g30049)
--	g24339 = OR(g23690, g18756)
--	g33973 = OR(g33840, g18344)
--	g29304 = OR(g28588, g18810)
--	g32262 = OR(g31186, g29710)
--	g23716 = OR(g9194, g20905)
--	g25673 = OR(g24727, g21830)
--	g32990 = OR(g32281, g18341)
--	I18417 = OR(g14444, g14414, g14392)
--	g24338 = OR(g23658, g18755)
--	g11370 = OR(g8807, g550)
--	g30452 = OR(g29891, g21861)
--	g34452 = OR(g34401, g18665)
--	g13858 = OR(g209, g10685)
--	g33732 = OR(g33104, g32011)
--	g30311 = OR(g28265, g27265)
--	g24968 = OR(g22360, g22409, g23389)
--	g25634 = OR(g24559, g18284)
--	g31761 = OR(g30009, g30028)
--	g33692 = OR(g32400, g33428)
--	g19475 = OR(g16930, g14126)
--	g27456 = OR(g25978, g24607)
--	g26396 = OR(g24762, g23062)
--	g28545 = OR(g27301, g26230)
--	g28078 = OR(g27140, g21880)
--	g33013 = OR(g32283, g18484)
--	g22669 = OR(g7763, g19525)
--	g32247 = OR(g31168, g29686)
--	I18543 = OR(g14568, g14540, g14516)
--	g28086 = OR(g27268, g18702)
--	g32389 = OR(g31496, g29966)
--	g30350 = OR(g30118, g18334)
--	g34350 = OR(g26048, g34106)
--	g33539 = OR(g33245, g18178)
--	g32388 = OR(g31495, g29962)
--	g33005 = OR(g32260, g18432)
--	g27596 = OR(g26207, g24775)
--	g11025 = OR(g2980, g7831)
--	g28817 = OR(g27548, g16845)
--	g33538 = OR(g33252, g18144)
--	g28322 = OR(g27117, g15809)
--	g27243 = OR(g25884, g24475)
--	g30396 = OR(g29856, g21755)
--	g32251 = OR(g30599, g29352)
--	g13540 = OR(g10822, g10827)
--	g27431 = OR(g24582, g25977)
--	g20202 = OR(g16211, g13507)
--	g34731 = OR(g34662, g18272)
--	g29484 = OR(g28124, g22191)
--	g24202 = OR(g22899, g18106)
--	g26929 = OR(g26635, g18543)
--	g24257 = OR(g22938, g18310)
--	g30413 = OR(g30001, g21772)
--	g24496 = OR(g24008, g21557)
--	g31241 = OR(g25959, g29510)
--	g26928 = OR(g26713, g18541)
--	g17488 = OR(g14361, g14335, g11954, I18417)
--	g25592 = OR(g24672, g21706)
--	g25756 = OR(g25112, g22103)
--	g28561 = OR(g27312, g26250)
--	g28295 = OR(g27094, g15783)
--	g28680 = OR(g27427, g16633)
--	g32997 = OR(g32269, g18378)
--	g30405 = OR(g29767, g21764)
--	g16173 = OR(g8796, g13464)
--	g34405 = OR(g34183, g25103)
--	g33235 = OR(g32040, g30982)
--	g23317 = OR(g19715, g16191)
--	I22852 = OR(g21459, g21350, g21339)
--	g29813 = OR(g26020, g28261)
--	g22679 = OR(g19145, g15701)
--	g23129 = OR(g19500, g15863)
--	g13699 = OR(g10921, g10947)
--	g34020 = OR(g33904, g18514)
--	g25731 = OR(g25128, g22014)
--	g28631 = OR(g27372, g16534)
--	I28567 = OR(g29204, g29205, g29206, g29207)
--	I24117 = OR(g23088, g23154, g23172)
--	g32360 = OR(g29868, g31299)
--	g16506 = OR(g13294, g10966)
--	g15789 = OR(g10819, g13211)
--	I30261 = OR(g29385, g31376, g30735, g30825)
--	g34046 = OR(g33906, g33908)
--	g31882 = OR(g31115, g21776)
--	g33991 = OR(g33885, g18400)
--	g14078 = OR(g10776, g8703)
--	g20196 = OR(g16207, g13497)
--	g25691 = OR(g24536, g21890)
--	g27487 = OR(g25990, g24629)
--	g34282 = OR(g26838, g34214)
--	g23298 = OR(g19693, g16179)
--	g30357 = OR(g30107, g18366)
--	g28309 = OR(g27106, g15796)
--	g32220 = OR(g31139, g29633)
--	g26881 = OR(g26629, g24187)
--	g16927 = OR(g13524, g11126)
--	g25929 = OR(g24395, g22193)
--	g28308 = OR(g27105, g15795)
--	g27278 = OR(g15786, g25921)
--	g29692 = OR(g28197, g10873)
--	g24457 = OR(g10902, g22400)
--	g14977 = OR(g10776, g8703)
--	g25583 = OR(g21666, g24153)
--	g33584 = OR(g33406, g18449)
--	g34640 = OR(g34487, g18723)
--	g19274 = OR(g17753, g14791)
--	g19593 = OR(g17145, g14210)
--	g34803 = OR(g34758, g18590)
--	g28816 = OR(g27547, g16843)
--	g20077 = OR(g16025, g13320)
--	g23261 = OR(g19660, g16125)
--	g26890 = OR(g26630, g24196)
--	g28687 = OR(g27434, g16638)
--	g29539 = OR(g2864, g28220)
--	g32355 = OR(g29855, g31286)
--	g34881 = OR(g34866, g18187)
--	g24256 = OR(g22873, g18309)
--	g32370 = OR(g29882, g31312)
--	g28374 = OR(g27181, g15850)
--	g24280 = OR(g23292, g15109)
--	g25743 = OR(g25110, g22058)
--	g28643 = OR(g27386, g16592)
--	g27937 = OR(g14506, g26793)
--	g32996 = OR(g32256, g18377)
--	g34027 = OR(g33718, g18683)
--	g29241 = OR(g28638, g18332)
--	g13385 = OR(g11967, g9479)
--	
--	g11980 = NAND(I14817, I14818)
--	g13889 = NAND(g11566, g11435)
--	g13980 = NAND(g10295, g11435)
--	g12169 = NAND(g9804, g5448)
--	I22761 = NAND(g11939, I22760)
--	I13443 = NAND(g262, I13442)
--	I14185 = NAND(g8442, g3470)
--	g16719 = NAND(g3243, g13700, g3310, g11350)
--	I14518 = NAND(g661, I14516)
--	g10224 = NAND(g6661, g6704, g6675, g6697)
--	g17595 = NAND(g8616, g14367)
--	g22984 = NAND(g20114, g2868)
--	I12346 = NAND(g3111, I12344)
--	g12478 = NAND(I15299, I15300)
--	g21432 = NAND(g17790, g14820, g17761, g14780)
--	g28830 = NAND(g27886, g7451, g7369)
--	I14883 = NAND(g9500, g5489)
--	g19474 = NAND(g11609, g17794)
--	g11426 = NAND(g8742, g4878)
--	g11190 = NAND(g8539, g3447)
--	g9852 = NAND(g3684, g4871)
--	g23342 = NAND(g6928, g21163)
--	g27223 = NAND(I25908, I25909)
--	I15089 = NAND(g2393, I15087)
--	g22853 = NAND(g20219, g2922)
--	g25003 = NAND(g21353, g23462)
--	I15088 = NAND(g9832, I15087)
--	g24916 = NAND(g19450, g23154)
--	g25779 = NAND(g19694, g24362)
--	g12084 = NAND(g2342, g8211)
--	g28270 = NAND(g10504, g26105, g26987)
--	g22836 = NAND(g18918, g2852)
--	g21330 = NAND(g11401, g17157)
--	g20076 = NAND(g13795, g16521)
--	g21365 = NAND(g15744, g13119, g15730, g13100)
--	g23132 = NAND(g8155, g19932)
--	I22683 = NAND(g11893, g21434)
--	g28938 = NAND(g27796, g8205)
--	g9825 = NAND(I13391, I13392)
--	g7201 = NAND(I11865, I11866)
--	g15719 = NAND(g5256, g14490, g5335, g9780)
--	g27654 = NAND(g164, g26598, g23042)
--	g22864 = NAND(g7780, g21156)
--	I20165 = NAND(g16246, g990)
--	g14489 = NAND(g12126, g5084)
--	g29082 = NAND(g27837, g9694)
--	g25233 = NAND(g20838, g23623)
--	g24942 = NAND(g20039, g23172)
--	I26459 = NAND(g26576, g14306)
--	g15832 = NAND(g7903, g7479, g13256)
--	g14830 = NAND(g6605, g12211, g6723, g12721)
--	I32431 = NAND(g34056, g34051)
--	g9972 = NAND(I13510, I13511)
--	I20222 = NAND(g16272, I20221)
--	g17748 = NAND(g562, g14708, g12323)
--	g11969 = NAND(g7252, g1636)
--	g20734 = NAND(g14408, g17312)
--	g28837 = NAND(g27800, g7374, g2197)
--	I25244 = NAND(g24744, I25242)
--	g11968 = NAND(g837, g9334, g9086)
--	g13968 = NAND(g3913, g11255, g4031, g11631)
--	g15045 = NAND(g12716, g7142)
--	g12423 = NAND(I15242, I15243)
--	g27587 = NAND(g24917, g25018, g24918, g26857)
--	g20838 = NAND(g5041, g17284)
--	g13855 = NAND(g4944, g11804)
--	g19483 = NAND(g15969, g10841, g10922)
--	g10610 = NAND(g7462, g7490)
--	g11411 = NAND(g9713, g3625)
--	I13110 = NAND(g5808, I13109)
--	g22642 = NAND(g7870, g19560)
--	g12587 = NAND(g7497, g6315)
--	g13870 = NAND(g11773, g4732)
--	g13527 = NAND(g182, g168, g203, g12812)
--	g23810 = NAND(I22973, I22974)
--	g20619 = NAND(g14317, g17217)
--	g16628 = NAND(g3602, g11207, g3618, g13902)
--	I23119 = NAND(g20076, I23118)
--	g10124 = NAND(g5276, g5320, g5290, g5313)
--	g12000 = NAND(g8418, g2610)
--	I23118 = NAND(g20076, g417)
--	g22874 = NAND(g18918, g2844)
--	g10939 = NAND(g7352, g1459)
--	g13867 = NAND(g11312, g8449)
--	g14686 = NAND(g5268, g12059, g5276, g12239)
--	I12840 = NAND(g4222, g4235)
--	g29049 = NAND(g9640, g27779)
--	g16776 = NAND(g3945, g13772, g4012, g11419)
--	g13315 = NAND(g1459, g10715)
--	g11707 = NAND(g8718, g4864)
--	I18530 = NAND(g1811, I18529)
--	g20039 = NAND(g11250, g17794)
--	I14609 = NAND(g8993, g8678)
--	I13334 = NAND(g1687, g1691)
--	g13257 = NAND(g1389, g10544)
--	g29004 = NAND(g27933, g8330)
--	g21459 = NAND(g17814, g14854, g17605, g17581)
--	g11979 = NAND(g9861, g5452)
--	g13496 = NAND(g1351, g11336, g11815)
--	g11590 = NAND(g6928, g3990, g4049)
--	g12639 = NAND(g10194, g6682, g6732)
--	g22712 = NAND(g18957, g2864)
--	g23010 = NAND(g20516, g2984)
--	g7897 = NAND(I12288, I12289)
--	g24601 = NAND(g22957, g2965)
--	g13986 = NAND(g10323, g11747)
--	g12293 = NAND(g7436, g5283)
--	g24677 = NAND(g22957, g2975)
--	g12638 = NAND(g7514, g6661)
--	g24975 = NAND(g21388, g23363)
--	g10160 = NAND(g5623, g5666, g5637, g5659)
--	g17712 = NAND(g5599, g14425, g5666, g12301)
--	g12416 = NAND(g10133, g7064, g10166)
--	g14160 = NAND(g11626, g8958)
--	g28853 = NAND(g27742, g1636, g7252)
--	g13067 = NAND(g5240, g12059, g5331, g9780)
--	g28167 = NAND(g925, g27046)
--	I18635 = NAND(g14713, I18633)
--	g10617 = NAND(g10151, g9909)
--	g16319 = NAND(g8224, g8170, g13736)
--	I32187 = NAND(g33661, I32185)
--	I12252 = NAND(g1124, I12251)
--	g14915 = NAND(g12553, g10266)
--	g22941 = NAND(g20219, g2970)
--	I17406 = NAND(g1472, I17404)
--	g12578 = NAND(g7791, g10341)
--	g27586 = NAND(g24924, g24916, g24905, g26863)
--	g12014 = NAND(g7197, g703)
--	g14075 = NAND(g11658, g11527)
--	g15591 = NAND(g4332, g4322, g13202)
--	g28864 = NAND(g27886, g7411, g1996)
--	g10623 = NAND(g10181, g9976)
--	g17675 = NAND(g5252, g14399, g5320, g12239)
--	g23656 = NAND(I22800, I22801)
--	g21353 = NAND(g11467, g17157)
--	I13751 = NAND(g4584, I13749)
--	g14782 = NAND(g12755, g10491)
--	I14400 = NAND(g3654, I14398)
--	g12116 = NAND(g2051, g8255)
--	g14984 = NAND(g7812, g12680)
--	g13866 = NAND(g3239, g11194, g3321, g11519)
--	I18537 = NAND(g2236, I18536)
--	g16281 = NAND(g4754, g13937, g12054)
--	g28900 = NAND(g27886, g7451, g2040)
--	g14822 = NAND(g12755, g12632)
--	g14170 = NAND(g11715, g11537)
--	g15844 = NAND(g14714, g9340, g12378)
--	I22972 = NAND(g9657, g19638)
--	g21364 = NAND(g15787, g15781, g15753, g13131)
--	I13391 = NAND(g1821, I13390)
--	g13256 = NAND(g11846, g11294, g11812)
--	I13510 = NAND(g2089, I13509)
--	g11923 = NAND(I14734, I14735)
--	g12340 = NAND(g4888, g8984)
--	g12035 = NAND(g10000, g6144)
--	g13923 = NAND(g11692, g11527)
--	I15300 = NAND(g1982, I15298)
--	g9830 = NAND(I13402, I13403)
--	g20186 = NAND(g16926, g8177)
--	g20676 = NAND(g14379, g17287)
--	g21289 = NAND(g14616, g17493)
--	I12205 = NAND(g1135, I12203)
--	g13102 = NAND(g7523, g10759)
--	g25429 = NAND(g22417, g1917, g8302)
--	g23309 = NAND(g6905, g21024)
--	g28874 = NAND(g27907, g7424, g2421)
--	g29121 = NAND(g9755, g27886)
--	g21288 = NAND(g14616, g17492)
--	g7582 = NAND(g1361, g1373)
--	I13442 = NAND(g262, g239)
--	g13066 = NAND(g4430, g7178, g10590)
--	g24936 = NAND(g20186, g20173, g23379, g14029)
--	g31262 = NAND(g767, g29916, g11679)
--	g10022 = NAND(g6474, g6466)
--	g14864 = NAND(g7791, g10421)
--	g8769 = NAND(g691, g714)
--	g7227 = NAND(g4584, g4593)
--	I32186 = NAND(g33665, I32185)
--	g12523 = NAND(g7563, g6346)
--	g28892 = NAND(g27779, g1772, g7275)
--	g13854 = NAND(g4765, g11797)
--	g11511 = NAND(I14481, I14482)
--	I14991 = NAND(g9685, g6527)
--	g8967 = NAND(g4264, g4258)
--	g13511 = NAND(g182, g174, g203, g12812)
--	g20216 = NAND(I20487, I20488)
--	g14254 = NAND(g11968, g11933, g11951)
--	g28914 = NAND(g27937, g7462, g2555)
--	g29134 = NAND(g9762, g27907)
--	g28907 = NAND(g27858, g2361, g2287)
--	g12222 = NAND(g8310, g2028)
--	g29028 = NAND(g27933, g8381)
--	g22852 = NAND(g18957, g2856)
--	g14101 = NAND(g11653, g11729)
--	g25002 = NAND(g19474, g23154)
--	I29297 = NAND(g12117, I29295)
--	g14177 = NAND(g11741, g11721, g753)
--	g11480 = NAND(g10323, g8906)
--	I26460 = NAND(g26576, I26459)
--	I22946 = NAND(g19620, I22944)
--	I18536 = NAND(g2236, g14642)
--	I15287 = NAND(g10061, g6697)
--	I14206 = NAND(g3821, I14204)
--	g16956 = NAND(g3925, g13824, g4019, g11631)
--	I26093 = NAND(g26055, g13539)
--	I15307 = NAND(g10116, I15306)
--	g23195 = NAND(g20136, g37)
--	g13307 = NAND(g1116, g10695)
--	I15243 = NAND(g6351, I15241)
--	g16181 = NAND(g13475, g13495, g13057, g13459)
--	g12351 = NAND(I15194, I15195)
--	g24814 = NAND(g20011, g23167)
--	g22312 = NAND(g907, g19063)
--	g28935 = NAND(g27800, g2227, g7328)
--	g24807 = NAND(I23979, I23980)
--	I15341 = NAND(g10154, I15340)
--	g14665 = NAND(g12604, g12798)
--	g24974 = NAND(g21301, g23363)
--	g31997 = NAND(g22306, g30580)
--	g14008 = NAND(g11610, g11435)
--	I14399 = NAND(g8542, I14398)
--	I22760 = NAND(g11939, g21434)
--	g9258 = NAND(I13044, I13045)
--	g22921 = NAND(g20219, g2950)
--	g15715 = NAND(g336, g305, g13385)
--	g17312 = NAND(g7297, g14248)
--	g25995 = NAND(g24621, g22853)
--	g14892 = NAND(g12700, g12515)
--	g17608 = NAND(g5953, g12067, g5969, g14701)
--	I14398 = NAND(g8542, g3654)
--	g15572 = NAND(g12969, g7219)
--	I18634 = NAND(g2504, I18633)
--	I15335 = NAND(g2116, I15333)
--	g34056 = NAND(I31984, I31985)
--	g14570 = NAND(g3933, g11255, g4023, g8595)
--	g11993 = NAND(g1894, g8302)
--	g13993 = NAND(g3961, g11255, g3969, g11419)
--	I23963 = NAND(g13631, I23961)
--	g9975 = NAND(I13519, I13520)
--	g21124 = NAND(g5731, g17393)
--	I14332 = NAND(g9966, I14330)
--	g13667 = NAND(g3723, g11119)
--	g13131 = NAND(g6243, g12101, g6377, g10003)
--	g10567 = NAND(g1862, g7405)
--	g20007 = NAND(g11512, g17794)
--	I23585 = NAND(g22409, g4332)
--	g28349 = NAND(g27074, g24770, g27187, g19644)
--	g29719 = NAND(g28406, g13739)
--	g21294 = NAND(g11324, g17157)
--	g25498 = NAND(g22498, g2610, g8418)
--	g28906 = NAND(g27796, g8150)
--	g13210 = NAND(g7479, g10521)
--	g34650 = NAND(I32757, I32758)
--	g16625 = NAND(g3203, g13700, g3274, g11519)
--	g17732 = NAND(g3937, g13824, g4012, g13933)
--	g10185 = NAND(g5969, g6012, g5983, g6005)
--	g11443 = NAND(g9916, g3649)
--	g12436 = NAND(I15263, I15264)
--	g11279 = NAND(g8504, g3443)
--	g14519 = NAND(g3889, g11225, g4000, g8595)
--	I29296 = NAND(g29495, I29295)
--	g14675 = NAND(g12317, g9898)
--	I25219 = NAND(g482, g24718)
--	g27593 = NAND(g24972, g24950, g24906, g26861)
--	I26419 = NAND(g14247, I26417)
--	I22755 = NAND(g21434, I22753)
--	g12073 = NAND(g10058, g6490)
--	g14154 = NAND(g11669, g8958)
--	g17761 = NAND(g6291, g14529, g6358, g12423)
--	I26418 = NAND(g26519, I26417)
--	g13469 = NAND(g4983, g10862)
--	g25432 = NAND(g12374, g22384)
--	g10935 = NAND(g1459, g7352)
--	g14637 = NAND(g12255, g9815)
--	I15306 = NAND(g10116, g2407)
--	g16296 = NAND(g9360, g13501)
--	g25271 = NAND(I24462, I24463)
--	g7133 = NAND(I11825, I11826)
--	g12464 = NAND(g10169, g7087, g10191)
--	g7846 = NAND(g4843, g4878)
--	g12797 = NAND(g10275, g7655, g7643, g7627)
--	I22794 = NAND(g21434, I22792)
--	I22845 = NAND(g12113, I22844)
--	g7803 = NAND(I12204, I12205)
--	g31950 = NAND(g7285, g30573)
--	g12292 = NAND(g4698, g8933)
--	g9461 = NAND(I13140, I13141)
--	g12153 = NAND(g2610, g8330)
--	g25199 = NAND(I24364, I24365)
--	I22899 = NAND(g12193, g21228)
--	g8829 = NAND(g5011, g4836)
--	g11975 = NAND(g8267, g8316)
--	I12204 = NAND(g1094, I12203)
--	g19513 = NAND(g15969, g10841, g10922)
--	g23617 = NAND(I22761, I22762)
--	g15024 = NAND(g12780, g10421)
--	I20205 = NAND(g11147, I20203)
--	g12136 = NAND(I14992, I14993)
--	I22719 = NAND(g21434, I22717)
--	g9904 = NAND(I13443, I13444)
--	g13143 = NAND(g10695, g7661, g979, g1061)
--	I13453 = NAND(g1955, I13452)
--	I22718 = NAND(g11916, I22717)
--	g33394 = NAND(g10159, g4474, g32426)
--	g11169 = NAND(I14229, I14230)
--	I29315 = NAND(g12154, I29313)
--	I15168 = NAND(g9823, I15166)
--	g13884 = NAND(g11797, g4727)
--	g11410 = NAND(g6875, g6895, g8696)
--	g23623 = NAND(g9364, g20717)
--	g9391 = NAND(I13110, I13111)
--	I15363 = NAND(g10182, g2675)
--	g8124 = NAND(I12402, I12403)
--	g24362 = NAND(g21370, g22136)
--	g11479 = NAND(g6875, g3288, g3347)
--	g23782 = NAND(g2741, g21062)
--	g13666 = NAND(g11190, g8441)
--	g13479 = NAND(g12686, g12639, g12590, g12526)
--	g8069 = NAND(I12373, I12374)
--	I32517 = NAND(g34424, I32516)
--	g13217 = NAND(g4082, g10808)
--	g10622 = NAND(g10178, g9973)
--	g10566 = NAND(g7315, g7356)
--	g13478 = NAND(g12511, g12460, g12414, g12344)
--	I13565 = NAND(g2648, I13564)
--	I13464 = NAND(g2384, I13462)
--	g13486 = NAND(g10862, g4983, g4966)
--	g25258 = NAND(I24439, I24440)
--	g23266 = NAND(g18918, g2894)
--	g13580 = NAND(g11849, g7503, g7922, g10544)
--	g10653 = NAND(g10204, g10042)
--	g14139 = NAND(g11626, g11584)
--	g16741 = NAND(g3207, g13765, g3303, g11519)
--	I14789 = NAND(g9891, I14788)
--	g23167 = NAND(g8219, g19981)
--	g13084 = NAND(g5587, g12093, g5677, g9864)
--	g28973 = NAND(g27907, g2465, g7387)
--	g14636 = NAND(g5595, g12029, g5677, g12563)
--	I14788 = NAND(g9891, g6167)
--	g14333 = NAND(g12042, g12014, g11990, g11892)
--	I17462 = NAND(g1300, I17460)
--	g21401 = NAND(g17755, g14730, g17712, g14695)
--	g27796 = NAND(g21228, g25263, g26424, g26171)
--	g20236 = NAND(g16875, g14014, g16625, g16604)
--	g12796 = NAND(g4467, g6961)
--	g9654 = NAND(g2485, g2453)
--	g15867 = NAND(g14714, g9417, g9340)
--	g25337 = NAND(g22342, g1648, g8187)
--	g28934 = NAND(g27882, g14641)
--	g14664 = NAND(g5220, g12059, g5339, g12497)
--	g16196 = NAND(g13496, g13513, g13079, g13476)
--	g11676 = NAND(g358, g8944, g376, g385)
--	g34545 = NAND(g11679, g794, g34354)
--	I22871 = NAND(g12150, g21228)
--	g11953 = NAND(g8195, g8241)
--	g13676 = NAND(g11834, g11283)
--	g23616 = NAND(I22754, I22755)
--	g29355 = NAND(g24383, g28109)
--	g15581 = NAND(g7232, g12999)
--	g10585 = NAND(g1996, g7451)
--	g9595 = NAND(g2351, g2319)
--	g23748 = NAND(I22872, I22873)
--	I14291 = NAND(g3835, I14289)
--	g11936 = NAND(g8241, g1783)
--	I15334 = NAND(g10152, I15333)
--	g12192 = NAND(g8267, g2319)
--	g10609 = NAND(g10111, g9826)
--	I13109 = NAND(g5808, g5813)
--	g22940 = NAND(g18918, g2860)
--	I12097 = NAND(g1339, I12096)
--	g25425 = NAND(g20081, g23172)
--	g12522 = NAND(g10133, g5990, g6040)
--	g23809 = NAND(I22966, I22967)
--	g17744 = NAND(g6303, g14529, g6373, g12672)
--	I17447 = NAND(g13336, I17446)
--	g28207 = NAND(g12546, g26131, g27977)
--	g17399 = NAND(g9626, g9574, g14535)
--	g14921 = NAND(g12492, g10266)
--	g15741 = NAND(g5244, g14490, g5320, g14631)
--	I32516 = NAND(g34424, g34422)
--	g9629 = NAND(g6462, g6466)
--	I13750 = NAND(g4608, I13749)
--	g14813 = NAND(g7766, g12824)
--	g11543 = NAND(g9714, g3969)
--	I12850 = NAND(g4277, I12848)
--	g13909 = NAND(g11396, g8847, g11674, g8803)
--	g23733 = NAND(g20751, g11178)
--	g15735 = NAND(g5547, g14425, g5659, g9864)
--	g15877 = NAND(g14833, g9340, g12543)
--	g9800 = NAND(g5436, g5428)
--	g14674 = NAND(g5941, g12067, g6023, g12614)
--	g11117 = NAND(g8087, g8186, g8239)
--	g29025 = NAND(g27937, g2629, g7462)
--	g13000 = NAND(g7228, g10598)
--	I22754 = NAND(g11937, I22753)
--	g29540 = NAND(g28336, g13464)
--	g23630 = NAND(g20739, g11123)
--	g22833 = NAND(g1193, g19560, g10666)
--	g15695 = NAND(g1266, g13125)
--	g25532 = NAND(g21360, g23363)
--	g15018 = NAND(g12739, g12515)
--	I13390 = NAND(g1821, g1825)
--	g14732 = NAND(g12662, g12515)
--	g24905 = NAND(g534, g23088)
--	I15242 = NAND(g10003, I15241)
--	g19857 = NAND(g13628, g16296)
--	g17500 = NAND(g14573, g14548)
--	I15123 = NAND(g2102, I15121)
--	g14761 = NAND(g12651, g10281)
--	I22844 = NAND(g12113, g21228)
--	g21555 = NAND(g17846, g14946, g17686, g17650)
--	g16854 = NAND(g3965, g13824, g3976, g8595)
--	g11974 = NAND(g2185, g8259)
--	g31671 = NAND(I29262, I29263)
--	g27933 = NAND(g21228, g25356, g26424, g26236)
--	g19549 = NAND(g15969, g10841, g10899)
--	g8806 = NAND(g358, g370, g376, g385)
--	g11639 = NAND(g8933, g4722)
--	g9823 = NAND(I13383, I13384)
--	g12933 = NAND(g7150, g10515)
--	I25907 = NAND(g26256, g24782)
--	g10207 = NAND(g6315, g6358, g6329, g6351)
--	I20204 = NAND(g16246, I20203)
--	g26752 = NAND(g9397, g25189)
--	g14005 = NAND(g11514, g11729)
--	g16660 = NAND(g3953, g11225, g3969, g13933)
--	I26439 = NAND(g26549, I26438)
--	g17605 = NAND(g5559, g14425, g5630, g12563)
--	g11992 = NAND(g7275, g1772)
--	I29314 = NAND(g29501, I29313)
--	I26438 = NAND(g26549, g14271)
--	I12096 = NAND(g1339, g1322)
--	I23962 = NAND(g23184, I23961)
--	I17446 = NAND(g13336, g956)
--	g28206 = NAND(g12546, g26105, g27985)
--	g25309 = NAND(g22384, g12021)
--	I13564 = NAND(g2648, g2652)
--	I12730 = NAND(g4287, I12728)
--	g7857 = NAND(I12241, I12242)
--	g28758 = NAND(g27779, g7356, g7275)
--	I29269 = NAND(g29486, g12050)
--	g14771 = NAND(g5961, g12129, g5969, g12351)
--	g8913 = NAND(I12877, I12878)
--	g11442 = NAND(g8644, g3288, g3343)
--	I13183 = NAND(g6500, I13182)
--	g14683 = NAND(g12553, g12443)
--	g17514 = NAND(g3917, g13772, g4019, g8595)
--	g25495 = NAND(g12483, g22472)
--	g12592 = NAND(I15364, I15365)
--	I13509 = NAND(g2089, g2093)
--	I14247 = NAND(g1322, g8091)
--	I15041 = NAND(g9752, g1834)
--	g10515 = NAND(g10337, g5022)
--	I13851 = NAND(g862, I13850)
--	g25985 = NAND(g24631, g23956)
--	g14882 = NAND(g12558, g12453)
--	g34424 = NAND(I32440, I32441)
--	g14407 = NAND(g12008, g9807)
--	g19856 = NAND(g13626, g16278, g8105)
--	I23951 = NAND(g13603, I23949)
--	I15340 = NAND(g10154, g2541)
--	g26255 = NAND(g8075, g24779)
--	g12152 = NAND(g2485, g8324)
--	g22325 = NAND(g1252, g19140)
--	g13983 = NAND(g11658, g8906)
--	g16694 = NAND(g3905, g13772, g3976, g11631)
--	g17788 = NAND(g5232, g14490, g5327, g12497)
--	g12413 = NAND(g7521, g5654)
--	g10584 = NAND(g7362, g7405)
--	g28406 = NAND(g27064, g13675)
--	I13452 = NAND(g1955, g1959)
--	g28962 = NAND(g27886, g2040, g7369)
--	I29279 = NAND(g12081, I29277)
--	g28500 = NAND(g590, g27629, g12323)
--	g10759 = NAND(g7537, g324)
--	g15721 = NAND(g7564, g311, g13385)
--	I29278 = NAND(g29488, I29277)
--	I14766 = NAND(g5821, I14764)
--	I15130 = NAND(g2527, I15128)
--	I15193 = NAND(g9935, g6005)
--	I29286 = NAND(g12085, I29284)
--	g14758 = NAND(g7704, g12405)
--	g11130 = NAND(g1221, g7918)
--	g14082 = NAND(g11697, g11537)
--	g11193 = NAND(I14258, I14259)
--	g13130 = NAND(g1351, g11815, g11336)
--	g14107 = NAND(g11571, g11527)
--	g16278 = NAND(g8102, g8057, g13664)
--	g12020 = NAND(g2028, g8365)
--	g19611 = NAND(g1070, g1199, g15995)
--	g23139 = NAND(g21163, g10756)
--	g16306 = NAND(g4944, g13971, g12088)
--	I12261 = NAND(g1454, g1448)
--	g14940 = NAND(g12744, g12581)
--	I18627 = NAND(g14712, I18625)
--	g13475 = NAND(g1008, g11294, g11786)
--	g14848 = NAND(g12651, g12453)
--	g27282 = NAND(g11192, g26269, g26248, g479)
--	g21415 = NAND(g17773, g14771, g17740, g14739)
--	g16815 = NAND(g3909, g13824, g4005, g11631)
--	g13727 = NAND(g174, g203, g168, g12812)
--	g15734 = NAND(g5228, g12059, g5290, g14631)
--	g14804 = NAND(g12651, g12798)
--	g25255 = NAND(g20979, g23659)
--	I13731 = NAND(g4537, I13729)
--	g12357 = NAND(g7439, g6329)
--	g31978 = NAND(g30580, g15591)
--	I22824 = NAND(g21434, I22822)
--	I15253 = NAND(g10078, g1848)
--	g24621 = NAND(g22957, g2927)
--	I18681 = NAND(g2638, I18680)
--	g14962 = NAND(g12558, g10281)
--	g13600 = NAND(g3021, g11039)
--	I22931 = NAND(g21228, I22929)
--	g9645 = NAND(g2060, g2028)
--	g23576 = NAND(I22718, I22719)
--	g19764 = NAND(I20166, I20167)
--	g11952 = NAND(g1624, g8187)
--	I15175 = NAND(g9977, I15174)
--	I32757 = NAND(g34469, I32756)
--	I14370 = NAND(g3303, I14368)
--	g26782 = NAND(g9467, g25203)
--	g13821 = NAND(g11251, g8340)
--	g14048 = NAND(g11658, g11483)
--	I15264 = NAND(g2273, I15262)
--	g22755 = NAND(g20136, g18984)
--	g28421 = NAND(g27074, g13715)
--	g26352 = NAND(g744, g24875, g11679)
--	I12271 = NAND(g956, I12269)
--	g13264 = NAND(g11869, g11336, g11849)
--	g24933 = NAND(g19466, g23154)
--	g13137 = NAND(g10699, g7675, g1322, g1404)
--	g13516 = NAND(g11533, g11490, g11444, g11412)
--	g15039 = NAND(g12755, g7142)
--	g29060 = NAND(g9649, g27800)
--	g17755 = NAND(g5619, g14522, g5630, g9864)
--	g13873 = NAND(g11566, g11729)
--	I31974 = NAND(g33631, I31972)
--	g14947 = NAND(g12785, g10491)
--	g10605 = NAND(g2555, g7490)
--	g12482 = NAND(I15307, I15308)
--	g25470 = NAND(g22457, g2051, g8365)
--	g13834 = NAND(g4754, g11773)
--	g16321 = NAND(g4955, g13996, g12088)
--	g10951 = NAND(g7845, g7868)
--	g28920 = NAND(g27779, g1802, g7315)
--	g24574 = NAND(g22709, g22687)
--	g14234 = NAND(g9177, g11881)
--	g31706 = NAND(I29270, I29271)
--	I18626 = NAND(g2079, I18625)
--	g28946 = NAND(g27907, g2495, g2421)
--	g25467 = NAND(g12432, g22417)
--	g23761 = NAND(I22893, I22894)
--	g23692 = NAND(g9501, g20995)
--	g27380 = NAND(I26071, I26072)
--	g12356 = NAND(g7438, g6012)
--	g9591 = NAND(g1926, g1894)
--	g12999 = NAND(g4392, g10476, g4401)
--	g11320 = NAND(g4633, g4621, g7202)
--	g25984 = NAND(g24567, g22668)
--	g19886 = NAND(g11403, g17794)
--	I15122 = NAND(g9910, I15121)
--	g13346 = NAND(g4854, g11012)
--	g19792 = NAND(I20204, I20205)
--	I14957 = NAND(g6181, I14955)
--	g26053 = NAND(g22875, g24677, g22941)
--	g13464 = NAND(g10831, g4793, g4776)
--	g13797 = NAND(g8102, g11273)
--	g11292 = NAND(I14331, I14332)
--	I32756 = NAND(g34469, g25779)
--	g11153 = NAND(I14205, I14206)
--	g29094 = NAND(g27858, g9700)
--	g12449 = NAND(g7004, g5297, g5352)
--	I14290 = NAND(g8282, I14289)
--	g11409 = NAND(g9842, g3298)
--	I22894 = NAND(g21228, I22892)
--	I14427 = NAND(g8595, g4005)
--	g14829 = NAND(g6621, g12137, g6675, g12471)
--	I31983 = NAND(g33653, g33648)
--	g14434 = NAND(g6415, g11945)
--	g29018 = NAND(g9586, g27742)
--	I12878 = NAND(g4180, I12876)
--	g10946 = NAND(g1489, g7876)
--	g28927 = NAND(g27837, g1906, g7322)
--	g14946 = NAND(g6247, g12173, g6346, g12672)
--	g9750 = NAND(I13335, I13336)
--	I11826 = NAND(g4601, I11824)
--	g14344 = NAND(g5377, g11885)
--	g24583 = NAND(g22753, g22711)
--	I13182 = NAND(g6500, g6505)
--	I17496 = NAND(g1448, I17494)
--	g28903 = NAND(g27800, g2197, g7280)
--	g14682 = NAND(g4933, g11780)
--	g12149 = NAND(g8205, g2185)
--	I14481 = NAND(g10074, I14480)
--	g28755 = NAND(g27742, g7268, g1592)
--	g12148 = NAND(g2060, g8310)
--	g13109 = NAND(g6279, g12173, g6369, g10003)
--	g16772 = NAND(g3558, g13799, g3654, g11576)
--	g24787 = NAND(g3391, g23079)
--	g29001 = NAND(g27937, g2599, g7431)
--	g13108 = NAND(g5551, g12029, g5685, g9864)
--	g12343 = NAND(g7470, g5630)
--	g13283 = NAND(g12440, g12399, g9843)
--	I22801 = NAND(g21434, I22799)
--	g11492 = NAND(g6928, g6941, g8756)
--	g12971 = NAND(g9024, g8977, g10664)
--	I12545 = NAND(g191, I12544)
--	g9528 = NAND(I13183, I13184)
--	g12369 = NAND(g9049, g637)
--	g28395 = NAND(g27074, g13655)
--	I14956 = NAND(g9620, I14955)
--	g11381 = NAND(g9660, g3274)
--	g28899 = NAND(g27833, g14612)
--	I18529 = NAND(g1811, g14640)
--	g28990 = NAND(g27882, g8310)
--	g17220 = NAND(g9369, g9298, g14376)
--	I15174 = NAND(g9977, g2661)
--	g29157 = NAND(g9835, g27937)
--	g17246 = NAND(g9439, g9379, g14405)
--	g12412 = NAND(g10044, g5297, g5348)
--	I26049 = NAND(g25997, g13500)
--	g26382 = NAND(g577, g24953, g12323)
--	g33930 = NAND(g33394, g12767, g9848)
--	g22754 = NAND(g20114, g19376)
--	g33838 = NAND(g33083, g4369)
--	g14927 = NAND(g12695, g10281)
--	g16586 = NAND(g13851, g13823)
--	I22866 = NAND(g21228, I22864)
--	g21345 = NAND(g11429, g17157)
--	g27582 = NAND(g10857, g26131, g26105)
--	g9372 = NAND(g5080, g5084)
--	g28861 = NAND(g27837, g7405, g1906)
--	I20461 = NAND(g17515, I20460)
--	g25476 = NAND(g22472, g2476, g8373)
--	g8359 = NAND(I12545, I12546)
--	g24662 = NAND(g22957, g2955)
--	I24461 = NAND(g23796, g14437)
--	g10604 = NAND(g7424, g7456)
--	g15751 = NAND(g5591, g14522, g5666, g14669)
--	g10755 = NAND(g7352, g7675, g1322, g1404)
--	g24890 = NAND(g13852, g22929)
--	g14755 = NAND(g12593, g12772)
--	g19495 = NAND(g15969, g10841, g7781)
--	g27925 = NAND(I26439, I26440)
--	I22923 = NAND(g21284, I22921)
--	g29660 = NAND(g28448, g9582)
--	g20248 = NAND(g17056, g14146, g14123)
--	g16275 = NAND(g9291, g13480)
--	g14981 = NAND(g12785, g12632)
--	I14211 = NAND(g9252, g9295)
--	g9334 = NAND(g827, g832)
--	g12112 = NAND(g8139, g1624)
--	I17923 = NAND(g13378, g1478)
--	g33306 = NAND(g776, g32212, g11679)
--	g11326 = NAND(g8993, g376, g365, g370)
--	g20081 = NAND(g11325, g17794)
--	g14794 = NAND(g12492, g12772)
--	g14845 = NAND(g12558, g12798)
--	I14497 = NAND(g9020, g8737)
--	I24365 = NAND(g14320, I24363)
--	I13850 = NAND(g862, g7397)
--	g13040 = NAND(g5196, g12002, g5308, g9780)
--	g13948 = NAND(g11610, g8864)
--	g14899 = NAND(g12744, g10421)
--	g29085 = NAND(g9694, g27837)
--	g28997 = NAND(g27903, g8324)
--	g25382 = NAND(g12333, g22342)
--	I12289 = NAND(g1300, I12287)
--	g14898 = NAND(g5901, g12129, g6000, g12614)
--	I32204 = NAND(g33670, I32202)
--	I23950 = NAND(g23162, I23949)
--	g15014 = NAND(g12785, g12680)
--	I12288 = NAND(g1484, I12287)
--	g24380 = NAND(I23601, I23602)
--	g12429 = NAND(g7473, g6675)
--	g14521 = NAND(g12170, g5428)
--	I25221 = NAND(g24718, I25219)
--	g12428 = NAND(g7472, g6358)
--	g28871 = NAND(g27858, g7418, g2331)
--	I17885 = NAND(g1135, I17883)
--	g9908 = NAND(I13453, I13454)
--	g22902 = NAND(g18957, g2848)
--	I16780 = NAND(g12332, I16778)
--	g10573 = NAND(g7992, g8179)
--	g9567 = NAND(g6116, g6120)
--	g14861 = NAND(g12744, g10341)
--	g14573 = NAND(g9506, g12249)
--	g24932 = NAND(g19886, g23172)
--	g15720 = NAND(g5917, g14497, g6019, g9935)
--	g11933 = NAND(g837, g9334, g7197)
--	I14855 = NAND(g5142, I14853)
--	g14045 = NAND(g11571, g11747)
--	g29335 = NAND(g25540, g28131)
--	g13634 = NAND(g11797, g11261)
--	g13851 = NAND(g8224, g11360)
--	g27317 = NAND(g24793, g26255)
--	I12374 = NAND(g3462, I12372)
--	g25215 = NAND(I24384, I24385)
--	g7850 = NAND(g554, g807)
--	g12317 = NAND(g10026, g6486)
--	g29694 = NAND(g28391, g13709)
--	g14098 = NAND(g11566, g8864)
--	g17699 = NAND(I18681, I18682)
--	g25439 = NAND(g22498, g12122)
--	g28911 = NAND(g27907, g7456, g2465)
--	g23972 = NAND(g7097, g20751)
--	g17290 = NAND(g9506, g9449, g14431)
--	I29253 = NAND(g29482, g12017)
--	g29131 = NAND(g27907, g9762)
--	I15213 = NAND(g10035, I15212)
--	I12842 = NAND(g4235, I12840)
--	g25349 = NAND(g22432, g12051)
--	g12245 = NAND(g7344, g5637)
--	g12323 = NAND(g9480, g640)
--	I14714 = NAND(g5128, I14712)
--	g22661 = NAND(g20136, g94)
--	I13730 = NAND(g4534, I13729)
--	g27775 = NAND(g21228, g25262, g26424, g26166)
--	g16236 = NAND(g13573, g13554, g13058)
--	I14257 = NAND(g8154, g3133)
--	g28950 = NAND(g27937, g7490, g2599)
--	I15051 = NAND(g9759, g2259)
--	I14818 = NAND(g6513, I14816)
--	g9724 = NAND(g5092, g5084)
--	g22715 = NAND(g20114, g2999)
--	I23120 = NAND(g417, I23118)
--	g24620 = NAND(g22902, g22874)
--	g14871 = NAND(g6653, g12211, g6661, g12471)
--	I12544 = NAND(g191, g194)
--	g13756 = NAND(g203, g12812)
--	I18680 = NAND(g2638, g14752)
--	g12232 = NAND(g8804, g4878)
--	g16264 = NAND(g518, g9158, g13223)
--	g19875 = NAND(g13667, g16316)
--	I22930 = NAND(g12223, I22929)
--	g26052 = NAND(g22714, g24662, g22921)
--	g26745 = NAND(g6856, g25317)
--	g17572 = NAND(g3598, g13799, g3676, g8542)
--	g11350 = NAND(I14369, I14370)
--	I22965 = NAND(g12288, g21228)
--	I32433 = NAND(g34051, I32431)
--	g24369 = NAND(I23586, I23587)
--	g12512 = NAND(g7766, g10312)
--	g21359 = NAND(g11509, g17157)
--	g13846 = NAND(g1116, g10649)
--	g10472 = NAND(I13851, I13852)
--	g11396 = NAND(g8713, g4688)
--	I12270 = NAND(g1141, I12269)
--	I14735 = NAND(g5475, I14733)
--	g19455 = NAND(g15969, g10841, g7781)
--	g20133 = NAND(g17668, g17634, g17597, g14569)
--	g17297 = NAND(g2729, g14291)
--	g21344 = NAND(g11428, g17157)
--	g11405 = NAND(g2741, g2735, g6856, g2748)
--	g15781 = NAND(g6267, g12173, g6329, g14745)
--	g20011 = NAND(g3731, g16476)
--	g14776 = NAND(g12780, g12622)
--	g28203 = NAND(g12546, g27985, g27977)
--	g10754 = NAND(g7936, g7913, g8411)
--	g29015 = NAND(g27742, g9586)
--	g13929 = NAND(g11669, g11763)
--	I12219 = NAND(g1478, I12217)
--	g25200 = NAND(g5742, g23642)
--	g14825 = NAND(g12806, g12680)
--	g14950 = NAND(g7812, g12632)
--	g11020 = NAND(g9187, g9040)
--	g12080 = NAND(g1917, g8201)
--	g13928 = NAND(g3562, g11238, g3680, g11576)
--	I12218 = NAND(g1437, I12217)
--	g14858 = NAND(g7766, g12515)
--	g19782 = NAND(I20188, I20189)
--	g29556 = NAND(g28349, g13486)
--	g31747 = NAND(I29296, I29297)
--	g14151 = NAND(g11692, g11483)
--	g14996 = NAND(g12662, g10312)
--	g24925 = NAND(g20092, g23154)
--	g24958 = NAND(g21330, g23462)
--	g17520 = NAND(g5260, g12002, g5276, g14631)
--	g12461 = NAND(g7536, g6000)
--	I24364 = NAND(g23687, I24363)
--	g12342 = NAND(g7004, g7018, g10129)
--	I22937 = NAND(g12226, I22936)
--	I26395 = NAND(g14227, I26393)
--	I14923 = NAND(g9558, g5835)
--	g12145 = NAND(g8195, g1760)
--	g11302 = NAND(g9496, g3281)
--	I15105 = NAND(g9780, g5313)
--	I23980 = NAND(g13670, I23978)
--	g24944 = NAND(g21354, g23363)
--	g13105 = NAND(g10671, g7675, g1322, g1404)
--	I16779 = NAND(g11292, I16778)
--	I12470 = NAND(g392, I12468)
--	g9092 = NAND(g3004, g3050)
--	I16778 = NAND(g11292, g12332)
--	g19589 = NAND(g15969, g10841, g10884)
--	I12277 = NAND(g1467, g1472)
--	I13499 = NAND(g232, I13497)
--	I17884 = NAND(g13336, I17883)
--	g15021 = NAND(g12711, g10341)
--	I12075 = NAND(g996, I12074)
--	g27365 = NAND(I26050, I26051)
--	g24802 = NAND(I23970, I23971)
--	g29186 = NAND(g27051, g4507)
--	g29676 = NAND(g28381, g13676)
--	g7690 = NAND(g4669, g4659, g4653)
--	g15726 = NAND(g6263, g14529, g6365, g10003)
--	I13498 = NAND(g255, I13497)
--	g24793 = NAND(g3742, g23124)
--	g26235 = NAND(g8016, g24766)
--	g14058 = NAND(g7121, g11537)
--	I26440 = NAND(g14271, I26438)
--	g28895 = NAND(g27775, g8146)
--	I14885 = NAND(g5489, I14883)
--	g11881 = NAND(g9060, g3361)
--	I14854 = NAND(g9433, I14853)
--	g25400 = NAND(g22472, g12086)
--	g12225 = NAND(g8324, g2453)
--	g14902 = NAND(g7791, g12581)
--	g12471 = NAND(I15288, I15289)
--	I29303 = NAND(g29496, I29302)
--	g12087 = NAND(g7431, g2599)
--	g14120 = NAND(g11780, g4907)
--	g14739 = NAND(g5929, g12067, g5983, g12351)
--	g10738 = NAND(g6961, g10308)
--	I22922 = NAND(g14677, I22921)
--	I25845 = NAND(g26212, g24799)
--	g14146 = NAND(g11020, g691)
--	g32072 = NAND(g31009, g13301)
--	g19466 = NAND(g11562, g17794)
--	I15003 = NAND(g9691, I15002)
--	g12244 = NAND(g7343, g5320)
--	g13248 = NAND(g9985, g12399, g9843)
--	I14480 = NAND(g10074, g655)
--	g28376 = NAND(g27064, g13620)
--	g13779 = NAND(g11804, g11283)
--	I22685 = NAND(g21434, I22683)
--	g27955 = NAND(I26460, I26461)
--	g28980 = NAND(g27933, g14680)
--	I23987 = NAND(g482, I23985)
--	g23719 = NAND(I22845, I22846)
--	I12401 = NAND(g3808, g3813)
--	g28888 = NAND(g27738, g8139)
--	g28824 = NAND(g27779, g7356, g1772)
--	I20488 = NAND(g16757, I20486)
--	I22800 = NAND(g11960, I22799)
--	I22936 = NAND(g12226, g21228)
--	g11356 = NAND(g9552, g3632)
--	g8691 = NAND(g3267, g3310, g3281, g3303)
--	g13945 = NAND(g691, g11740)
--	g19874 = NAND(g13665, g16299, g8163)
--	g17581 = NAND(g5607, g12029, g5623, g14669)
--	g17315 = NAND(g9564, g9516, g14503)
--	g28931 = NAND(g27886, g2070, g1996)
--	I23969 = NAND(g22202, g490)
--	g14547 = NAND(g9439, g12201)
--	g14895 = NAND(g7766, g12571)
--	g11998 = NAND(g8324, g8373)
--	I22762 = NAND(g21434, I22760)
--	g13672 = NAND(g8933, g11261)
--	g12459 = NAND(g7437, g5623)
--	g16663 = NAND(g13854, g13834, g14655, g12292)
--	g10551 = NAND(g1728, g7356)
--	g21388 = NAND(g11608, g17157)
--	g24880 = NAND(g23281, g23266, g22839)
--	g23324 = NAND(g703, g20181)
--	g14572 = NAND(g12169, g9678)
--	I14734 = NAND(g9732, I14733)
--	I20189 = NAND(g1333, I20187)
--	g21272 = NAND(g11268, g17157)
--	I13043 = NAND(g5115, g5120)
--	I14993 = NAND(g6527, I14991)
--	I20188 = NAND(g16272, I20187)
--	g13513 = NAND(g1351, g11815, g8002)
--	g14127 = NAND(g11653, g11435)
--	g21462 = NAND(g17816, g14871, g17779, g14829)
--	g11961 = NAND(g9777, g5105)
--	g12079 = NAND(g1792, g8195)
--	g28860 = NAND(g27775, g14586)
--	g13897 = NAND(g3211, g11217, g3329, g11519)
--	I20460 = NAND(g17515, g14187)
--	I24383 = NAND(g23721, g14347)
--	g12078 = NAND(g8187, g8093)
--	I26071 = NAND(g26026, I26070)
--	I15212 = NAND(g10035, g1714)
--	g14956 = NAND(g12604, g10281)
--	I11879 = NAND(g4430, I11877)
--	g14889 = NAND(g12609, g12824)
--	g16757 = NAND(g13911, g13886, g14120, g11675)
--	I11878 = NAND(g4388, I11877)
--	g28987 = NAND(g27886, g2070, g7411)
--	g25435 = NAND(g22432, g2342, g8316)
--	I23979 = NAND(g23198, I23978)
--	g24989 = NAND(g21345, g23363)
--	g12159 = NAND(g8765, g4864)
--	g12125 = NAND(g9728, g5101)
--	I21978 = NAND(g19620, I21976)
--	I22974 = NAND(g19638, I22972)
--	I23978 = NAND(g23198, g13670)
--	g24988 = NAND(g546, g23088)
--	g24924 = NAND(g20007, g23172)
--	I15149 = NAND(g5659, I15147)
--	g21360 = NAND(g11510, g17157)
--	I23986 = NAND(g22182, I23985)
--	g27295 = NAND(g24776, g26208)
--	g20271 = NAND(g16925, g14054, g16657, g16628)
--	g11149 = NAND(g1564, g7948)
--	I15148 = NAND(g9864, I15147)
--	g28969 = NAND(g27854, g8267)
--	I26367 = NAND(g26400, I26366)
--	I26394 = NAND(g26488, I26393)
--	g12144 = NAND(I15003, I15004)
--	g9543 = NAND(g2217, g2185)
--	g13097 = NAND(g5204, g12002, g5339, g9780)
--	g10520 = NAND(g7195, g7115)
--	g13104 = NAND(g1404, g10794)
--	g12336 = NAND(I15175, I15176)
--	g14520 = NAND(g9369, g12163)
--	I14187 = NAND(g3470, I14185)
--	g7150 = NAND(g5016, g5062)
--	I25220 = NAND(g482, I25219)
--	g20199 = NAND(g16815, g13968, g16749, g13907)
--	g11971 = NAND(g8249, g8302)
--	g28870 = NAND(g27796, g14588)
--	g34048 = NAND(g33669, g10583, g7442)
--	I13079 = NAND(g5467, I13077)
--	I13444 = NAND(g239, I13442)
--	I32432 = NAND(g34056, I32431)
--	g14546 = NAND(g12125, g9613)
--	g14089 = NAND(g11755, g4717)
--	g22688 = NAND(g20219, g2936)
--	g20198 = NAND(g16813, g13958, g16745, g13927)
--	g17706 = NAND(g3921, g11255, g3983, g13933)
--	g17597 = NAND(g3191, g13700, g3303, g8481)
--	I12074 = NAND(g996, g979)
--	I13078 = NAND(g5462, I13077)
--	g14088 = NAND(g3901, g11255, g4000, g11631)
--	g14024 = NAND(g7121, g11763)
--	g17689 = NAND(g6645, g12137, g6661, g14786)
--	I18589 = NAND(g14679, I18587)
--	g24528 = NAND(g4098, g22654)
--	g17624 = NAND(I18588, I18589)
--	g28867 = NAND(g27800, g2227, g2153)
--	I18588 = NAND(g2370, I18587)
--	g7836 = NAND(g4653, g4688)
--	I20467 = NAND(g16663, g16728)
--	I14169 = NAND(g8389, g3119)
--	I14884 = NAND(g9500, I14883)
--	g11412 = NAND(g8666, g6918, g8697)
--	g15702 = NAND(g13066, g7293)
--	g13850 = NAND(g11279, g8396)
--	g15904 = NAND(I17380, I17381)
--	g25049 = NAND(g21344, g23462)
--	g12289 = NAND(g9978, g9766, g9708)
--	g14659 = NAND(g12646, g12443)
--	g14625 = NAND(g3897, g11225, g4031, g8595)
--	g14987 = NAND(g6593, g12211, g6692, g12721)
--	g20161 = NAND(g17732, g17706, g17670, g14625)
--	g22885 = NAND(g9104, g20154)
--	g12023 = NAND(g2453, g8373)
--	g28910 = NAND(g27854, g14614)
--	g13896 = NAND(g3227, g11194, g3281, g11350)
--	I23917 = NAND(g23975, g9333)
--	g25048 = NAND(g542, g23088)
--	g12224 = NAND(I15088, I15089)
--	g14943 = NAND(g7791, g12622)
--	I13336 = NAND(g1691, I13334)
--	g27687 = NAND(g25200, g26714)
--	g14968 = NAND(g12739, g10312)
--	g11959 = NAND(g8316, g2342)
--	g13627 = NAND(g11172, g8388)
--	I22684 = NAND(g11893, I22683)
--	I20167 = NAND(g990, I20165)
--	g14855 = NAND(g12700, g12824)
--	I12729 = NAND(g4291, I12728)
--	g13050 = NAND(g5543, g12029, g5654, g9864)
--	g13958 = NAND(g3610, g11238, g3618, g11389)
--	I12728 = NAND(g4291, g4287)
--	g28877 = NAND(g27937, g7490, g7431)
--	g20068 = NAND(g11293, g17794)
--	I26366 = NAND(g26400, g14211)
--	I14531 = NAND(g8840, I14530)
--	g13742 = NAND(g11780, g11283)
--	g11944 = NAND(I14765, I14766)
--	g7620 = NAND(I12097, I12098)
--	g8010 = NAND(I12345, I12346)
--	I14186 = NAND(g8442, I14185)
--	g17287 = NAND(g7262, g14228)
--	g12195 = NAND(g2619, g8381)
--	g17596 = NAND(g8686, g14367)
--	g25514 = NAND(g12540, g22498)
--	g24792 = NAND(I23950, I23951)
--	g17243 = NAND(g7247, g14212)
--	g12525 = NAND(g7522, g6668)
--	g12016 = NAND(g1648, g8093)
--	g23281 = NAND(g18957, g2898)
--	g21301 = NAND(g11371, g17157)
--	g21377 = NAND(g11560, g17157)
--	g14055 = NAND(g11697, g11763)
--	g17773 = NAND(g5965, g14549, g5976, g9935)
--	I18485 = NAND(g1677, g14611)
--	g14978 = NAND(g12716, g10491)
--	g15780 = NAND(g5937, g14549, g6012, g14701)
--	I17475 = NAND(g13336, I17474)
--	g14590 = NAND(g3546, g11207, g3680, g8542)
--	g24918 = NAND(g136, g23088)
--	g17670 = NAND(g3893, g13772, g4005, g8595)
--	g22839 = NAND(g20114, g2988)
--	g23699 = NAND(g21012, g11160)
--	I29302 = NAND(g29496, g12121)
--	g25473 = NAND(g12437, g22432)
--	g14741 = NAND(g12711, g10421)
--	g27705 = NAND(g25237, g26782)
--	g22838 = NAND(g20219, g2960)
--	g17734 = NAND(g5272, g14490, g5283, g9780)
--	g28923 = NAND(g27775, g8195)
--	g16282 = NAND(g4933, g13939, g12088)
--	g9442 = NAND(g5424, g5428)
--	g27679 = NAND(g25186, g26685)
--	I15129 = NAND(g9914, I15128)
--	g12042 = NAND(g9086, g703)
--	I15002 = NAND(g9691, g1700)
--	I26095 = NAND(g13539, I26093)
--	g12255 = NAND(g9958, g6140)
--	g11002 = NAND(g7475, g862)
--	I15128 = NAND(g9914, g2527)
--	g13057 = NAND(g969, g11294)
--	g14735 = NAND(g12739, g12571)
--	g12188 = NAND(g8249, g1894)
--	g12124 = NAND(g8741, g4674)
--	I13392 = NAND(g1825, I13390)
--	g11245 = NAND(g7636, g7733, g7697)
--	I15299 = NAND(g10112, I15298)
--	g12460 = NAND(g10093, g5644, g5694)
--	g12686 = NAND(g7097, g6682, g6736)
--	I20166 = NAND(g16246, I20165)
--	g11323 = NAND(I14351, I14352)
--	g14695 = NAND(g5583, g12029, g5637, g12301)
--	g14018 = NAND(g10323, g11483)
--	I15298 = NAND(g10112, g1982)
--	g11533 = NAND(g6905, g3639, g3698)
--	g21403 = NAND(g11652, g17157)
--	g20783 = NAND(g14616, g17225)
--	g12294 = NAND(g10044, g7018, g10090)
--	g17618 = NAND(I18580, I18581)
--	g28885 = NAND(g27742, g1668, g7268)
--	g22306 = NAND(g4584, g4616, g13202, g19071)
--	I22873 = NAND(g21228, I22871)
--	I11865 = NAND(g4434, I11864)
--	I14230 = NAND(g8055, I14228)
--	g17468 = NAND(g3215, g13700, g3317, g8481)
--	I21993 = NAND(g7670, I21992)
--	g15787 = NAND(g6283, g14575, g6358, g14745)
--	g14706 = NAND(g6287, g12101, g6369, g12672)
--	I14992 = NAND(g9685, I14991)
--	g21385 = NAND(g17736, g14696, g17679, g14636)
--	I14510 = NAND(g8721, I14508)
--	g15743 = NAND(g5893, g14497, g6005, g9935)
--	g21354 = NAND(g11468, g17157)
--	g14688 = NAND(g12604, g12453)
--	g28287 = NAND(g10504, g26131, g26973)
--	g12915 = NAND(g12806, g12632)
--	I13383 = NAND(g269, I13382)
--	g11445 = NAND(g9771, g3976)
--	g14157 = NAND(g11715, g11763)
--	g22666 = NAND(g18957, g2878)
--	g13499 = NAND(g11479, g11442, g11410, g11382)
--	I13065 = NAND(g4308, g4304)
--	g14066 = NAND(g11514, g11473)
--	g13498 = NAND(g12577, g12522, g12462, g12416)
--	I15080 = NAND(g1968, I15078)
--	g17363 = NAND(g8635, g14367)
--	g28942 = NAND(g27858, g2331, g7335)
--	g17217 = NAND(g7239, g14194)
--	g21190 = NAND(g6077, g17420)
--	g14876 = NAND(g12492, g12443)
--	g14885 = NAND(g12651, g12505)
--	g14854 = NAND(g5555, g12093, g5654, g12563)
--	g10511 = NAND(g4628, g7202, g4621)
--	g11432 = NAND(g10295, g8864)
--	I23601 = NAND(g22360, I23600)
--	g13432 = NAND(g4793, g10831)
--	I14275 = NAND(g8218, g3484)
--	g12155 = NAND(g7753, g7717)
--	g12822 = NAND(g6978, g7236, g7224, g7163)
--	g15027 = NAND(g12667, g10341)
--	I15342 = NAND(g2541, I15340)
--	g28930 = NAND(g27833, g8201)
--	I24439 = NAND(g23771, I24438)
--	g28965 = NAND(g27882, g8255)
--	g30573 = NAND(g29355, g19666)
--	I24438 = NAND(g23771, g14411)
--	g15710 = NAND(g319, g13385)
--	g9715 = NAND(g5011, g4836)
--	g28131 = NAND(g27051, g25838)
--	g31509 = NAND(g599, g29933, g12323)
--	g10916 = NAND(g1146, g7854)
--	I12241 = NAND(g1111, I12240)
--	g33933 = NAND(g33394, g12491, g12819, g12796)
--	g12589 = NAND(g7591, g6692)
--	g12194 = NAND(g8373, g8273)
--	g10550 = NAND(g7268, g7308)
--	g13529 = NAND(g11590, g11544, g11492, g11446)
--	I14517 = NAND(g10147, I14516)
--	g12588 = NAND(g10169, g6336, g6386)
--	g27401 = NAND(I26094, I26095)
--	g12524 = NAND(g7074, g7087, g10212)
--	g23659 = NAND(g9434, g20854)
--	g11330 = NAND(g9483, g1193)
--	g13528 = NAND(g11294, g7549, g1008)
--	g13330 = NAND(g4664, g11006)
--	g10307 = NAND(I13730, I13731)
--	I15365 = NAND(g2675, I15363)
--	g14085 = NAND(g7121, g11584)
--	g17740 = NAND(g5945, g14497, g6012, g12351)
--	g13764 = NAND(g11252, g3072)
--	g8238 = NAND(I12469, I12470)
--	g14596 = NAND(g12196, g9775, g12124, g9663)
--	g12119 = NAND(g2351, g8267)
--	g14054 = NAND(g3550, g11238, g3649, g11576)
--	I22711 = NAND(g11915, I22710)
--	g7701 = NAND(g4859, g4849, g4843)
--	g21339 = NAND(g15725, g13084, g15713, g13050)
--	g13960 = NAND(g11669, g11537)
--	g32057 = NAND(g31003, g13297)
--	g12118 = NAND(g8259, g8150)
--	g12022 = NAND(g7335, g2331)
--	g21338 = NAND(g15741, g15734, g15728, g13097)
--	I26070 = NAND(g26026, g13517)
--	I17474 = NAND(g13336, g1105)
--	g16723 = NAND(g3606, g13730, g3676, g11576)
--	g14773 = NAND(g12711, g12581)
--	g24544 = NAND(g22666, g22661, g22651)
--	g13709 = NAND(g11755, g11261)
--	g25389 = NAND(g22457, g12082)
--	g12285 = NAND(I15122, I15123)
--	I15087 = NAND(g9832, g2393)
--	g14655 = NAND(g4743, g11755)
--	g11708 = NAND(g10147, g10110)
--	g13708 = NAND(g11200, g8507)
--	g12053 = NAND(g2587, g8418)
--	g16097 = NAND(g13319, g10998)
--	I26094 = NAND(g26055, I26093)
--	I24415 = NAND(g23751, I24414)
--	I15043 = NAND(g1834, I15041)
--	g13043 = NAND(g10521, g969)
--	g14930 = NAND(g12609, g12515)
--	g14993 = NAND(g12695, g12453)
--	I17381 = NAND(g1129, I17379)
--	g24678 = NAND(g22994, g23010)
--	g14838 = NAND(g12492, g12405)
--	g14965 = NAND(g12609, g12571)
--	g22908 = NAND(g9104, g20175)
--	g13069 = NAND(g5889, g12067, g6000, g9935)
--	g29702 = NAND(g28395, g13712)
--	g34162 = NAND(g785, g33823, g11679)
--	g15717 = NAND(g10754, g13092)
--	I13401 = NAND(g2246, g2250)
--	g11955 = NAND(g8302, g1917)
--	g13955 = NAND(g11621, g11527)
--	g11970 = NAND(g1760, g8241)
--	g28410 = NAND(g27074, g13679)
--	g19962 = NAND(g11470, g17794)
--	g10618 = NAND(g10153, g9913)
--	I14351 = NAND(g8890, I14350)
--	g27693 = NAND(g25216, g26752)
--	I11864 = NAND(g4434, g4401)
--	g34220 = NAND(I32186, I32187)
--	g28363 = NAND(g27064, g13593)
--	g17568 = NAND(I18486, I18487)
--	g14279 = NAND(g12111, g9246)
--	g7887 = NAND(I12278, I12279)
--	I13749 = NAND(g4608, g4584)
--	g13886 = NAND(g11804, g4922)
--	g7228 = NAND(g6398, g6444)
--	g11994 = NAND(g8310, g8365)
--	g15723 = NAND(g10775, g13104)
--	g23978 = NAND(g572, g21389, g12323)
--	g13967 = NAND(g3929, g11225, g3983, g11419)
--	I12345 = NAND(g3106, I12344)
--	I14790 = NAND(g6167, I14788)
--	I14516 = NAND(g10147, g661)
--	g23590 = NAND(g20682, g11111)
--	I12849 = NAND(g4281, I12848)
--	g12008 = NAND(g9932, g5798)
--	g17814 = NAND(g5579, g14522, g5673, g12563)
--	g22638 = NAND(g18957, g2886)
--	I12848 = NAND(g4281, g4277)
--	g12476 = NAND(g7498, g6704)
--	g13459 = NAND(g7479, g11294, g11846)
--	g21384 = NAND(g17734, g14686, g17675, g14663)
--	I23587 = NAND(g4332, I23585)
--	g8889 = NAND(g3684, g4871)
--	g14038 = NAND(g11514, g11435)
--	g23067 = NAND(g20887, g10721)
--	g10601 = NAND(g896, g7397)
--	g13918 = NAND(g3259, g11217, g3267, g11350)
--	g16925 = NAND(g3574, g13799, g3668, g11576)
--	g14601 = NAND(g12318, g6466)
--	I18538 = NAND(g14642, I18536)
--	g8871 = NAND(I12841, I12842)
--	I15079 = NAND(g9827, I15078)
--	g14677 = NAND(I16779, I16780)
--	I12263 = NAND(g1448, I12261)
--	g11545 = NAND(I14498, I14499)
--	g11444 = NAND(g6905, g6918, g8733)
--	g13079 = NAND(g1312, g11336)
--	I15078 = NAND(g9827, g1968)
--	g12239 = NAND(I15106, I15107)
--	g20201 = NAND(I20468, I20469)
--	g8500 = NAND(g3431, g3423)
--	g14937 = NAND(g12667, g10421)
--	g26025 = NAND(g22405, g24631)
--	g13086 = NAND(g6235, g12101, g6346, g10003)
--	g16681 = NAND(I17884, I17885)
--	g17578 = NAND(g5212, g14399, g5283, g12497)
--	g12941 = NAND(g7167, g10537)
--	g19795 = NAND(g13600, g16275)
--	g12185 = NAND(g9905, g799)
--	g21402 = NAND(g17757, g14740, g17716, g14674)
--	g17586 = NAND(g14638, g14601)
--	g11977 = NAND(g8373, g2476)
--	g13977 = NAND(g11610, g11729)
--	I14530 = NAND(g8840, g8873)
--	g8737 = NAND(I12729, I12730)
--	g15011 = NAND(g12716, g12632)
--	g34227 = NAND(I32203, I32204)
--	g14015 = NAND(g11658, g11747)
--	g11561 = NAND(I14517, I14518)
--	g25172 = NAND(g5052, g23560)
--	I22872 = NAND(g12150, I22871)
--	g25996 = NAND(g24601, g22838)
--	g20170 = NAND(g16741, g13897, g16687, g13866)
--	g10556 = NAND(g7971, g8133)
--	g13823 = NAND(g11313, g3774)
--	I13454 = NAND(g1959, I13452)
--	I21992 = NAND(g7670, g19638)
--	g14223 = NAND(g9092, g11858)
--	g17493 = NAND(g8659, g14367)
--	g15959 = NAND(I17405, I17406)
--	g27577 = NAND(g25019, g25002, g24988, g25765)
--	I15364 = NAND(g10182, I15363)
--	g12577 = NAND(g7051, g5990, g6044)
--	g14110 = NAND(g11692, g8906)
--	g9246 = NAND(g847, g812)
--	g15742 = NAND(g5575, g12093, g5637, g14669)
--	I23586 = NAND(g22409, I23585)
--	g9203 = NAND(g3706, g3752)
--	g14740 = NAND(g5913, g12129, g6031, g12614)
--	I13382 = NAND(g269, g246)
--	I15289 = NAND(g6697, I15287)
--	g19358 = NAND(g15723, g1399)
--	I13519 = NAND(g2514, I13518)
--	g16299 = NAND(g8160, g8112, g13706)
--	g31003 = NAND(g27163, g29497, g19644)
--	g14953 = NAND(g12646, g12405)
--	I15288 = NAND(g10061, I15287)
--	I13518 = NAND(g2514, g2518)
--	g12083 = NAND(g2217, g8205)
--	I15308 = NAND(g2407, I15306)
--	g11224 = NAND(I14290, I14291)
--	g13288 = NAND(g10946, g1442)
--	g15730 = NAND(g6609, g14556, g6711, g10061)
--	g14800 = NAND(g7704, g12443)
--	I24414 = NAND(g23751, g14382)
--	g29046 = NAND(g27779, g9640)
--	g13495 = NAND(g1008, g11786, g7972)
--	I29261 = NAND(g29485, g12046)
--	g24809 = NAND(g19965, g23132)
--	I22846 = NAND(g21228, I22844)
--	g24808 = NAND(I23986, I23987)
--	I13729 = NAND(g4534, g4537)
--	g10587 = NAND(g2421, g7456)
--	g11374 = NAND(g9536, g1536)
--	g28391 = NAND(g27064, g13637)
--	g12415 = NAND(g7496, g5976)
--	g21287 = NAND(g14616, g17571)
--	g19506 = NAND(g4087, g15825)
--	g10909 = NAND(g7304, g1116)
--	g20733 = NAND(g14406, g17290, g9509)
--	g21307 = NAND(g15719, g13067, g15709, g13040)
--	g15002 = NAND(g12609, g10312)
--	I25243 = NAND(g490, I25242)
--	g13260 = NAND(g1116, g10666)
--	g14908 = NAND(g7812, g10491)
--	g10569 = NAND(g2287, g7418)
--	I22929 = NAND(g12223, g21228)
--	I15195 = NAND(g6005, I15193)
--	I17405 = NAND(g13378, I17404)
--	I12344 = NAND(g3106, g3111)
--	g14569 = NAND(g3195, g11194, g3329, g8481)
--	g11489 = NAND(g9661, g3618)
--	g10568 = NAND(g7328, g7374)
--	g25895 = NAND(g1259, g24453)
--	g16316 = NAND(g9429, g13518)
--	g11559 = NAND(I14509, I14510)
--	g11424 = NAND(g9662, g4012)
--	I13566 = NAND(g2652, I13564)
--	g23655 = NAND(I22793, I22794)
--	I29271 = NAND(g12050, I29269)
--	g9883 = NAND(g5782, g5774)
--	g14123 = NAND(g10685, g10928)
--	g15737 = NAND(g13240, g13115, g7903, g13210)
--	g14807 = NAND(g7738, g12453)
--	g19903 = NAND(g13707, g16319, g8227)
--	g12115 = NAND(g1926, g8249)
--	g14974 = NAND(g12744, g12622)
--	g17790 = NAND(g6311, g14575, g6322, g10003)
--	g17137 = NAND(g13727, g13511, g13527)
--	I13139 = NAND(g6154, g6159)
--	g11544 = NAND(g8700, g3990, g4045)
--	g13544 = NAND(g7972, g10521, g7549, g1008)
--	g24570 = NAND(g22957, g2941)
--	g12052 = NAND(g7387, g2465)
--	g14638 = NAND(g9626, g12361)
--	I15042 = NAND(g9752, I15041)
--	I15255 = NAND(g1848, I15253)
--	I13852 = NAND(g7397, I13850)
--	g14841 = NAND(g12593, g12443)
--	g25385 = NAND(g22369, g1783, g8241)
--	g24567 = NAND(g22957, g2917)
--	g11189 = NAND(I14248, I14249)
--	g11679 = NAND(g8836, g802)
--	I23600 = NAND(g22360, g4322)
--	g29778 = NAND(g294, g28444, g23204)
--	g13124 = NAND(g10666, g7661, g979, g1061)
--	g25888 = NAND(g914, g24439)
--	g31971 = NAND(g30573, g10511)
--	g23210 = NAND(g18957, g2882)
--	g16696 = NAND(g13871, g13855, g14682, g12340)
--	g20185 = NAND(g16772, g13928, g16723, g13882)
--	g10578 = NAND(g7174, g6058)
--	g20675 = NAND(g14377, g17246, g9442)
--	g20092 = NAND(g11373, g17794)
--	g14014 = NAND(g3199, g11217, g3298, g11519)
--	g11938 = NAND(g8259, g2208)
--	g10586 = NAND(g7380, g7418)
--	g13093 = NAND(g10649, g7661, g979, g1061)
--	g8873 = NAND(I12849, I12850)
--	g8632 = NAND(g1514, g1500)
--	g9538 = NAND(g1792, g1760)
--	I20221 = NAND(g16272, g11170)
--	I12240 = NAND(g1111, g1105)
--	g9509 = NAND(g5770, g5774)
--	g23286 = NAND(g6875, g20887)
--	g25426 = NAND(g12371, g22369)
--	g29672 = NAND(g28376, g13672)
--	g17593 = NAND(I18537, I18538)
--	g14116 = NAND(g11697, g11584)
--	I32185 = NAND(g33665, g33661)
--	I14509 = NAND(g370, I14508)
--	g10041 = NAND(I13565, I13566)
--	g14720 = NAND(g12593, g10266)
--	I32518 = NAND(g34422, I32516)
--	g16259 = NAND(g4743, g13908, g12054)
--	I14508 = NAND(g370, g8721)
--	g16225 = NAND(g13544, g13528, g13043)
--	g14041 = NAND(g11610, g11473)
--	g21187 = NAND(g14616, g17364)
--	I22710 = NAND(g11915, g21434)
--	g12207 = NAND(g9887, g5794)
--	g23975 = NAND(I23119, I23120)
--	g12539 = NAND(I15341, I15342)
--	I24463 = NAND(g14437, I24461)
--	g15753 = NAND(g6239, g14529, g6351, g10003)
--	g12538 = NAND(I15334, I15335)
--	I12262 = NAND(g1454, I12261)
--	I13184 = NAND(g6505, I13182)
--	I14213 = NAND(g9295, I14211)
--	g15736 = NAND(g6295, g14575, g6373, g10003)
--	g17635 = NAND(g3542, g13730, g3654, g8542)
--	g16069 = NAND(I17447, I17448)
--	g13915 = NAND(g11566, g11473)
--	I22945 = NAND(g9492, I22944)
--	g14142 = NAND(g11715, g8958)
--	g33925 = NAND(g33394, g4462, g4467)
--	g16657 = NAND(g3554, g13730, g3625, g11576)
--	I14205 = NAND(g8508, I14204)
--	g15843 = NAND(g7922, g7503, g13264)
--	g14517 = NAND(g3231, g11217, g3321, g8481)
--	g24906 = NAND(g8743, g23088)
--	g26714 = NAND(g9316, g25175)
--	g23666 = NAND(g20875, g11139)
--	I26417 = NAND(g26519, g14247)
--	g21363 = NAND(g17708, g14664, g17640, g14598)
--	I32439 = NAND(g34227, g34220)
--	g12100 = NAND(I14956, I14957)
--	I17380 = NAND(g13336, I17379)
--	g24566 = NAND(g22755, g22713)
--	g22711 = NAND(g19581, g7888)
--	g14130 = NAND(g11621, g8906)
--	I18682 = NAND(g14752, I18680)
--	g17474 = NAND(g14547, g14521)
--	g28516 = NAND(g10857, g26105, g27155)
--	g11419 = NAND(I14428, I14429)
--	g29097 = NAND(g9700, g27858)
--	g15709 = NAND(g5224, g14399, g5327, g9780)
--	g27882 = NAND(g21228, g25307, g26424, g26213)
--	g11155 = NAND(g4776, g7892, g9030)
--	I14350 = NAND(g8890, g8848)
--	g15708 = NAND(g7340, g13083)
--	g12414 = NAND(g7028, g7041, g10165)
--	g13822 = NAND(g8160, g11306)
--	g13266 = NAND(g12440, g9920, g9843)
--	g25527 = NAND(g21294, g23462)
--	I12098 = NAND(g1322, I12096)
--	g14727 = NAND(g12604, g12505)
--	I12251 = NAND(g1124, g1129)
--	I22717 = NAND(g11916, g21434)
--	g17492 = NAND(g8655, g14367)
--	I17448 = NAND(g956, I17446)
--	I15167 = NAND(g9904, I15166)
--	I15194 = NAND(g9935, I15193)
--	I17404 = NAND(g13378, g1472)
--	I31985 = NAND(g33648, I31983)
--	g21186 = NAND(g14616, g17363)
--	g23685 = NAND(I22823, I22824)
--	g7223 = NAND(I11878, I11879)
--	g14600 = NAND(g9564, g12311)
--	g14781 = NAND(g6259, g12173, g6377, g12672)
--	g24576 = NAND(g22957, g2902)
--	g13119 = NAND(g6625, g12211, g6715, g10061)
--	g21417 = NAND(g11677, g17157)
--	g11118 = NAND(I14170, I14171)
--	g12114 = NAND(g8241, g8146)
--	g13118 = NAND(g5897, g12067, g6031, g9935)
--	g21334 = NAND(g14616, g17596)
--	g24609 = NAND(g22850, g22650)
--	g20200 = NAND(I20461, I20462)
--	I29295 = NAND(g29495, g12117)
--	g22663 = NAND(I21977, I21978)
--	g33299 = NAND(g608, g32296, g12323)
--	g23762 = NAND(I22900, I22901)
--	I15053 = NAND(g2259, I15051)
--	I15254 = NAND(g10078, I15253)
--	g27141 = NAND(I25846, I25847)
--	I25909 = NAND(g24782, I25907)
--	g24798 = NAND(I23962, I23963)
--	g14422 = NAND(g3187, g11194, g3298, g8481)
--	g24973 = NAND(g21272, g23462)
--	g20184 = NAND(g16770, g13918, g16719, g13896)
--	g23909 = NAND(g7028, g20739)
--	I25908 = NAND(g26256, I25907)
--	g22757 = NAND(g20114, g7891)
--	g12332 = NAND(I15167, I15168)
--	g25019 = NAND(g20055, g23172)
--	g25018 = NAND(g20107, g23154)
--	I18633 = NAND(g2504, g14713)
--	g14542 = NAND(g3582, g11238, g3672, g8542)
--	g14021 = NAND(g11697, g8958)
--	g24934 = NAND(g21283, g23462)
--	I25242 = NAND(g490, g24744)
--	g17757 = NAND(g5909, g14549, g6005, g12614)
--	g10726 = NAND(g7304, g7661, g979, g1061)
--	g23747 = NAND(I22865, I22866)
--	g10614 = NAND(g9024, g8977, g8928)
--	g27833 = NAND(g21228, g25282, g26424, g26190)
--	g12049 = NAND(g2208, g8150)
--	g10905 = NAND(g1116, g7304)
--	I15166 = NAND(g9904, g9823)
--	g14905 = NAND(g12785, g7142)
--	g12048 = NAND(g7369, g2040)
--	g20214 = NAND(g16854, g13993, g16776, g13967)
--	g28109 = NAND(g27051, g25783)
--	g12221 = NAND(I15079, I15080)
--	g27613 = NAND(g24942, g24933, g25048, g26871)
--	g11892 = NAND(g7777, g9086)
--	g13892 = NAND(g11653, g11473)
--	g13476 = NAND(g7503, g11336, g11869)
--	g21416 = NAND(g17775, g14781, g17744, g14706)
--	I13141 = NAND(g6159, I13139)
--	I14249 = NAND(g8091, I14247)
--	I17379 = NAND(g13336, g1129)
--	I17925 = NAND(g1478, I17923)
--	I23949 = NAND(g23162, g13603)
--	g14797 = NAND(g12593, g12405)
--	g27273 = NAND(g10504, g26131, g26105)
--	I14482 = NAND(g655, I14480)
--	g16687 = NAND(g3255, g13700, g3325, g11519)
--	g13712 = NAND(g8984, g11283)
--	g17634 = NAND(g3219, g11217, g3281, g13877)
--	g11914 = NAND(g8187, g1648)
--	g17872 = NAND(g6617, g14602, g6711, g12721)
--	g12947 = NAND(g7184, g10561)
--	I14248 = NAND(g1322, I14247)
--	I22944 = NAND(g9492, g19620)
--	g8728 = NAND(g3618, g3661, g3632, g3654)
--	I14204 = NAND(g8508, g3821)
--	g25300 = NAND(g22369, g12018)
--	g27463 = NAND(g287, g26330, g23204)
--	g13907 = NAND(g3941, g11225, g4023, g11631)
--	g28381 = NAND(g27074, g13621)
--	g29057 = NAND(g27800, g9649)
--	g12463 = NAND(g7513, g6322)
--	g14136 = NAND(g11571, g8906)
--	g14408 = NAND(g6069, g11924)
--	g12972 = NAND(g7209, g10578)
--	g28174 = NAND(g1270, g27059)
--	g28796 = NAND(g27858, g7418, g7335)
--	g31753 = NAND(I29314, I29315)
--	I22793 = NAND(g11956, I22792)
--	g16260 = NAND(g4888, g13910, g12088)
--	g7823 = NAND(I12218, I12219)
--	g28840 = NAND(g27858, g7380, g2287)
--	g11382 = NAND(g8644, g6895, g8663)
--	I15176 = NAND(g2661, I15174)
--	I12203 = NAND(g1094, g1135)
--	g19632 = NAND(g1413, g1542, g16047)
--	I24440 = NAND(g14411, I24438)
--	g11675 = NAND(g8984, g4912)
--	g13176 = NAND(g10715, g7675, g1322, g1404)
--	g13092 = NAND(g1061, g10761)
--	g26269 = NAND(I25243, I25244)
--	g34550 = NAND(g626, g34359, g12323)
--	g11154 = NAND(I14212, I14213)
--	g29737 = NAND(g28421, g13779)
--	g28522 = NAND(g10857, g26131, g27142)
--	g8678 = NAND(g376, g358)
--	g17592 = NAND(I18530, I18531)
--	g16893 = NAND(g10685, g13252, g703)
--	g10537 = NAND(g7138, g5366)
--	I14331 = NAND(g225, I14330)
--	g8105 = NAND(g3068, g3072)
--	I31984 = NAND(g33653, I31983)
--	g16713 = NAND(I17924, I17925)
--	I20462 = NAND(g14187, I20460)
--	I29255 = NAND(g12017, I29253)
--	I24462 = NAND(g23796, I24461)
--	g17820 = NAND(g5925, g14549, g6019, g12614)
--	g31709 = NAND(I29285, I29286)
--	g15752 = NAND(g5921, g12129, g5983, g14701)
--	I29270 = NAND(g29486, I29269)
--	g28949 = NAND(g27903, g14643)
--	I13463 = NAND(g2380, I13462)
--	g31708 = NAND(I29278, I29279)
--	g17846 = NAND(g6271, g14575, g6365, g12672)
--	g17396 = NAND(g7345, g14272)
--	g14750 = NAND(g6633, g12137, g6715, g12721)
--	g24584 = NAND(g22852, g22836, g22715)
--	I14212 = NAND(g9252, I14211)
--	g7167 = NAND(g5360, g5406)
--	g10796 = NAND(g7537, g7523)
--	g20107 = NAND(g11404, g17794)
--	g11906 = NAND(I14713, I14714)
--	I12403 = NAND(g3813, I12401)
--	g16093 = NAND(I17461, I17462)
--	g12344 = NAND(g10093, g7041, g10130)
--	g13083 = NAND(g4392, g10590, g4434)
--	I32441 = NAND(g34220, I32439)
--	g13284 = NAND(g10695, g1157)
--	g7549 = NAND(g1018, g1030)
--	g25341 = NAND(g22417, g12047)
--	g29722 = NAND(g28410, g13742)
--	g25268 = NAND(g21124, g23692)
--	g16875 = NAND(g3223, g13765, g3317, g11519)
--	g7598 = NAND(I12075, I12076)
--	I32758 = NAND(g25779, I32756)
--	g14663 = NAND(g5236, g12002, g5290, g12239)
--	g24804 = NAND(g19916, g23105)
--	g24652 = NAND(g22712, g22940, g22757)
--	g13139 = NAND(g6589, g12137, g6723, g10061)
--	g15713 = NAND(g5571, g14425, g5673, g9864)
--	I14369 = NAND(g8481, I14368)
--	g34469 = NAND(I32517, I32518)
--	I15333 = NAND(g10152, g2116)
--	g19546 = NAND(g15969, g10841, g10884)
--	g8227 = NAND(g3770, g3774)
--	I14368 = NAND(g8481, g3303)
--	g12028 = NAND(I14884, I14885)
--	g15042 = NAND(g12806, g10491)
--	g21253 = NAND(g6423, g17482)
--	I29277 = NAND(g29488, g12081)
--	g23781 = NAND(I22937, I22938)
--	g13963 = NAND(g11715, g11584)
--	g17640 = NAND(g5264, g14399, g5335, g12497)
--	I14229 = NAND(g979, I14228)
--	g21351 = NAND(g15729, g13098, g15720, g13069)
--	g26666 = NAND(g9229, g25144)
--	I14228 = NAND(g979, g8055)
--	g15030 = NAND(g12716, g12680)
--	g27903 = NAND(g21228, g25316, g26424, g26218)
--	g13554 = NAND(g11336, g7582, g1351)
--	I17924 = NAND(g13378, I17923)
--	g12491 = NAND(g7285, g4462, g6961)
--	g28780 = NAND(g27742, g7308, g1636)
--	I22753 = NAND(g11937, g21434)
--	g11312 = NAND(g8565, g3794)
--	g11200 = NAND(g8592, g3798)
--	g25038 = NAND(g21331, g23363)
--	g13115 = NAND(g1008, g11786, g11294)
--	I15052 = NAND(g9759, I15051)
--	g14933 = NAND(g12700, g12571)
--	I14925 = NAND(g5835, I14923)
--	g16155 = NAND(I17495, I17496)
--	g17662 = NAND(I18634, I18635)
--	g28820 = NAND(g27742, g1668, g1592)
--	I12546 = NAND(g194, I12544)
--	I17461 = NAND(g13378, I17460)
--	g14851 = NAND(g7738, g12505)
--	g27767 = NAND(I26367, I26368)
--	g9775 = NAND(g4831, g4681)
--	g20371 = NAND(g16956, g14088, g16694, g16660)
--	g24951 = NAND(g199, g23088)
--	g24972 = NAND(g19962, g23172)
--	g12767 = NAND(g4467, g6961)
--	g13798 = NAND(g11280, g3423)
--	g11973 = NAND(g8365, g2051)
--	g30580 = NAND(g29335, g19666)
--	g29657 = NAND(g28363, g13634)
--	g17779 = NAND(g6637, g14556, g6704, g12471)
--	g11674 = NAND(g8676, g4674)
--	g7879 = NAND(I12262, I12263)
--	g23726 = NAND(g9559, g21140)
--	I20203 = NAND(g16246, g11147)
--	g16524 = NAND(g13822, g13798)
--	g26685 = NAND(g9264, g25160)
--	I14429 = NAND(g4005, I14427)
--	g14574 = NAND(g12256, g6120)
--	g12191 = NAND(I15052, I15053)
--	g14452 = NAND(g3538, g11207, g3649, g8542)
--	g11934 = NAND(g8139, g8187)
--	g16119 = NAND(I17475, I17476)
--	I14428 = NAND(g8595, I14427)
--	g12521 = NAND(g7471, g5969)
--	g17647 = NAND(g5905, g14497, g5976, g12614)
--	I29313 = NAND(g29501, g12154)
--	g8609 = NAND(g1171, g1157)
--	g19450 = NAND(g11471, g17794)
--	I14765 = NAND(g9808, I14764)
--	g11761 = NAND(I14610, I14611)
--	g22651 = NAND(g20114, g2873)
--	I29285 = NAND(g29489, I29284)
--	g14051 = NAND(g10323, g11527)
--	g14072 = NAND(g11571, g11483)
--	g16749 = NAND(g3957, g13772, g4027, g11631)
--	g20163 = NAND(g16663, g13938)
--	g15782 = NAND(g6585, g14556, g6697, g10061)
--	I29254 = NAND(g29482, I29253)
--	I15214 = NAND(g1714, I15212)
--	g14780 = NAND(g6275, g12101, g6329, g12423)
--	g12045 = NAND(g1783, g8146)
--	g10820 = NAND(g9985, g9920, g9843)
--	g14820 = NAND(g6307, g12173, g6315, g12423)
--	g17513 = NAND(g3247, g13765, g3325, g8481)
--	g28827 = NAND(g27837, g7362, g1862)
--	g25531 = NAND(g22763, g2868)
--	g15853 = NAND(g14714, g9417, g12337)
--	I15241 = NAND(g10003, g6351)
--	g12462 = NAND(g7051, g7064, g10190)
--	g13241 = NAND(g7503, g10544)
--	g25186 = NAND(g5396, g23602)
--	g14691 = NAND(g12695, g12505)
--	g25953 = NAND(g22756, g24570, g22688)
--	g8803 = NAND(g128, g4646)
--	g9954 = NAND(g6128, g6120)
--	I22792 = NAND(g11956, g21434)
--	I22967 = NAND(g21228, I22965)
--	g13100 = NAND(g6581, g12137, g6692, g10061)
--	g23575 = NAND(I22711, I22712)
--	g20173 = NAND(g16696, g13972)
--	g10929 = NAND(g1099, g7854)
--	g31669 = NAND(I29254, I29255)
--	g15864 = NAND(g14833, g12543, g12487)
--	g33669 = NAND(g33378, g862)
--	g25334 = NAND(g21253, g23756)
--	g17723 = NAND(g6597, g14556, g6668, g12721)
--	g10583 = NAND(g7475, g862)
--	g10928 = NAND(g8181, g8137, g417)
--	g15748 = NAND(g13257, g13130, g7922, g13241)
--	g21283 = NAND(g11291, g17157)
--	g9912 = NAND(I13463, I13464)
--	I13045 = NAND(g5120, I13043)
--	g20134 = NAND(g17572, g14542, g17495, g14452)
--	g13515 = NAND(g12628, g12588, g12524, g12464)
--	g13882 = NAND(g3590, g11207, g3672, g11576)
--	g24760 = NAND(I23918, I23919)
--	I23961 = NAND(g23184, g13631)
--	g25216 = NAND(g6088, g23678)
--	g14113 = NAND(g11626, g11537)
--	I24385 = NAND(g14347, I24383)
--	g15036 = NAND(g12780, g12581)
--	g19597 = NAND(g1199, g15995)
--	g12629 = NAND(g7812, g7142)
--	I12877 = NAND(g4200, I12876)
--	I13462 = NAND(g2380, g2384)
--	g8847 = NAND(g4831, g4681)
--	g12628 = NAND(g7074, g6336, g6390)
--	g22850 = NAND(g1536, g19581, g10699)
--	g11441 = NAND(g9599, g3267)
--	I13140 = NAND(g6154, I13139)
--	I22901 = NAND(g21228, I22899)
--	g28786 = NAND(g27837, g7405, g7322)
--	g11206 = NAND(I14276, I14277)
--	g16238 = NAND(g4698, g13883, g12054)
--	I14499 = NAND(g8737, I14497)
--	g17412 = NAND(g14520, g14489)
--	I18625 = NAND(g2079, g14712)
--	g14768 = NAND(g12662, g12571)
--	g28945 = NAND(g27854, g8211)
--	g14803 = NAND(g5208, g12059, g5308, g12497)
--	I14498 = NAND(g9020, I14497)
--	g33679 = NAND(g33394, g10737, g10308)
--	g12147 = NAND(g8302, g8201)
--	I12402 = NAND(g3808, I12401)
--	I15107 = NAND(g5313, I15105)
--	I22823 = NAND(g11978, I22822)
--	I14611 = NAND(g8678, I14609)
--	I14924 = NAND(g9558, I14923)
--	g12370 = NAND(I15213, I15214)
--	g25974 = NAND(g24576, g22837)
--	g17716 = NAND(g5957, g14497, g6027, g12614)
--	g15008 = NAND(g12780, g10341)
--	I23971 = NAND(g490, I23969)
--	g25293 = NAND(g21190, g23726)
--	g12151 = NAND(g8316, g8211)
--	g19854 = NAND(I20222, I20223)
--	g13940 = NAND(g11426, g8889, g11707, g8829)
--	I22966 = NAND(g12288, I22965)
--	g23949 = NAND(g7074, g21012)
--	g28448 = NAND(g23975, g27377)
--	I15263 = NAND(g10081, I15262)
--	g10552 = NAND(g2153, g7374)
--	g8751 = NAND(g3969, g4012, g3983, g4005)
--	g15907 = NAND(g14833, g9417, g12487)
--	g22681 = NAND(I21993, I21994)
--	g11135 = NAND(I14186, I14187)
--	I14330 = NAND(g225, g9966)
--	g19916 = NAND(g3029, g16313)
--	g16728 = NAND(g13884, g13870, g14089, g11639)
--	g12227 = NAND(g8418, g8330)
--	I14764 = NAND(g9808, g5821)
--	g11962 = NAND(I14789, I14790)
--	I29284 = NAND(g29489, g12085)
--	I31973 = NAND(g33641, I31972)
--	I29304 = NAND(g12121, I29302)
--	I18581 = NAND(g14678, I18579)
--	I26051 = NAND(g13500, I26049)
--	I25847 = NAND(g24799, I25845)
--	I26072 = NAND(g13517, I26070)
--	I11825 = NAND(g4593, I11824)
--	I12876 = NAND(g4200, g4180)
--	g14999 = NAND(g12739, g12824)
--	g16304 = NAND(g4765, g13970, g12054)
--	g12044 = NAND(g1657, g8139)
--	I15004 = NAND(g1700, I15002)
--	g21509 = NAND(g17820, g14898, g17647, g17608)
--	g17765 = NAND(g6649, g14556, g6719, g12721)
--	I14259 = NAND(g3133, I14257)
--	I17495 = NAND(g13378, I17494)
--	g27377 = NAND(g10685, g25930)
--	g24926 = NAND(g20172, g20163, g23357, g13995)
--	g25275 = NAND(g22342, g11991)
--	g12301 = NAND(I15148, I15149)
--	I14258 = NAND(g8154, I14257)
--	g12120 = NAND(g2476, g8273)
--	g27738 = NAND(g21228, g25243, g26424, g26148)
--	I32440 = NAND(g34227, I32439)
--	g25237 = NAND(g6434, g23711)
--	I15106 = NAND(g9780, I15105)
--	g13273 = NAND(g1459, g10699)
--	g19335 = NAND(g15717, g1056)
--	g10961 = NAND(g1442, g7876)
--	g29679 = NAND(g153, g28353, g23042)
--	g15729 = NAND(g5949, g14549, g6027, g9935)
--	g14505 = NAND(g12073, g9961)
--	I12287 = NAND(g1484, g1300)
--	I14955 = NAND(g9620, g6181)
--	g19965 = NAND(g3380, g16424)
--	g11951 = NAND(g9166, g847, g703)
--	g15728 = NAND(g5200, g14399, g5313, g9780)
--	g13951 = NAND(g10295, g11729)
--	I12076 = NAND(g979, I12074)
--	g23047 = NAND(g482, g20000)
--	g13795 = NAND(g11216, g401)
--	g28896 = NAND(g27837, g1936, g1862)
--	I14171 = NAND(g3119, I14169)
--	g20871 = NAND(g14434, g17396)
--	I22893 = NAND(g12189, I22892)
--	I12269 = NAND(g1141, g956)
--	I13044 = NAND(g5115, I13043)
--	g17775 = NAND(g6255, g14575, g6351, g12672)
--	I22865 = NAND(g12146, I22864)
--	g23756 = NAND(g9621, g21206)
--	g14723 = NAND(g7704, g12772)
--	g23780 = NAND(I22930, I22931)
--	g14433 = NAND(g12035, g9890)
--	I24384 = NAND(g23721, I24383)
--	g21350 = NAND(g15751, g15742, g15735, g13108)
--	g16312 = NAND(g13580, g13574)
--	g14104 = NAND(g11514, g8864)
--	I25846 = NAND(g26212, I25845)
--	g14343 = NAND(g11961, g9670)
--	g10971 = NAND(g7867, g7886)
--	g28958 = NAND(g27833, g8249)
--	g14971 = NAND(g12667, g12581)
--	g16745 = NAND(g3594, g13730, g3661, g11389)
--	g31748 = NAND(I29303, I29304)
--	g26208 = NAND(g7975, g24751)
--	g16813 = NAND(g3614, g13799, g3625, g8542)
--	I22938 = NAND(g21228, I22936)
--	g27824 = NAND(I26394, I26395)
--	g13920 = NAND(g11621, g11483)
--	I17460 = NAND(g13378, g1300)
--	g24591 = NAND(g22833, g22642)
--	g24776 = NAND(g3040, g23052)
--	I14817 = NAND(g9962, I14816)
--	g25236 = NAND(I24415, I24416)
--	I15121 = NAND(g9910, g2102)
--	g34422 = NAND(I32432, I32433)
--	g28857 = NAND(g27779, g1802, g1728)
--	g14133 = NAND(g11692, g11747)
--	I12279 = NAND(g1472, I12277)
--	I14532 = NAND(g8873, I14530)
--	g13121 = NAND(g11117, g8411)
--	g28793 = NAND(g27800, g7328, g2153)
--	I13403 = NAND(g2250, I13401)
--	I12278 = NAND(g1467, I12277)
--	g24950 = NAND(g19442, g23154)
--	I12469 = NAND(g405, I12468)
--	g27931 = NAND(g25425, g25381, g25780)
--	g28765 = NAND(g27800, g7374, g7280)
--	g7611 = NAND(g4057, g4064)
--	g14011 = NAND(g10295, g11473)
--	g20151 = NAND(g17598, g14570, g17514, g14519)
--	g20172 = NAND(g16876, g8131)
--	I12468 = NAND(g405, g392)
--	g13291 = NAND(g10715, g1500)
--	g11173 = NAND(g4966, g7898, g9064)
--	g12190 = NAND(g8365, g8255)
--	g22753 = NAND(g1536, g19632)
--	g28504 = NAND(g758, g27528, g11679)
--	g21357 = NAND(g15736, g13109, g15726, g13086)
--	g31009 = NAND(g27187, g29503, g19644)
--	g14627 = NAND(g12553, g12772)
--	g23357 = NAND(g20201, g11231)
--	g14959 = NAND(g12695, g12798)
--	g14379 = NAND(g5723, g11907)
--	g22650 = NAND(g7888, g19581)
--	g11134 = NAND(g8138, g8240, g8301)
--	g23105 = NAND(g8097, g19887)
--	g13134 = NAND(g11134, g8470)
--	g14378 = NAND(g11979, g9731)
--	g7209 = NAND(g6052, g6098)
--	g12024 = NAND(g8381, g8418)
--	g17650 = NAND(g6299, g12101, g6315, g14745)
--	g10603 = NAND(g10077, g9751)
--	g17736 = NAND(g5563, g14522, g5659, g12563)
--	g15798 = NAND(g6629, g14602, g6704, g14786)
--	g25021 = NAND(g21417, g23363)
--	I11824 = NAND(g4593, g4601)
--	g15674 = NAND(g921, g13110)
--	g9310 = NAND(I13078, I13079)
--	I14289 = NAND(g8282, g3835)
--	g28298 = NAND(g10533, g26131, g26990)
--	g9663 = NAND(g128, g4646)
--	g13927 = NAND(g3578, g11207, g3632, g11389)
--	I17494 = NAND(g13378, g1448)
--	g29118 = NAND(g27886, g9755)
--	I12217 = NAND(g1437, g1478)
--	g14730 = NAND(g5615, g12093, g5623, g12301)
--	g22709 = NAND(g1193, g19611)
--	I22822 = NAND(g11978, g21434)
--	g13240 = NAND(g1046, g10521)
--	g24957 = NAND(g21359, g23462)
--	g11491 = NAND(g9982, g4000)
--	g12644 = NAND(g10233, g4531)
--	g11903 = NAND(g9099, g3712)
--	I14816 = NAND(g9962, g6513)
--	I32203 = NAND(g33937, I32202)
--	g23890 = NAND(g7004, g20682)
--	g12969 = NAND(g4388, g7178, g10476)
--	I13520 = NAND(g2518, I13518)
--	g20645 = NAND(g14344, g17243)
--	g28856 = NAND(g27738, g8093)
--	g14548 = NAND(g12208, g5774)
--	g17225 = NAND(g8612, g14367)
--	g17708 = NAND(g5216, g14490, g5313, g12497)
--	g12197 = NAND(g7296, g5290)
--	g8434 = NAND(g3080, g3072)
--	g28512 = NAND(g10857, g27155, g27142)
--	g23552 = NAND(I22684, I22685)
--	g15005 = NAND(g12667, g12622)
--	g14317 = NAND(g5033, g11862)
--	g12411 = NAND(g7393, g5276)
--	g8347 = NAND(g4358, g4349, g4340)
--	I15262 = NAND(g10081, g2273)
--	g23778 = NAND(I22922, I22923)
--	g11395 = NAND(g9601, g3983)
--	I13497 = NAND(g255, g232)
--	g11990 = NAND(g9166, g703)
--	g13990 = NAND(g11669, g11584)
--	g23786 = NAND(I22945, I22946)
--	I18487 = NAND(g14611, I18485)
--	g13898 = NAND(g11621, g11747)
--	I22864 = NAND(g12146, g21228)
--	g21356 = NAND(g15780, g15752, g15743, g13118)
--	I12373 = NAND(g3457, I12372)
--	g14626 = NAND(g12232, g9852, g12159, g9715)
--	g24661 = NAND(g23210, g23195, g22984)
--	g24547 = NAND(g22638, g22643, g22754)
--	I31972 = NAND(g33641, g33631)
--	g12450 = NAND(g7738, g10281)
--	g10775 = NAND(g7960, g7943, g8470)
--	g9295 = NAND(I13066, I13067)
--	g12819 = NAND(g9848, g6961)
--	g12910 = NAND(g11002, g10601)
--	g34174 = NAND(g617, g33851, g12323)
--	g17792 = NAND(g6601, g14602, g6697, g12721)
--	I22900 = NAND(g12193, I22899)
--	g10737 = NAND(g6961, g9848)
--	g25537 = NAND(g22763, g2873)
--	g12111 = NAND(g847, g9166)
--	g28271 = NAND(g10533, g27004, g26990)
--	g13861 = NAND(g1459, g10671)
--	g21331 = NAND(g11402, g17157)
--	g13573 = NAND(g8002, g10544, g7582, g1351)
--	g23932 = NAND(g7051, g20875)
--	I14713 = NAND(g9671, I14712)
--	g12590 = NAND(g7097, g7110, g10229)
--	g33083 = NAND(g7805, g32118)
--	g11389 = NAND(I14399, I14400)
--	g25492 = NAND(g12479, g22457)
--	g14697 = NAND(g12662, g12824)
--	g9966 = NAND(I13498, I13499)
--	g7184 = NAND(g5706, g5752)
--	g9705 = NAND(g2619, g2587)
--	I14610 = NAND(g8993, I14609)
--	I26368 = NAND(g14211, I26366)
--	I29263 = NAND(g12046, I29261)
--	g11534 = NAND(g7121, g8958)
--	I23602 = NAND(g4322, I23600)
--	g20784 = NAND(g14616, g17595)
--	g28736 = NAND(g27742, g7308, g7252)
--	g19265 = NAND(g15721, g15715, g13091, g15710)
--	g13098 = NAND(g5933, g12129, g6023, g9935)
--	I20487 = NAND(g16696, I20486)
--	g11251 = NAND(g8438, g3092)
--	g25381 = NAND(g538, g23088)
--	I23970 = NAND(g22202, I23969)
--	g13462 = NAND(g12449, g12412, g12342, g12294)
--	g28843 = NAND(g27907, g7456, g7387)
--	g19510 = NAND(g15969, g10841, g10899)
--	g20181 = NAND(g13252, g16846)
--	g12019 = NAND(g7322, g1906)
--	g17598 = NAND(g3949, g13824, g4027, g8595)
--	g12196 = NAND(g8764, g4688)
--	g11997 = NAND(g2319, g8316)
--	I20469 = NAND(g16728, I20467)
--	I21994 = NAND(g19638, I21992)
--	I12242 = NAND(g1105, I12240)
--	g12526 = NAND(g10194, g7110, g10213)
--	g15725 = NAND(g5603, g14522, g5681, g9864)
--	I20468 = NAND(g16663, I20467)
--	g29154 = NAND(g27937, g9835)
--	g21433 = NAND(g17792, g14830, g17765, g14750)
--	I22892 = NAND(g12189, g21228)
--	g19442 = NAND(g11431, g17794)
--	g12402 = NAND(g7704, g10266)
--	g10611 = NAND(g10115, g9831)
--	I13111 = NAND(g5813, I13109)
--	g13871 = NAND(g4955, g11834)
--	I23919 = NAND(g9333, I23917)
--	I18486 = NAND(g1677, I18485)
--	g28259 = NAND(g10504, g26987, g26973)
--	g14924 = NAND(g12558, g12505)
--	I22712 = NAND(g21434, I22710)
--	g17656 = NAND(I18626, I18627)
--	I20187 = NAND(g16272, g1333)
--	g15744 = NAND(g6641, g14602, g6719, g10061)
--	I17476 = NAND(g1105, I17474)
--	I23918 = NAND(g23975, I23917)
--	I18580 = NAND(g1945, I18579)
--	I26050 = NAND(g25997, I26049)
--	I13384 = NAND(g246, I13382)
--	g12001 = NAND(I14854, I14855)
--	I13067 = NAND(g4304, I13065)
--	I12841 = NAND(g4222, I12840)
--	I11877 = NAND(g4388, g4430)
--	g10529 = NAND(g1592, g7308)
--	g13628 = NAND(g3372, g11107)
--	g23850 = NAND(g12185, g19462)
--	g13911 = NAND(g11834, g4917)
--	I18531 = NAND(g14640, I18529)
--	g17364 = NAND(g8639, g14367)
--	g28955 = NAND(g27837, g1936, g7362)
--	I14277 = NAND(g3484, I14275)
--	I21977 = NAND(g7680, I21976)
--	g14696 = NAND(g5567, g12093, g5685, g12563)
--	I24363 = NAND(g23687, g14320)
--	g8163 = NAND(g3419, g3423)
--	g15962 = NAND(g14833, g9417, g9340)
--	g14764 = NAND(g7738, g12798)
--	g11591 = NAND(I14531, I14532)
--	g21011 = NAND(g14504, g17399, g9629)
--	I15147 = NAND(g9864, g5659)
--	g12066 = NAND(I14924, I14925)
--	I20486 = NAND(g16696, g16757)
--	g24943 = NAND(g20068, g23172)
--	g20644 = NAND(g14342, g17220, g9372)
--	g27876 = NAND(I26418, I26419)
--	g15833 = NAND(g14714, g12378, g12337)
--	I13402 = NAND(g2246, I13401)
--	g11355 = NAND(g9551, g3310)
--	g28994 = NAND(g27907, g2495, g7424)
--	g14868 = NAND(g12755, g12680)
--	g17571 = NAND(g8579, g14367)
--	I11866 = NAND(g4401, I11864)
--	g27854 = NAND(g21228, g25283, g26424, g26195)
--	g25062 = NAND(g21403, g23363)
--	I20223 = NAND(g11170, I20221)
--	g16507 = NAND(g13797, g13764)
--	g11858 = NAND(g9014, g3010)
--	I14352 = NAND(g8848, I14350)
--	I17883 = NAND(g13336, g1135)
--	g11172 = NAND(g8478, g3096)
--	g12511 = NAND(g7028, g5644, g5698)
--	g22687 = NAND(g19560, g7870)
--	g7885 = NAND(I12270, I12271)
--	g11996 = NAND(g7280, g2197)
--	g17495 = NAND(g3566, g13730, g3668, g8542)
--	g23379 = NAND(g20216, g11248)
--	I14170 = NAND(g8389, I14169)
--	I13077 = NAND(g5462, g5467)
--	g23112 = NAND(g21024, g10733)
--	g20870 = NAND(g14432, g17315, g9567)
--	g17816 = NAND(g6657, g14602, g6668, g10061)
--	g14258 = NAND(g9203, g11903)
--	g11394 = NAND(g9600, g3661)
--	g22643 = NAND(g20136, g18954)
--	g34051 = NAND(I31973, I31974)
--	g21386 = NAND(g15798, g15788, g15782, g13139)
--	I18587 = NAND(g2370, g14679)
--	g21603 = NAND(g17872, g14987, g17723, g17689)
--	I14853 = NAND(g9433, g5142)
--	g27550 = NAND(g24943, g25772)
--	g9485 = NAND(g1657, g1624)
--	g14069 = NAND(g11653, g8864)
--	g22668 = NAND(g20219, g2912)
--	g10602 = NAND(g7411, g7451)
--	g11446 = NAND(g8700, g6941, g8734)
--	g14810 = NAND(g12700, g10312)
--	g15033 = NAND(g12806, g7142)
--	g12287 = NAND(g8381, g2587)
--	g21429 = NAND(g17788, g14803, g17578, g17520)
--	g17669 = NAND(g3570, g11238, g3632, g13902)
--	g12307 = NAND(g7395, g5983)
--	g14879 = NAND(g12646, g10266)
--	I13066 = NAND(g4308, I13065)
--	g17668 = NAND(g3235, g13765, g3310, g13877)
--	g23428 = NAND(g13945, g20522)
--	g13058 = NAND(g10544, g1312)
--	g28977 = NAND(g27937, g2629, g2555)
--	g12431 = NAND(I15254, I15255)
--	g20979 = NAND(g5385, g17309)
--	g28783 = NAND(g27779, g7315, g1728)
--	g20055 = NAND(g11269, g17794)
--	g20111 = NAND(g17513, g14517, g17468, g14422)
--	g17525 = NAND(g14600, g14574)
--	I13511 = NAND(g2093, I13509)
--	g12341 = NAND(g7512, g5308)
--	g28823 = NAND(g27738, g14565)
--	I14276 = NAND(g8218, I14275)
--	I21976 = NAND(g7680, g19620)
--	g16291 = NAND(g13551, g13545)
--	I23985 = NAND(g22182, g482)
--	g13281 = NAND(g10916, g1099)
--	g27670 = NAND(g25172, g26666)
--	g22713 = NAND(g20114, g2890)
--	g11957 = NAND(g8205, g8259)
--	g28336 = NAND(g27064, g24756, g27163, g19644)
--	I32202 = NAND(g33937, g33670)
--	g13739 = NAND(g11773, g11261)
--	g25396 = NAND(g22384, g2208, g8259)
--	g28966 = NAND(g27858, g2361, g7380)
--	g14918 = NAND(g12646, g12772)
--	g20150 = NAND(g17705, g17669, g17635, g14590)
--	g14079 = NAND(g11626, g11763)
--	g17705 = NAND(g3586, g13799, g3661, g13902)
--	g8292 = NAND(g218, g215)
--	g14599 = NAND(g12207, g9739)
--	I12253 = NAND(g1129, I12251)
--	g17679 = NAND(g5611, g14425, g5681, g12563)
--	g7869 = NAND(I12252, I12253)
--	g10598 = NAND(g7191, g6404)
--	g15788 = NAND(g6613, g12211, g6675, g14786)
--	I18579 = NAND(g1945, g14678)
--	g14598 = NAND(g5248, g12002, g5331, g12497)
--	I14733 = NAND(g9732, g5475)
--	g15829 = NAND(g4112, g13831)
--	g17686 = NAND(g6251, g14529, g6322, g12672)
--	I12372 = NAND(g3457, g3462)
--	g14817 = NAND(g12711, g12622)
--	g28288 = NAND(g10533, g26105, g27004)
--	g19913 = NAND(g11430, g17794)
--	g19614 = NAND(g1542, g16047)
--	g22875 = NAND(g20516, g2980)
--	g25020 = NAND(g21377, g23462)
--	g7442 = NAND(g896, g890)
--	g24917 = NAND(g19913, g23172)
--	g10561 = NAND(g7157, g5712)
--	g27468 = NAND(g24951, g24932, g24925, g26852)
--	I22921 = NAND(g14677, g21284)
--	g27306 = NAND(g24787, g26235)
--	g19530 = NAND(g15829, g10841)
--	g12286 = NAND(I15129, I15130)
--	g14656 = NAND(g12553, g12405)
--	g9177 = NAND(g3355, g3401)
--	g22837 = NAND(g20219, g2907)
--	g12306 = NAND(g7394, g5666)
--	I26461 = NAND(g14306, I26459)
--	I24416 = NAND(g14382, I24414)
--	g16604 = NAND(g3251, g11194, g3267, g13877)
--	I22799 = NAND(g11960, g21434)
--	g13551 = NAND(g11812, g7479, g7903, g10521)
--	g10336 = NAND(I13750, I13751)
--	g28976 = NAND(g27903, g8273)
--	I14712 = NAND(g9671, g5128)
--	I13335 = NAND(g1687, I13334)
--	g16770 = NAND(g3263, g13765, g3274, g8481)
--	g8561 = NAND(g3782, g3774)
--	I22973 = NAND(g9657, I22972)
--	g26248 = NAND(I25220, I25221)
--	g12187 = NAND(I15042, I15043)
--	I29262 = NAND(g29485, I29261)
--	g11490 = NAND(g8666, g3639, g3694)
--	I26393 = NAND(g26488, g14227)
--	
--	g30249 = NOR(g5297, g28982)
--	g33141 = NOR(g32099, g8400)
--	g13824 = NOR(g8623, g11702)
--	g27479 = NOR(g9056, g26616)
--	g12479 = NOR(g2028, g8310)
--	g20854 = NOR(g5381, g17243)
--	g33135 = NOR(g32090, g8350)
--	g7675 = NOR(g1554, g1559, g1564, g1548)
--	g12486 = NOR(g9055, g9013, g8957, g8905)
--	g9694 = NOR(g1936, g1862)
--	g8906 = NOR(g3530, g3522)
--	g14816 = NOR(g10166, g12252)
--	g12223 = NOR(g2051, g8365)
--	g14687 = NOR(g5352, g12166)
--	g14752 = NOR(g12540, g10040)
--	g16272 = NOR(g13580, g11189)
--	g22524 = NOR(g19720, g1361)
--	g25778 = NOR(g25459, g25420)
--	g26212 = NOR(g23837, g25408)
--	g17194 = NOR(g11039, g13480)
--	g14392 = NOR(g12114, g9537)
--	g13700 = NOR(g3288, g11615)
--	g11658 = NOR(g8021, g3506)
--	g15718 = NOR(g13858, g11330)
--	g10488 = NOR(g4616, g7133, g10336)
--	g29107 = NOR(g6203, g7791, g26977)
--	g10893 = NOR(g1189, g7715, g7749)
--	g25932 = NOR(g7680, g24528)
--	g29141 = NOR(g9374, g27999)
--	g14713 = NOR(g12483, g9974)
--	g31507 = NOR(g9064, g29556)
--	g15099 = NOR(g13191, g12869)
--	g11527 = NOR(g8165, g8114)
--	g32715 = NOR(g31327, I30261, I30262)
--	g15098 = NOR(g13191, g6927)
--	g30148 = NOR(g28799, g7335)
--	g23602 = NOR(g9672, g20979)
--	g28470 = NOR(g8021, g27617)
--	g16220 = NOR(g13499, g4939)
--	g14679 = NOR(g12437, g9911)
--	g23955 = NOR(g2823, g18890)
--	g33163 = NOR(g32099, g7809)
--	g24619 = NOR(g23554, g23581)
--	g14188 = NOR(g9162, g12259)
--	g14124 = NOR(g8830, g11083)
--	g14678 = NOR(g12432, g9907)
--	g16246 = NOR(g13551, g11169)
--	g12117 = NOR(g10113, g9755)
--	g29361 = NOR(g7553, g28174)
--	g15140 = NOR(g12887, g13680)
--	g14093 = NOR(g8833, g11083)
--	g15061 = NOR(g6815, g13394)
--	g13910 = NOR(g4899, g4975, g11173)
--	g13202 = NOR(g8347, g10511)
--	g12123 = NOR(g6856, g2748)
--	g27772 = NOR(g7297, g25839)
--	g12772 = NOR(g5188, g9300)
--	g31121 = NOR(g4776, g29540)
--	g23918 = NOR(g2799, g21382)
--	g15162 = NOR(g13809, g12904)
--	g11384 = NOR(g8538, g8540)
--	g23079 = NOR(g8390, g19965)
--	g29106 = NOR(g9451, g28020)
--	g13094 = NOR(g7487, g10762)
--	g26603 = NOR(g24908, g24900)
--	g29033 = NOR(g5511, g7738, g28010)
--	g15628 = NOR(g11907, g14228)
--	g32520 = NOR(g31554, I30054, I30055)
--	g17239 = NOR(g11119, g13518)
--	g31134 = NOR(g8033, g29679, g24732)
--	g33134 = NOR(g7686, g32057)
--	g16227 = NOR(g1554, g13574)
--	g27007 = NOR(g5706, g25821)
--	g31506 = NOR(g4793, g29540)
--	g15071 = NOR(g6831, g13416)
--	g15147 = NOR(g13716, g12892)
--	g15754 = NOR(g341, g7440, g13385)
--	g14037 = NOR(g8748, g11083)
--	g15825 = NOR(g7666, g13217)
--	g16044 = NOR(g10961, g13861)
--	g27720 = NOR(g9253, g25791)
--	g14419 = NOR(g12152, g9546)
--	g29012 = NOR(g5863, g28020)
--	g15151 = NOR(g13745, g7027)
--	g14418 = NOR(g12151, g9594)
--	g10266 = NOR(g5188, g5180)
--	g25958 = NOR(g7779, g24609)
--	g32296 = NOR(g9044, g31509, g12259)
--	g31491 = NOR(g8938, g29725)
--	g11280 = NOR(g8647, g3408)
--	g25944 = NOR(g7716, g24591)
--	g29359 = NOR(g7528, g28167)
--	g12806 = NOR(g9472, g9407)
--	g14194 = NOR(g5029, g10515)
--	g19413 = NOR(g17151, g14221)
--	g24953 = NOR(g10262, g23978, g12259)
--	g15059 = NOR(g12839, g13350)
--	g26298 = NOR(g8297, g24825)
--	g30129 = NOR(g28739, g14537)
--	g15058 = NOR(g12838, g13350)
--	g11231 = NOR(g7928, g4801, g4793)
--	g17284 = NOR(g9253, g14317)
--	g12193 = NOR(g2342, g8316)
--	g11885 = NOR(g7153, g7167)
--	g29173 = NOR(g9259, g27999, g7704)
--	g14313 = NOR(g12016, g9250)
--	g28476 = NOR(g27627, g26547)
--	g16226 = NOR(g8052, g13545)
--	g11763 = NOR(g3881, g8172)
--	g25504 = NOR(g22550, g7222)
--	g15120 = NOR(g12873, g13605)
--	g32910 = NOR(g31327, I30468, I30469)
--	g25317 = NOR(g9766, g23782)
--	g10808 = NOR(g8509, g7611)
--	g15146 = NOR(g13716, g7003)
--	g14036 = NOR(g8725, g11083)
--	g34737 = NOR(g34706, g30003)
--	g12437 = NOR(g2319, g8267)
--	g27703 = NOR(g9607, g25791)
--	g20000 = NOR(g13661, g16264)
--	g13480 = NOR(g3017, g11858)
--	g14642 = NOR(g12374, g9829)
--	g12347 = NOR(g9321, g9274)
--	g14064 = NOR(g9214, g12259)
--	g13076 = NOR(g7443, g10741)
--	g33098 = NOR(g31997, g4616)
--	g28519 = NOR(g8011, g27602, g10295)
--	g12821 = NOR(g7132, g10223, g7149, g10261)
--	g27063 = NOR(g26485, g26516)
--	g24751 = NOR(g3034, g23105)
--	g29903 = NOR(g6928, g28484)
--	g11773 = NOR(g8883, g4785)
--	g27516 = NOR(g9180, g26657)
--	g33140 = NOR(g7693, g32072)
--	g13341 = NOR(g7863, g10762)
--	g12137 = NOR(g6682, g7097)
--	g13670 = NOR(g8123, g10756)
--	g10555 = NOR(g7227, g4601, g4608)
--	g20841 = NOR(g17847, g12027)
--	g23042 = NOR(g16581, g19462, g10685)
--	g14712 = NOR(g12479, g9971)
--	g13335 = NOR(g7851, g10741)
--	g19890 = NOR(g16987, g8058)
--	g14914 = NOR(g12822, g12797)
--	g24391 = NOR(g22190, g14645)
--	g15127 = NOR(g12879, g13605)
--	g30271 = NOR(g7041, g29008)
--	g23124 = NOR(g8443, g20011)
--	g23678 = NOR(g9809, g21190)
--	g16024 = NOR(g14216, g11890)
--	g12208 = NOR(g10096, g5759)
--	g33447 = NOR(g31978, g7643)
--	g26330 = NOR(g8631, g24825)
--	g23686 = NOR(g2767, g21066)
--	g20014 = NOR(g17096, g11244)
--	g33162 = NOR(g4859, g32072)
--	g29898 = NOR(g6895, g28458)
--	g12453 = NOR(g9444, g5527)
--	g15095 = NOR(g13177, g12866)
--	g29191 = NOR(g7738, g28010)
--	g19778 = NOR(g16268, g1061)
--	g11618 = NOR(g8114, g8070)
--	g14382 = NOR(g9390, g11139)
--	g14176 = NOR(g9044, g12259)
--	g14092 = NOR(g8774, g11083)
--	g19999 = NOR(g16232, g13742)
--	g22400 = NOR(g19345, g15718)
--	g20720 = NOR(g17847, g9299)
--	g11469 = NOR(g650, g9903, g645)
--	g12593 = NOR(g9234, g5164)
--	g12346 = NOR(g9931, g9933)
--	g24720 = NOR(g1322, g23051, g19793)
--	g11039 = NOR(g9056, g9092)
--	g11306 = NOR(g3412, g8647)
--	g30132 = NOR(g28789, g7362)
--	g22539 = NOR(g1030, g19699)
--	g8958 = NOR(g3881, g3873)
--	g33147 = NOR(g32090, g7788)
--	g9061 = NOR(g3401, g3361)
--	g19932 = NOR(g3376, g16296)
--	g25887 = NOR(g24984, g11706)
--	g15089 = NOR(g13144, g12861)
--	g15088 = NOR(g13144, g6874)
--	g13937 = NOR(g8883, g4785, g11155)
--	g21277 = NOR(g9417, g9340, g17467)
--	g29032 = NOR(g9300, g27999)
--	g15126 = NOR(g12878, g13605)
--	g11666 = NOR(g8172, g8125)
--	g16581 = NOR(g13756, g8086)
--	g11363 = NOR(g8626, g8751)
--	g11217 = NOR(g8531, g6875)
--	g31318 = NOR(g4785, g29697)
--	g12711 = NOR(g6209, g9326)
--	g8177 = NOR(g4966, g4991, g4983)
--	g30171 = NOR(g28880, g7431)
--	g17515 = NOR(g13221, g10828)
--	g15060 = NOR(g13350, g6814)
--	g12492 = NOR(g7704, g5170, g5164)
--	g26545 = NOR(g24881, g24855)
--	g27982 = NOR(g7212, g25856)
--	g27381 = NOR(g8075, g26657)
--	g14415 = NOR(g12147, g9590)
--	g13110 = NOR(g7841, g10741)
--	g26598 = NOR(g8990, g13756, g24732)
--	g33146 = NOR(g4669, g32057)
--	g29071 = NOR(g5873, g28020)
--	g29370 = NOR(g28585, g28599)
--	g33427 = NOR(g10278, g31950)
--	g22399 = NOR(g1367, g19720)
--	g10312 = NOR(g5881, g5873)
--	g15055 = NOR(g6808, g13350)
--	g15070 = NOR(g6829, g13416)
--	g30159 = NOR(g28799, g14589)
--	g23560 = NOR(g9607, g20838)
--	g12483 = NOR(g2453, g8324)
--	g11216 = NOR(g7998, g8037)
--	g10799 = NOR(g347, g7541)
--	g12553 = NOR(g5170, g9206)
--	g23642 = NOR(g9733, g21124)
--	g15067 = NOR(g12842, g13394)
--	g15094 = NOR(g13177, g12865)
--	g30144 = NOR(g28789, g7322)
--	g24453 = NOR(g7446, g22325)
--	g15150 = NOR(g12895, g13745)
--	g31127 = NOR(g4966, g29556)
--	g13908 = NOR(g4709, g8796, g11155)
--	g12252 = NOR(g9995, g10185)
--	g26309 = NOR(g8575, g24825)
--	g11747 = NOR(g3530, g8114)
--	g13568 = NOR(g8046, g12527)
--	g16066 = NOR(g10929, g13307)
--	g16231 = NOR(g13515, g4771)
--	g33103 = NOR(g32176, g31212)
--	g19793 = NOR(g16292, g1404)
--	g33095 = NOR(g31997, g7236)
--	g12847 = NOR(g6838, g10430)
--	g25144 = NOR(g5046, g23623)
--	g13772 = NOR(g3990, g11702)
--	g28515 = NOR(g3881, g27635)
--	g28414 = NOR(g27467, g26347)
--	g30288 = NOR(g7087, g29073)
--	g26976 = NOR(g5016, g25791)
--	g29146 = NOR(g6565, g26994)
--	g12851 = NOR(g6846, g10430)
--	g14539 = NOR(g11977, g9833)
--	g9649 = NOR(g2227, g2153)
--	g14538 = NOR(g11973, g9828)
--	g28584 = NOR(g7121, g27635)
--	g16287 = NOR(g13622, g11144)
--	g33089 = NOR(g31978, g4322)
--	g15102 = NOR(g14591, g6954)
--	g15157 = NOR(g13782, g12900)
--	g33088 = NOR(g31997, g7224)
--	g22514 = NOR(g19699, g1018)
--	g12311 = NOR(g6109, g10136)
--	g15066 = NOR(g12841, g13394)
--	g24575 = NOR(g23498, g23514)
--	g30260 = NOR(g7018, g28982)
--	g23883 = NOR(g2779, g21067)
--	g26865 = NOR(g25328, g25290)
--	g31126 = NOR(g7928, g29540)
--	g16268 = NOR(g7913, g13121)
--	g12780 = NOR(g9402, g9326)
--	g14515 = NOR(g12225, g9761)
--	g14414 = NOR(g12145, g9639)
--	g11493 = NOR(g8964, g8967)
--	g25954 = NOR(g7750, g24591)
--	g23729 = NOR(g17482, g21206)
--	g20982 = NOR(g17929, g12065)
--	g19880 = NOR(g16201, g13634)
--	g27731 = NOR(g9229, g25791)
--	g12846 = NOR(g6837, g10430)
--	g22535 = NOR(g19699, g1030)
--	g13806 = NOR(g11245, g4076)
--	g29889 = NOR(g6905, g28471)
--	g26686 = NOR(g23678, g25189)
--	g13517 = NOR(g8541, g12692)
--	g20390 = NOR(g17182, g14257)
--	g29181 = NOR(g6573, g26994)
--	g21284 = NOR(g16646, g9690)
--	g26267 = NOR(g8033, g24732)
--	g12405 = NOR(g9374, g5180)
--	g16210 = NOR(g13479, g4894)
--	g15054 = NOR(g12837, g13350)
--	g27046 = NOR(g7544, g25888)
--	g15156 = NOR(g13782, g7050)
--	g30294 = NOR(g7110, g29110)
--	g12046 = NOR(g10036, g9640)
--	g14399 = NOR(g5297, g12598)
--	g11006 = NOR(g7686, g7836)
--	g12113 = NOR(g1648, g8187)
--	g28106 = NOR(g7812, g26994)
--	g25189 = NOR(g6082, g23726)
--	g27827 = NOR(g9456, g25839)
--	g9586 = NOR(g1668, g1592)
--	g19887 = NOR(g3025, g16275)
--	g29497 = NOR(g22763, g28241)
--	g27769 = NOR(g9434, g25805)
--	g15131 = NOR(g12881, g13638)
--	g27768 = NOR(g9264, g25805)
--	g30160 = NOR(g28846, g7387)
--	g33094 = NOR(g31950, g4639)
--	g14361 = NOR(g12079, g9413)
--	g20183 = NOR(g17152, g14222)
--	g28514 = NOR(g8165, g27617)
--	g22491 = NOR(g1361, g19720)
--	g16479 = NOR(g14719, g12490)
--	g27027 = NOR(g26398, g26484)
--	g24508 = NOR(g23577, g23618)
--	g23052 = NOR(g8334, g19916)
--	g12662 = NOR(g5863, g9274)
--	g25160 = NOR(g5390, g23659)
--	g12249 = NOR(g5763, g10096)
--	g11834 = NOR(g8938, g8822)
--	g12204 = NOR(g9927, g10160)
--	g15143 = NOR(g6998, g13680)
--	g30170 = NOR(g28846, g14615)
--	g29503 = NOR(g22763, g28250)
--	g14033 = NOR(g8808, g12259)
--	g12081 = NOR(g10079, g9694)
--	g13021 = NOR(g7544, g10741)
--	g22521 = NOR(g1036, g19699)
--	g27647 = NOR(g3004, g26616)
--	g11913 = NOR(g7197, g9166)
--	g13913 = NOR(g8859, g11083)
--	g27356 = NOR(g9429, g26657)
--	g7601 = NOR(g1322, g1333)
--	g15168 = NOR(g13835, g12909)
--	g27826 = NOR(g9501, g25821)
--	g29910 = NOR(g3990, g28484)
--	g11607 = NOR(g8848, g8993, g376)
--	g14514 = NOR(g11959, g9760)
--	g11346 = NOR(g7980, g7964)
--	g29070 = NOR(g5857, g7766, g28020)
--	g12651 = NOR(g9269, g5511)
--	g10421 = NOR(g6227, g9518)
--	g30119 = NOR(g28761, g7315)
--	g14163 = NOR(g8997, g12259)
--	g11797 = NOR(g8883, g8796)
--	g19919 = NOR(g16987, g11205)
--	g30276 = NOR(g7074, g29073)
--	g30285 = NOR(g7097, g29110)
--	g19444 = NOR(g17192, g14295)
--	g12505 = NOR(g9444, g9381)
--	g27717 = NOR(g9492, g26745)
--	g9100 = NOR(g3752, g3712)
--	g12026 = NOR(g9417, g9340)
--	g8984 = NOR(g4899, g4975)
--	g14121 = NOR(g8891, g12259)
--	g25022 = NOR(g714, g23324)
--	g11891 = NOR(g812, g9166)
--	g16242 = NOR(g13529, g4961)
--	g28491 = NOR(g8114, g27617)
--	g33085 = NOR(g31978, g4311)
--	g14291 = NOR(g9839, g12155)
--	g11537 = NOR(g8229, g3873)
--	g27343 = NOR(g8005, g26616)
--	g28981 = NOR(g9234, g27999)
--	g29077 = NOR(g6555, g26994)
--	g12646 = NOR(g9234, g9206)
--	g11283 = NOR(g7953, g4991, g9064)
--	g10760 = NOR(g1046, g7479)
--	g11303 = NOR(g8497, g8500)
--	g31942 = NOR(g8977, g30583)
--	g27368 = NOR(g8119, g26657)
--	g21206 = NOR(g6419, g17396)
--	g12850 = NOR(g10430, g6845)
--	g13796 = NOR(g9158, g12527)
--	g28521 = NOR(g27649, g26604)
--	g31965 = NOR(g30583, g4358)
--	g33131 = NOR(g4659, g32057)
--	g12228 = NOR(g10222, g10206, g10184, g10335)
--	g10649 = NOR(g1183, g8407)
--	g12716 = NOR(g7812, g6555, g6549)
--	g15123 = NOR(g6975, g13605)
--	g10491 = NOR(g6573, g9576)
--	g20027 = NOR(g16242, g13779)
--	g21652 = NOR(g17619, g17663)
--	g27379 = NOR(g8492, g26636)
--	g11483 = NOR(g8165, g3522)
--	g31469 = NOR(g8822, g29725)
--	g11862 = NOR(g7134, g7150)
--	g12050 = NOR(g10038, g9649)
--	g24779 = NOR(g3736, g23167)
--	g16237 = NOR(g8088, g13574)
--	g29916 = NOR(g8681, g28504, g11083)
--	g23135 = NOR(g16476, g19981)
--	g15992 = NOR(g10929, g13846)
--	g28462 = NOR(g3512, g27617)
--	g13326 = NOR(g10929, g10905)
--	g14767 = NOR(g10130, g12204)
--	g14395 = NOR(g12118, g9542)
--	g17420 = NOR(g9456, g14408)
--	g10899 = NOR(g4064, g8451)
--	g22540 = NOR(g19720, g1373)
--	g11252 = NOR(g8620, g3057)
--	g11621 = NOR(g3512, g7985)
--	g15578 = NOR(g7216, g14279)
--	g20998 = NOR(g18065, g9450)
--	g33143 = NOR(g32293, g31518)
--	g7661 = NOR(g1211, g1216, g1221, g1205)
--	g29180 = NOR(g9569, g26977)
--	g14247 = NOR(g9934, g10869)
--	g13872 = NOR(g8745, g11083)
--	g25501 = NOR(g23918, g14645)
--	g20717 = NOR(g5037, g17217)
--	g14272 = NOR(g6411, g10598)
--	g12129 = NOR(g9992, g7051)
--	g12002 = NOR(g5297, g7004)
--	g11213 = NOR(g4776, g7892, g9030)
--	g15142 = NOR(g13680, g12889)
--	g33084 = NOR(g31978, g7655)
--	g20149 = NOR(g17091, g14185)
--	g26609 = NOR(g146, g24732)
--	g15130 = NOR(g13638, g6985)
--	g24148 = NOR(g19268, g19338)
--	g15165 = NOR(g12907, g13835)
--	g31373 = NOR(g4975, g29725)
--	g11780 = NOR(g4899, g8822)
--	g14360 = NOR(g12078, g9484)
--	g9835 = NOR(g2629, g2555)
--	g14447 = NOR(g11938, g9698)
--	g12856 = NOR(g10430, g6855)
--	g29187 = NOR(g7704, g27999)
--	g11846 = NOR(g7635, g7518, g7548)
--	g16209 = NOR(g13478, g4749)
--	g14911 = NOR(g10213, g12364)
--	g27499 = NOR(g9095, g26636)
--	g28540 = NOR(g8125, g27635, g7121)
--	g15372 = NOR(g817, g14279)
--	g14754 = NOR(g12821, g2988)
--	g27722 = NOR(g7247, g25805)
--	g31117 = NOR(g4991, g29556)
--	g27924 = NOR(g9946, g25839)
--	g33117 = NOR(g31261, g32205)
--	g22190 = NOR(g2827, g18949)
--	g8720 = NOR(g358, g365)
--	g15063 = NOR(g6818, g13394)
--	g30934 = NOR(g29836, g29850)
--	g19984 = NOR(g17096, g8171)
--	g15137 = NOR(g6992, g13680)
--	g12432 = NOR(g1894, g8249)
--	g24959 = NOR(g8858, g23324)
--	g17190 = NOR(g723, g14279)
--	g14394 = NOR(g12116, g9414)
--	g14367 = NOR(g9547, g12289)
--	g16292 = NOR(g7943, g13134)
--	g11357 = NOR(g8558, g8561)
--	g29179 = NOR(g9311, g28010, g7738)
--	g14420 = NOR(g12153, g9490)
--	g12198 = NOR(g9797, g9800)
--	g19853 = NOR(g15746, g1052)
--	g27528 = NOR(g8770, g26352, g11083)
--	g10318 = NOR(g25, g22)
--	g14446 = NOR(g12190, g9644)
--	g14227 = NOR(g9863, g10838)
--	g20857 = NOR(g17929, g9380)
--	g27960 = NOR(g7134, g25791)
--	g14540 = NOR(g12287, g9834)
--	g19401 = NOR(g17193, g14296)
--	g17700 = NOR(g14792, g12983)
--	g17625 = NOR(g14541, g12123)
--	g15073 = NOR(g12844, g13416)
--	g28481 = NOR(g3506, g10323, g27617)
--	g10281 = NOR(g5535, g5527)
--	g15122 = NOR(g6959, g13605)
--	g26515 = NOR(g24843, g24822)
--	g12708 = NOR(g9518, g9462)
--	g25005 = NOR(g6811, g23324)
--	g10699 = NOR(g8526, g1514)
--	g15153 = NOR(g13745, g12897)
--	g31116 = NOR(g7892, g29540)
--	g11248 = NOR(g7953, g4991, g4983)
--	g32780 = NOR(g31327, I30330, I30331)
--	g15136 = NOR(g13680, g12885)
--	g29908 = NOR(g6918, g28471)
--	g27879 = NOR(g9523, g25856)
--	g22450 = NOR(g19345, g15724)
--	g12970 = NOR(g10555, g10510, g10488)
--	g27878 = NOR(g9559, g25839)
--	g27337 = NOR(g8334, g26616)
--	g15164 = NOR(g13835, g12906)
--	g11945 = NOR(g7212, g7228)
--	g11999 = NOR(g9654, g7423)
--	g10715 = NOR(g8526, g8466)
--	g21389 = NOR(g10143, g17748, g12259)
--	g20995 = NOR(g5727, g17287)
--	g28520 = NOR(g8229, g27635)
--	g25407 = NOR(g23871, g14645)
--	g27010 = NOR(g6052, g25839)
--	g11932 = NOR(g843, g9166)
--	g33130 = NOR(g32265, g31497)
--	g11448 = NOR(g4191, g8790)
--	g14490 = NOR(g9853, g12598)
--	g19907 = NOR(g16210, g13676)
--	g21140 = NOR(g6073, g17312)
--	g15091 = NOR(g13177, g12863)
--	g33437 = NOR(g31997, g10275)
--	g29007 = NOR(g9269, g28010)
--	g10671 = NOR(g1526, g8466)
--	g14181 = NOR(g9083, g12259)
--	g23871 = NOR(g2811, g21348)
--	g27353 = NOR(g8097, g26616)
--	g16183 = NOR(g9223, g13545)
--	g27823 = NOR(g9792, g25805)
--	g11148 = NOR(g8052, g9197, g9174, g9050)
--	g12680 = NOR(g9631, g9576)
--	g19935 = NOR(g17062, g8113)
--	g31372 = NOR(g8796, g29697)
--	g25141 = NOR(g22228, g10334)
--	g33175 = NOR(g32099, g7828)
--	g24145 = NOR(g19402, g19422)
--	g27966 = NOR(g7153, g25805)
--	g13971 = NOR(g8938, g4975, g11173)
--	g29035 = NOR(g9321, g28020)
--	g14211 = NOR(g9779, g10823)
--	g27364 = NOR(g8426, g26616)
--	g33137 = NOR(g4849, g32072)
--	g12017 = NOR(g9969, g9586)
--	g12364 = NOR(g10102, g10224)
--	g30613 = NOR(g4507, g29365)
--	g29142 = NOR(g5535, g28010)
--	g14497 = NOR(g5990, g12705)
--	g30273 = NOR(g5990, g29036)
--	g30106 = NOR(g28739, g7268)
--	g12288 = NOR(g2610, g8418)
--	g29193 = NOR(g9529, g26994, g7812)
--	g19906 = NOR(g16209, g13672)
--	g12571 = NOR(g9511, g9451)
--	g12308 = NOR(g9951, g9954)
--	g25004 = NOR(g676, g23324)
--	g28496 = NOR(g3179, g27602)
--	g29165 = NOR(g5881, g28020)
--	g14339 = NOR(g12289, g2735)
--	g16072 = NOR(g10961, g13273)
--	g10338 = NOR(g5062, g5022)
--	g15062 = NOR(g6817, g13394)
--	g28986 = NOR(g5517, g28010)
--	g29006 = NOR(g5180, g27999)
--	g25947 = NOR(g1199, g24591)
--	g15508 = NOR(g10320, g14279)
--	g13959 = NOR(g3698, g11309)
--	g27954 = NOR(g10014, g25856)
--	g12752 = NOR(g9576, g9529)
--	g11958 = NOR(g9543, g7327)
--	g12374 = NOR(g2185, g8205)
--	g13378 = NOR(g11374, g11017)
--	g14411 = NOR(g9460, g11160)
--	g13603 = NOR(g8009, g10721)
--	g13944 = NOR(g10262, g12259)
--	g14867 = NOR(g10191, g12314)
--	g14450 = NOR(g12195, g9598)
--	g29175 = NOR(g6227, g26977)
--	g10819 = NOR(g7479, g1041)
--	g13730 = NOR(g3639, g11663)
--	g34359 = NOR(g9162, g34174, g12259)
--	g14707 = NOR(g10143, g12259)
--	g28457 = NOR(g7980, g27602)
--	g32212 = NOR(g8859, g31262, g11083)
--	g12558 = NOR(g7738, g5517, g5511)
--	g13765 = NOR(g8531, g11615)
--	g15051 = NOR(g6801, g13350)
--	g15072 = NOR(g13416, g12843)
--	g7192 = NOR(g6444, g6404)
--	g29873 = NOR(g6875, g28458)
--	g17180 = NOR(g1559, g13574)
--	g22993 = NOR(g1322, g16292, g19873)
--	g14094 = NOR(g8770, g11083)
--	g15152 = NOR(g13745, g12896)
--	g33109 = NOR(g31997, g4584)
--	g12189 = NOR(g1917, g8302)
--	g13129 = NOR(g7553, g10762)
--	g10801 = NOR(g1041, g7479)
--	g17694 = NOR(g12435, g12955)
--	g33108 = NOR(g32183, g31228)
--	g30134 = NOR(g28768, g7280)
--	g11626 = NOR(g7121, g3863, g3857)
--	g10695 = NOR(g8462, g8407)
--	g27093 = NOR(g26712, g26749)
--	g17619 = NOR(g10179, g12955)
--	g12093 = NOR(g9924, g7028)
--	g26649 = NOR(g9037, g24732)
--	g27875 = NOR(g9875, g25821)
--	g33174 = NOR(g8714, g32072)
--	g11232 = NOR(g4966, g7898, g9064)
--	g29034 = NOR(g5527, g28010)
--	g19400 = NOR(g17139, g14206)
--	g21127 = NOR(g18065, g12099)
--	g11697 = NOR(g8080, g3857)
--	g11995 = NOR(g9645, g7410)
--	g16027 = NOR(g10929, g13260)
--	g11261 = NOR(g7928, g4801, g9030)
--	g14001 = NOR(g739, g11083)
--	g30240 = NOR(g7004, g28982)
--	g24631 = NOR(g20516, g20436, g20219, g22957)
--	g12160 = NOR(g9721, g9724)
--	g13512 = NOR(g9077, g12527)
--	g28480 = NOR(g8059, g27602)
--	g23956 = NOR(g18957, g18918, g20136, g20114)
--	g8933 = NOR(g4709, g4785)
--	g31483 = NOR(g4899, g29725)
--	g13831 = NOR(g11245, g7666)
--	g12201 = NOR(g5417, g10047)
--	g29164 = NOR(g9444, g28010)
--	g12467 = NOR(g9472, g9407)
--	g30262 = NOR(g5644, g29008)
--	g13989 = NOR(g8697, g11309)
--	g13056 = NOR(g7400, g10741)
--	g16090 = NOR(g10961, g13315)
--	g26573 = NOR(g24897, g24884)
--	g11924 = NOR(g7187, g7209)
--	g29109 = NOR(g9472, g26994)
--	g27352 = NOR(g7975, g26616)
--	g26247 = NOR(g7995, g24732)
--	g7781 = NOR(g4064, g4057)
--	g12419 = NOR(g9402, g9326)
--	g25770 = NOR(g25417, g25377)
--	g29108 = NOR(g6219, g26977)
--	g24976 = NOR(g671, g23324)
--	g12418 = NOR(g9999, g10001)
--	g12170 = NOR(g10047, g5413)
--	g26098 = NOR(g9073, g24732)
--	g23024 = NOR(g7936, g19407)
--	g13342 = NOR(g10961, g10935)
--	g13031 = NOR(g7301, g10741)
--	g12853 = NOR(g6848, g10430)
--	g33851 = NOR(g8854, g33299, g12259)
--	g29174 = NOR(g9511, g28020)
--	g21250 = NOR(g9417, g9340, g17494)
--	g21658 = NOR(g17694, g17727)
--	g22654 = NOR(g7733, g19506)
--	g25521 = NOR(g23955, g14645)
--	g11869 = NOR(g7649, g7534, g7581)
--	g15647 = NOR(g11924, g14248)
--	g28469 = NOR(g3171, g27602)
--	g15090 = NOR(g13144, g12862)
--	g28468 = NOR(g3155, g10295, g27602)
--	g10341 = NOR(g6227, g6219)
--	g25247 = NOR(g23763, g14645)
--	g27704 = NOR(g7239, g25791)
--	g11225 = NOR(g3990, g6928)
--	g26162 = NOR(g23052, g24751)
--	g16646 = NOR(g13437, g11020, g11372)
--	g12466 = NOR(g10057, g10059)
--	g25777 = NOR(g25482, g25456)
--	g14335 = NOR(g12045, g9283)
--	g12101 = NOR(g6336, g7074)
--	g26628 = NOR(g8990, g24732)
--	g29040 = NOR(g6209, g26977)
--	g30162 = NOR(g28880, g7462)
--	g8864 = NOR(g3179, g3171)
--	g24383 = NOR(g22409, g22360)
--	g27733 = NOR(g9305, g25805)
--	g13970 = NOR(g8883, g8796, g11155)
--	g11171 = NOR(g8088, g9226, g9200, g9091)
--	g29183 = NOR(g9392, g28020, g7766)
--	g24875 = NOR(g8725, g23850, g11083)
--	g12166 = NOR(g9856, g10124)
--	g14278 = NOR(g562, g12259, g9217)
--	g13994 = NOR(g4049, g11363)
--	g15149 = NOR(g13745, g12894)
--	g25447 = NOR(g23883, g14645)
--	g14306 = NOR(g10060, g10887)
--	g29933 = NOR(g8808, g28500, g12259)
--	g15148 = NOR(g13716, g12893)
--	g15097 = NOR(g12868, g13191)
--	g30147 = NOR(g28768, g14567)
--	g13919 = NOR(g3347, g11276)
--	g9755 = NOR(g2070, g1996)
--	g13078 = NOR(g7446, g10762)
--	g23695 = NOR(g17420, g21140)
--	g19951 = NOR(g16219, g13709)
--	g25776 = NOR(g7166, g24380, g24369)
--	g25785 = NOR(g25488, g25462)
--	g10884 = NOR(g7650, g8451)
--	g27382 = NOR(g8219, g26657)
--	g28953 = NOR(g5170, g27999)
--	g24494 = NOR(g23513, g23532)
--	g15133 = NOR(g12883, g13638)
--	g32650 = NOR(g31579, I30192, I30193)
--	g13125 = NOR(g7863, g10762)
--	g10666 = NOR(g8462, g1171)
--	g25950 = NOR(g1070, g24591)
--	g7142 = NOR(g6573, g6565)
--	g12154 = NOR(g10155, g9835)
--	g29072 = NOR(g9402, g26977)
--	g9602 = NOR(g4688, g4681, g4674, g4646)
--	g14556 = NOR(g6682, g12790)
--	g26645 = NOR(g23602, g25160)
--	g13336 = NOR(g11330, g11011)
--	g21256 = NOR(g15483, g12179)
--	g22983 = NOR(g979, g16268, g19853)
--	g9015 = NOR(g3050, g3010)
--	g15050 = NOR(g12834, g13350)
--	g12729 = NOR(g1657, g8139)
--	g13631 = NOR(g8068, g10733)
--	g10922 = NOR(g7650, g4057)
--	g25446 = NOR(g23686, g14645)
--	g22517 = NOR(g19720, g1345)
--	g10179 = NOR(g2098, g1964, g1830, g1696)
--	g9664 = NOR(g4878, g4871, g4864, g4836)
--	g15096 = NOR(g13191, g12867)
--	g30146 = NOR(g28833, g7411)
--	g25540 = NOR(g22409, g22360)
--	g14178 = NOR(g8899, g11083)
--	g31482 = NOR(g8883, g29697)
--	g30290 = NOR(g6682, g29110)
--	g28568 = NOR(g10323, g27617)
--	g25203 = NOR(g6428, g23756)
--	g11309 = NOR(g8587, g8728)
--	g11571 = NOR(g10323, g3512, g3506)
--	g22523 = NOR(g1345, g19720)
--	g14417 = NOR(g12149, g9648)
--	g12622 = NOR(g9569, g9518)
--	g26715 = NOR(g23711, g25203)
--	g23763 = NOR(g2795, g21276)
--	g14334 = NOR(g12044, g9337)
--	g16232 = NOR(g13516, g4950)
--	g11976 = NOR(g9595, g7379)
--	g33090 = NOR(g31997, g4593)
--	g31233 = NOR(g8522, g29778, g24825)
--	g17727 = NOR(g12486, g12983)
--	g11954 = NOR(g9538, g7314)
--	g13954 = NOR(g8663, g11276)
--	g28510 = NOR(g3530, g27617)
--	g12333 = NOR(g1624, g8139)
--	g26297 = NOR(g8519, g24825)
--	g15129 = NOR(g6984, g13638)
--	g12852 = NOR(g6847, g10430)
--	g15057 = NOR(g6810, g13350)
--	g11669 = NOR(g3863, g8026)
--	g15128 = NOR(g13638, g12880)
--	g14000 = NOR(g8766, g12259)
--	g33449 = NOR(g10311, g31950)
--	g33448 = NOR(g7785, g31950)
--	g14568 = NOR(g12000, g9915)
--	g17175 = NOR(g1216, g13545)
--	g10123 = NOR(g4294, g4297)
--	g21655 = NOR(g17657, g17700)
--	g34354 = NOR(g9003, g34162, g11083)
--	g12609 = NOR(g7766, g5863, g5857)
--	g14751 = NOR(g10622, g10617, g10609, g10603)
--	g14772 = NOR(g6044, g12252)
--	g8182 = NOR(g405, g392)
--	g28493 = NOR(g3873, g27635)
--	g26546 = NOR(g24858, g24846)
--	g19981 = NOR(g3727, g16316)
--	g28340 = NOR(g27439, g26339)
--	g14416 = NOR(g12148, g9541)
--	g11610 = NOR(g7980, g3155)
--	g25784 = NOR(g25507, g25485)
--	g27973 = NOR(g7187, g25839)
--	g33148 = NOR(g4854, g32072)
--	g25956 = NOR(g1413, g24609)
--	g11255 = NOR(g8623, g6928)
--	g33097 = NOR(g31950, g4628)
--	g14391 = NOR(g12112, g9585)
--	g12798 = NOR(g5535, g9381)
--	g10510 = NOR(g7183, g4593, g4584)
--	g11270 = NOR(g8431, g8434)
--	g16198 = NOR(g9247, g13574)
--	g7352 = NOR(g1526, g1514)
--	g26625 = NOR(g23560, g25144)
--	g27732 = NOR(g9364, g25791)
--	g13939 = NOR(g4899, g8822, g11173)
--	g32017 = NOR(g31504, g23475)
--	g26296 = NOR(g8287, g24732)
--	g26338 = NOR(g8458, g24825)
--	g15056 = NOR(g6809, g13350)
--	g27400 = NOR(g8553, g26657)
--	g10615 = NOR(g1636, g7308)
--	g31133 = NOR(g7953, g29556)
--	g33133 = NOR(g32278, g31503)
--	g28475 = NOR(g3863, g27635)
--	g21143 = NOR(g15348, g9517)
--	g19388 = NOR(g17181, g14256)
--	g15145 = NOR(g12891, g13716)
--	g24439 = NOR(g7400, g22312)
--	g9700 = NOR(g2361, g2287)
--	g11201 = NOR(g4125, g7765)
--	g33112 = NOR(g31240, g32194)
--	g27771 = NOR(g9809, g25839)
--	g19140 = NOR(g7939, g15695)
--	g19997 = NOR(g16231, g13739)
--	g15132 = NOR(g12882, g13638)
--	g12235 = NOR(g9234, g9206)
--	g33096 = NOR(g31997, g4608)
--	g14362 = NOR(g12080, g9338)
--	g22537 = NOR(g19720, g1367)
--	g15161 = NOR(g13809, g7073)
--	g14165 = NOR(g8951, g11083)
--	g29104 = NOR(g5188, g27999)
--	g12515 = NOR(g9511, g5873)
--	g15087 = NOR(g12860, g13144)
--	g32424 = NOR(g8721, g31294)
--	g34496 = NOR(g34370, g27648)
--	g14437 = NOR(g9527, g11178)
--	g11194 = NOR(g3288, g6875)
--	g15069 = NOR(g6828, g13416)
--	g14347 = NOR(g9309, g11123)
--	g14253 = NOR(g10032, g12259, g9217)
--	g15068 = NOR(g6826, g13416)
--	g17174 = NOR(g9194, g14279)
--	g34067 = NOR(g33859, g11772)
--	g11119 = NOR(g9180, g9203)
--	g30150 = NOR(g28846, g7424)
--	g33129 = NOR(g8630, g32072)
--	g10821 = NOR(g7503, g1384)
--	g12435 = NOR(g9012, g8956, g8904, g8863)
--	g33128 = NOR(g4653, g32057)
--	g14821 = NOR(g6390, g12314)
--	g22522 = NOR(g19699, g1024)
--	g11313 = NOR(g8669, g3759)
--	g27345 = NOR(g9360, g26636)
--	g12744 = NOR(g9402, g6203)
--	g14516 = NOR(g12227, g9704)
--	g11276 = NOR(g8534, g8691)
--	g12849 = NOR(g6840, g10430)
--	g17663 = NOR(g10205, g12983)
--	g12848 = NOR(g6839, g10430)
--	g27652 = NOR(g3355, g26636)
--	g26256 = NOR(g23873, g25479)
--	g22536 = NOR(g1379, g19720)
--	g15086 = NOR(g13144, g12859)
--	g12361 = NOR(g6455, g10172)
--	g14726 = NOR(g10090, g12166)
--	g30280 = NOR(g7064, g29036)
--	g32455 = NOR(g31566, I29985, I29986)
--	g15159 = NOR(g13809, g12902)
--	g16288 = NOR(g13794, g417)
--	g14320 = NOR(g9257, g11111)
--	g15158 = NOR(g13782, g12901)
--	g30157 = NOR(g28833, g7369)
--	g14122 = NOR(g8895, g12259)
--	g15144 = NOR(g13716, g12890)
--	g31498 = NOR(g9030, g29540)
--	g28492 = NOR(g3857, g7121, g27635)
--	g8086 = NOR(g168, g174, g182)
--	g11907 = NOR(g7170, g7184)
--	g33432 = NOR(g31997, g6978)
--	g26314 = NOR(g24808, g24802)
--	g12371 = NOR(g1760, g8195)
--	g23835 = NOR(g2791, g21303)
--	g11238 = NOR(g8584, g6905)
--	g17213 = NOR(g11107, g13501)
--	g12234 = NOR(g9776, g9778)
--	g23586 = NOR(g17284, g20717)
--	g33145 = NOR(g8677, g32072)
--	g14164 = NOR(g9000, g12259)
--	g11185 = NOR(g8038, g8183, g6804)
--	g13518 = NOR(g3719, g11903)
--	g16488 = NOR(g13697, g13656)
--	g16424 = NOR(g8064, g13628)
--	g26268 = NOR(g283, g24825)
--	g14575 = NOR(g10050, g12749)
--	g11935 = NOR(g9485, g7267)
--	g8131 = NOR(g4776, g4801, g4793)
--	g27012 = NOR(g6398, g25856)
--	g13883 = NOR(g4709, g4785, g11155)
--	g33132 = NOR(g4843, g32072)
--	g12163 = NOR(g5073, g9989)
--	g28483 = NOR(g8080, g27635)
--	g26993 = NOR(g5360, g25805)
--	g33161 = NOR(g32090, g7806)
--	g26667 = NOR(g23642, g25175)
--	g30156 = NOR(g28789, g14587)
--	g11729 = NOR(g3179, g8059)
--	g13501 = NOR(g3368, g11881)
--	g27829 = NOR(g7345, g25856)
--	g14091 = NOR(g8854, g12259)
--	g27828 = NOR(g9892, g25856)
--	g22405 = NOR(g18957, g20136, g20114)
--	g15669 = NOR(g11945, g14272)
--	g12358 = NOR(g10019, g10022)
--	g27344 = NOR(g8390, g26636)
--	g12121 = NOR(g10117, g9762)
--	g21193 = NOR(g15348, g12135)
--	g22929 = NOR(g19773, g12970)
--	g31068 = NOR(g4801, g29540)
--	g11566 = NOR(g3161, g7964)
--	g13622 = NOR(g278, g11166)
--	g31970 = NOR(g9024, g30583)
--	g12173 = NOR(g10050, g7074)
--	g28509 = NOR(g8107, g27602)
--	g16219 = NOR(g13498, g4760)
--	g14522 = NOR(g9924, g12656)
--	g11653 = NOR(g7980, g7964)
--	g22357 = NOR(g1024, g19699)
--	g29145 = NOR(g6549, g7812, g26994)
--	g12029 = NOR(g5644, g7028)
--	g10862 = NOR(g7701, g7840)
--	g11415 = NOR(g8080, g8026)
--	g29198 = NOR(g7766, g28020)
--	g13852 = NOR(g11320, g8347)
--	g30601 = NOR(g16279, g29718)
--	g28452 = NOR(g3161, g27602)
--	g27927 = NOR(g9621, g25856)
--	g16201 = NOR(g13462, g4704)
--	g15093 = NOR(g13177, g6904)
--	g30143 = NOR(g28761, g14566)
--	g23063 = NOR(g16313, g19887)
--	g15065 = NOR(g13394, g12840)
--	g30169 = NOR(g28833, g14613)
--	g14397 = NOR(g12120, g9416)
--	g12604 = NOR(g5517, g9239)
--	g27770 = NOR(g9386, g25821)
--	g19338 = NOR(g16031, g1306)
--	g12755 = NOR(g6555, g9407)
--	g33125 = NOR(g8606, g32057)
--	g21209 = NOR(g15483, g9575)
--	g14872 = NOR(g6736, g12364)
--	g19968 = NOR(g17062, g11223)
--	g23208 = NOR(g20035, g16324)
--	g15160 = NOR(g12903, g13809)
--	g13799 = NOR(g8584, g11663)
--	g17482 = NOR(g9523, g14434)
--	g33144 = NOR(g4664, g32057)
--	g33823 = NOR(g8774, g33306, g11083)
--	g20234 = NOR(g17140, g14207)
--	g29069 = NOR(g9381, g28010)
--	g11184 = NOR(g513, g9040)
--	g7158 = NOR(g5752, g5712)
--	g10205 = NOR(g2657, g2523, g2389, g2255)
--	g24514 = NOR(g23619, g23657)
--	g30922 = NOR(g16662, g29810)
--	g29886 = NOR(g3288, g28458)
--	g11692 = NOR(g8021, g7985)
--	g16313 = NOR(g8005, g13600)
--	g27926 = NOR(g9467, g25856)
--	g13013 = NOR(g7957, g10762)
--	g19070 = NOR(g16957, g11720)
--	g22513 = NOR(g1002, g19699)
--	g15155 = NOR(g12899, g13782)
--	g11207 = NOR(g3639, g6905)
--	g15170 = NOR(g7118, g14279)
--	g22448 = NOR(g1018, g19699)
--	g13539 = NOR(g8594, g12735)
--	g13005 = NOR(g7939, g10762)
--	g25321 = NOR(g23835, g14645)
--	g14396 = NOR(g12119, g9489)
--	g14731 = NOR(g5698, g12204)
--	g15167 = NOR(g13835, g12908)
--	g14413 = NOR(g11914, g9638)
--	g28803 = NOR(g27730, g22763)
--	g11771 = NOR(g8921, g4185)
--	g25800 = NOR(g25518, g25510)
--	g27766 = NOR(g9716, g25791)
--	g23711 = NOR(g9892, g21253)
--	g30117 = NOR(g28739, g7252)
--	g29144 = NOR(g9518, g26977)
--	g19402 = NOR(g15979, g13133)
--	g23108 = NOR(g16424, g19932)
--	g17148 = NOR(g827, g14279)
--	g11414 = NOR(g8591, g8593)
--	g16476 = NOR(g8119, g13667)
--	g32585 = NOR(g31542, I30123, I30124)
--	g15053 = NOR(g12836, g13350)
--	g28482 = NOR(g3522, g27617)
--	g30123 = NOR(g28768, g7328)
--	g27629 = NOR(g8891, g26382, g12259)
--	g28552 = NOR(g10295, g27602)
--	g15101 = NOR(g12871, g14591)
--	g12246 = NOR(g9880, g9883)
--	g11584 = NOR(g8229, g8172)
--	g30265 = NOR(g7051, g29036)
--	g14640 = NOR(g12371, g9824)
--	g15064 = NOR(g6820, g13394)
--	g10803 = NOR(g1384, g7503)
--	g12591 = NOR(g504, g9040)
--	g12785 = NOR(g9472, g6549)
--	g27355 = NOR(g8443, g26657)
--	g13114 = NOR(g7528, g10741)
--	g27825 = NOR(g9316, g25821)
--	g11435 = NOR(g8107, g3171)
--	g11107 = NOR(g9095, g9177)
--	g15166 = NOR(g13835, g7096)
--	g12858 = NOR(g10365, g10430)
--	g11345 = NOR(g8477, g8479)
--	g33093 = NOR(g31997, g4601)
--	g31294 = NOR(g11326, g29660)
--	g11940 = NOR(g2712, g10084)
--	g27367 = NOR(g8155, g26636)
--	g14027 = NOR(g8734, g11363)
--	g11804 = NOR(g8938, g4975)
--	g15570 = NOR(g822, g14279)
--	g14248 = NOR(g6065, g10578)
--	g16215 = NOR(g1211, g13545)
--	g24990 = NOR(g8898, g23324)
--	g14003 = NOR(g9003, g11083)
--	g15074 = NOR(g12845, g13416)
--	g12318 = NOR(g10172, g6451)
--	g27059 = NOR(g7577, g25895)
--	g15594 = NOR(g10614, g13026, g7285)
--	g12059 = NOR(g9853, g7004)
--	g12025 = NOR(g9705, g7461)
--	g33160 = NOR(g8672, g32057)
--	g12540 = NOR(g2587, g8381)
--	g13500 = NOR(g8480, g12641)
--	g15092 = NOR(g12864, g13177)
--	g28149 = NOR(g27598, g27612)
--	g15154 = NOR(g13782, g12898)
--	g21062 = NOR(g9547, g17297)
--	g14090 = NOR(g8851, g12259)
--	g13004 = NOR(g7933, g10741)
--	g33075 = NOR(g31997, g7163)
--	g19268 = NOR(g15979, g962)
--	g12377 = NOR(g6856, g2748, g9708)
--	g12739 = NOR(g9321, g9274)
--	g30130 = NOR(g28761, g7275)
--	g24701 = NOR(g979, g23024, g19778)
--	g12146 = NOR(g1783, g8241)
--	g12645 = NOR(g4467, g6961)
--	g13947 = NOR(g8948, g11083)
--	g11273 = NOR(g3061, g8620)
--	g14513 = NOR(g12222, g9754)
--	g29705 = NOR(g28399, g8284, g8404)
--	g14449 = NOR(g12194, g9653)
--	g29189 = NOR(g9462, g26977, g7791)
--	g33419 = NOR(g31978, g7627)
--	g14448 = NOR(g12192, g9699)
--	g11972 = NOR(g9591, g7361)
--	g27366 = NOR(g8016, g26636)
--	g7567 = NOR(g979, g990)
--	g14212 = NOR(g5373, g10537)
--	g12632 = NOR(g9631, g6565)
--	g24766 = NOR(g3385, g23132)
--	g23051 = NOR(g7960, g19427)
--	g34703 = NOR(g8899, g34545, g11083)
--	g11514 = NOR(g10295, g3161, g3155)
--	g12226 = NOR(g2476, g8373)
--	g31119 = NOR(g7898, g29556)
--	g26873 = NOR(g25374, g25331)
--	g11012 = NOR(g7693, g7846)
--	g15139 = NOR(g12886, g13680)
--	g26209 = NOR(g23124, g24779)
--	g15138 = NOR(g13680, g6993)
--	g11473 = NOR(g8107, g8059)
--	g29915 = NOR(g6941, g28484)
--	g27354 = NOR(g8064, g26636)
--	g12297 = NOR(g9269, g9239)
--	g13325 = NOR(g7841, g10741)
--	g12980 = NOR(g7909, g10741)
--	g12824 = NOR(g5881, g9451)
--	g25952 = NOR(g1542, g24609)
--	g13946 = NOR(g8651, g11083)
--	g25175 = NOR(g5736, g23692)
--	g14228 = NOR(g5719, g10561)
--	g15585 = NOR(g11862, g14194)
--	g26346 = NOR(g8522, g24825)
--	g15608 = NOR(g11885, g14212)
--	g15052 = NOR(g12835, g13350)
--	g12211 = NOR(g10099, g7097)
--	g31008 = NOR(g30004, g30026)
--	g31476 = NOR(g4709, g29697)
--	g29167 = NOR(g9576, g26994)
--	g17198 = NOR(g9282, g14279)
--	g27659 = NOR(g3706, g26657)
--	g17393 = NOR(g9386, g14379)
--	g12700 = NOR(g9321, g5857)
--	g12659 = NOR(g9451, g9392)
--	g12126 = NOR(g9989, g5069)
--	g30136 = NOR(g28799, g7380)
--	g19953 = NOR(g16220, g13712)
--	g10793 = NOR(g1389, g7503)
--	g14793 = NOR(g2988, g12228)
--	g27338 = NOR(g9291, g26616)
--	g12296 = NOR(g9860, g9862)
--	g9762 = NOR(g2495, g2421)
--	g23662 = NOR(g17393, g20995)
--	g27969 = NOR(g7170, g25821)
--	g14549 = NOR(g9992, g12705)
--	g11755 = NOR(g4709, g8796)
--	g29900 = NOR(g3639, g28471)
--	g33092 = NOR(g31978, g4332)
--	g11563 = NOR(g8059, g8011)
--	g12855 = NOR(g10430, g6854)
--	g31935 = NOR(g30583, g4349)
--	g23204 = NOR(g10685, g19462, g16488)
--	g14002 = NOR(g8681, g11083)
--	g17657 = NOR(g14751, g12955)
--	g11191 = NOR(g4776, g4801, g9030)
--	g28498 = NOR(g8172, g27635)
--	g15100 = NOR(g13191, g12870)
--	g12581 = NOR(g9569, g6219)
--	g33439 = NOR(g31950, g4633)
--	g7175 = NOR(g6098, g6058)
--	g33438 = NOR(g31950, g4621)
--	g7139 = NOR(g5406, g5366)
--	g22545 = NOR(g1373, g19720)
--	g28031 = NOR(g21209, I26522, I26523)
--	g12067 = NOR(g5990, g7051)
--	g14512 = NOR(g11955, g9753)
--	g27735 = NOR(g7262, g25821)
--	g27877 = NOR(g9397, g25839)
--	g28529 = NOR(g8070, g27617, g10323)
--	g12150 = NOR(g2208, g8259)
--	g33139 = NOR(g8650, g32057)
--	g10831 = NOR(g7690, g7827)
--	g13032 = NOR(g7577, g10762)
--	g33138 = NOR(g32287, g31514)
--	g14445 = NOR(g12188, g9693)
--	g12695 = NOR(g9269, g9239)
--	g29675 = NOR(g28380, g8236, g8354)
--	g26183 = NOR(g23079, g24766)
--	g30252 = NOR(g7028, g29008)
--	g7304 = NOR(g1183, g1171)
--	g14611 = NOR(g12333, g9749)
--	g7499 = NOR(g333, g355)
--	g14988 = NOR(g10816, g10812, g10805)
--	g11360 = NOR(g3763, g8669)
--	g26872 = NOR(g25411, g25371)
--	g14271 = NOR(g10002, g10874)
--	g30183 = NOR(g28880, g14644)
--	g19430 = NOR(g17150, g14220)
--	g15141 = NOR(g12888, g13680)
--	g14145 = NOR(g8945, g12259)
--	g12256 = NOR(g10136, g6105)
--	g25948 = NOR(g7752, g24609)
--	g24497 = NOR(g23533, g23553)
--	g14529 = NOR(g6336, g12749)
--	g27102 = NOR(g26750, g26779)
--	g15135 = NOR(g6990, g13638)
--	g26574 = NOR(g24887, g24861)
--	g14393 = NOR(g12115, g9488)
--	g14365 = NOR(g12084, g9339)
--	g32845 = NOR(g30673, I30399, I30400)
--	g17309 = NOR(g9305, g14344)
--	g15049 = NOR(g13350, g6799)
--	g11950 = NOR(g9220, g9166)
--	g10709 = NOR(g7499, g351)
--	g27511 = NOR(g22137, g26866, g20277)
--	g12854 = NOR(g6849, g10430)
--	g28425 = NOR(g27493, g26351)
--	g34912 = NOR(g34883, g20277, g20242, g21370)
--	g25851 = NOR(g4311, g24380, g24369)
--	g13996 = NOR(g8938, g8822, g11173)
--	g28444 = NOR(g8575, g27463, g24825)
--	g15106 = NOR(g12872, g10430)
--	g17954 = NOR(g832, g14279)
--	g12550 = NOR(g9300, g9259)
--	g12314 = NOR(g10053, g10207)
--	g14602 = NOR(g10099, g12790)
--	g27721 = NOR(g9672, g25805)
--	g12085 = NOR(g10082, g9700)
--	g22488 = NOR(g19699, g1002)
--	g14337 = NOR(g12049, g9284)
--	g11203 = NOR(g4966, g4991, g9064)
--	g13044 = NOR(g7349, g10762)
--	g14792 = NOR(g10653, g10623, g10618, g10611)
--	g28353 = NOR(g9073, g27654, g24732)
--	g29200 = NOR(g7791, g26977)
--	g9640 = NOR(g1802, g1728)
--	g19063 = NOR(g7909, g15674)
--	g33100 = NOR(g32172, g31188)
--	g13377 = NOR(g7873, g10762)
--	g14425 = NOR(g5644, g12656)
--	g27734 = NOR(g9733, g25821)
--	g15163 = NOR(g13809, g12905)
--	g30929 = NOR(g29803, g29835)
--	g19873 = NOR(g15755, g1395)
--	g10918 = NOR(g1532, g7751, g7778)
--	g19422 = NOR(g16031, g13141)
--	g14444 = NOR(g11936, g9692)
--	g12667 = NOR(g7791, g6209, g6203)
--	g19209 = NOR(g12971, g15614, g11320)
--	g13698 = NOR(g528, g12527, g11185)
--	g31515 = NOR(g4983, g29556)
--	g29184 = NOR(g9631, g26994)
--	g23626 = NOR(g17309, g20854)
--	g15724 = NOR(g13858, g11374)
--	g24018 = NOR(I23162, I23163)
--	g30282 = NOR(g6336, g29073)
--	g19453 = NOR(g17199, g14316)
--	g15121 = NOR(g12874, g13605)
--	g12443 = NOR(g9374, g9300)
--	g19436 = NOR(g17176, g14233)
--	g13661 = NOR(g528, g11185)
--	g11715 = NOR(g8080, g8026)
--	g29005 = NOR(g5164, g7704, g27999)
--	g33107 = NOR(g32180, g31223)
--	g12601 = NOR(g9381, g9311)
--	g15134 = NOR(g13638, g12884)
--	g14364 = NOR(g12083, g9415)
--	g25769 = NOR(g25453, g25414)
--	g11385 = NOR(g8021, g7985)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s38584 is
	port (
		CLK: in std_logic;
		G5: in std_logic;
		G35: in std_logic;
		G36: in std_logic;
		G44: in std_logic;
		G53: in std_logic;
		G54: in std_logic;
		G56: in std_logic;
		G57: in std_logic;
		G64: in std_logic;
		G72: in std_logic;
		G73: in std_logic;
		G84: in std_logic;
		G90: in std_logic;
		G91: in std_logic;
		G92: in std_logic;
		G99: in std_logic;
		G100: in std_logic;
		G113: in std_logic;
		G114: in std_logic;
		G115: in std_logic;
		G116: in std_logic;
		G120: in std_logic;
		G124: in std_logic;
		G125: in std_logic;
		G126: in std_logic;
		G127: in std_logic;
		G134: in std_logic;
		G135: in std_logic;
		G6744: in std_logic;
		G6745: in std_logic;
		G6746: in std_logic;
		G6747: in std_logic;
		G6748: in std_logic;
		G6749: in std_logic;
		G6750: in std_logic;
		G6751: in std_logic;
		G6752: in std_logic;
		G6753: in std_logic;
		G7243: out std_logic;
		G7245: out std_logic;
		G7257: out std_logic;
		G7260: out std_logic;
		G7540: out std_logic;
		G7916: out std_logic;
		G7946: out std_logic;
		G8132: out std_logic;
		G8178: out std_logic;
		G8215: out std_logic;
		G8235: out std_logic;
		G8277: out std_logic;
		G8279: out std_logic;
		G8283: out std_logic;
		G8291: out std_logic;
		G8342: out std_logic;
		G8344: out std_logic;
		G8353: out std_logic;
		G8358: out std_logic;
		G8398: out std_logic;
		G8403: out std_logic;
		G8416: out std_logic;
		G8475: out std_logic;
		G8719: out std_logic;
		G8783: out std_logic;
		G8784: out std_logic;
		G8785: out std_logic;
		G8786: out std_logic;
		G8787: out std_logic;
		G8788: out std_logic;
		G8789: out std_logic;
		G8839: out std_logic;
		G8870: out std_logic;
		G8915: out std_logic;
		G8916: out std_logic;
		G8917: out std_logic;
		G8918: out std_logic;
		G8919: out std_logic;
		G8920: out std_logic;
		G9019: out std_logic;
		G9048: out std_logic;
		G9251: out std_logic;
		G9497: out std_logic;
		G9553: out std_logic;
		G9555: out std_logic;
		G9615: out std_logic;
		G9617: out std_logic;
		G9680: out std_logic;
		G9682: out std_logic;
		G9741: out std_logic;
		G9743: out std_logic;
		G9817: out std_logic;
		G10122: out std_logic;
		G10306: out std_logic;
		G10500: out std_logic;
		G10527: out std_logic;
		G11349: out std_logic;
		G11388: out std_logic;
		G11418: out std_logic;
		G11447: out std_logic;
		G11678: out std_logic;
		G11770: out std_logic;
		G12184: out std_logic;
		G12238: out std_logic;
		G12300: out std_logic;
		G12350: out std_logic;
		G12368: out std_logic;
		G12422: out std_logic;
		G12470: out std_logic;
		G12832: out std_logic;
		G12833: out std_logic;
		G12919: out std_logic;
		G12923: out std_logic;
		G13039: out std_logic;
		G13049: out std_logic;
		G13068: out std_logic;
		G13085: out std_logic;
		G13099: out std_logic;
		G13259: out std_logic;
		G13272: out std_logic;
		G13865: out std_logic;
		G13881: out std_logic;
		G13895: out std_logic;
		G13906: out std_logic;
		G13926: out std_logic;
		G13966: out std_logic;
		G14096: out std_logic;
		G14125: out std_logic;
		G14147: out std_logic;
		G14167: out std_logic;
		G14189: out std_logic;
		G14201: out std_logic;
		G14217: out std_logic;
		G14421: out std_logic;
		G14451: out std_logic;
		G14518: out std_logic;
		G14597: out std_logic;
		G14635: out std_logic;
		G14662: out std_logic;
		G14673: out std_logic;
		G14694: out std_logic;
		G14705: out std_logic;
		G14738: out std_logic;
		G14749: out std_logic;
		G14779: out std_logic;
		G14828: out std_logic;
		G16603: out std_logic;
		G16624: out std_logic;
		G16627: out std_logic;
		G16656: out std_logic;
		G16659: out std_logic;
		G16686: out std_logic;
		G16693: out std_logic;
		G16718: out std_logic;
		G16722: out std_logic;
		G16744: out std_logic;
		G16748: out std_logic;
		G16775: out std_logic;
		G16874: out std_logic;
		G16924: out std_logic;
		G16955: out std_logic;
		G17291: out std_logic;
		G17316: out std_logic;
		G17320: out std_logic;
		G17400: out std_logic;
		G17404: out std_logic;
		G17423: out std_logic;
		G17519: out std_logic;
		G17577: out std_logic;
		G17580: out std_logic;
		G17604: out std_logic;
		G17607: out std_logic;
		G17639: out std_logic;
		G17646: out std_logic;
		G17649: out std_logic;
		G17674: out std_logic;
		G17678: out std_logic;
		G17685: out std_logic;
		G17688: out std_logic;
		G17711: out std_logic;
		G17715: out std_logic;
		G17722: out std_logic;
		G17739: out std_logic;
		G17743: out std_logic;
		G17760: out std_logic;
		G17764: out std_logic;
		G17778: out std_logic;
		G17787: out std_logic;
		G17813: out std_logic;
		G17819: out std_logic;
		G17845: out std_logic;
		G17871: out std_logic;
		G18092: out std_logic;
		G18094: out std_logic;
		G18095: out std_logic;
		G18096: out std_logic;
		G18097: out std_logic;
		G18098: out std_logic;
		G18099: out std_logic;
		G18100: out std_logic;
		G18101: out std_logic;
		G18881: out std_logic;
		G19334: out std_logic;
		G19357: out std_logic;
		G20049: out std_logic;
		G20557: out std_logic;
		G20652: out std_logic;
		G20654: out std_logic;
		G20763: out std_logic;
		G20899: out std_logic;
		G20901: out std_logic;
		G21176: out std_logic;
		G21245: out std_logic;
		G21270: out std_logic;
		G21292: out std_logic;
		G21698: out std_logic;
		G21727: out std_logic;
		G23002: out std_logic;
		G23190: out std_logic;
		G23612: out std_logic;
		G23652: out std_logic;
		G23683: out std_logic;
		G23759: out std_logic;
		G24151: out std_logic;
		G24161: out std_logic;
		G24162: out std_logic;
		G24163: out std_logic;
		G24164: out std_logic;
		G24165: out std_logic;
		G24166: out std_logic;
		G24167: out std_logic;
		G24168: out std_logic;
		G24169: out std_logic;
		G24170: out std_logic;
		G24171: out std_logic;
		G24172: out std_logic;
		G24173: out std_logic;
		G24174: out std_logic;
		G24175: out std_logic;
		G24176: out std_logic;
		G24177: out std_logic;
		G24178: out std_logic;
		G24179: out std_logic;
		G24180: out std_logic;
		G24181: out std_logic;
		G24182: out std_logic;
		G24183: out std_logic;
		G24184: out std_logic;
		G24185: out std_logic;
		G25114: out std_logic;
		G25167: out std_logic;
		G25219: out std_logic;
		G25259: out std_logic;
		G25582: out std_logic;
		G25583: out std_logic;
		G25584: out std_logic;
		G25585: out std_logic;
		G25586: out std_logic;
		G25587: out std_logic;
		G25588: out std_logic;
		G25589: out std_logic;
		G25590: out std_logic;
		G26801: out std_logic;
		G26875: out std_logic;
		G26876: out std_logic;
		G26877: out std_logic;
		G27831: out std_logic;
		G28030: out std_logic;
		G28041: out std_logic;
		G28042: out std_logic;
		G28753: out std_logic;
		G29210: out std_logic;
		G29211: out std_logic;
		G29212: out std_logic;
		G29213: out std_logic;
		G29214: out std_logic;
		G29215: out std_logic;
		G29216: out std_logic;
		G29217: out std_logic;
		G29218: out std_logic;
		G29219: out std_logic;
		G29220: out std_logic;
		G29221: out std_logic;
		G30327: out std_logic;
		G30329: out std_logic;
		G30330: out std_logic;
		G30331: out std_logic;
		G30332: out std_logic;
		G31521: out std_logic;
		G31656: out std_logic;
		G31665: out std_logic;
		G31793: out std_logic;
		G31860: out std_logic;
		G31861: out std_logic;
		G31862: out std_logic;
		G31863: out std_logic;
		G32185: out std_logic;
		G32429: out std_logic;
		G32454: out std_logic;
		G32975: out std_logic;
		G33079: out std_logic;
		G33435: out std_logic;
		G33533: out std_logic;
		G33636: out std_logic;
		G33659: out std_logic;
		G33874: out std_logic;
		G33894: out std_logic;
		G33935: out std_logic;
		G33945: out std_logic;
		G33946: out std_logic;
		G33947: out std_logic;
		G33948: out std_logic;
		G33949: out std_logic;
		G33950: out std_logic;
		G33959: out std_logic;
		G34201: out std_logic;
		G34221: out std_logic;
		G34232: out std_logic;
		G34233: out std_logic;
		G34234: out std_logic;
		G34235: out std_logic;
		G34236: out std_logic;
		G34237: out std_logic;
		G34238: out std_logic;
		G34239: out std_logic;
		G34240: out std_logic;
		G34383: out std_logic;
		G34425: out std_logic;
		G34435: out std_logic;
		G34436: out std_logic;
		G34437: out std_logic;
		G34597: out std_logic;
		G34788: out std_logic;
		G34839: out std_logic;
		G34913: out std_logic;
		G34915: out std_logic;
		G34917: out std_logic;
		G34919: out std_logic;
		G34921: out std_logic;
		G34923: out std_logic;
		G34925: out std_logic;
		G34927: out std_logic;
		G34956: out std_logic;
		G34972: out std_logic
	);
end entity;

architecture RTL of s38584 is
	attribute dont_touch: boolean;

	signal G1: std_logic; attribute dont_touch of G1: signal is true;
	signal G6: std_logic; attribute dont_touch of G6: signal is true;
	signal G7: std_logic; attribute dont_touch of G7: signal is true;
	signal G8: std_logic; attribute dont_touch of G8: signal is true;
	signal G9: std_logic; attribute dont_touch of G9: signal is true;
	signal G12: std_logic; attribute dont_touch of G12: signal is true;
	signal G16: std_logic; attribute dont_touch of G16: signal is true;
	signal G19: std_logic; attribute dont_touch of G19: signal is true;
	signal G22: std_logic; attribute dont_touch of G22: signal is true;
	signal G25: std_logic; attribute dont_touch of G25: signal is true;
	signal G28: std_logic; attribute dont_touch of G28: signal is true;
	signal G31: std_logic; attribute dont_touch of G31: signal is true;
	signal G34: std_logic; attribute dont_touch of G34: signal is true;
	signal G37: std_logic; attribute dont_touch of G37: signal is true;
	signal G43: std_logic; attribute dont_touch of G43: signal is true;
	signal G45: std_logic; attribute dont_touch of G45: signal is true;
	signal G46: std_logic; attribute dont_touch of G46: signal is true;
	signal G47: std_logic; attribute dont_touch of G47: signal is true;
	signal G48: std_logic; attribute dont_touch of G48: signal is true;
	signal G49: std_logic; attribute dont_touch of G49: signal is true;
	signal G50: std_logic; attribute dont_touch of G50: signal is true;
	signal G51: std_logic; attribute dont_touch of G51: signal is true;
	signal G52: std_logic; attribute dont_touch of G52: signal is true;
	signal G55: std_logic; attribute dont_touch of G55: signal is true;
	signal G58: std_logic; attribute dont_touch of G58: signal is true;
	signal G59: std_logic; attribute dont_touch of G59: signal is true;
	signal G63: std_logic; attribute dont_touch of G63: signal is true;
	signal G65: std_logic; attribute dont_touch of G65: signal is true;
	signal G66: std_logic; attribute dont_touch of G66: signal is true;
	signal G70: std_logic; attribute dont_touch of G70: signal is true;
	signal G71: std_logic; attribute dont_touch of G71: signal is true;
	signal G74: std_logic; attribute dont_touch of G74: signal is true;
	signal G79: std_logic; attribute dont_touch of G79: signal is true;
	signal G85: std_logic; attribute dont_touch of G85: signal is true;
	signal G86: std_logic; attribute dont_touch of G86: signal is true;
	signal G93: std_logic; attribute dont_touch of G93: signal is true;
	signal G94: std_logic; attribute dont_touch of G94: signal is true;
	signal G101: std_logic; attribute dont_touch of G101: signal is true;
	signal G102: std_logic; attribute dont_touch of G102: signal is true;
	signal G106: std_logic; attribute dont_touch of G106: signal is true;
	signal G110: std_logic; attribute dont_touch of G110: signal is true;
	signal G111: std_logic; attribute dont_touch of G111: signal is true;
	signal G112: std_logic; attribute dont_touch of G112: signal is true;
	signal G117: std_logic; attribute dont_touch of G117: signal is true;
	signal G121: std_logic; attribute dont_touch of G121: signal is true;
	signal G128: std_logic; attribute dont_touch of G128: signal is true;
	signal G136: std_logic; attribute dont_touch of G136: signal is true;
	signal G142: std_logic; attribute dont_touch of G142: signal is true;
	signal G146: std_logic; attribute dont_touch of G146: signal is true;
	signal G150: std_logic; attribute dont_touch of G150: signal is true;
	signal G153: std_logic; attribute dont_touch of G153: signal is true;
	signal G157: std_logic; attribute dont_touch of G157: signal is true;
	signal G160: std_logic; attribute dont_touch of G160: signal is true;
	signal G164: std_logic; attribute dont_touch of G164: signal is true;
	signal G168: std_logic; attribute dont_touch of G168: signal is true;
	signal G174: std_logic; attribute dont_touch of G174: signal is true;
	signal G182: std_logic; attribute dont_touch of G182: signal is true;
	signal G191: std_logic; attribute dont_touch of G191: signal is true;
	signal G194: std_logic; attribute dont_touch of G194: signal is true;
	signal G199: std_logic; attribute dont_touch of G199: signal is true;
	signal G203: std_logic; attribute dont_touch of G203: signal is true;
	signal G209: std_logic; attribute dont_touch of G209: signal is true;
	signal G215: std_logic; attribute dont_touch of G215: signal is true;
	signal G218: std_logic; attribute dont_touch of G218: signal is true;
	signal G222: std_logic; attribute dont_touch of G222: signal is true;
	signal G225: std_logic; attribute dont_touch of G225: signal is true;
	signal G232: std_logic; attribute dont_touch of G232: signal is true;
	signal G239: std_logic; attribute dont_touch of G239: signal is true;
	signal G246: std_logic; attribute dont_touch of G246: signal is true;
	signal G255: std_logic; attribute dont_touch of G255: signal is true;
	signal G262: std_logic; attribute dont_touch of G262: signal is true;
	signal G269: std_logic; attribute dont_touch of G269: signal is true;
	signal G278: std_logic; attribute dont_touch of G278: signal is true;
	signal G283: std_logic; attribute dont_touch of G283: signal is true;
	signal G287: std_logic; attribute dont_touch of G287: signal is true;
	signal G291: std_logic; attribute dont_touch of G291: signal is true;
	signal G294: std_logic; attribute dont_touch of G294: signal is true;
	signal G298: std_logic; attribute dont_touch of G298: signal is true;
	signal G301: std_logic; attribute dont_touch of G301: signal is true;
	signal G305: std_logic; attribute dont_touch of G305: signal is true;
	signal G311: std_logic; attribute dont_touch of G311: signal is true;
	signal G316: std_logic; attribute dont_touch of G316: signal is true;
	signal G319: std_logic; attribute dont_touch of G319: signal is true;
	signal G324: std_logic; attribute dont_touch of G324: signal is true;
	signal G329: std_logic; attribute dont_touch of G329: signal is true;
	signal G333: std_logic; attribute dont_touch of G333: signal is true;
	signal G336: std_logic; attribute dont_touch of G336: signal is true;
	signal G341: std_logic; attribute dont_touch of G341: signal is true;
	signal G344: std_logic; attribute dont_touch of G344: signal is true;
	signal G347: std_logic; attribute dont_touch of G347: signal is true;
	signal G351: std_logic; attribute dont_touch of G351: signal is true;
	signal G355: std_logic; attribute dont_touch of G355: signal is true;
	signal G358: std_logic; attribute dont_touch of G358: signal is true;
	signal G365: std_logic; attribute dont_touch of G365: signal is true;
	signal G370: std_logic; attribute dont_touch of G370: signal is true;
	signal G376: std_logic; attribute dont_touch of G376: signal is true;
	signal G385: std_logic; attribute dont_touch of G385: signal is true;
	signal G391: std_logic; attribute dont_touch of G391: signal is true;
	signal G392: std_logic; attribute dont_touch of G392: signal is true;
	signal G401: std_logic; attribute dont_touch of G401: signal is true;
	signal G405: std_logic; attribute dont_touch of G405: signal is true;
	signal G411: std_logic; attribute dont_touch of G411: signal is true;
	signal G417: std_logic; attribute dont_touch of G417: signal is true;
	signal G424: std_logic; attribute dont_touch of G424: signal is true;
	signal G429: std_logic; attribute dont_touch of G429: signal is true;
	signal G433: std_logic; attribute dont_touch of G433: signal is true;
	signal G437: std_logic; attribute dont_touch of G437: signal is true;
	signal G441: std_logic; attribute dont_touch of G441: signal is true;
	signal G446: std_logic; attribute dont_touch of G446: signal is true;
	signal G452: std_logic; attribute dont_touch of G452: signal is true;
	signal G457: std_logic; attribute dont_touch of G457: signal is true;
	signal G460: std_logic; attribute dont_touch of G460: signal is true;
	signal G464: std_logic; attribute dont_touch of G464: signal is true;
	signal G468: std_logic; attribute dont_touch of G468: signal is true;
	signal G471: std_logic; attribute dont_touch of G471: signal is true;
	signal G475: std_logic; attribute dont_touch of G475: signal is true;
	signal G479: std_logic; attribute dont_touch of G479: signal is true;
	signal G482: std_logic; attribute dont_touch of G482: signal is true;
	signal G490: std_logic; attribute dont_touch of G490: signal is true;
	signal G496: std_logic; attribute dont_touch of G496: signal is true;
	signal G499: std_logic; attribute dont_touch of G499: signal is true;
	signal G504: std_logic; attribute dont_touch of G504: signal is true;
	signal G513: std_logic; attribute dont_touch of G513: signal is true;
	signal G518: std_logic; attribute dont_touch of G518: signal is true;
	signal G528: std_logic; attribute dont_touch of G528: signal is true;
	signal G534: std_logic; attribute dont_touch of G534: signal is true;
	signal G538: std_logic; attribute dont_touch of G538: signal is true;
	signal G542: std_logic; attribute dont_touch of G542: signal is true;
	signal G546: std_logic; attribute dont_touch of G546: signal is true;
	signal G550: std_logic; attribute dont_touch of G550: signal is true;
	signal G554: std_logic; attribute dont_touch of G554: signal is true;
	signal G559: std_logic; attribute dont_touch of G559: signal is true;
	signal G562: std_logic; attribute dont_touch of G562: signal is true;
	signal G568: std_logic; attribute dont_touch of G568: signal is true;
	signal G572: std_logic; attribute dont_touch of G572: signal is true;
	signal G577: std_logic; attribute dont_touch of G577: signal is true;
	signal G582: std_logic; attribute dont_touch of G582: signal is true;
	signal G586: std_logic; attribute dont_touch of G586: signal is true;
	signal G590: std_logic; attribute dont_touch of G590: signal is true;
	signal G595: std_logic; attribute dont_touch of G595: signal is true;
	signal G599: std_logic; attribute dont_touch of G599: signal is true;
	signal G604: std_logic; attribute dont_touch of G604: signal is true;
	signal G608: std_logic; attribute dont_touch of G608: signal is true;
	signal G613: std_logic; attribute dont_touch of G613: signal is true;
	signal G617: std_logic; attribute dont_touch of G617: signal is true;
	signal G622: std_logic; attribute dont_touch of G622: signal is true;
	signal G626: std_logic; attribute dont_touch of G626: signal is true;
	signal G632: std_logic; attribute dont_touch of G632: signal is true;
	signal G637: std_logic; attribute dont_touch of G637: signal is true;
	signal G640: std_logic; attribute dont_touch of G640: signal is true;
	signal G645: std_logic; attribute dont_touch of G645: signal is true;
	signal G650: std_logic; attribute dont_touch of G650: signal is true;
	signal G655: std_logic; attribute dont_touch of G655: signal is true;
	signal G661: std_logic; attribute dont_touch of G661: signal is true;
	signal G667: std_logic; attribute dont_touch of G667: signal is true;
	signal G671: std_logic; attribute dont_touch of G671: signal is true;
	signal G676: std_logic; attribute dont_touch of G676: signal is true;
	signal G681: std_logic; attribute dont_touch of G681: signal is true;
	signal G686: std_logic; attribute dont_touch of G686: signal is true;
	signal G691: std_logic; attribute dont_touch of G691: signal is true;
	signal G699: std_logic; attribute dont_touch of G699: signal is true;
	signal G703: std_logic; attribute dont_touch of G703: signal is true;
	signal G714: std_logic; attribute dont_touch of G714: signal is true;
	signal G718: std_logic; attribute dont_touch of G718: signal is true;
	signal G723: std_logic; attribute dont_touch of G723: signal is true;
	signal G728: std_logic; attribute dont_touch of G728: signal is true;
	signal G732: std_logic; attribute dont_touch of G732: signal is true;
	signal G736: std_logic; attribute dont_touch of G736: signal is true;
	signal G739: std_logic; attribute dont_touch of G739: signal is true;
	signal G744: std_logic; attribute dont_touch of G744: signal is true;
	signal G749: std_logic; attribute dont_touch of G749: signal is true;
	signal G753: std_logic; attribute dont_touch of G753: signal is true;
	signal G758: std_logic; attribute dont_touch of G758: signal is true;
	signal G763: std_logic; attribute dont_touch of G763: signal is true;
	signal G767: std_logic; attribute dont_touch of G767: signal is true;
	signal G772: std_logic; attribute dont_touch of G772: signal is true;
	signal G776: std_logic; attribute dont_touch of G776: signal is true;
	signal G781: std_logic; attribute dont_touch of G781: signal is true;
	signal G785: std_logic; attribute dont_touch of G785: signal is true;
	signal G790: std_logic; attribute dont_touch of G790: signal is true;
	signal G794: std_logic; attribute dont_touch of G794: signal is true;
	signal G799: std_logic; attribute dont_touch of G799: signal is true;
	signal G802: std_logic; attribute dont_touch of G802: signal is true;
	signal G807: std_logic; attribute dont_touch of G807: signal is true;
	signal G812: std_logic; attribute dont_touch of G812: signal is true;
	signal G817: std_logic; attribute dont_touch of G817: signal is true;
	signal G822: std_logic; attribute dont_touch of G822: signal is true;
	signal G827: std_logic; attribute dont_touch of G827: signal is true;
	signal G832: std_logic; attribute dont_touch of G832: signal is true;
	signal G837: std_logic; attribute dont_touch of G837: signal is true;
	signal G843: std_logic; attribute dont_touch of G843: signal is true;
	signal G847: std_logic; attribute dont_touch of G847: signal is true;
	signal G854: std_logic; attribute dont_touch of G854: signal is true;
	signal G859: std_logic; attribute dont_touch of G859: signal is true;
	signal G862: std_logic; attribute dont_touch of G862: signal is true;
	signal G869: std_logic; attribute dont_touch of G869: signal is true;
	signal G872: std_logic; attribute dont_touch of G872: signal is true;
	signal G875: std_logic; attribute dont_touch of G875: signal is true;
	signal G878: std_logic; attribute dont_touch of G878: signal is true;
	signal G881: std_logic; attribute dont_touch of G881: signal is true;
	signal G884: std_logic; attribute dont_touch of G884: signal is true;
	signal G887: std_logic; attribute dont_touch of G887: signal is true;
	signal G890: std_logic; attribute dont_touch of G890: signal is true;
	signal G896: std_logic; attribute dont_touch of G896: signal is true;
	signal G901: std_logic; attribute dont_touch of G901: signal is true;
	signal G904: std_logic; attribute dont_touch of G904: signal is true;
	signal G907: std_logic; attribute dont_touch of G907: signal is true;
	signal G911: std_logic; attribute dont_touch of G911: signal is true;
	signal G914: std_logic; attribute dont_touch of G914: signal is true;
	signal G918: std_logic; attribute dont_touch of G918: signal is true;
	signal G921: std_logic; attribute dont_touch of G921: signal is true;
	signal G925: std_logic; attribute dont_touch of G925: signal is true;
	signal G929: std_logic; attribute dont_touch of G929: signal is true;
	signal G930: std_logic; attribute dont_touch of G930: signal is true;
	signal G933: std_logic; attribute dont_touch of G933: signal is true;
	signal G936: std_logic; attribute dont_touch of G936: signal is true;
	signal G939: std_logic; attribute dont_touch of G939: signal is true;
	signal G943: std_logic; attribute dont_touch of G943: signal is true;
	signal G947: std_logic; attribute dont_touch of G947: signal is true;
	signal G952: std_logic; attribute dont_touch of G952: signal is true;
	signal G956: std_logic; attribute dont_touch of G956: signal is true;
	signal G962: std_logic; attribute dont_touch of G962: signal is true;
	signal G967: std_logic; attribute dont_touch of G967: signal is true;
	signal G968: std_logic; attribute dont_touch of G968: signal is true;
	signal G969: std_logic; attribute dont_touch of G969: signal is true;
	signal G976: std_logic; attribute dont_touch of G976: signal is true;
	signal G979: std_logic; attribute dont_touch of G979: signal is true;
	signal G990: std_logic; attribute dont_touch of G990: signal is true;
	signal G996: std_logic; attribute dont_touch of G996: signal is true;
	signal G1002: std_logic; attribute dont_touch of G1002: signal is true;
	signal G1008: std_logic; attribute dont_touch of G1008: signal is true;
	signal G1018: std_logic; attribute dont_touch of G1018: signal is true;
	signal G1024: std_logic; attribute dont_touch of G1024: signal is true;
	signal G1030: std_logic; attribute dont_touch of G1030: signal is true;
	signal G1036: std_logic; attribute dont_touch of G1036: signal is true;
	signal G1041: std_logic; attribute dont_touch of G1041: signal is true;
	signal G1046: std_logic; attribute dont_touch of G1046: signal is true;
	signal G1052: std_logic; attribute dont_touch of G1052: signal is true;
	signal G1056: std_logic; attribute dont_touch of G1056: signal is true;
	signal G1061: std_logic; attribute dont_touch of G1061: signal is true;
	signal G1070: std_logic; attribute dont_touch of G1070: signal is true;
	signal G1075: std_logic; attribute dont_touch of G1075: signal is true;
	signal G1079: std_logic; attribute dont_touch of G1079: signal is true;
	signal G1083: std_logic; attribute dont_touch of G1083: signal is true;
	signal G1087: std_logic; attribute dont_touch of G1087: signal is true;
	signal G1094: std_logic; attribute dont_touch of G1094: signal is true;
	signal G1099: std_logic; attribute dont_touch of G1099: signal is true;
	signal G1105: std_logic; attribute dont_touch of G1105: signal is true;
	signal G1111: std_logic; attribute dont_touch of G1111: signal is true;
	signal G1116: std_logic; attribute dont_touch of G1116: signal is true;
	signal G1124: std_logic; attribute dont_touch of G1124: signal is true;
	signal G1129: std_logic; attribute dont_touch of G1129: signal is true;
	signal G1135: std_logic; attribute dont_touch of G1135: signal is true;
	signal G1141: std_logic; attribute dont_touch of G1141: signal is true;
	signal G1146: std_logic; attribute dont_touch of G1146: signal is true;
	signal G1152: std_logic; attribute dont_touch of G1152: signal is true;
	signal G1157: std_logic; attribute dont_touch of G1157: signal is true;
	signal G1171: std_logic; attribute dont_touch of G1171: signal is true;
	signal G1178: std_logic; attribute dont_touch of G1178: signal is true;
	signal G1183: std_logic; attribute dont_touch of G1183: signal is true;
	signal G1189: std_logic; attribute dont_touch of G1189: signal is true;
	signal G1193: std_logic; attribute dont_touch of G1193: signal is true;
	signal G1199: std_logic; attribute dont_touch of G1199: signal is true;
	signal G1205: std_logic; attribute dont_touch of G1205: signal is true;
	signal G1211: std_logic; attribute dont_touch of G1211: signal is true;
	signal G1216: std_logic; attribute dont_touch of G1216: signal is true;
	signal G1221: std_logic; attribute dont_touch of G1221: signal is true;
	signal G1227: std_logic; attribute dont_touch of G1227: signal is true;
	signal G1233: std_logic; attribute dont_touch of G1233: signal is true;
	signal G1236: std_logic; attribute dont_touch of G1236: signal is true;
	signal G1239: std_logic; attribute dont_touch of G1239: signal is true;
	signal G1242: std_logic; attribute dont_touch of G1242: signal is true;
	signal G1246: std_logic; attribute dont_touch of G1246: signal is true;
	signal G1249: std_logic; attribute dont_touch of G1249: signal is true;
	signal G1252: std_logic; attribute dont_touch of G1252: signal is true;
	signal G1256: std_logic; attribute dont_touch of G1256: signal is true;
	signal G1259: std_logic; attribute dont_touch of G1259: signal is true;
	signal G1263: std_logic; attribute dont_touch of G1263: signal is true;
	signal G1266: std_logic; attribute dont_touch of G1266: signal is true;
	signal G1270: std_logic; attribute dont_touch of G1270: signal is true;
	signal G1274: std_logic; attribute dont_touch of G1274: signal is true;
	signal G1277: std_logic; attribute dont_touch of G1277: signal is true;
	signal G1280: std_logic; attribute dont_touch of G1280: signal is true;
	signal G1283: std_logic; attribute dont_touch of G1283: signal is true;
	signal G1287: std_logic; attribute dont_touch of G1287: signal is true;
	signal G1291: std_logic; attribute dont_touch of G1291: signal is true;
	signal G1296: std_logic; attribute dont_touch of G1296: signal is true;
	signal G1300: std_logic; attribute dont_touch of G1300: signal is true;
	signal G1306: std_logic; attribute dont_touch of G1306: signal is true;
	signal G1311: std_logic; attribute dont_touch of G1311: signal is true;
	signal G1312: std_logic; attribute dont_touch of G1312: signal is true;
	signal G1319: std_logic; attribute dont_touch of G1319: signal is true;
	signal G1322: std_logic; attribute dont_touch of G1322: signal is true;
	signal G1333: std_logic; attribute dont_touch of G1333: signal is true;
	signal G1339: std_logic; attribute dont_touch of G1339: signal is true;
	signal G1345: std_logic; attribute dont_touch of G1345: signal is true;
	signal G1351: std_logic; attribute dont_touch of G1351: signal is true;
	signal G1361: std_logic; attribute dont_touch of G1361: signal is true;
	signal G1367: std_logic; attribute dont_touch of G1367: signal is true;
	signal G1373: std_logic; attribute dont_touch of G1373: signal is true;
	signal G1379: std_logic; attribute dont_touch of G1379: signal is true;
	signal G1384: std_logic; attribute dont_touch of G1384: signal is true;
	signal G1389: std_logic; attribute dont_touch of G1389: signal is true;
	signal G1395: std_logic; attribute dont_touch of G1395: signal is true;
	signal G1399: std_logic; attribute dont_touch of G1399: signal is true;
	signal G1404: std_logic; attribute dont_touch of G1404: signal is true;
	signal G1413: std_logic; attribute dont_touch of G1413: signal is true;
	signal G1418: std_logic; attribute dont_touch of G1418: signal is true;
	signal G1422: std_logic; attribute dont_touch of G1422: signal is true;
	signal G1426: std_logic; attribute dont_touch of G1426: signal is true;
	signal G1430: std_logic; attribute dont_touch of G1430: signal is true;
	signal G1437: std_logic; attribute dont_touch of G1437: signal is true;
	signal G1442: std_logic; attribute dont_touch of G1442: signal is true;
	signal G1448: std_logic; attribute dont_touch of G1448: signal is true;
	signal G1454: std_logic; attribute dont_touch of G1454: signal is true;
	signal G1459: std_logic; attribute dont_touch of G1459: signal is true;
	signal G1467: std_logic; attribute dont_touch of G1467: signal is true;
	signal G1472: std_logic; attribute dont_touch of G1472: signal is true;
	signal G1478: std_logic; attribute dont_touch of G1478: signal is true;
	signal G1484: std_logic; attribute dont_touch of G1484: signal is true;
	signal G1489: std_logic; attribute dont_touch of G1489: signal is true;
	signal G1495: std_logic; attribute dont_touch of G1495: signal is true;
	signal G1500: std_logic; attribute dont_touch of G1500: signal is true;
	signal G1514: std_logic; attribute dont_touch of G1514: signal is true;
	signal G1521: std_logic; attribute dont_touch of G1521: signal is true;
	signal G1526: std_logic; attribute dont_touch of G1526: signal is true;
	signal G1532: std_logic; attribute dont_touch of G1532: signal is true;
	signal G1536: std_logic; attribute dont_touch of G1536: signal is true;
	signal G1542: std_logic; attribute dont_touch of G1542: signal is true;
	signal G1548: std_logic; attribute dont_touch of G1548: signal is true;
	signal G1554: std_logic; attribute dont_touch of G1554: signal is true;
	signal G1559: std_logic; attribute dont_touch of G1559: signal is true;
	signal G1564: std_logic; attribute dont_touch of G1564: signal is true;
	signal G1570: std_logic; attribute dont_touch of G1570: signal is true;
	signal G1576: std_logic; attribute dont_touch of G1576: signal is true;
	signal G1579: std_logic; attribute dont_touch of G1579: signal is true;
	signal G1582: std_logic; attribute dont_touch of G1582: signal is true;
	signal G1585: std_logic; attribute dont_touch of G1585: signal is true;
	signal G1589: std_logic; attribute dont_touch of G1589: signal is true;
	signal G1592: std_logic; attribute dont_touch of G1592: signal is true;
	signal G1600: std_logic; attribute dont_touch of G1600: signal is true;
	signal G1604: std_logic; attribute dont_touch of G1604: signal is true;
	signal G1608: std_logic; attribute dont_touch of G1608: signal is true;
	signal G1612: std_logic; attribute dont_touch of G1612: signal is true;
	signal G1616: std_logic; attribute dont_touch of G1616: signal is true;
	signal G1620: std_logic; attribute dont_touch of G1620: signal is true;
	signal G1624: std_logic; attribute dont_touch of G1624: signal is true;
	signal G1632: std_logic; attribute dont_touch of G1632: signal is true;
	signal G1636: std_logic; attribute dont_touch of G1636: signal is true;
	signal G1644: std_logic; attribute dont_touch of G1644: signal is true;
	signal G1648: std_logic; attribute dont_touch of G1648: signal is true;
	signal G1657: std_logic; attribute dont_touch of G1657: signal is true;
	signal G1664: std_logic; attribute dont_touch of G1664: signal is true;
	signal G1668: std_logic; attribute dont_touch of G1668: signal is true;
	signal G1677: std_logic; attribute dont_touch of G1677: signal is true;
	signal G1682: std_logic; attribute dont_touch of G1682: signal is true;
	signal G1687: std_logic; attribute dont_touch of G1687: signal is true;
	signal G1691: std_logic; attribute dont_touch of G1691: signal is true;
	signal G1696: std_logic; attribute dont_touch of G1696: signal is true;
	signal G1700: std_logic; attribute dont_touch of G1700: signal is true;
	signal G1706: std_logic; attribute dont_touch of G1706: signal is true;
	signal G1710: std_logic; attribute dont_touch of G1710: signal is true;
	signal G1714: std_logic; attribute dont_touch of G1714: signal is true;
	signal G1720: std_logic; attribute dont_touch of G1720: signal is true;
	signal G1724: std_logic; attribute dont_touch of G1724: signal is true;
	signal G1728: std_logic; attribute dont_touch of G1728: signal is true;
	signal G1736: std_logic; attribute dont_touch of G1736: signal is true;
	signal G1740: std_logic; attribute dont_touch of G1740: signal is true;
	signal G1744: std_logic; attribute dont_touch of G1744: signal is true;
	signal G1748: std_logic; attribute dont_touch of G1748: signal is true;
	signal G1752: std_logic; attribute dont_touch of G1752: signal is true;
	signal G1756: std_logic; attribute dont_touch of G1756: signal is true;
	signal G1760: std_logic; attribute dont_touch of G1760: signal is true;
	signal G1768: std_logic; attribute dont_touch of G1768: signal is true;
	signal G1772: std_logic; attribute dont_touch of G1772: signal is true;
	signal G1779: std_logic; attribute dont_touch of G1779: signal is true;
	signal G1783: std_logic; attribute dont_touch of G1783: signal is true;
	signal G1792: std_logic; attribute dont_touch of G1792: signal is true;
	signal G1798: std_logic; attribute dont_touch of G1798: signal is true;
	signal G1802: std_logic; attribute dont_touch of G1802: signal is true;
	signal G1811: std_logic; attribute dont_touch of G1811: signal is true;
	signal G1816: std_logic; attribute dont_touch of G1816: signal is true;
	signal G1821: std_logic; attribute dont_touch of G1821: signal is true;
	signal G1825: std_logic; attribute dont_touch of G1825: signal is true;
	signal G1830: std_logic; attribute dont_touch of G1830: signal is true;
	signal G1834: std_logic; attribute dont_touch of G1834: signal is true;
	signal G1840: std_logic; attribute dont_touch of G1840: signal is true;
	signal G1844: std_logic; attribute dont_touch of G1844: signal is true;
	signal G1848: std_logic; attribute dont_touch of G1848: signal is true;
	signal G1854: std_logic; attribute dont_touch of G1854: signal is true;
	signal G1858: std_logic; attribute dont_touch of G1858: signal is true;
	signal G1862: std_logic; attribute dont_touch of G1862: signal is true;
	signal G1870: std_logic; attribute dont_touch of G1870: signal is true;
	signal G1874: std_logic; attribute dont_touch of G1874: signal is true;
	signal G1878: std_logic; attribute dont_touch of G1878: signal is true;
	signal G1882: std_logic; attribute dont_touch of G1882: signal is true;
	signal G1886: std_logic; attribute dont_touch of G1886: signal is true;
	signal G1890: std_logic; attribute dont_touch of G1890: signal is true;
	signal G1894: std_logic; attribute dont_touch of G1894: signal is true;
	signal G1902: std_logic; attribute dont_touch of G1902: signal is true;
	signal G1906: std_logic; attribute dont_touch of G1906: signal is true;
	signal G1913: std_logic; attribute dont_touch of G1913: signal is true;
	signal G1917: std_logic; attribute dont_touch of G1917: signal is true;
	signal G1926: std_logic; attribute dont_touch of G1926: signal is true;
	signal G1932: std_logic; attribute dont_touch of G1932: signal is true;
	signal G1936: std_logic; attribute dont_touch of G1936: signal is true;
	signal G1945: std_logic; attribute dont_touch of G1945: signal is true;
	signal G1950: std_logic; attribute dont_touch of G1950: signal is true;
	signal G1955: std_logic; attribute dont_touch of G1955: signal is true;
	signal G1959: std_logic; attribute dont_touch of G1959: signal is true;
	signal G1964: std_logic; attribute dont_touch of G1964: signal is true;
	signal G1968: std_logic; attribute dont_touch of G1968: signal is true;
	signal G1974: std_logic; attribute dont_touch of G1974: signal is true;
	signal G1978: std_logic; attribute dont_touch of G1978: signal is true;
	signal G1982: std_logic; attribute dont_touch of G1982: signal is true;
	signal G1988: std_logic; attribute dont_touch of G1988: signal is true;
	signal G1992: std_logic; attribute dont_touch of G1992: signal is true;
	signal G1996: std_logic; attribute dont_touch of G1996: signal is true;
	signal G2004: std_logic; attribute dont_touch of G2004: signal is true;
	signal G2008: std_logic; attribute dont_touch of G2008: signal is true;
	signal G2012: std_logic; attribute dont_touch of G2012: signal is true;
	signal G2016: std_logic; attribute dont_touch of G2016: signal is true;
	signal G2020: std_logic; attribute dont_touch of G2020: signal is true;
	signal G2024: std_logic; attribute dont_touch of G2024: signal is true;
	signal G2028: std_logic; attribute dont_touch of G2028: signal is true;
	signal G2036: std_logic; attribute dont_touch of G2036: signal is true;
	signal G2040: std_logic; attribute dont_touch of G2040: signal is true;
	signal G2047: std_logic; attribute dont_touch of G2047: signal is true;
	signal G2051: std_logic; attribute dont_touch of G2051: signal is true;
	signal G2060: std_logic; attribute dont_touch of G2060: signal is true;
	signal G2066: std_logic; attribute dont_touch of G2066: signal is true;
	signal G2070: std_logic; attribute dont_touch of G2070: signal is true;
	signal G2079: std_logic; attribute dont_touch of G2079: signal is true;
	signal G2084: std_logic; attribute dont_touch of G2084: signal is true;
	signal G2089: std_logic; attribute dont_touch of G2089: signal is true;
	signal G2093: std_logic; attribute dont_touch of G2093: signal is true;
	signal G2098: std_logic; attribute dont_touch of G2098: signal is true;
	signal G2102: std_logic; attribute dont_touch of G2102: signal is true;
	signal G2108: std_logic; attribute dont_touch of G2108: signal is true;
	signal G2112: std_logic; attribute dont_touch of G2112: signal is true;
	signal G2116: std_logic; attribute dont_touch of G2116: signal is true;
	signal G2122: std_logic; attribute dont_touch of G2122: signal is true;
	signal G2126: std_logic; attribute dont_touch of G2126: signal is true;
	signal G2130: std_logic; attribute dont_touch of G2130: signal is true;
	signal G2138: std_logic; attribute dont_touch of G2138: signal is true;
	signal G2145: std_logic; attribute dont_touch of G2145: signal is true;
	signal G2151: std_logic; attribute dont_touch of G2151: signal is true;
	signal G2152: std_logic; attribute dont_touch of G2152: signal is true;
	signal G2153: std_logic; attribute dont_touch of G2153: signal is true;
	signal G2161: std_logic; attribute dont_touch of G2161: signal is true;
	signal G2165: std_logic; attribute dont_touch of G2165: signal is true;
	signal G2169: std_logic; attribute dont_touch of G2169: signal is true;
	signal G2173: std_logic; attribute dont_touch of G2173: signal is true;
	signal G2177: std_logic; attribute dont_touch of G2177: signal is true;
	signal G2181: std_logic; attribute dont_touch of G2181: signal is true;
	signal G2185: std_logic; attribute dont_touch of G2185: signal is true;
	signal G2193: std_logic; attribute dont_touch of G2193: signal is true;
	signal G2197: std_logic; attribute dont_touch of G2197: signal is true;
	signal G2204: std_logic; attribute dont_touch of G2204: signal is true;
	signal G2208: std_logic; attribute dont_touch of G2208: signal is true;
	signal G2217: std_logic; attribute dont_touch of G2217: signal is true;
	signal G2223: std_logic; attribute dont_touch of G2223: signal is true;
	signal G2227: std_logic; attribute dont_touch of G2227: signal is true;
	signal G2236: std_logic; attribute dont_touch of G2236: signal is true;
	signal G2241: std_logic; attribute dont_touch of G2241: signal is true;
	signal G2246: std_logic; attribute dont_touch of G2246: signal is true;
	signal G2250: std_logic; attribute dont_touch of G2250: signal is true;
	signal G2255: std_logic; attribute dont_touch of G2255: signal is true;
	signal G2259: std_logic; attribute dont_touch of G2259: signal is true;
	signal G2265: std_logic; attribute dont_touch of G2265: signal is true;
	signal G2269: std_logic; attribute dont_touch of G2269: signal is true;
	signal G2273: std_logic; attribute dont_touch of G2273: signal is true;
	signal G2279: std_logic; attribute dont_touch of G2279: signal is true;
	signal G2283: std_logic; attribute dont_touch of G2283: signal is true;
	signal G2287: std_logic; attribute dont_touch of G2287: signal is true;
	signal G2295: std_logic; attribute dont_touch of G2295: signal is true;
	signal G2299: std_logic; attribute dont_touch of G2299: signal is true;
	signal G2303: std_logic; attribute dont_touch of G2303: signal is true;
	signal G2307: std_logic; attribute dont_touch of G2307: signal is true;
	signal G2311: std_logic; attribute dont_touch of G2311: signal is true;
	signal G2315: std_logic; attribute dont_touch of G2315: signal is true;
	signal G2319: std_logic; attribute dont_touch of G2319: signal is true;
	signal G2327: std_logic; attribute dont_touch of G2327: signal is true;
	signal G2331: std_logic; attribute dont_touch of G2331: signal is true;
	signal G2338: std_logic; attribute dont_touch of G2338: signal is true;
	signal G2342: std_logic; attribute dont_touch of G2342: signal is true;
	signal G2351: std_logic; attribute dont_touch of G2351: signal is true;
	signal G2357: std_logic; attribute dont_touch of G2357: signal is true;
	signal G2361: std_logic; attribute dont_touch of G2361: signal is true;
	signal G2370: std_logic; attribute dont_touch of G2370: signal is true;
	signal G2375: std_logic; attribute dont_touch of G2375: signal is true;
	signal G2380: std_logic; attribute dont_touch of G2380: signal is true;
	signal G2384: std_logic; attribute dont_touch of G2384: signal is true;
	signal G2389: std_logic; attribute dont_touch of G2389: signal is true;
	signal G2393: std_logic; attribute dont_touch of G2393: signal is true;
	signal G2399: std_logic; attribute dont_touch of G2399: signal is true;
	signal G2403: std_logic; attribute dont_touch of G2403: signal is true;
	signal G2407: std_logic; attribute dont_touch of G2407: signal is true;
	signal G2413: std_logic; attribute dont_touch of G2413: signal is true;
	signal G2417: std_logic; attribute dont_touch of G2417: signal is true;
	signal G2421: std_logic; attribute dont_touch of G2421: signal is true;
	signal G2429: std_logic; attribute dont_touch of G2429: signal is true;
	signal G2433: std_logic; attribute dont_touch of G2433: signal is true;
	signal G2437: std_logic; attribute dont_touch of G2437: signal is true;
	signal G2441: std_logic; attribute dont_touch of G2441: signal is true;
	signal G2445: std_logic; attribute dont_touch of G2445: signal is true;
	signal G2449: std_logic; attribute dont_touch of G2449: signal is true;
	signal G2453: std_logic; attribute dont_touch of G2453: signal is true;
	signal G2461: std_logic; attribute dont_touch of G2461: signal is true;
	signal G2465: std_logic; attribute dont_touch of G2465: signal is true;
	signal G2472: std_logic; attribute dont_touch of G2472: signal is true;
	signal G2476: std_logic; attribute dont_touch of G2476: signal is true;
	signal G2485: std_logic; attribute dont_touch of G2485: signal is true;
	signal G2491: std_logic; attribute dont_touch of G2491: signal is true;
	signal G2495: std_logic; attribute dont_touch of G2495: signal is true;
	signal G2504: std_logic; attribute dont_touch of G2504: signal is true;
	signal G2509: std_logic; attribute dont_touch of G2509: signal is true;
	signal G2514: std_logic; attribute dont_touch of G2514: signal is true;
	signal G2518: std_logic; attribute dont_touch of G2518: signal is true;
	signal G2523: std_logic; attribute dont_touch of G2523: signal is true;
	signal G2527: std_logic; attribute dont_touch of G2527: signal is true;
	signal G2533: std_logic; attribute dont_touch of G2533: signal is true;
	signal G2537: std_logic; attribute dont_touch of G2537: signal is true;
	signal G2541: std_logic; attribute dont_touch of G2541: signal is true;
	signal G2547: std_logic; attribute dont_touch of G2547: signal is true;
	signal G2551: std_logic; attribute dont_touch of G2551: signal is true;
	signal G2555: std_logic; attribute dont_touch of G2555: signal is true;
	signal G2563: std_logic; attribute dont_touch of G2563: signal is true;
	signal G2567: std_logic; attribute dont_touch of G2567: signal is true;
	signal G2571: std_logic; attribute dont_touch of G2571: signal is true;
	signal G2575: std_logic; attribute dont_touch of G2575: signal is true;
	signal G2579: std_logic; attribute dont_touch of G2579: signal is true;
	signal G2583: std_logic; attribute dont_touch of G2583: signal is true;
	signal G2587: std_logic; attribute dont_touch of G2587: signal is true;
	signal G2595: std_logic; attribute dont_touch of G2595: signal is true;
	signal G2599: std_logic; attribute dont_touch of G2599: signal is true;
	signal G2606: std_logic; attribute dont_touch of G2606: signal is true;
	signal G2610: std_logic; attribute dont_touch of G2610: signal is true;
	signal G2619: std_logic; attribute dont_touch of G2619: signal is true;
	signal G2625: std_logic; attribute dont_touch of G2625: signal is true;
	signal G2629: std_logic; attribute dont_touch of G2629: signal is true;
	signal G2638: std_logic; attribute dont_touch of G2638: signal is true;
	signal G2643: std_logic; attribute dont_touch of G2643: signal is true;
	signal G2648: std_logic; attribute dont_touch of G2648: signal is true;
	signal G2652: std_logic; attribute dont_touch of G2652: signal is true;
	signal G2657: std_logic; attribute dont_touch of G2657: signal is true;
	signal G2661: std_logic; attribute dont_touch of G2661: signal is true;
	signal G2667: std_logic; attribute dont_touch of G2667: signal is true;
	signal G2671: std_logic; attribute dont_touch of G2671: signal is true;
	signal G2675: std_logic; attribute dont_touch of G2675: signal is true;
	signal G2681: std_logic; attribute dont_touch of G2681: signal is true;
	signal G2685: std_logic; attribute dont_touch of G2685: signal is true;
	signal G2689: std_logic; attribute dont_touch of G2689: signal is true;
	signal G2697: std_logic; attribute dont_touch of G2697: signal is true;
	signal G2704: std_logic; attribute dont_touch of G2704: signal is true;
	signal G2710: std_logic; attribute dont_touch of G2710: signal is true;
	signal G2711: std_logic; attribute dont_touch of G2711: signal is true;
	signal G2712: std_logic; attribute dont_touch of G2712: signal is true;
	signal G2715: std_logic; attribute dont_touch of G2715: signal is true;
	signal G2719: std_logic; attribute dont_touch of G2719: signal is true;
	signal G2724: std_logic; attribute dont_touch of G2724: signal is true;
	signal G2729: std_logic; attribute dont_touch of G2729: signal is true;
	signal G2735: std_logic; attribute dont_touch of G2735: signal is true;
	signal G2741: std_logic; attribute dont_touch of G2741: signal is true;
	signal G2748: std_logic; attribute dont_touch of G2748: signal is true;
	signal G2756: std_logic; attribute dont_touch of G2756: signal is true;
	signal G2759: std_logic; attribute dont_touch of G2759: signal is true;
	signal G2763: std_logic; attribute dont_touch of G2763: signal is true;
	signal G2767: std_logic; attribute dont_touch of G2767: signal is true;
	signal G2771: std_logic; attribute dont_touch of G2771: signal is true;
	signal G2775: std_logic; attribute dont_touch of G2775: signal is true;
	signal G2779: std_logic; attribute dont_touch of G2779: signal is true;
	signal G2783: std_logic; attribute dont_touch of G2783: signal is true;
	signal G2787: std_logic; attribute dont_touch of G2787: signal is true;
	signal G2791: std_logic; attribute dont_touch of G2791: signal is true;
	signal G2795: std_logic; attribute dont_touch of G2795: signal is true;
	signal G2799: std_logic; attribute dont_touch of G2799: signal is true;
	signal G2803: std_logic; attribute dont_touch of G2803: signal is true;
	signal G2807: std_logic; attribute dont_touch of G2807: signal is true;
	signal G2811: std_logic; attribute dont_touch of G2811: signal is true;
	signal G2815: std_logic; attribute dont_touch of G2815: signal is true;
	signal G2819: std_logic; attribute dont_touch of G2819: signal is true;
	signal G2823: std_logic; attribute dont_touch of G2823: signal is true;
	signal G2827: std_logic; attribute dont_touch of G2827: signal is true;
	signal G2831: std_logic; attribute dont_touch of G2831: signal is true;
	signal G2834: std_logic; attribute dont_touch of G2834: signal is true;
	signal G2837: std_logic; attribute dont_touch of G2837: signal is true;
	signal G2841: std_logic; attribute dont_touch of G2841: signal is true;
	signal G2844: std_logic; attribute dont_touch of G2844: signal is true;
	signal G2848: std_logic; attribute dont_touch of G2848: signal is true;
	signal G2852: std_logic; attribute dont_touch of G2852: signal is true;
	signal G2856: std_logic; attribute dont_touch of G2856: signal is true;
	signal G2860: std_logic; attribute dont_touch of G2860: signal is true;
	signal G2864: std_logic; attribute dont_touch of G2864: signal is true;
	signal G2868: std_logic; attribute dont_touch of G2868: signal is true;
	signal G2873: std_logic; attribute dont_touch of G2873: signal is true;
	signal G2878: std_logic; attribute dont_touch of G2878: signal is true;
	signal G2882: std_logic; attribute dont_touch of G2882: signal is true;
	signal G2886: std_logic; attribute dont_touch of G2886: signal is true;
	signal G2890: std_logic; attribute dont_touch of G2890: signal is true;
	signal G2894: std_logic; attribute dont_touch of G2894: signal is true;
	signal G2898: std_logic; attribute dont_touch of G2898: signal is true;
	signal G2902: std_logic; attribute dont_touch of G2902: signal is true;
	signal G2907: std_logic; attribute dont_touch of G2907: signal is true;
	signal G2912: std_logic; attribute dont_touch of G2912: signal is true;
	signal G2917: std_logic; attribute dont_touch of G2917: signal is true;
	signal G2922: std_logic; attribute dont_touch of G2922: signal is true;
	signal G2927: std_logic; attribute dont_touch of G2927: signal is true;
	signal G2932: std_logic; attribute dont_touch of G2932: signal is true;
	signal G2936: std_logic; attribute dont_touch of G2936: signal is true;
	signal G2941: std_logic; attribute dont_touch of G2941: signal is true;
	signal G2946: std_logic; attribute dont_touch of G2946: signal is true;
	signal G2950: std_logic; attribute dont_touch of G2950: signal is true;
	signal G2955: std_logic; attribute dont_touch of G2955: signal is true;
	signal G2960: std_logic; attribute dont_touch of G2960: signal is true;
	signal G2965: std_logic; attribute dont_touch of G2965: signal is true;
	signal G2970: std_logic; attribute dont_touch of G2970: signal is true;
	signal G2975: std_logic; attribute dont_touch of G2975: signal is true;
	signal G2980: std_logic; attribute dont_touch of G2980: signal is true;
	signal G2984: std_logic; attribute dont_touch of G2984: signal is true;
	signal G2988: std_logic; attribute dont_touch of G2988: signal is true;
	signal G2994: std_logic; attribute dont_touch of G2994: signal is true;
	signal G2999: std_logic; attribute dont_touch of G2999: signal is true;
	signal G3003: std_logic; attribute dont_touch of G3003: signal is true;
	signal G3004: std_logic; attribute dont_touch of G3004: signal is true;
	signal G3010: std_logic; attribute dont_touch of G3010: signal is true;
	signal G3017: std_logic; attribute dont_touch of G3017: signal is true;
	signal G3021: std_logic; attribute dont_touch of G3021: signal is true;
	signal G3025: std_logic; attribute dont_touch of G3025: signal is true;
	signal G3029: std_logic; attribute dont_touch of G3029: signal is true;
	signal G3034: std_logic; attribute dont_touch of G3034: signal is true;
	signal G3040: std_logic; attribute dont_touch of G3040: signal is true;
	signal G3045: std_logic; attribute dont_touch of G3045: signal is true;
	signal G3050: std_logic; attribute dont_touch of G3050: signal is true;
	signal G3057: std_logic; attribute dont_touch of G3057: signal is true;
	signal G3061: std_logic; attribute dont_touch of G3061: signal is true;
	signal G3065: std_logic; attribute dont_touch of G3065: signal is true;
	signal G3068: std_logic; attribute dont_touch of G3068: signal is true;
	signal G3072: std_logic; attribute dont_touch of G3072: signal is true;
	signal G3080: std_logic; attribute dont_touch of G3080: signal is true;
	signal G3085: std_logic; attribute dont_touch of G3085: signal is true;
	signal G3089: std_logic; attribute dont_touch of G3089: signal is true;
	signal G3092: std_logic; attribute dont_touch of G3092: signal is true;
	signal G3096: std_logic; attribute dont_touch of G3096: signal is true;
	signal G3100: std_logic; attribute dont_touch of G3100: signal is true;
	signal G3103: std_logic; attribute dont_touch of G3103: signal is true;
	signal G3106: std_logic; attribute dont_touch of G3106: signal is true;
	signal G3111: std_logic; attribute dont_touch of G3111: signal is true;
	signal G3115: std_logic; attribute dont_touch of G3115: signal is true;
	signal G3119: std_logic; attribute dont_touch of G3119: signal is true;
	signal G3125: std_logic; attribute dont_touch of G3125: signal is true;
	signal G3129: std_logic; attribute dont_touch of G3129: signal is true;
	signal G3133: std_logic; attribute dont_touch of G3133: signal is true;
	signal G3139: std_logic; attribute dont_touch of G3139: signal is true;
	signal G3143: std_logic; attribute dont_touch of G3143: signal is true;
	signal G3147: std_logic; attribute dont_touch of G3147: signal is true;
	signal G3151: std_logic; attribute dont_touch of G3151: signal is true;
	signal G3155: std_logic; attribute dont_touch of G3155: signal is true;
	signal G3161: std_logic; attribute dont_touch of G3161: signal is true;
	signal G3167: std_logic; attribute dont_touch of G3167: signal is true;
	signal G3171: std_logic; attribute dont_touch of G3171: signal is true;
	signal G3179: std_logic; attribute dont_touch of G3179: signal is true;
	signal G3187: std_logic; attribute dont_touch of G3187: signal is true;
	signal G3191: std_logic; attribute dont_touch of G3191: signal is true;
	signal G3195: std_logic; attribute dont_touch of G3195: signal is true;
	signal G3199: std_logic; attribute dont_touch of G3199: signal is true;
	signal G3203: std_logic; attribute dont_touch of G3203: signal is true;
	signal G3207: std_logic; attribute dont_touch of G3207: signal is true;
	signal G3211: std_logic; attribute dont_touch of G3211: signal is true;
	signal G3215: std_logic; attribute dont_touch of G3215: signal is true;
	signal G3219: std_logic; attribute dont_touch of G3219: signal is true;
	signal G3223: std_logic; attribute dont_touch of G3223: signal is true;
	signal G3227: std_logic; attribute dont_touch of G3227: signal is true;
	signal G3231: std_logic; attribute dont_touch of G3231: signal is true;
	signal G3235: std_logic; attribute dont_touch of G3235: signal is true;
	signal G3239: std_logic; attribute dont_touch of G3239: signal is true;
	signal G3243: std_logic; attribute dont_touch of G3243: signal is true;
	signal G3247: std_logic; attribute dont_touch of G3247: signal is true;
	signal G3251: std_logic; attribute dont_touch of G3251: signal is true;
	signal G3255: std_logic; attribute dont_touch of G3255: signal is true;
	signal G3259: std_logic; attribute dont_touch of G3259: signal is true;
	signal G3263: std_logic; attribute dont_touch of G3263: signal is true;
	signal G3267: std_logic; attribute dont_touch of G3267: signal is true;
	signal G3274: std_logic; attribute dont_touch of G3274: signal is true;
	signal G3281: std_logic; attribute dont_touch of G3281: signal is true;
	signal G3288: std_logic; attribute dont_touch of G3288: signal is true;
	signal G3298: std_logic; attribute dont_touch of G3298: signal is true;
	signal G3303: std_logic; attribute dont_touch of G3303: signal is true;
	signal G3310: std_logic; attribute dont_touch of G3310: signal is true;
	signal G3317: std_logic; attribute dont_touch of G3317: signal is true;
	signal G3321: std_logic; attribute dont_touch of G3321: signal is true;
	signal G3325: std_logic; attribute dont_touch of G3325: signal is true;
	signal G3329: std_logic; attribute dont_touch of G3329: signal is true;
	signal G3333: std_logic; attribute dont_touch of G3333: signal is true;
	signal G3338: std_logic; attribute dont_touch of G3338: signal is true;
	signal G3343: std_logic; attribute dont_touch of G3343: signal is true;
	signal G3347: std_logic; attribute dont_touch of G3347: signal is true;
	signal G3352: std_logic; attribute dont_touch of G3352: signal is true;
	signal G3355: std_logic; attribute dont_touch of G3355: signal is true;
	signal G3361: std_logic; attribute dont_touch of G3361: signal is true;
	signal G3368: std_logic; attribute dont_touch of G3368: signal is true;
	signal G3372: std_logic; attribute dont_touch of G3372: signal is true;
	signal G3376: std_logic; attribute dont_touch of G3376: signal is true;
	signal G3380: std_logic; attribute dont_touch of G3380: signal is true;
	signal G3385: std_logic; attribute dont_touch of G3385: signal is true;
	signal G3391: std_logic; attribute dont_touch of G3391: signal is true;
	signal G3396: std_logic; attribute dont_touch of G3396: signal is true;
	signal G3401: std_logic; attribute dont_touch of G3401: signal is true;
	signal G3408: std_logic; attribute dont_touch of G3408: signal is true;
	signal G3412: std_logic; attribute dont_touch of G3412: signal is true;
	signal G3416: std_logic; attribute dont_touch of G3416: signal is true;
	signal G3419: std_logic; attribute dont_touch of G3419: signal is true;
	signal G3423: std_logic; attribute dont_touch of G3423: signal is true;
	signal G3431: std_logic; attribute dont_touch of G3431: signal is true;
	signal G3436: std_logic; attribute dont_touch of G3436: signal is true;
	signal G3440: std_logic; attribute dont_touch of G3440: signal is true;
	signal G3443: std_logic; attribute dont_touch of G3443: signal is true;
	signal G3447: std_logic; attribute dont_touch of G3447: signal is true;
	signal G3451: std_logic; attribute dont_touch of G3451: signal is true;
	signal G3454: std_logic; attribute dont_touch of G3454: signal is true;
	signal G3457: std_logic; attribute dont_touch of G3457: signal is true;
	signal G3462: std_logic; attribute dont_touch of G3462: signal is true;
	signal G3466: std_logic; attribute dont_touch of G3466: signal is true;
	signal G3470: std_logic; attribute dont_touch of G3470: signal is true;
	signal G3476: std_logic; attribute dont_touch of G3476: signal is true;
	signal G3480: std_logic; attribute dont_touch of G3480: signal is true;
	signal G3484: std_logic; attribute dont_touch of G3484: signal is true;
	signal G3490: std_logic; attribute dont_touch of G3490: signal is true;
	signal G3494: std_logic; attribute dont_touch of G3494: signal is true;
	signal G3498: std_logic; attribute dont_touch of G3498: signal is true;
	signal G3502: std_logic; attribute dont_touch of G3502: signal is true;
	signal G3506: std_logic; attribute dont_touch of G3506: signal is true;
	signal G3512: std_logic; attribute dont_touch of G3512: signal is true;
	signal G3518: std_logic; attribute dont_touch of G3518: signal is true;
	signal G3522: std_logic; attribute dont_touch of G3522: signal is true;
	signal G3530: std_logic; attribute dont_touch of G3530: signal is true;
	signal G3538: std_logic; attribute dont_touch of G3538: signal is true;
	signal G3542: std_logic; attribute dont_touch of G3542: signal is true;
	signal G3546: std_logic; attribute dont_touch of G3546: signal is true;
	signal G3550: std_logic; attribute dont_touch of G3550: signal is true;
	signal G3554: std_logic; attribute dont_touch of G3554: signal is true;
	signal G3558: std_logic; attribute dont_touch of G3558: signal is true;
	signal G3562: std_logic; attribute dont_touch of G3562: signal is true;
	signal G3566: std_logic; attribute dont_touch of G3566: signal is true;
	signal G3570: std_logic; attribute dont_touch of G3570: signal is true;
	signal G3574: std_logic; attribute dont_touch of G3574: signal is true;
	signal G3578: std_logic; attribute dont_touch of G3578: signal is true;
	signal G3582: std_logic; attribute dont_touch of G3582: signal is true;
	signal G3586: std_logic; attribute dont_touch of G3586: signal is true;
	signal G3590: std_logic; attribute dont_touch of G3590: signal is true;
	signal G3594: std_logic; attribute dont_touch of G3594: signal is true;
	signal G3598: std_logic; attribute dont_touch of G3598: signal is true;
	signal G3602: std_logic; attribute dont_touch of G3602: signal is true;
	signal G3606: std_logic; attribute dont_touch of G3606: signal is true;
	signal G3610: std_logic; attribute dont_touch of G3610: signal is true;
	signal G3614: std_logic; attribute dont_touch of G3614: signal is true;
	signal G3618: std_logic; attribute dont_touch of G3618: signal is true;
	signal G3625: std_logic; attribute dont_touch of G3625: signal is true;
	signal G3632: std_logic; attribute dont_touch of G3632: signal is true;
	signal G3639: std_logic; attribute dont_touch of G3639: signal is true;
	signal G3649: std_logic; attribute dont_touch of G3649: signal is true;
	signal G3654: std_logic; attribute dont_touch of G3654: signal is true;
	signal G3661: std_logic; attribute dont_touch of G3661: signal is true;
	signal G3668: std_logic; attribute dont_touch of G3668: signal is true;
	signal G3672: std_logic; attribute dont_touch of G3672: signal is true;
	signal G3676: std_logic; attribute dont_touch of G3676: signal is true;
	signal G3680: std_logic; attribute dont_touch of G3680: signal is true;
	signal G3684: std_logic; attribute dont_touch of G3684: signal is true;
	signal G3689: std_logic; attribute dont_touch of G3689: signal is true;
	signal G3694: std_logic; attribute dont_touch of G3694: signal is true;
	signal G3698: std_logic; attribute dont_touch of G3698: signal is true;
	signal G3703: std_logic; attribute dont_touch of G3703: signal is true;
	signal G3706: std_logic; attribute dont_touch of G3706: signal is true;
	signal G3712: std_logic; attribute dont_touch of G3712: signal is true;
	signal G3719: std_logic; attribute dont_touch of G3719: signal is true;
	signal G3723: std_logic; attribute dont_touch of G3723: signal is true;
	signal G3727: std_logic; attribute dont_touch of G3727: signal is true;
	signal G3731: std_logic; attribute dont_touch of G3731: signal is true;
	signal G3736: std_logic; attribute dont_touch of G3736: signal is true;
	signal G3742: std_logic; attribute dont_touch of G3742: signal is true;
	signal G3747: std_logic; attribute dont_touch of G3747: signal is true;
	signal G3752: std_logic; attribute dont_touch of G3752: signal is true;
	signal G3759: std_logic; attribute dont_touch of G3759: signal is true;
	signal G3763: std_logic; attribute dont_touch of G3763: signal is true;
	signal G3767: std_logic; attribute dont_touch of G3767: signal is true;
	signal G3770: std_logic; attribute dont_touch of G3770: signal is true;
	signal G3774: std_logic; attribute dont_touch of G3774: signal is true;
	signal G3782: std_logic; attribute dont_touch of G3782: signal is true;
	signal G3787: std_logic; attribute dont_touch of G3787: signal is true;
	signal G3791: std_logic; attribute dont_touch of G3791: signal is true;
	signal G3794: std_logic; attribute dont_touch of G3794: signal is true;
	signal G3798: std_logic; attribute dont_touch of G3798: signal is true;
	signal G3802: std_logic; attribute dont_touch of G3802: signal is true;
	signal G3805: std_logic; attribute dont_touch of G3805: signal is true;
	signal G3808: std_logic; attribute dont_touch of G3808: signal is true;
	signal G3813: std_logic; attribute dont_touch of G3813: signal is true;
	signal G3817: std_logic; attribute dont_touch of G3817: signal is true;
	signal G3821: std_logic; attribute dont_touch of G3821: signal is true;
	signal G3827: std_logic; attribute dont_touch of G3827: signal is true;
	signal G3831: std_logic; attribute dont_touch of G3831: signal is true;
	signal G3835: std_logic; attribute dont_touch of G3835: signal is true;
	signal G3841: std_logic; attribute dont_touch of G3841: signal is true;
	signal G3845: std_logic; attribute dont_touch of G3845: signal is true;
	signal G3849: std_logic; attribute dont_touch of G3849: signal is true;
	signal G3853: std_logic; attribute dont_touch of G3853: signal is true;
	signal G3857: std_logic; attribute dont_touch of G3857: signal is true;
	signal G3863: std_logic; attribute dont_touch of G3863: signal is true;
	signal G3869: std_logic; attribute dont_touch of G3869: signal is true;
	signal G3873: std_logic; attribute dont_touch of G3873: signal is true;
	signal G3881: std_logic; attribute dont_touch of G3881: signal is true;
	signal G3889: std_logic; attribute dont_touch of G3889: signal is true;
	signal G3893: std_logic; attribute dont_touch of G3893: signal is true;
	signal G3897: std_logic; attribute dont_touch of G3897: signal is true;
	signal G3901: std_logic; attribute dont_touch of G3901: signal is true;
	signal G3905: std_logic; attribute dont_touch of G3905: signal is true;
	signal G3909: std_logic; attribute dont_touch of G3909: signal is true;
	signal G3913: std_logic; attribute dont_touch of G3913: signal is true;
	signal G3917: std_logic; attribute dont_touch of G3917: signal is true;
	signal G3921: std_logic; attribute dont_touch of G3921: signal is true;
	signal G3925: std_logic; attribute dont_touch of G3925: signal is true;
	signal G3929: std_logic; attribute dont_touch of G3929: signal is true;
	signal G3933: std_logic; attribute dont_touch of G3933: signal is true;
	signal G3937: std_logic; attribute dont_touch of G3937: signal is true;
	signal G3941: std_logic; attribute dont_touch of G3941: signal is true;
	signal G3945: std_logic; attribute dont_touch of G3945: signal is true;
	signal G3949: std_logic; attribute dont_touch of G3949: signal is true;
	signal G3953: std_logic; attribute dont_touch of G3953: signal is true;
	signal G3957: std_logic; attribute dont_touch of G3957: signal is true;
	signal G3961: std_logic; attribute dont_touch of G3961: signal is true;
	signal G3965: std_logic; attribute dont_touch of G3965: signal is true;
	signal G3969: std_logic; attribute dont_touch of G3969: signal is true;
	signal G3976: std_logic; attribute dont_touch of G3976: signal is true;
	signal G3983: std_logic; attribute dont_touch of G3983: signal is true;
	signal G3990: std_logic; attribute dont_touch of G3990: signal is true;
	signal G4000: std_logic; attribute dont_touch of G4000: signal is true;
	signal G4005: std_logic; attribute dont_touch of G4005: signal is true;
	signal G4012: std_logic; attribute dont_touch of G4012: signal is true;
	signal G4019: std_logic; attribute dont_touch of G4019: signal is true;
	signal G4023: std_logic; attribute dont_touch of G4023: signal is true;
	signal G4027: std_logic; attribute dont_touch of G4027: signal is true;
	signal G4031: std_logic; attribute dont_touch of G4031: signal is true;
	signal G4035: std_logic; attribute dont_touch of G4035: signal is true;
	signal G4040: std_logic; attribute dont_touch of G4040: signal is true;
	signal G4045: std_logic; attribute dont_touch of G4045: signal is true;
	signal G4049: std_logic; attribute dont_touch of G4049: signal is true;
	signal G4054: std_logic; attribute dont_touch of G4054: signal is true;
	signal G4057: std_logic; attribute dont_touch of G4057: signal is true;
	signal G4064: std_logic; attribute dont_touch of G4064: signal is true;
	signal G4072: std_logic; attribute dont_touch of G4072: signal is true;
	signal G4076: std_logic; attribute dont_touch of G4076: signal is true;
	signal G4082: std_logic; attribute dont_touch of G4082: signal is true;
	signal G4087: std_logic; attribute dont_touch of G4087: signal is true;
	signal G4093: std_logic; attribute dont_touch of G4093: signal is true;
	signal G4098: std_logic; attribute dont_touch of G4098: signal is true;
	signal G4104: std_logic; attribute dont_touch of G4104: signal is true;
	signal G4108: std_logic; attribute dont_touch of G4108: signal is true;
	signal G4112: std_logic; attribute dont_touch of G4112: signal is true;
	signal G4116: std_logic; attribute dont_touch of G4116: signal is true;
	signal G4119: std_logic; attribute dont_touch of G4119: signal is true;
	signal G4122: std_logic; attribute dont_touch of G4122: signal is true;
	signal G4125: std_logic; attribute dont_touch of G4125: signal is true;
	signal G4129: std_logic; attribute dont_touch of G4129: signal is true;
	signal G4132: std_logic; attribute dont_touch of G4132: signal is true;
	signal G4135: std_logic; attribute dont_touch of G4135: signal is true;
	signal G4138: std_logic; attribute dont_touch of G4138: signal is true;
	signal G4141: std_logic; attribute dont_touch of G4141: signal is true;
	signal G4145: std_logic; attribute dont_touch of G4145: signal is true;
	signal G4146: std_logic; attribute dont_touch of G4146: signal is true;
	signal G4153: std_logic; attribute dont_touch of G4153: signal is true;
	signal G4157: std_logic; attribute dont_touch of G4157: signal is true;
	signal G4164: std_logic; attribute dont_touch of G4164: signal is true;
	signal G4165: std_logic; attribute dont_touch of G4165: signal is true;
	signal G4169: std_logic; attribute dont_touch of G4169: signal is true;
	signal G4172: std_logic; attribute dont_touch of G4172: signal is true;
	signal G4176: std_logic; attribute dont_touch of G4176: signal is true;
	signal G4180: std_logic; attribute dont_touch of G4180: signal is true;
	signal G4185: std_logic; attribute dont_touch of G4185: signal is true;
	signal G4188: std_logic; attribute dont_touch of G4188: signal is true;
	signal G4191: std_logic; attribute dont_touch of G4191: signal is true;
	signal G4194: std_logic; attribute dont_touch of G4194: signal is true;
	signal G4197: std_logic; attribute dont_touch of G4197: signal is true;
	signal G4200: std_logic; attribute dont_touch of G4200: signal is true;
	signal G4204: std_logic; attribute dont_touch of G4204: signal is true;
	signal G4207: std_logic; attribute dont_touch of G4207: signal is true;
	signal G4210: std_logic; attribute dont_touch of G4210: signal is true;
	signal G4213: std_logic; attribute dont_touch of G4213: signal is true;
	signal G4216: std_logic; attribute dont_touch of G4216: signal is true;
	signal G4219: std_logic; attribute dont_touch of G4219: signal is true;
	signal G4222: std_logic; attribute dont_touch of G4222: signal is true;
	signal G4226: std_logic; attribute dont_touch of G4226: signal is true;
	signal G4229: std_logic; attribute dont_touch of G4229: signal is true;
	signal G4232: std_logic; attribute dont_touch of G4232: signal is true;
	signal G4235: std_logic; attribute dont_touch of G4235: signal is true;
	signal G4239: std_logic; attribute dont_touch of G4239: signal is true;
	signal G4242: std_logic; attribute dont_touch of G4242: signal is true;
	signal G4245: std_logic; attribute dont_touch of G4245: signal is true;
	signal G4249: std_logic; attribute dont_touch of G4249: signal is true;
	signal G4253: std_logic; attribute dont_touch of G4253: signal is true;
	signal G4258: std_logic; attribute dont_touch of G4258: signal is true;
	signal G4264: std_logic; attribute dont_touch of G4264: signal is true;
	signal G4269: std_logic; attribute dont_touch of G4269: signal is true;
	signal G4273: std_logic; attribute dont_touch of G4273: signal is true;
	signal G4277: std_logic; attribute dont_touch of G4277: signal is true;
	signal G4281: std_logic; attribute dont_touch of G4281: signal is true;
	signal G4284: std_logic; attribute dont_touch of G4284: signal is true;
	signal G4287: std_logic; attribute dont_touch of G4287: signal is true;
	signal G4291: std_logic; attribute dont_touch of G4291: signal is true;
	signal G4294: std_logic; attribute dont_touch of G4294: signal is true;
	signal G4297: std_logic; attribute dont_touch of G4297: signal is true;
	signal G4300: std_logic; attribute dont_touch of G4300: signal is true;
	signal G4304: std_logic; attribute dont_touch of G4304: signal is true;
	signal G4308: std_logic; attribute dont_touch of G4308: signal is true;
	signal G4311: std_logic; attribute dont_touch of G4311: signal is true;
	signal G4322: std_logic; attribute dont_touch of G4322: signal is true;
	signal G4332: std_logic; attribute dont_touch of G4332: signal is true;
	signal G4340: std_logic; attribute dont_touch of G4340: signal is true;
	signal G4349: std_logic; attribute dont_touch of G4349: signal is true;
	signal G4358: std_logic; attribute dont_touch of G4358: signal is true;
	signal G4366: std_logic; attribute dont_touch of G4366: signal is true;
	signal G4369: std_logic; attribute dont_touch of G4369: signal is true;
	signal G4372: std_logic; attribute dont_touch of G4372: signal is true;
	signal G4375: std_logic; attribute dont_touch of G4375: signal is true;
	signal G4382: std_logic; attribute dont_touch of G4382: signal is true;
	signal G4388: std_logic; attribute dont_touch of G4388: signal is true;
	signal G4392: std_logic; attribute dont_touch of G4392: signal is true;
	signal G4401: std_logic; attribute dont_touch of G4401: signal is true;
	signal G4405: std_logic; attribute dont_touch of G4405: signal is true;
	signal G4408: std_logic; attribute dont_touch of G4408: signal is true;
	signal G4411: std_logic; attribute dont_touch of G4411: signal is true;
	signal G4414: std_logic; attribute dont_touch of G4414: signal is true;
	signal G4417: std_logic; attribute dont_touch of G4417: signal is true;
	signal G4420: std_logic; attribute dont_touch of G4420: signal is true;
	signal G4423: std_logic; attribute dont_touch of G4423: signal is true;
	signal G4427: std_logic; attribute dont_touch of G4427: signal is true;
	signal G4430: std_logic; attribute dont_touch of G4430: signal is true;
	signal G4434: std_logic; attribute dont_touch of G4434: signal is true;
	signal G4438: std_logic; attribute dont_touch of G4438: signal is true;
	signal G4443: std_logic; attribute dont_touch of G4443: signal is true;
	signal G4446: std_logic; attribute dont_touch of G4446: signal is true;
	signal G4449: std_logic; attribute dont_touch of G4449: signal is true;
	signal G4452: std_logic; attribute dont_touch of G4452: signal is true;
	signal G4455: std_logic; attribute dont_touch of G4455: signal is true;
	signal G4456: std_logic; attribute dont_touch of G4456: signal is true;
	signal G4459: std_logic; attribute dont_touch of G4459: signal is true;
	signal G4462: std_logic; attribute dont_touch of G4462: signal is true;
	signal G4467: std_logic; attribute dont_touch of G4467: signal is true;
	signal G4473: std_logic; attribute dont_touch of G4473: signal is true;
	signal G4474: std_logic; attribute dont_touch of G4474: signal is true;
	signal G4477: std_logic; attribute dont_touch of G4477: signal is true;
	signal G4480: std_logic; attribute dont_touch of G4480: signal is true;
	signal G4483: std_logic; attribute dont_touch of G4483: signal is true;
	signal G4486: std_logic; attribute dont_touch of G4486: signal is true;
	signal G4489: std_logic; attribute dont_touch of G4489: signal is true;
	signal G4492: std_logic; attribute dont_touch of G4492: signal is true;
	signal G4495: std_logic; attribute dont_touch of G4495: signal is true;
	signal G4498: std_logic; attribute dont_touch of G4498: signal is true;
	signal G4501: std_logic; attribute dont_touch of G4501: signal is true;
	signal G4504: std_logic; attribute dont_touch of G4504: signal is true;
	signal G4507: std_logic; attribute dont_touch of G4507: signal is true;
	signal G4512: std_logic; attribute dont_touch of G4512: signal is true;
	signal G4515: std_logic; attribute dont_touch of G4515: signal is true;
	signal G4519: std_logic; attribute dont_touch of G4519: signal is true;
	signal G4520: std_logic; attribute dont_touch of G4520: signal is true;
	signal G4521: std_logic; attribute dont_touch of G4521: signal is true;
	signal G4527: std_logic; attribute dont_touch of G4527: signal is true;
	signal G4531: std_logic; attribute dont_touch of G4531: signal is true;
	signal G4534: std_logic; attribute dont_touch of G4534: signal is true;
	signal G4537: std_logic; attribute dont_touch of G4537: signal is true;
	signal G4540: std_logic; attribute dont_touch of G4540: signal is true;
	signal G4543: std_logic; attribute dont_touch of G4543: signal is true;
	signal G4546: std_logic; attribute dont_touch of G4546: signal is true;
	signal G4549: std_logic; attribute dont_touch of G4549: signal is true;
	signal G4552: std_logic; attribute dont_touch of G4552: signal is true;
	signal G4555: std_logic; attribute dont_touch of G4555: signal is true;
	signal G4558: std_logic; attribute dont_touch of G4558: signal is true;
	signal G4561: std_logic; attribute dont_touch of G4561: signal is true;
	signal G4564: std_logic; attribute dont_touch of G4564: signal is true;
	signal G4567: std_logic; attribute dont_touch of G4567: signal is true;
	signal G4570: std_logic; attribute dont_touch of G4570: signal is true;
	signal G4571: std_logic; attribute dont_touch of G4571: signal is true;
	signal G4572: std_logic; attribute dont_touch of G4572: signal is true;
	signal G4575: std_logic; attribute dont_touch of G4575: signal is true;
	signal G4578: std_logic; attribute dont_touch of G4578: signal is true;
	signal G4581: std_logic; attribute dont_touch of G4581: signal is true;
	signal G4584: std_logic; attribute dont_touch of G4584: signal is true;
	signal G4593: std_logic; attribute dont_touch of G4593: signal is true;
	signal G4601: std_logic; attribute dont_touch of G4601: signal is true;
	signal G4608: std_logic; attribute dont_touch of G4608: signal is true;
	signal G4616: std_logic; attribute dont_touch of G4616: signal is true;
	signal G4621: std_logic; attribute dont_touch of G4621: signal is true;
	signal G4628: std_logic; attribute dont_touch of G4628: signal is true;
	signal G4633: std_logic; attribute dont_touch of G4633: signal is true;
	signal G4639: std_logic; attribute dont_touch of G4639: signal is true;
	signal G4643: std_logic; attribute dont_touch of G4643: signal is true;
	signal G4646: std_logic; attribute dont_touch of G4646: signal is true;
	signal G4653: std_logic; attribute dont_touch of G4653: signal is true;
	signal G4659: std_logic; attribute dont_touch of G4659: signal is true;
	signal G4664: std_logic; attribute dont_touch of G4664: signal is true;
	signal G4669: std_logic; attribute dont_touch of G4669: signal is true;
	signal G4674: std_logic; attribute dont_touch of G4674: signal is true;
	signal G4681: std_logic; attribute dont_touch of G4681: signal is true;
	signal G4688: std_logic; attribute dont_touch of G4688: signal is true;
	signal G4698: std_logic; attribute dont_touch of G4698: signal is true;
	signal G4704: std_logic; attribute dont_touch of G4704: signal is true;
	signal G4709: std_logic; attribute dont_touch of G4709: signal is true;
	signal G4717: std_logic; attribute dont_touch of G4717: signal is true;
	signal G4722: std_logic; attribute dont_touch of G4722: signal is true;
	signal G4727: std_logic; attribute dont_touch of G4727: signal is true;
	signal G4732: std_logic; attribute dont_touch of G4732: signal is true;
	signal G4737: std_logic; attribute dont_touch of G4737: signal is true;
	signal G4741: std_logic; attribute dont_touch of G4741: signal is true;
	signal G4742: std_logic; attribute dont_touch of G4742: signal is true;
	signal G4743: std_logic; attribute dont_touch of G4743: signal is true;
	signal G4749: std_logic; attribute dont_touch of G4749: signal is true;
	signal G4754: std_logic; attribute dont_touch of G4754: signal is true;
	signal G4760: std_logic; attribute dont_touch of G4760: signal is true;
	signal G4765: std_logic; attribute dont_touch of G4765: signal is true;
	signal G4771: std_logic; attribute dont_touch of G4771: signal is true;
	signal G4776: std_logic; attribute dont_touch of G4776: signal is true;
	signal G4785: std_logic; attribute dont_touch of G4785: signal is true;
	signal G4793: std_logic; attribute dont_touch of G4793: signal is true;
	signal G4801: std_logic; attribute dont_touch of G4801: signal is true;
	signal G4809: std_logic; attribute dont_touch of G4809: signal is true;
	signal G4812: std_logic; attribute dont_touch of G4812: signal is true;
	signal G4815: std_logic; attribute dont_touch of G4815: signal is true;
	signal G4818: std_logic; attribute dont_touch of G4818: signal is true;
	signal G4821: std_logic; attribute dont_touch of G4821: signal is true;
	signal G4826: std_logic; attribute dont_touch of G4826: signal is true;
	signal G4831: std_logic; attribute dont_touch of G4831: signal is true;
	signal G4836: std_logic; attribute dont_touch of G4836: signal is true;
	signal G4843: std_logic; attribute dont_touch of G4843: signal is true;
	signal G4849: std_logic; attribute dont_touch of G4849: signal is true;
	signal G4854: std_logic; attribute dont_touch of G4854: signal is true;
	signal G4859: std_logic; attribute dont_touch of G4859: signal is true;
	signal G4864: std_logic; attribute dont_touch of G4864: signal is true;
	signal G4871: std_logic; attribute dont_touch of G4871: signal is true;
	signal G4878: std_logic; attribute dont_touch of G4878: signal is true;
	signal G4888: std_logic; attribute dont_touch of G4888: signal is true;
	signal G4894: std_logic; attribute dont_touch of G4894: signal is true;
	signal G4899: std_logic; attribute dont_touch of G4899: signal is true;
	signal G4907: std_logic; attribute dont_touch of G4907: signal is true;
	signal G4912: std_logic; attribute dont_touch of G4912: signal is true;
	signal G4917: std_logic; attribute dont_touch of G4917: signal is true;
	signal G4922: std_logic; attribute dont_touch of G4922: signal is true;
	signal G4927: std_logic; attribute dont_touch of G4927: signal is true;
	signal G4931: std_logic; attribute dont_touch of G4931: signal is true;
	signal G4932: std_logic; attribute dont_touch of G4932: signal is true;
	signal G4933: std_logic; attribute dont_touch of G4933: signal is true;
	signal G4939: std_logic; attribute dont_touch of G4939: signal is true;
	signal G4944: std_logic; attribute dont_touch of G4944: signal is true;
	signal G4950: std_logic; attribute dont_touch of G4950: signal is true;
	signal G4955: std_logic; attribute dont_touch of G4955: signal is true;
	signal G4961: std_logic; attribute dont_touch of G4961: signal is true;
	signal G4966: std_logic; attribute dont_touch of G4966: signal is true;
	signal G4975: std_logic; attribute dont_touch of G4975: signal is true;
	signal G4983: std_logic; attribute dont_touch of G4983: signal is true;
	signal G4991: std_logic; attribute dont_touch of G4991: signal is true;
	signal G4999: std_logic; attribute dont_touch of G4999: signal is true;
	signal G5002: std_logic; attribute dont_touch of G5002: signal is true;
	signal G5005: std_logic; attribute dont_touch of G5005: signal is true;
	signal G5008: std_logic; attribute dont_touch of G5008: signal is true;
	signal G5011: std_logic; attribute dont_touch of G5011: signal is true;
	signal G5016: std_logic; attribute dont_touch of G5016: signal is true;
	signal G5022: std_logic; attribute dont_touch of G5022: signal is true;
	signal G5029: std_logic; attribute dont_touch of G5029: signal is true;
	signal G5033: std_logic; attribute dont_touch of G5033: signal is true;
	signal G5037: std_logic; attribute dont_touch of G5037: signal is true;
	signal G5041: std_logic; attribute dont_touch of G5041: signal is true;
	signal G5046: std_logic; attribute dont_touch of G5046: signal is true;
	signal G5052: std_logic; attribute dont_touch of G5052: signal is true;
	signal G5057: std_logic; attribute dont_touch of G5057: signal is true;
	signal G5062: std_logic; attribute dont_touch of G5062: signal is true;
	signal G5069: std_logic; attribute dont_touch of G5069: signal is true;
	signal G5073: std_logic; attribute dont_touch of G5073: signal is true;
	signal G5077: std_logic; attribute dont_touch of G5077: signal is true;
	signal G5080: std_logic; attribute dont_touch of G5080: signal is true;
	signal G5084: std_logic; attribute dont_touch of G5084: signal is true;
	signal G5092: std_logic; attribute dont_touch of G5092: signal is true;
	signal G5097: std_logic; attribute dont_touch of G5097: signal is true;
	signal G5101: std_logic; attribute dont_touch of G5101: signal is true;
	signal G5105: std_logic; attribute dont_touch of G5105: signal is true;
	signal G5109: std_logic; attribute dont_touch of G5109: signal is true;
	signal G5112: std_logic; attribute dont_touch of G5112: signal is true;
	signal G5115: std_logic; attribute dont_touch of G5115: signal is true;
	signal G5120: std_logic; attribute dont_touch of G5120: signal is true;
	signal G5124: std_logic; attribute dont_touch of G5124: signal is true;
	signal G5128: std_logic; attribute dont_touch of G5128: signal is true;
	signal G5134: std_logic; attribute dont_touch of G5134: signal is true;
	signal G5138: std_logic; attribute dont_touch of G5138: signal is true;
	signal G5142: std_logic; attribute dont_touch of G5142: signal is true;
	signal G5148: std_logic; attribute dont_touch of G5148: signal is true;
	signal G5152: std_logic; attribute dont_touch of G5152: signal is true;
	signal G5156: std_logic; attribute dont_touch of G5156: signal is true;
	signal G5160: std_logic; attribute dont_touch of G5160: signal is true;
	signal G5164: std_logic; attribute dont_touch of G5164: signal is true;
	signal G5170: std_logic; attribute dont_touch of G5170: signal is true;
	signal G5176: std_logic; attribute dont_touch of G5176: signal is true;
	signal G5180: std_logic; attribute dont_touch of G5180: signal is true;
	signal G5188: std_logic; attribute dont_touch of G5188: signal is true;
	signal G5196: std_logic; attribute dont_touch of G5196: signal is true;
	signal G5200: std_logic; attribute dont_touch of G5200: signal is true;
	signal G5204: std_logic; attribute dont_touch of G5204: signal is true;
	signal G5208: std_logic; attribute dont_touch of G5208: signal is true;
	signal G5212: std_logic; attribute dont_touch of G5212: signal is true;
	signal G5216: std_logic; attribute dont_touch of G5216: signal is true;
	signal G5220: std_logic; attribute dont_touch of G5220: signal is true;
	signal G5224: std_logic; attribute dont_touch of G5224: signal is true;
	signal G5228: std_logic; attribute dont_touch of G5228: signal is true;
	signal G5232: std_logic; attribute dont_touch of G5232: signal is true;
	signal G5236: std_logic; attribute dont_touch of G5236: signal is true;
	signal G5240: std_logic; attribute dont_touch of G5240: signal is true;
	signal G5244: std_logic; attribute dont_touch of G5244: signal is true;
	signal G5248: std_logic; attribute dont_touch of G5248: signal is true;
	signal G5252: std_logic; attribute dont_touch of G5252: signal is true;
	signal G5256: std_logic; attribute dont_touch of G5256: signal is true;
	signal G5260: std_logic; attribute dont_touch of G5260: signal is true;
	signal G5264: std_logic; attribute dont_touch of G5264: signal is true;
	signal G5268: std_logic; attribute dont_touch of G5268: signal is true;
	signal G5272: std_logic; attribute dont_touch of G5272: signal is true;
	signal G5276: std_logic; attribute dont_touch of G5276: signal is true;
	signal G5283: std_logic; attribute dont_touch of G5283: signal is true;
	signal G5290: std_logic; attribute dont_touch of G5290: signal is true;
	signal G5297: std_logic; attribute dont_touch of G5297: signal is true;
	signal G5308: std_logic; attribute dont_touch of G5308: signal is true;
	signal G5313: std_logic; attribute dont_touch of G5313: signal is true;
	signal G5320: std_logic; attribute dont_touch of G5320: signal is true;
	signal G5327: std_logic; attribute dont_touch of G5327: signal is true;
	signal G5331: std_logic; attribute dont_touch of G5331: signal is true;
	signal G5335: std_logic; attribute dont_touch of G5335: signal is true;
	signal G5339: std_logic; attribute dont_touch of G5339: signal is true;
	signal G5343: std_logic; attribute dont_touch of G5343: signal is true;
	signal G5348: std_logic; attribute dont_touch of G5348: signal is true;
	signal G5352: std_logic; attribute dont_touch of G5352: signal is true;
	signal G5357: std_logic; attribute dont_touch of G5357: signal is true;
	signal G5360: std_logic; attribute dont_touch of G5360: signal is true;
	signal G5366: std_logic; attribute dont_touch of G5366: signal is true;
	signal G5373: std_logic; attribute dont_touch of G5373: signal is true;
	signal G5377: std_logic; attribute dont_touch of G5377: signal is true;
	signal G5381: std_logic; attribute dont_touch of G5381: signal is true;
	signal G5385: std_logic; attribute dont_touch of G5385: signal is true;
	signal G5390: std_logic; attribute dont_touch of G5390: signal is true;
	signal G5396: std_logic; attribute dont_touch of G5396: signal is true;
	signal G5401: std_logic; attribute dont_touch of G5401: signal is true;
	signal G5406: std_logic; attribute dont_touch of G5406: signal is true;
	signal G5413: std_logic; attribute dont_touch of G5413: signal is true;
	signal G5417: std_logic; attribute dont_touch of G5417: signal is true;
	signal G5421: std_logic; attribute dont_touch of G5421: signal is true;
	signal G5424: std_logic; attribute dont_touch of G5424: signal is true;
	signal G5428: std_logic; attribute dont_touch of G5428: signal is true;
	signal G5436: std_logic; attribute dont_touch of G5436: signal is true;
	signal G5441: std_logic; attribute dont_touch of G5441: signal is true;
	signal G5445: std_logic; attribute dont_touch of G5445: signal is true;
	signal G5448: std_logic; attribute dont_touch of G5448: signal is true;
	signal G5452: std_logic; attribute dont_touch of G5452: signal is true;
	signal G5456: std_logic; attribute dont_touch of G5456: signal is true;
	signal G5459: std_logic; attribute dont_touch of G5459: signal is true;
	signal G5462: std_logic; attribute dont_touch of G5462: signal is true;
	signal G5467: std_logic; attribute dont_touch of G5467: signal is true;
	signal G5471: std_logic; attribute dont_touch of G5471: signal is true;
	signal G5475: std_logic; attribute dont_touch of G5475: signal is true;
	signal G5481: std_logic; attribute dont_touch of G5481: signal is true;
	signal G5485: std_logic; attribute dont_touch of G5485: signal is true;
	signal G5489: std_logic; attribute dont_touch of G5489: signal is true;
	signal G5495: std_logic; attribute dont_touch of G5495: signal is true;
	signal G5499: std_logic; attribute dont_touch of G5499: signal is true;
	signal G5503: std_logic; attribute dont_touch of G5503: signal is true;
	signal G5507: std_logic; attribute dont_touch of G5507: signal is true;
	signal G5511: std_logic; attribute dont_touch of G5511: signal is true;
	signal G5517: std_logic; attribute dont_touch of G5517: signal is true;
	signal G5523: std_logic; attribute dont_touch of G5523: signal is true;
	signal G5527: std_logic; attribute dont_touch of G5527: signal is true;
	signal G5535: std_logic; attribute dont_touch of G5535: signal is true;
	signal G5543: std_logic; attribute dont_touch of G5543: signal is true;
	signal G5547: std_logic; attribute dont_touch of G5547: signal is true;
	signal G5551: std_logic; attribute dont_touch of G5551: signal is true;
	signal G5555: std_logic; attribute dont_touch of G5555: signal is true;
	signal G5559: std_logic; attribute dont_touch of G5559: signal is true;
	signal G5563: std_logic; attribute dont_touch of G5563: signal is true;
	signal G5567: std_logic; attribute dont_touch of G5567: signal is true;
	signal G5571: std_logic; attribute dont_touch of G5571: signal is true;
	signal G5575: std_logic; attribute dont_touch of G5575: signal is true;
	signal G5579: std_logic; attribute dont_touch of G5579: signal is true;
	signal G5583: std_logic; attribute dont_touch of G5583: signal is true;
	signal G5587: std_logic; attribute dont_touch of G5587: signal is true;
	signal G5591: std_logic; attribute dont_touch of G5591: signal is true;
	signal G5595: std_logic; attribute dont_touch of G5595: signal is true;
	signal G5599: std_logic; attribute dont_touch of G5599: signal is true;
	signal G5603: std_logic; attribute dont_touch of G5603: signal is true;
	signal G5607: std_logic; attribute dont_touch of G5607: signal is true;
	signal G5611: std_logic; attribute dont_touch of G5611: signal is true;
	signal G5615: std_logic; attribute dont_touch of G5615: signal is true;
	signal G5619: std_logic; attribute dont_touch of G5619: signal is true;
	signal G5623: std_logic; attribute dont_touch of G5623: signal is true;
	signal G5630: std_logic; attribute dont_touch of G5630: signal is true;
	signal G5637: std_logic; attribute dont_touch of G5637: signal is true;
	signal G5644: std_logic; attribute dont_touch of G5644: signal is true;
	signal G5654: std_logic; attribute dont_touch of G5654: signal is true;
	signal G5659: std_logic; attribute dont_touch of G5659: signal is true;
	signal G5666: std_logic; attribute dont_touch of G5666: signal is true;
	signal G5673: std_logic; attribute dont_touch of G5673: signal is true;
	signal G5677: std_logic; attribute dont_touch of G5677: signal is true;
	signal G5681: std_logic; attribute dont_touch of G5681: signal is true;
	signal G5685: std_logic; attribute dont_touch of G5685: signal is true;
	signal G5689: std_logic; attribute dont_touch of G5689: signal is true;
	signal G5694: std_logic; attribute dont_touch of G5694: signal is true;
	signal G5698: std_logic; attribute dont_touch of G5698: signal is true;
	signal G5703: std_logic; attribute dont_touch of G5703: signal is true;
	signal G5706: std_logic; attribute dont_touch of G5706: signal is true;
	signal G5712: std_logic; attribute dont_touch of G5712: signal is true;
	signal G5719: std_logic; attribute dont_touch of G5719: signal is true;
	signal G5723: std_logic; attribute dont_touch of G5723: signal is true;
	signal G5727: std_logic; attribute dont_touch of G5727: signal is true;
	signal G5731: std_logic; attribute dont_touch of G5731: signal is true;
	signal G5736: std_logic; attribute dont_touch of G5736: signal is true;
	signal G5742: std_logic; attribute dont_touch of G5742: signal is true;
	signal G5747: std_logic; attribute dont_touch of G5747: signal is true;
	signal G5752: std_logic; attribute dont_touch of G5752: signal is true;
	signal G5759: std_logic; attribute dont_touch of G5759: signal is true;
	signal G5763: std_logic; attribute dont_touch of G5763: signal is true;
	signal G5767: std_logic; attribute dont_touch of G5767: signal is true;
	signal G5770: std_logic; attribute dont_touch of G5770: signal is true;
	signal G5774: std_logic; attribute dont_touch of G5774: signal is true;
	signal G5782: std_logic; attribute dont_touch of G5782: signal is true;
	signal G5787: std_logic; attribute dont_touch of G5787: signal is true;
	signal G5791: std_logic; attribute dont_touch of G5791: signal is true;
	signal G5794: std_logic; attribute dont_touch of G5794: signal is true;
	signal G5798: std_logic; attribute dont_touch of G5798: signal is true;
	signal G5802: std_logic; attribute dont_touch of G5802: signal is true;
	signal G5805: std_logic; attribute dont_touch of G5805: signal is true;
	signal G5808: std_logic; attribute dont_touch of G5808: signal is true;
	signal G5813: std_logic; attribute dont_touch of G5813: signal is true;
	signal G5817: std_logic; attribute dont_touch of G5817: signal is true;
	signal G5821: std_logic; attribute dont_touch of G5821: signal is true;
	signal G5827: std_logic; attribute dont_touch of G5827: signal is true;
	signal G5831: std_logic; attribute dont_touch of G5831: signal is true;
	signal G5835: std_logic; attribute dont_touch of G5835: signal is true;
	signal G5841: std_logic; attribute dont_touch of G5841: signal is true;
	signal G5845: std_logic; attribute dont_touch of G5845: signal is true;
	signal G5849: std_logic; attribute dont_touch of G5849: signal is true;
	signal G5853: std_logic; attribute dont_touch of G5853: signal is true;
	signal G5857: std_logic; attribute dont_touch of G5857: signal is true;
	signal G5863: std_logic; attribute dont_touch of G5863: signal is true;
	signal G5869: std_logic; attribute dont_touch of G5869: signal is true;
	signal G5873: std_logic; attribute dont_touch of G5873: signal is true;
	signal G5881: std_logic; attribute dont_touch of G5881: signal is true;
	signal G5889: std_logic; attribute dont_touch of G5889: signal is true;
	signal G5893: std_logic; attribute dont_touch of G5893: signal is true;
	signal G5897: std_logic; attribute dont_touch of G5897: signal is true;
	signal G5901: std_logic; attribute dont_touch of G5901: signal is true;
	signal G5905: std_logic; attribute dont_touch of G5905: signal is true;
	signal G5909: std_logic; attribute dont_touch of G5909: signal is true;
	signal G5913: std_logic; attribute dont_touch of G5913: signal is true;
	signal G5917: std_logic; attribute dont_touch of G5917: signal is true;
	signal G5921: std_logic; attribute dont_touch of G5921: signal is true;
	signal G5925: std_logic; attribute dont_touch of G5925: signal is true;
	signal G5929: std_logic; attribute dont_touch of G5929: signal is true;
	signal G5933: std_logic; attribute dont_touch of G5933: signal is true;
	signal G5937: std_logic; attribute dont_touch of G5937: signal is true;
	signal G5941: std_logic; attribute dont_touch of G5941: signal is true;
	signal G5945: std_logic; attribute dont_touch of G5945: signal is true;
	signal G5949: std_logic; attribute dont_touch of G5949: signal is true;
	signal G5953: std_logic; attribute dont_touch of G5953: signal is true;
	signal G5957: std_logic; attribute dont_touch of G5957: signal is true;
	signal G5961: std_logic; attribute dont_touch of G5961: signal is true;
	signal G5965: std_logic; attribute dont_touch of G5965: signal is true;
	signal G5969: std_logic; attribute dont_touch of G5969: signal is true;
	signal G5976: std_logic; attribute dont_touch of G5976: signal is true;
	signal G5983: std_logic; attribute dont_touch of G5983: signal is true;
	signal G5990: std_logic; attribute dont_touch of G5990: signal is true;
	signal G6000: std_logic; attribute dont_touch of G6000: signal is true;
	signal G6005: std_logic; attribute dont_touch of G6005: signal is true;
	signal G6012: std_logic; attribute dont_touch of G6012: signal is true;
	signal G6019: std_logic; attribute dont_touch of G6019: signal is true;
	signal G6023: std_logic; attribute dont_touch of G6023: signal is true;
	signal G6027: std_logic; attribute dont_touch of G6027: signal is true;
	signal G6031: std_logic; attribute dont_touch of G6031: signal is true;
	signal G6035: std_logic; attribute dont_touch of G6035: signal is true;
	signal G6040: std_logic; attribute dont_touch of G6040: signal is true;
	signal G6044: std_logic; attribute dont_touch of G6044: signal is true;
	signal G6049: std_logic; attribute dont_touch of G6049: signal is true;
	signal G6052: std_logic; attribute dont_touch of G6052: signal is true;
	signal G6058: std_logic; attribute dont_touch of G6058: signal is true;
	signal G6065: std_logic; attribute dont_touch of G6065: signal is true;
	signal G6069: std_logic; attribute dont_touch of G6069: signal is true;
	signal G6073: std_logic; attribute dont_touch of G6073: signal is true;
	signal G6077: std_logic; attribute dont_touch of G6077: signal is true;
	signal G6082: std_logic; attribute dont_touch of G6082: signal is true;
	signal G6088: std_logic; attribute dont_touch of G6088: signal is true;
	signal G6093: std_logic; attribute dont_touch of G6093: signal is true;
	signal G6098: std_logic; attribute dont_touch of G6098: signal is true;
	signal G6105: std_logic; attribute dont_touch of G6105: signal is true;
	signal G6109: std_logic; attribute dont_touch of G6109: signal is true;
	signal G6113: std_logic; attribute dont_touch of G6113: signal is true;
	signal G6116: std_logic; attribute dont_touch of G6116: signal is true;
	signal G6120: std_logic; attribute dont_touch of G6120: signal is true;
	signal G6128: std_logic; attribute dont_touch of G6128: signal is true;
	signal G6133: std_logic; attribute dont_touch of G6133: signal is true;
	signal G6137: std_logic; attribute dont_touch of G6137: signal is true;
	signal G6140: std_logic; attribute dont_touch of G6140: signal is true;
	signal G6144: std_logic; attribute dont_touch of G6144: signal is true;
	signal G6148: std_logic; attribute dont_touch of G6148: signal is true;
	signal G6151: std_logic; attribute dont_touch of G6151: signal is true;
	signal G6154: std_logic; attribute dont_touch of G6154: signal is true;
	signal G6159: std_logic; attribute dont_touch of G6159: signal is true;
	signal G6163: std_logic; attribute dont_touch of G6163: signal is true;
	signal G6167: std_logic; attribute dont_touch of G6167: signal is true;
	signal G6173: std_logic; attribute dont_touch of G6173: signal is true;
	signal G6177: std_logic; attribute dont_touch of G6177: signal is true;
	signal G6181: std_logic; attribute dont_touch of G6181: signal is true;
	signal G6187: std_logic; attribute dont_touch of G6187: signal is true;
	signal G6191: std_logic; attribute dont_touch of G6191: signal is true;
	signal G6195: std_logic; attribute dont_touch of G6195: signal is true;
	signal G6199: std_logic; attribute dont_touch of G6199: signal is true;
	signal G6203: std_logic; attribute dont_touch of G6203: signal is true;
	signal G6209: std_logic; attribute dont_touch of G6209: signal is true;
	signal G6215: std_logic; attribute dont_touch of G6215: signal is true;
	signal G6219: std_logic; attribute dont_touch of G6219: signal is true;
	signal G6227: std_logic; attribute dont_touch of G6227: signal is true;
	signal G6235: std_logic; attribute dont_touch of G6235: signal is true;
	signal G6239: std_logic; attribute dont_touch of G6239: signal is true;
	signal G6243: std_logic; attribute dont_touch of G6243: signal is true;
	signal G6247: std_logic; attribute dont_touch of G6247: signal is true;
	signal G6251: std_logic; attribute dont_touch of G6251: signal is true;
	signal G6255: std_logic; attribute dont_touch of G6255: signal is true;
	signal G6259: std_logic; attribute dont_touch of G6259: signal is true;
	signal G6263: std_logic; attribute dont_touch of G6263: signal is true;
	signal G6267: std_logic; attribute dont_touch of G6267: signal is true;
	signal G6271: std_logic; attribute dont_touch of G6271: signal is true;
	signal G6275: std_logic; attribute dont_touch of G6275: signal is true;
	signal G6279: std_logic; attribute dont_touch of G6279: signal is true;
	signal G6283: std_logic; attribute dont_touch of G6283: signal is true;
	signal G6287: std_logic; attribute dont_touch of G6287: signal is true;
	signal G6291: std_logic; attribute dont_touch of G6291: signal is true;
	signal G6295: std_logic; attribute dont_touch of G6295: signal is true;
	signal G6299: std_logic; attribute dont_touch of G6299: signal is true;
	signal G6303: std_logic; attribute dont_touch of G6303: signal is true;
	signal G6307: std_logic; attribute dont_touch of G6307: signal is true;
	signal G6311: std_logic; attribute dont_touch of G6311: signal is true;
	signal G6315: std_logic; attribute dont_touch of G6315: signal is true;
	signal G6322: std_logic; attribute dont_touch of G6322: signal is true;
	signal G6329: std_logic; attribute dont_touch of G6329: signal is true;
	signal G6336: std_logic; attribute dont_touch of G6336: signal is true;
	signal G6346: std_logic; attribute dont_touch of G6346: signal is true;
	signal G6351: std_logic; attribute dont_touch of G6351: signal is true;
	signal G6358: std_logic; attribute dont_touch of G6358: signal is true;
	signal G6365: std_logic; attribute dont_touch of G6365: signal is true;
	signal G6369: std_logic; attribute dont_touch of G6369: signal is true;
	signal G6373: std_logic; attribute dont_touch of G6373: signal is true;
	signal G6377: std_logic; attribute dont_touch of G6377: signal is true;
	signal G6381: std_logic; attribute dont_touch of G6381: signal is true;
	signal G6386: std_logic; attribute dont_touch of G6386: signal is true;
	signal G6390: std_logic; attribute dont_touch of G6390: signal is true;
	signal G6395: std_logic; attribute dont_touch of G6395: signal is true;
	signal G6398: std_logic; attribute dont_touch of G6398: signal is true;
	signal G6404: std_logic; attribute dont_touch of G6404: signal is true;
	signal G6411: std_logic; attribute dont_touch of G6411: signal is true;
	signal G6415: std_logic; attribute dont_touch of G6415: signal is true;
	signal G6419: std_logic; attribute dont_touch of G6419: signal is true;
	signal G6423: std_logic; attribute dont_touch of G6423: signal is true;
	signal G6428: std_logic; attribute dont_touch of G6428: signal is true;
	signal G6434: std_logic; attribute dont_touch of G6434: signal is true;
	signal G6439: std_logic; attribute dont_touch of G6439: signal is true;
	signal G6444: std_logic; attribute dont_touch of G6444: signal is true;
	signal G6451: std_logic; attribute dont_touch of G6451: signal is true;
	signal G6455: std_logic; attribute dont_touch of G6455: signal is true;
	signal G6459: std_logic; attribute dont_touch of G6459: signal is true;
	signal G6462: std_logic; attribute dont_touch of G6462: signal is true;
	signal G6466: std_logic; attribute dont_touch of G6466: signal is true;
	signal G6474: std_logic; attribute dont_touch of G6474: signal is true;
	signal G6479: std_logic; attribute dont_touch of G6479: signal is true;
	signal G6483: std_logic; attribute dont_touch of G6483: signal is true;
	signal G6486: std_logic; attribute dont_touch of G6486: signal is true;
	signal G6490: std_logic; attribute dont_touch of G6490: signal is true;
	signal G6494: std_logic; attribute dont_touch of G6494: signal is true;
	signal G6497: std_logic; attribute dont_touch of G6497: signal is true;
	signal G6500: std_logic; attribute dont_touch of G6500: signal is true;
	signal G6505: std_logic; attribute dont_touch of G6505: signal is true;
	signal G6509: std_logic; attribute dont_touch of G6509: signal is true;
	signal G6513: std_logic; attribute dont_touch of G6513: signal is true;
	signal G6519: std_logic; attribute dont_touch of G6519: signal is true;
	signal G6523: std_logic; attribute dont_touch of G6523: signal is true;
	signal G6527: std_logic; attribute dont_touch of G6527: signal is true;
	signal G6533: std_logic; attribute dont_touch of G6533: signal is true;
	signal G6537: std_logic; attribute dont_touch of G6537: signal is true;
	signal G6541: std_logic; attribute dont_touch of G6541: signal is true;
	signal G6545: std_logic; attribute dont_touch of G6545: signal is true;
	signal G6549: std_logic; attribute dont_touch of G6549: signal is true;
	signal G6555: std_logic; attribute dont_touch of G6555: signal is true;
	signal G6561: std_logic; attribute dont_touch of G6561: signal is true;
	signal G6565: std_logic; attribute dont_touch of G6565: signal is true;
	signal G6573: std_logic; attribute dont_touch of G6573: signal is true;
	signal G6581: std_logic; attribute dont_touch of G6581: signal is true;
	signal G6585: std_logic; attribute dont_touch of G6585: signal is true;
	signal G6589: std_logic; attribute dont_touch of G6589: signal is true;
	signal G6593: std_logic; attribute dont_touch of G6593: signal is true;
	signal G6597: std_logic; attribute dont_touch of G6597: signal is true;
	signal G6601: std_logic; attribute dont_touch of G6601: signal is true;
	signal G6605: std_logic; attribute dont_touch of G6605: signal is true;
	signal G6609: std_logic; attribute dont_touch of G6609: signal is true;
	signal G6613: std_logic; attribute dont_touch of G6613: signal is true;
	signal G6617: std_logic; attribute dont_touch of G6617: signal is true;
	signal G6621: std_logic; attribute dont_touch of G6621: signal is true;
	signal G6625: std_logic; attribute dont_touch of G6625: signal is true;
	signal G6629: std_logic; attribute dont_touch of G6629: signal is true;
	signal G6633: std_logic; attribute dont_touch of G6633: signal is true;
	signal G6637: std_logic; attribute dont_touch of G6637: signal is true;
	signal G6641: std_logic; attribute dont_touch of G6641: signal is true;
	signal G6645: std_logic; attribute dont_touch of G6645: signal is true;
	signal G6649: std_logic; attribute dont_touch of G6649: signal is true;
	signal G6653: std_logic; attribute dont_touch of G6653: signal is true;
	signal G6657: std_logic; attribute dont_touch of G6657: signal is true;
	signal G6661: std_logic; attribute dont_touch of G6661: signal is true;
	signal G6668: std_logic; attribute dont_touch of G6668: signal is true;
	signal G6675: std_logic; attribute dont_touch of G6675: signal is true;
	signal G6682: std_logic; attribute dont_touch of G6682: signal is true;
	signal G6692: std_logic; attribute dont_touch of G6692: signal is true;
	signal G6697: std_logic; attribute dont_touch of G6697: signal is true;
	signal G6704: std_logic; attribute dont_touch of G6704: signal is true;
	signal G6711: std_logic; attribute dont_touch of G6711: signal is true;
	signal G6715: std_logic; attribute dont_touch of G6715: signal is true;
	signal G6719: std_logic; attribute dont_touch of G6719: signal is true;
	signal G6723: std_logic; attribute dont_touch of G6723: signal is true;
	signal G6727: std_logic; attribute dont_touch of G6727: signal is true;
	signal G6732: std_logic; attribute dont_touch of G6732: signal is true;
	signal G6736: std_logic; attribute dont_touch of G6736: signal is true;
	signal G6741: std_logic; attribute dont_touch of G6741: signal is true;
	signal G6754: std_logic; attribute dont_touch of G6754: signal is true;
	signal G6755: std_logic; attribute dont_touch of G6755: signal is true;
	signal G6756: std_logic; attribute dont_touch of G6756: signal is true;
	signal G6767: std_logic; attribute dont_touch of G6767: signal is true;
	signal G6772: std_logic; attribute dont_touch of G6772: signal is true;
	signal G6782: std_logic; attribute dont_touch of G6782: signal is true;
	signal G6789: std_logic; attribute dont_touch of G6789: signal is true;
	signal G6799: std_logic; attribute dont_touch of G6799: signal is true;
	signal G6800: std_logic; attribute dont_touch of G6800: signal is true;
	signal G6801: std_logic; attribute dont_touch of G6801: signal is true;
	signal G6802: std_logic; attribute dont_touch of G6802: signal is true;
	signal G6803: std_logic; attribute dont_touch of G6803: signal is true;
	signal G6804: std_logic; attribute dont_touch of G6804: signal is true;
	signal G6808: std_logic; attribute dont_touch of G6808: signal is true;
	signal G6809: std_logic; attribute dont_touch of G6809: signal is true;
	signal G6810: std_logic; attribute dont_touch of G6810: signal is true;
	signal G6811: std_logic; attribute dont_touch of G6811: signal is true;
	signal G6814: std_logic; attribute dont_touch of G6814: signal is true;
	signal G6815: std_logic; attribute dont_touch of G6815: signal is true;
	signal G6816: std_logic; attribute dont_touch of G6816: signal is true;
	signal G6817: std_logic; attribute dont_touch of G6817: signal is true;
	signal G6818: std_logic; attribute dont_touch of G6818: signal is true;
	signal G6819: std_logic; attribute dont_touch of G6819: signal is true;
	signal G6820: std_logic; attribute dont_touch of G6820: signal is true;
	signal G6821: std_logic; attribute dont_touch of G6821: signal is true;
	signal G6825: std_logic; attribute dont_touch of G6825: signal is true;
	signal G6826: std_logic; attribute dont_touch of G6826: signal is true;
	signal G6827: std_logic; attribute dont_touch of G6827: signal is true;
	signal G6828: std_logic; attribute dont_touch of G6828: signal is true;
	signal G6829: std_logic; attribute dont_touch of G6829: signal is true;
	signal G6830: std_logic; attribute dont_touch of G6830: signal is true;
	signal G6831: std_logic; attribute dont_touch of G6831: signal is true;
	signal G6832: std_logic; attribute dont_touch of G6832: signal is true;
	signal G6836: std_logic; attribute dont_touch of G6836: signal is true;
	signal G6837: std_logic; attribute dont_touch of G6837: signal is true;
	signal G6838: std_logic; attribute dont_touch of G6838: signal is true;
	signal G6839: std_logic; attribute dont_touch of G6839: signal is true;
	signal G6840: std_logic; attribute dont_touch of G6840: signal is true;
	signal G6841: std_logic; attribute dont_touch of G6841: signal is true;
	signal G6845: std_logic; attribute dont_touch of G6845: signal is true;
	signal G6846: std_logic; attribute dont_touch of G6846: signal is true;
	signal G6847: std_logic; attribute dont_touch of G6847: signal is true;
	signal G6848: std_logic; attribute dont_touch of G6848: signal is true;
	signal G6849: std_logic; attribute dont_touch of G6849: signal is true;
	signal G6850: std_logic; attribute dont_touch of G6850: signal is true;
	signal G6854: std_logic; attribute dont_touch of G6854: signal is true;
	signal G6855: std_logic; attribute dont_touch of G6855: signal is true;
	signal G6856: std_logic; attribute dont_touch of G6856: signal is true;
	signal G6867: std_logic; attribute dont_touch of G6867: signal is true;
	signal G6868: std_logic; attribute dont_touch of G6868: signal is true;
	signal G6869: std_logic; attribute dont_touch of G6869: signal is true;
	signal G6870: std_logic; attribute dont_touch of G6870: signal is true;
	signal G6873: std_logic; attribute dont_touch of G6873: signal is true;
	signal G6874: std_logic; attribute dont_touch of G6874: signal is true;
	signal G6875: std_logic; attribute dont_touch of G6875: signal is true;
	signal G6887: std_logic; attribute dont_touch of G6887: signal is true;
	signal G6888: std_logic; attribute dont_touch of G6888: signal is true;
	signal G6895: std_logic; attribute dont_touch of G6895: signal is true;
	signal G6900: std_logic; attribute dont_touch of G6900: signal is true;
	signal G6903: std_logic; attribute dont_touch of G6903: signal is true;
	signal G6904: std_logic; attribute dont_touch of G6904: signal is true;
	signal G6905: std_logic; attribute dont_touch of G6905: signal is true;
	signal G6917: std_logic; attribute dont_touch of G6917: signal is true;
	signal G6918: std_logic; attribute dont_touch of G6918: signal is true;
	signal G6923: std_logic; attribute dont_touch of G6923: signal is true;
	signal G6926: std_logic; attribute dont_touch of G6926: signal is true;
	signal G6927: std_logic; attribute dont_touch of G6927: signal is true;
	signal G6928: std_logic; attribute dont_touch of G6928: signal is true;
	signal G6940: std_logic; attribute dont_touch of G6940: signal is true;
	signal G6941: std_logic; attribute dont_touch of G6941: signal is true;
	signal G6946: std_logic; attribute dont_touch of G6946: signal is true;
	signal G6953: std_logic; attribute dont_touch of G6953: signal is true;
	signal G6954: std_logic; attribute dont_touch of G6954: signal is true;
	signal G6955: std_logic; attribute dont_touch of G6955: signal is true;
	signal G6956: std_logic; attribute dont_touch of G6956: signal is true;
	signal G6957: std_logic; attribute dont_touch of G6957: signal is true;
	signal G6958: std_logic; attribute dont_touch of G6958: signal is true;
	signal G6959: std_logic; attribute dont_touch of G6959: signal is true;
	signal G6960: std_logic; attribute dont_touch of G6960: signal is true;
	signal G6961: std_logic; attribute dont_touch of G6961: signal is true;
	signal G6971: std_logic; attribute dont_touch of G6971: signal is true;
	signal G6972: std_logic; attribute dont_touch of G6972: signal is true;
	signal G6973: std_logic; attribute dont_touch of G6973: signal is true;
	signal G6974: std_logic; attribute dont_touch of G6974: signal is true;
	signal G6975: std_logic; attribute dont_touch of G6975: signal is true;
	signal G6976: std_logic; attribute dont_touch of G6976: signal is true;
	signal G6977: std_logic; attribute dont_touch of G6977: signal is true;
	signal G6978: std_logic; attribute dont_touch of G6978: signal is true;
	signal G6982: std_logic; attribute dont_touch of G6982: signal is true;
	signal G6983: std_logic; attribute dont_touch of G6983: signal is true;
	signal G6984: std_logic; attribute dont_touch of G6984: signal is true;
	signal G6985: std_logic; attribute dont_touch of G6985: signal is true;
	signal G6986: std_logic; attribute dont_touch of G6986: signal is true;
	signal G6987: std_logic; attribute dont_touch of G6987: signal is true;
	signal G6988: std_logic; attribute dont_touch of G6988: signal is true;
	signal G6989: std_logic; attribute dont_touch of G6989: signal is true;
	signal G6990: std_logic; attribute dont_touch of G6990: signal is true;
	signal G6991: std_logic; attribute dont_touch of G6991: signal is true;
	signal G6992: std_logic; attribute dont_touch of G6992: signal is true;
	signal G6993: std_logic; attribute dont_touch of G6993: signal is true;
	signal G6994: std_logic; attribute dont_touch of G6994: signal is true;
	signal G6995: std_logic; attribute dont_touch of G6995: signal is true;
	signal G6996: std_logic; attribute dont_touch of G6996: signal is true;
	signal G6997: std_logic; attribute dont_touch of G6997: signal is true;
	signal G6998: std_logic; attribute dont_touch of G6998: signal is true;
	signal G6999: std_logic; attribute dont_touch of G6999: signal is true;
	signal G7002: std_logic; attribute dont_touch of G7002: signal is true;
	signal G7003: std_logic; attribute dont_touch of G7003: signal is true;
	signal G7004: std_logic; attribute dont_touch of G7004: signal is true;
	signal G7017: std_logic; attribute dont_touch of G7017: signal is true;
	signal G7018: std_logic; attribute dont_touch of G7018: signal is true;
	signal G7023: std_logic; attribute dont_touch of G7023: signal is true;
	signal G7026: std_logic; attribute dont_touch of G7026: signal is true;
	signal G7027: std_logic; attribute dont_touch of G7027: signal is true;
	signal G7028: std_logic; attribute dont_touch of G7028: signal is true;
	signal G7040: std_logic; attribute dont_touch of G7040: signal is true;
	signal G7041: std_logic; attribute dont_touch of G7041: signal is true;
	signal G7046: std_logic; attribute dont_touch of G7046: signal is true;
	signal G7049: std_logic; attribute dont_touch of G7049: signal is true;
	signal G7050: std_logic; attribute dont_touch of G7050: signal is true;
	signal G7051: std_logic; attribute dont_touch of G7051: signal is true;
	signal G7063: std_logic; attribute dont_touch of G7063: signal is true;
	signal G7064: std_logic; attribute dont_touch of G7064: signal is true;
	signal G7069: std_logic; attribute dont_touch of G7069: signal is true;
	signal G7072: std_logic; attribute dont_touch of G7072: signal is true;
	signal G7073: std_logic; attribute dont_touch of G7073: signal is true;
	signal G7074: std_logic; attribute dont_touch of G7074: signal is true;
	signal G7086: std_logic; attribute dont_touch of G7086: signal is true;
	signal G7087: std_logic; attribute dont_touch of G7087: signal is true;
	signal G7092: std_logic; attribute dont_touch of G7092: signal is true;
	signal G7095: std_logic; attribute dont_touch of G7095: signal is true;
	signal G7096: std_logic; attribute dont_touch of G7096: signal is true;
	signal G7097: std_logic; attribute dont_touch of G7097: signal is true;
	signal G7109: std_logic; attribute dont_touch of G7109: signal is true;
	signal G7110: std_logic; attribute dont_touch of G7110: signal is true;
	signal G7115: std_logic; attribute dont_touch of G7115: signal is true;
	signal G7116: std_logic; attribute dont_touch of G7116: signal is true;
	signal G7117: std_logic; attribute dont_touch of G7117: signal is true;
	signal G7118: std_logic; attribute dont_touch of G7118: signal is true;
	signal G7121: std_logic; attribute dont_touch of G7121: signal is true;
	signal G7132: std_logic; attribute dont_touch of G7132: signal is true;
	signal G7133: std_logic; attribute dont_touch of G7133: signal is true;
	signal G7134: std_logic; attribute dont_touch of G7134: signal is true;
	signal G7138: std_logic; attribute dont_touch of G7138: signal is true;
	signal G7139: std_logic; attribute dont_touch of G7139: signal is true;
	signal G7142: std_logic; attribute dont_touch of G7142: signal is true;
	signal G7148: std_logic; attribute dont_touch of G7148: signal is true;
	signal G7149: std_logic; attribute dont_touch of G7149: signal is true;
	signal G7150: std_logic; attribute dont_touch of G7150: signal is true;
	signal G7153: std_logic; attribute dont_touch of G7153: signal is true;
	signal G7157: std_logic; attribute dont_touch of G7157: signal is true;
	signal G7158: std_logic; attribute dont_touch of G7158: signal is true;
	signal G7161: std_logic; attribute dont_touch of G7161: signal is true;
	signal G7162: std_logic; attribute dont_touch of G7162: signal is true;
	signal G7163: std_logic; attribute dont_touch of G7163: signal is true;
	signal G7166: std_logic; attribute dont_touch of G7166: signal is true;
	signal G7167: std_logic; attribute dont_touch of G7167: signal is true;
	signal G7170: std_logic; attribute dont_touch of G7170: signal is true;
	signal G7174: std_logic; attribute dont_touch of G7174: signal is true;
	signal G7175: std_logic; attribute dont_touch of G7175: signal is true;
	signal G7178: std_logic; attribute dont_touch of G7178: signal is true;
	signal G7183: std_logic; attribute dont_touch of G7183: signal is true;
	signal G7184: std_logic; attribute dont_touch of G7184: signal is true;
	signal G7187: std_logic; attribute dont_touch of G7187: signal is true;
	signal G7191: std_logic; attribute dont_touch of G7191: signal is true;
	signal G7192: std_logic; attribute dont_touch of G7192: signal is true;
	signal G7195: std_logic; attribute dont_touch of G7195: signal is true;
	signal G7196: std_logic; attribute dont_touch of G7196: signal is true;
	signal G7197: std_logic; attribute dont_touch of G7197: signal is true;
	signal G7201: std_logic; attribute dont_touch of G7201: signal is true;
	signal G7202: std_logic; attribute dont_touch of G7202: signal is true;
	signal G7209: std_logic; attribute dont_touch of G7209: signal is true;
	signal G7212: std_logic; attribute dont_touch of G7212: signal is true;
	signal G7216: std_logic; attribute dont_touch of G7216: signal is true;
	signal G7219: std_logic; attribute dont_touch of G7219: signal is true;
	signal G7222: std_logic; attribute dont_touch of G7222: signal is true;
	signal G7223: std_logic; attribute dont_touch of G7223: signal is true;
	signal G7224: std_logic; attribute dont_touch of G7224: signal is true;
	signal G7227: std_logic; attribute dont_touch of G7227: signal is true;
	signal G7228: std_logic; attribute dont_touch of G7228: signal is true;
	signal G7231: std_logic; attribute dont_touch of G7231: signal is true;
	signal G7232: std_logic; attribute dont_touch of G7232: signal is true;
	signal G7235: std_logic; attribute dont_touch of G7235: signal is true;
	signal G7236: std_logic; attribute dont_touch of G7236: signal is true;
	signal G7239: std_logic; attribute dont_touch of G7239: signal is true;
	signal G7244: std_logic; attribute dont_touch of G7244: signal is true;
	signal G7246: std_logic; attribute dont_touch of G7246: signal is true;
	signal G7247: std_logic; attribute dont_touch of G7247: signal is true;
	signal G7251: std_logic; attribute dont_touch of G7251: signal is true;
	signal G7252: std_logic; attribute dont_touch of G7252: signal is true;
	signal G7258: std_logic; attribute dont_touch of G7258: signal is true;
	signal G7259: std_logic; attribute dont_touch of G7259: signal is true;
	signal G7261: std_logic; attribute dont_touch of G7261: signal is true;
	signal G7262: std_logic; attribute dont_touch of G7262: signal is true;
	signal G7266: std_logic; attribute dont_touch of G7266: signal is true;
	signal G7267: std_logic; attribute dont_touch of G7267: signal is true;
	signal G7268: std_logic; attribute dont_touch of G7268: signal is true;
	signal G7275: std_logic; attribute dont_touch of G7275: signal is true;
	signal G7280: std_logic; attribute dont_touch of G7280: signal is true;
	signal G7285: std_logic; attribute dont_touch of G7285: signal is true;
	signal G7289: std_logic; attribute dont_touch of G7289: signal is true;
	signal G7293: std_logic; attribute dont_touch of G7293: signal is true;
	signal G7296: std_logic; attribute dont_touch of G7296: signal is true;
	signal G7297: std_logic; attribute dont_touch of G7297: signal is true;
	signal G7301: std_logic; attribute dont_touch of G7301: signal is true;
	signal G7304: std_logic; attribute dont_touch of G7304: signal is true;
	signal G7308: std_logic; attribute dont_touch of G7308: signal is true;
	signal G7314: std_logic; attribute dont_touch of G7314: signal is true;
	signal G7315: std_logic; attribute dont_touch of G7315: signal is true;
	signal G7322: std_logic; attribute dont_touch of G7322: signal is true;
	signal G7327: std_logic; attribute dont_touch of G7327: signal is true;
	signal G7328: std_logic; attribute dont_touch of G7328: signal is true;
	signal G7335: std_logic; attribute dont_touch of G7335: signal is true;
	signal G7340: std_logic; attribute dont_touch of G7340: signal is true;
	signal G7343: std_logic; attribute dont_touch of G7343: signal is true;
	signal G7344: std_logic; attribute dont_touch of G7344: signal is true;
	signal G7345: std_logic; attribute dont_touch of G7345: signal is true;
	signal G7349: std_logic; attribute dont_touch of G7349: signal is true;
	signal G7352: std_logic; attribute dont_touch of G7352: signal is true;
	signal G7356: std_logic; attribute dont_touch of G7356: signal is true;
	signal G7361: std_logic; attribute dont_touch of G7361: signal is true;
	signal G7362: std_logic; attribute dont_touch of G7362: signal is true;
	signal G7369: std_logic; attribute dont_touch of G7369: signal is true;
	signal G7374: std_logic; attribute dont_touch of G7374: signal is true;
	signal G7379: std_logic; attribute dont_touch of G7379: signal is true;
	signal G7380: std_logic; attribute dont_touch of G7380: signal is true;
	signal G7387: std_logic; attribute dont_touch of G7387: signal is true;
	signal G7392: std_logic; attribute dont_touch of G7392: signal is true;
	signal G7393: std_logic; attribute dont_touch of G7393: signal is true;
	signal G7394: std_logic; attribute dont_touch of G7394: signal is true;
	signal G7395: std_logic; attribute dont_touch of G7395: signal is true;
	signal G7396: std_logic; attribute dont_touch of G7396: signal is true;
	signal G7397: std_logic; attribute dont_touch of G7397: signal is true;
	signal G7400: std_logic; attribute dont_touch of G7400: signal is true;
	signal G7404: std_logic; attribute dont_touch of G7404: signal is true;
	signal G7405: std_logic; attribute dont_touch of G7405: signal is true;
	signal G7410: std_logic; attribute dont_touch of G7410: signal is true;
	signal G7411: std_logic; attribute dont_touch of G7411: signal is true;
	signal G7418: std_logic; attribute dont_touch of G7418: signal is true;
	signal G7423: std_logic; attribute dont_touch of G7423: signal is true;
	signal G7424: std_logic; attribute dont_touch of G7424: signal is true;
	signal G7431: std_logic; attribute dont_touch of G7431: signal is true;
	signal G7436: std_logic; attribute dont_touch of G7436: signal is true;
	signal G7437: std_logic; attribute dont_touch of G7437: signal is true;
	signal G7438: std_logic; attribute dont_touch of G7438: signal is true;
	signal G7439: std_logic; attribute dont_touch of G7439: signal is true;
	signal G7440: std_logic; attribute dont_touch of G7440: signal is true;
	signal G7441: std_logic; attribute dont_touch of G7441: signal is true;
	signal G7442: std_logic; attribute dont_touch of G7442: signal is true;
	signal G7443: std_logic; attribute dont_touch of G7443: signal is true;
	signal G7446: std_logic; attribute dont_touch of G7446: signal is true;
	signal G7450: std_logic; attribute dont_touch of G7450: signal is true;
	signal G7451: std_logic; attribute dont_touch of G7451: signal is true;
	signal G7456: std_logic; attribute dont_touch of G7456: signal is true;
	signal G7461: std_logic; attribute dont_touch of G7461: signal is true;
	signal G7462: std_logic; attribute dont_touch of G7462: signal is true;
	signal G7469: std_logic; attribute dont_touch of G7469: signal is true;
	signal G7470: std_logic; attribute dont_touch of G7470: signal is true;
	signal G7471: std_logic; attribute dont_touch of G7471: signal is true;
	signal G7472: std_logic; attribute dont_touch of G7472: signal is true;
	signal G7473: std_logic; attribute dont_touch of G7473: signal is true;
	signal G7474: std_logic; attribute dont_touch of G7474: signal is true;
	signal G7475: std_logic; attribute dont_touch of G7475: signal is true;
	signal G7479: std_logic; attribute dont_touch of G7479: signal is true;
	signal G7487: std_logic; attribute dont_touch of G7487: signal is true;
	signal G7490: std_logic; attribute dont_touch of G7490: signal is true;
	signal G7495: std_logic; attribute dont_touch of G7495: signal is true;
	signal G7496: std_logic; attribute dont_touch of G7496: signal is true;
	signal G7497: std_logic; attribute dont_touch of G7497: signal is true;
	signal G7498: std_logic; attribute dont_touch of G7498: signal is true;
	signal G7499: std_logic; attribute dont_touch of G7499: signal is true;
	signal G7502: std_logic; attribute dont_touch of G7502: signal is true;
	signal G7503: std_logic; attribute dont_touch of G7503: signal is true;
	signal G7511: std_logic; attribute dont_touch of G7511: signal is true;
	signal G7512: std_logic; attribute dont_touch of G7512: signal is true;
	signal G7513: std_logic; attribute dont_touch of G7513: signal is true;
	signal G7514: std_logic; attribute dont_touch of G7514: signal is true;
	signal G7515: std_logic; attribute dont_touch of G7515: signal is true;
	signal G7516: std_logic; attribute dont_touch of G7516: signal is true;
	signal G7517: std_logic; attribute dont_touch of G7517: signal is true;
	signal G7518: std_logic; attribute dont_touch of G7518: signal is true;
	signal G7519: std_logic; attribute dont_touch of G7519: signal is true;
	signal G7520: std_logic; attribute dont_touch of G7520: signal is true;
	signal G7521: std_logic; attribute dont_touch of G7521: signal is true;
	signal G7522: std_logic; attribute dont_touch of G7522: signal is true;
	signal G7523: std_logic; attribute dont_touch of G7523: signal is true;
	signal G7526: std_logic; attribute dont_touch of G7526: signal is true;
	signal G7527: std_logic; attribute dont_touch of G7527: signal is true;
	signal G7528: std_logic; attribute dont_touch of G7528: signal is true;
	signal G7532: std_logic; attribute dont_touch of G7532: signal is true;
	signal G7533: std_logic; attribute dont_touch of G7533: signal is true;
	signal G7534: std_logic; attribute dont_touch of G7534: signal is true;
	signal G7535: std_logic; attribute dont_touch of G7535: signal is true;
	signal G7536: std_logic; attribute dont_touch of G7536: signal is true;
	signal G7537: std_logic; attribute dont_touch of G7537: signal is true;
	signal G7541: std_logic; attribute dont_touch of G7541: signal is true;
	signal G7542: std_logic; attribute dont_touch of G7542: signal is true;
	signal G7543: std_logic; attribute dont_touch of G7543: signal is true;
	signal G7544: std_logic; attribute dont_touch of G7544: signal is true;
	signal G7548: std_logic; attribute dont_touch of G7548: signal is true;
	signal G7549: std_logic; attribute dont_touch of G7549: signal is true;
	signal G7553: std_logic; attribute dont_touch of G7553: signal is true;
	signal G7557: std_logic; attribute dont_touch of G7557: signal is true;
	signal G7558: std_logic; attribute dont_touch of G7558: signal is true;
	signal G7563: std_logic; attribute dont_touch of G7563: signal is true;
	signal G7564: std_logic; attribute dont_touch of G7564: signal is true;
	signal G7565: std_logic; attribute dont_touch of G7565: signal is true;
	signal G7566: std_logic; attribute dont_touch of G7566: signal is true;
	signal G7567: std_logic; attribute dont_touch of G7567: signal is true;
	signal G7577: std_logic; attribute dont_touch of G7577: signal is true;
	signal G7581: std_logic; attribute dont_touch of G7581: signal is true;
	signal G7582: std_logic; attribute dont_touch of G7582: signal is true;
	signal G7586: std_logic; attribute dont_touch of G7586: signal is true;
	signal G7591: std_logic; attribute dont_touch of G7591: signal is true;
	signal G7592: std_logic; attribute dont_touch of G7592: signal is true;
	signal G7593: std_logic; attribute dont_touch of G7593: signal is true;
	signal G7594: std_logic; attribute dont_touch of G7594: signal is true;
	signal G7595: std_logic; attribute dont_touch of G7595: signal is true;
	signal G7596: std_logic; attribute dont_touch of G7596: signal is true;
	signal G7597: std_logic; attribute dont_touch of G7597: signal is true;
	signal G7598: std_logic; attribute dont_touch of G7598: signal is true;
	signal G7601: std_logic; attribute dont_touch of G7601: signal is true;
	signal G7611: std_logic; attribute dont_touch of G7611: signal is true;
	signal G7615: std_logic; attribute dont_touch of G7615: signal is true;
	signal G7616: std_logic; attribute dont_touch of G7616: signal is true;
	signal G7617: std_logic; attribute dont_touch of G7617: signal is true;
	signal G7618: std_logic; attribute dont_touch of G7618: signal is true;
	signal G7619: std_logic; attribute dont_touch of G7619: signal is true;
	signal G7620: std_logic; attribute dont_touch of G7620: signal is true;
	signal G7623: std_logic; attribute dont_touch of G7623: signal is true;
	signal G7624: std_logic; attribute dont_touch of G7624: signal is true;
	signal G7625: std_logic; attribute dont_touch of G7625: signal is true;
	signal G7626: std_logic; attribute dont_touch of G7626: signal is true;
	signal G7627: std_logic; attribute dont_touch of G7627: signal is true;
	signal G7631: std_logic; attribute dont_touch of G7631: signal is true;
	signal G7632: std_logic; attribute dont_touch of G7632: signal is true;
	signal G7633: std_logic; attribute dont_touch of G7633: signal is true;
	signal G7634: std_logic; attribute dont_touch of G7634: signal is true;
	signal G7635: std_logic; attribute dont_touch of G7635: signal is true;
	signal G7636: std_logic; attribute dont_touch of G7636: signal is true;
	signal G7640: std_logic; attribute dont_touch of G7640: signal is true;
	signal G7643: std_logic; attribute dont_touch of G7643: signal is true;
	signal G7647: std_logic; attribute dont_touch of G7647: signal is true;
	signal G7648: std_logic; attribute dont_touch of G7648: signal is true;
	signal G7649: std_logic; attribute dont_touch of G7649: signal is true;
	signal G7650: std_logic; attribute dont_touch of G7650: signal is true;
	signal G7655: std_logic; attribute dont_touch of G7655: signal is true;
	signal G7659: std_logic; attribute dont_touch of G7659: signal is true;
	signal G7660: std_logic; attribute dont_touch of G7660: signal is true;
	signal G7661: std_logic; attribute dont_touch of G7661: signal is true;
	signal G7666: std_logic; attribute dont_touch of G7666: signal is true;
	signal G7670: std_logic; attribute dont_touch of G7670: signal is true;
	signal G7673: std_logic; attribute dont_touch of G7673: signal is true;
	signal G7674: std_logic; attribute dont_touch of G7674: signal is true;
	signal G7675: std_logic; attribute dont_touch of G7675: signal is true;
	signal G7680: std_logic; attribute dont_touch of G7680: signal is true;
	signal G7684: std_logic; attribute dont_touch of G7684: signal is true;
	signal G7685: std_logic; attribute dont_touch of G7685: signal is true;
	signal G7686: std_logic; attribute dont_touch of G7686: signal is true;
	signal G7689: std_logic; attribute dont_touch of G7689: signal is true;
	signal G7690: std_logic; attribute dont_touch of G7690: signal is true;
	signal G7693: std_logic; attribute dont_touch of G7693: signal is true;
	signal G7696: std_logic; attribute dont_touch of G7696: signal is true;
	signal G7697: std_logic; attribute dont_touch of G7697: signal is true;
	signal G7701: std_logic; attribute dont_touch of G7701: signal is true;
	signal G7704: std_logic; attribute dont_touch of G7704: signal is true;
	signal G7715: std_logic; attribute dont_touch of G7715: signal is true;
	signal G7716: std_logic; attribute dont_touch of G7716: signal is true;
	signal G7717: std_logic; attribute dont_touch of G7717: signal is true;
	signal G7733: std_logic; attribute dont_touch of G7733: signal is true;
	signal G7738: std_logic; attribute dont_touch of G7738: signal is true;
	signal G7749: std_logic; attribute dont_touch of G7749: signal is true;
	signal G7750: std_logic; attribute dont_touch of G7750: signal is true;
	signal G7751: std_logic; attribute dont_touch of G7751: signal is true;
	signal G7752: std_logic; attribute dont_touch of G7752: signal is true;
	signal G7753: std_logic; attribute dont_touch of G7753: signal is true;
	signal G7763: std_logic; attribute dont_touch of G7763: signal is true;
	signal G7764: std_logic; attribute dont_touch of G7764: signal is true;
	signal G7765: std_logic; attribute dont_touch of G7765: signal is true;
	signal G7766: std_logic; attribute dont_touch of G7766: signal is true;
	signal G7777: std_logic; attribute dont_touch of G7777: signal is true;
	signal G7778: std_logic; attribute dont_touch of G7778: signal is true;
	signal G7779: std_logic; attribute dont_touch of G7779: signal is true;
	signal G7780: std_logic; attribute dont_touch of G7780: signal is true;
	signal G7781: std_logic; attribute dont_touch of G7781: signal is true;
	signal G7785: std_logic; attribute dont_touch of G7785: signal is true;
	signal G7788: std_logic; attribute dont_touch of G7788: signal is true;
	signal G7791: std_logic; attribute dont_touch of G7791: signal is true;
	signal G7802: std_logic; attribute dont_touch of G7802: signal is true;
	signal G7803: std_logic; attribute dont_touch of G7803: signal is true;
	signal G7804: std_logic; attribute dont_touch of G7804: signal is true;
	signal G7805: std_logic; attribute dont_touch of G7805: signal is true;
	signal G7806: std_logic; attribute dont_touch of G7806: signal is true;
	signal G7809: std_logic; attribute dont_touch of G7809: signal is true;
	signal G7812: std_logic; attribute dont_touch of G7812: signal is true;
	signal G7823: std_logic; attribute dont_touch of G7823: signal is true;
	signal G7824: std_logic; attribute dont_touch of G7824: signal is true;
	signal G7827: std_logic; attribute dont_touch of G7827: signal is true;
	signal G7828: std_logic; attribute dont_touch of G7828: signal is true;
	signal G7831: std_logic; attribute dont_touch of G7831: signal is true;
	signal G7834: std_logic; attribute dont_touch of G7834: signal is true;
	signal G7835: std_logic; attribute dont_touch of G7835: signal is true;
	signal G7836: std_logic; attribute dont_touch of G7836: signal is true;
	signal G7840: std_logic; attribute dont_touch of G7840: signal is true;
	signal G7841: std_logic; attribute dont_touch of G7841: signal is true;
	signal G7845: std_logic; attribute dont_touch of G7845: signal is true;
	signal G7846: std_logic; attribute dont_touch of G7846: signal is true;
	signal G7850: std_logic; attribute dont_touch of G7850: signal is true;
	signal G7851: std_logic; attribute dont_touch of G7851: signal is true;
	signal G7854: std_logic; attribute dont_touch of G7854: signal is true;
	signal G7857: std_logic; attribute dont_touch of G7857: signal is true;
	signal G7858: std_logic; attribute dont_touch of G7858: signal is true;
	signal G7863: std_logic; attribute dont_touch of G7863: signal is true;
	signal G7867: std_logic; attribute dont_touch of G7867: signal is true;
	signal G7868: std_logic; attribute dont_touch of G7868: signal is true;
	signal G7869: std_logic; attribute dont_touch of G7869: signal is true;
	signal G7870: std_logic; attribute dont_touch of G7870: signal is true;
	signal G7873: std_logic; attribute dont_touch of G7873: signal is true;
	signal G7876: std_logic; attribute dont_touch of G7876: signal is true;
	signal G7879: std_logic; attribute dont_touch of G7879: signal is true;
	signal G7880: std_logic; attribute dont_touch of G7880: signal is true;
	signal G7885: std_logic; attribute dont_touch of G7885: signal is true;
	signal G7886: std_logic; attribute dont_touch of G7886: signal is true;
	signal G7887: std_logic; attribute dont_touch of G7887: signal is true;
	signal G7888: std_logic; attribute dont_touch of G7888: signal is true;
	signal G7891: std_logic; attribute dont_touch of G7891: signal is true;
	signal G7892: std_logic; attribute dont_touch of G7892: signal is true;
	signal G7897: std_logic; attribute dont_touch of G7897: signal is true;
	signal G7898: std_logic; attribute dont_touch of G7898: signal is true;
	signal G7903: std_logic; attribute dont_touch of G7903: signal is true;
	signal G7907: std_logic; attribute dont_touch of G7907: signal is true;
	signal G7908: std_logic; attribute dont_touch of G7908: signal is true;
	signal G7909: std_logic; attribute dont_touch of G7909: signal is true;
	signal G7913: std_logic; attribute dont_touch of G7913: signal is true;
	signal G7917: std_logic; attribute dont_touch of G7917: signal is true;
	signal G7918: std_logic; attribute dont_touch of G7918: signal is true;
	signal G7922: std_logic; attribute dont_touch of G7922: signal is true;
	signal G7926: std_logic; attribute dont_touch of G7926: signal is true;
	signal G7927: std_logic; attribute dont_touch of G7927: signal is true;
	signal G7928: std_logic; attribute dont_touch of G7928: signal is true;
	signal G7932: std_logic; attribute dont_touch of G7932: signal is true;
	signal G7933: std_logic; attribute dont_touch of G7933: signal is true;
	signal G7936: std_logic; attribute dont_touch of G7936: signal is true;
	signal G7939: std_logic; attribute dont_touch of G7939: signal is true;
	signal G7943: std_logic; attribute dont_touch of G7943: signal is true;
	signal G7947: std_logic; attribute dont_touch of G7947: signal is true;
	signal G7948: std_logic; attribute dont_touch of G7948: signal is true;
	signal G7952: std_logic; attribute dont_touch of G7952: signal is true;
	signal G7953: std_logic; attribute dont_touch of G7953: signal is true;
	signal G7957: std_logic; attribute dont_touch of G7957: signal is true;
	signal G7960: std_logic; attribute dont_touch of G7960: signal is true;
	signal G7963: std_logic; attribute dont_touch of G7963: signal is true;
	signal G7964: std_logic; attribute dont_touch of G7964: signal is true;
	signal G7970: std_logic; attribute dont_touch of G7970: signal is true;
	signal G7971: std_logic; attribute dont_touch of G7971: signal is true;
	signal G7972: std_logic; attribute dont_touch of G7972: signal is true;
	signal G7975: std_logic; attribute dont_touch of G7975: signal is true;
	signal G7980: std_logic; attribute dont_touch of G7980: signal is true;
	signal G7985: std_logic; attribute dont_touch of G7985: signal is true;
	signal G7991: std_logic; attribute dont_touch of G7991: signal is true;
	signal G7992: std_logic; attribute dont_touch of G7992: signal is true;
	signal G7993: std_logic; attribute dont_touch of G7993: signal is true;
	signal G7994: std_logic; attribute dont_touch of G7994: signal is true;
	signal G7995: std_logic; attribute dont_touch of G7995: signal is true;
	signal G7998: std_logic; attribute dont_touch of G7998: signal is true;
	signal G8002: std_logic; attribute dont_touch of G8002: signal is true;
	signal G8005: std_logic; attribute dont_touch of G8005: signal is true;
	signal G8009: std_logic; attribute dont_touch of G8009: signal is true;
	signal G8010: std_logic; attribute dont_touch of G8010: signal is true;
	signal G8011: std_logic; attribute dont_touch of G8011: signal is true;
	signal G8016: std_logic; attribute dont_touch of G8016: signal is true;
	signal G8021: std_logic; attribute dont_touch of G8021: signal is true;
	signal G8026: std_logic; attribute dont_touch of G8026: signal is true;
	signal G8032: std_logic; attribute dont_touch of G8032: signal is true;
	signal G8033: std_logic; attribute dont_touch of G8033: signal is true;
	signal G8037: std_logic; attribute dont_touch of G8037: signal is true;
	signal G8038: std_logic; attribute dont_touch of G8038: signal is true;
	signal G8046: std_logic; attribute dont_touch of G8046: signal is true;
	signal G8052: std_logic; attribute dont_touch of G8052: signal is true;
	signal G8055: std_logic; attribute dont_touch of G8055: signal is true;
	signal G8056: std_logic; attribute dont_touch of G8056: signal is true;
	signal G8057: std_logic; attribute dont_touch of G8057: signal is true;
	signal G8058: std_logic; attribute dont_touch of G8058: signal is true;
	signal G8059: std_logic; attribute dont_touch of G8059: signal is true;
	signal G8064: std_logic; attribute dont_touch of G8064: signal is true;
	signal G8068: std_logic; attribute dont_touch of G8068: signal is true;
	signal G8069: std_logic; attribute dont_touch of G8069: signal is true;
	signal G8070: std_logic; attribute dont_touch of G8070: signal is true;
	signal G8075: std_logic; attribute dont_touch of G8075: signal is true;
	signal G8080: std_logic; attribute dont_touch of G8080: signal is true;
	signal G8085: std_logic; attribute dont_touch of G8085: signal is true;
	signal G8086: std_logic; attribute dont_touch of G8086: signal is true;
	signal G8087: std_logic; attribute dont_touch of G8087: signal is true;
	signal G8088: std_logic; attribute dont_touch of G8088: signal is true;
	signal G8091: std_logic; attribute dont_touch of G8091: signal is true;
	signal G8092: std_logic; attribute dont_touch of G8092: signal is true;
	signal G8093: std_logic; attribute dont_touch of G8093: signal is true;
	signal G8097: std_logic; attribute dont_touch of G8097: signal is true;
	signal G8102: std_logic; attribute dont_touch of G8102: signal is true;
	signal G8105: std_logic; attribute dont_touch of G8105: signal is true;
	signal G8106: std_logic; attribute dont_touch of G8106: signal is true;
	signal G8107: std_logic; attribute dont_touch of G8107: signal is true;
	signal G8112: std_logic; attribute dont_touch of G8112: signal is true;
	signal G8113: std_logic; attribute dont_touch of G8113: signal is true;
	signal G8114: std_logic; attribute dont_touch of G8114: signal is true;
	signal G8119: std_logic; attribute dont_touch of G8119: signal is true;
	signal G8123: std_logic; attribute dont_touch of G8123: signal is true;
	signal G8124: std_logic; attribute dont_touch of G8124: signal is true;
	signal G8125: std_logic; attribute dont_touch of G8125: signal is true;
	signal G8130: std_logic; attribute dont_touch of G8130: signal is true;
	signal G8131: std_logic; attribute dont_touch of G8131: signal is true;
	signal G8133: std_logic; attribute dont_touch of G8133: signal is true;
	signal G8134: std_logic; attribute dont_touch of G8134: signal is true;
	signal G8135: std_logic; attribute dont_touch of G8135: signal is true;
	signal G8136: std_logic; attribute dont_touch of G8136: signal is true;
	signal G8137: std_logic; attribute dont_touch of G8137: signal is true;
	signal G8138: std_logic; attribute dont_touch of G8138: signal is true;
	signal G8139: std_logic; attribute dont_touch of G8139: signal is true;
	signal G8146: std_logic; attribute dont_touch of G8146: signal is true;
	signal G8150: std_logic; attribute dont_touch of G8150: signal is true;
	signal G8154: std_logic; attribute dont_touch of G8154: signal is true;
	signal G8155: std_logic; attribute dont_touch of G8155: signal is true;
	signal G8160: std_logic; attribute dont_touch of G8160: signal is true;
	signal G8163: std_logic; attribute dont_touch of G8163: signal is true;
	signal G8164: std_logic; attribute dont_touch of G8164: signal is true;
	signal G8165: std_logic; attribute dont_touch of G8165: signal is true;
	signal G8170: std_logic; attribute dont_touch of G8170: signal is true;
	signal G8171: std_logic; attribute dont_touch of G8171: signal is true;
	signal G8172: std_logic; attribute dont_touch of G8172: signal is true;
	signal G8177: std_logic; attribute dont_touch of G8177: signal is true;
	signal G8179: std_logic; attribute dont_touch of G8179: signal is true;
	signal G8180: std_logic; attribute dont_touch of G8180: signal is true;
	signal G8181: std_logic; attribute dont_touch of G8181: signal is true;
	signal G8182: std_logic; attribute dont_touch of G8182: signal is true;
	signal G8183: std_logic; attribute dont_touch of G8183: signal is true;
	signal G8186: std_logic; attribute dont_touch of G8186: signal is true;
	signal G8187: std_logic; attribute dont_touch of G8187: signal is true;
	signal G8195: std_logic; attribute dont_touch of G8195: signal is true;
	signal G8201: std_logic; attribute dont_touch of G8201: signal is true;
	signal G8205: std_logic; attribute dont_touch of G8205: signal is true;
	signal G8211: std_logic; attribute dont_touch of G8211: signal is true;
	signal G8216: std_logic; attribute dont_touch of G8216: signal is true;
	signal G8217: std_logic; attribute dont_touch of G8217: signal is true;
	signal G8218: std_logic; attribute dont_touch of G8218: signal is true;
	signal G8219: std_logic; attribute dont_touch of G8219: signal is true;
	signal G8224: std_logic; attribute dont_touch of G8224: signal is true;
	signal G8227: std_logic; attribute dont_touch of G8227: signal is true;
	signal G8228: std_logic; attribute dont_touch of G8228: signal is true;
	signal G8229: std_logic; attribute dont_touch of G8229: signal is true;
	signal G8234: std_logic; attribute dont_touch of G8234: signal is true;
	signal G8236: std_logic; attribute dont_touch of G8236: signal is true;
	signal G8237: std_logic; attribute dont_touch of G8237: signal is true;
	signal G8238: std_logic; attribute dont_touch of G8238: signal is true;
	signal G8239: std_logic; attribute dont_touch of G8239: signal is true;
	signal G8240: std_logic; attribute dont_touch of G8240: signal is true;
	signal G8241: std_logic; attribute dont_touch of G8241: signal is true;
	signal G8249: std_logic; attribute dont_touch of G8249: signal is true;
	signal G8255: std_logic; attribute dont_touch of G8255: signal is true;
	signal G8259: std_logic; attribute dont_touch of G8259: signal is true;
	signal G8267: std_logic; attribute dont_touch of G8267: signal is true;
	signal G8273: std_logic; attribute dont_touch of G8273: signal is true;
	signal G8278: std_logic; attribute dont_touch of G8278: signal is true;
	signal G8280: std_logic; attribute dont_touch of G8280: signal is true;
	signal G8281: std_logic; attribute dont_touch of G8281: signal is true;
	signal G8282: std_logic; attribute dont_touch of G8282: signal is true;
	signal G8284: std_logic; attribute dont_touch of G8284: signal is true;
	signal G8285: std_logic; attribute dont_touch of G8285: signal is true;
	signal G8286: std_logic; attribute dont_touch of G8286: signal is true;
	signal G8287: std_logic; attribute dont_touch of G8287: signal is true;
	signal G8290: std_logic; attribute dont_touch of G8290: signal is true;
	signal G8292: std_logic; attribute dont_touch of G8292: signal is true;
	signal G8296: std_logic; attribute dont_touch of G8296: signal is true;
	signal G8297: std_logic; attribute dont_touch of G8297: signal is true;
	signal G8300: std_logic; attribute dont_touch of G8300: signal is true;
	signal G8301: std_logic; attribute dont_touch of G8301: signal is true;
	signal G8302: std_logic; attribute dont_touch of G8302: signal is true;
	signal G8310: std_logic; attribute dont_touch of G8310: signal is true;
	signal G8316: std_logic; attribute dont_touch of G8316: signal is true;
	signal G8324: std_logic; attribute dont_touch of G8324: signal is true;
	signal G8330: std_logic; attribute dont_touch of G8330: signal is true;
	signal G8334: std_logic; attribute dont_touch of G8334: signal is true;
	signal G8340: std_logic; attribute dont_touch of G8340: signal is true;
	signal G8341: std_logic; attribute dont_touch of G8341: signal is true;
	signal G8343: std_logic; attribute dont_touch of G8343: signal is true;
	signal G8345: std_logic; attribute dont_touch of G8345: signal is true;
	signal G8346: std_logic; attribute dont_touch of G8346: signal is true;
	signal G8347: std_logic; attribute dont_touch of G8347: signal is true;
	signal G8350: std_logic; attribute dont_touch of G8350: signal is true;
	signal G8354: std_logic; attribute dont_touch of G8354: signal is true;
	signal G8355: std_logic; attribute dont_touch of G8355: signal is true;
	signal G8356: std_logic; attribute dont_touch of G8356: signal is true;
	signal G8357: std_logic; attribute dont_touch of G8357: signal is true;
	signal G8359: std_logic; attribute dont_touch of G8359: signal is true;
	signal G8362: std_logic; attribute dont_touch of G8362: signal is true;
	signal G8363: std_logic; attribute dont_touch of G8363: signal is true;
	signal G8364: std_logic; attribute dont_touch of G8364: signal is true;
	signal G8365: std_logic; attribute dont_touch of G8365: signal is true;
	signal G8373: std_logic; attribute dont_touch of G8373: signal is true;
	signal G8381: std_logic; attribute dont_touch of G8381: signal is true;
	signal G8387: std_logic; attribute dont_touch of G8387: signal is true;
	signal G8388: std_logic; attribute dont_touch of G8388: signal is true;
	signal G8389: std_logic; attribute dont_touch of G8389: signal is true;
	signal G8390: std_logic; attribute dont_touch of G8390: signal is true;
	signal G8396: std_logic; attribute dont_touch of G8396: signal is true;
	signal G8397: std_logic; attribute dont_touch of G8397: signal is true;
	signal G8399: std_logic; attribute dont_touch of G8399: signal is true;
	signal G8400: std_logic; attribute dont_touch of G8400: signal is true;
	signal G8404: std_logic; attribute dont_touch of G8404: signal is true;
	signal G8405: std_logic; attribute dont_touch of G8405: signal is true;
	signal G8406: std_logic; attribute dont_touch of G8406: signal is true;
	signal G8407: std_logic; attribute dont_touch of G8407: signal is true;
	signal G8411: std_logic; attribute dont_touch of G8411: signal is true;
	signal G8417: std_logic; attribute dont_touch of G8417: signal is true;
	signal G8418: std_logic; attribute dont_touch of G8418: signal is true;
	signal G8426: std_logic; attribute dont_touch of G8426: signal is true;
	signal G8431: std_logic; attribute dont_touch of G8431: signal is true;
	signal G8434: std_logic; attribute dont_touch of G8434: signal is true;
	signal G8438: std_logic; attribute dont_touch of G8438: signal is true;
	signal G8439: std_logic; attribute dont_touch of G8439: signal is true;
	signal G8440: std_logic; attribute dont_touch of G8440: signal is true;
	signal G8441: std_logic; attribute dont_touch of G8441: signal is true;
	signal G8442: std_logic; attribute dont_touch of G8442: signal is true;
	signal G8443: std_logic; attribute dont_touch of G8443: signal is true;
	signal G8449: std_logic; attribute dont_touch of G8449: signal is true;
	signal G8450: std_logic; attribute dont_touch of G8450: signal is true;
	signal G8451: std_logic; attribute dont_touch of G8451: signal is true;
	signal G8456: std_logic; attribute dont_touch of G8456: signal is true;
	signal G8457: std_logic; attribute dont_touch of G8457: signal is true;
	signal G8458: std_logic; attribute dont_touch of G8458: signal is true;
	signal G8461: std_logic; attribute dont_touch of G8461: signal is true;
	signal G8462: std_logic; attribute dont_touch of G8462: signal is true;
	signal G8466: std_logic; attribute dont_touch of G8466: signal is true;
	signal G8470: std_logic; attribute dont_touch of G8470: signal is true;
	signal G8476: std_logic; attribute dont_touch of G8476: signal is true;
	signal G8477: std_logic; attribute dont_touch of G8477: signal is true;
	signal G8478: std_logic; attribute dont_touch of G8478: signal is true;
	signal G8479: std_logic; attribute dont_touch of G8479: signal is true;
	signal G8480: std_logic; attribute dont_touch of G8480: signal is true;
	signal G8481: std_logic; attribute dont_touch of G8481: signal is true;
	signal G8492: std_logic; attribute dont_touch of G8492: signal is true;
	signal G8497: std_logic; attribute dont_touch of G8497: signal is true;
	signal G8500: std_logic; attribute dont_touch of G8500: signal is true;
	signal G8504: std_logic; attribute dont_touch of G8504: signal is true;
	signal G8505: std_logic; attribute dont_touch of G8505: signal is true;
	signal G8506: std_logic; attribute dont_touch of G8506: signal is true;
	signal G8507: std_logic; attribute dont_touch of G8507: signal is true;
	signal G8508: std_logic; attribute dont_touch of G8508: signal is true;
	signal G8509: std_logic; attribute dont_touch of G8509: signal is true;
	signal G8514: std_logic; attribute dont_touch of G8514: signal is true;
	signal G8515: std_logic; attribute dont_touch of G8515: signal is true;
	signal G8519: std_logic; attribute dont_touch of G8519: signal is true;
	signal G8522: std_logic; attribute dont_touch of G8522: signal is true;
	signal G8526: std_logic; attribute dont_touch of G8526: signal is true;
	signal G8530: std_logic; attribute dont_touch of G8530: signal is true;
	signal G8531: std_logic; attribute dont_touch of G8531: signal is true;
	signal G8534: std_logic; attribute dont_touch of G8534: signal is true;
	signal G8538: std_logic; attribute dont_touch of G8538: signal is true;
	signal G8539: std_logic; attribute dont_touch of G8539: signal is true;
	signal G8540: std_logic; attribute dont_touch of G8540: signal is true;
	signal G8541: std_logic; attribute dont_touch of G8541: signal is true;
	signal G8542: std_logic; attribute dont_touch of G8542: signal is true;
	signal G8553: std_logic; attribute dont_touch of G8553: signal is true;
	signal G8558: std_logic; attribute dont_touch of G8558: signal is true;
	signal G8561: std_logic; attribute dont_touch of G8561: signal is true;
	signal G8565: std_logic; attribute dont_touch of G8565: signal is true;
	signal G8566: std_logic; attribute dont_touch of G8566: signal is true;
	signal G8567: std_logic; attribute dont_touch of G8567: signal is true;
	signal G8571: std_logic; attribute dont_touch of G8571: signal is true;
	signal G8572: std_logic; attribute dont_touch of G8572: signal is true;
	signal G8575: std_logic; attribute dont_touch of G8575: signal is true;
	signal G8579: std_logic; attribute dont_touch of G8579: signal is true;
	signal G8583: std_logic; attribute dont_touch of G8583: signal is true;
	signal G8584: std_logic; attribute dont_touch of G8584: signal is true;
	signal G8587: std_logic; attribute dont_touch of G8587: signal is true;
	signal G8591: std_logic; attribute dont_touch of G8591: signal is true;
	signal G8592: std_logic; attribute dont_touch of G8592: signal is true;
	signal G8593: std_logic; attribute dont_touch of G8593: signal is true;
	signal G8594: std_logic; attribute dont_touch of G8594: signal is true;
	signal G8595: std_logic; attribute dont_touch of G8595: signal is true;
	signal G8606: std_logic; attribute dont_touch of G8606: signal is true;
	signal G8607: std_logic; attribute dont_touch of G8607: signal is true;
	signal G8608: std_logic; attribute dont_touch of G8608: signal is true;
	signal G8609: std_logic; attribute dont_touch of G8609: signal is true;
	signal G8612: std_logic; attribute dont_touch of G8612: signal is true;
	signal G8616: std_logic; attribute dont_touch of G8616: signal is true;
	signal G8620: std_logic; attribute dont_touch of G8620: signal is true;
	signal G8623: std_logic; attribute dont_touch of G8623: signal is true;
	signal G8626: std_logic; attribute dont_touch of G8626: signal is true;
	signal G8630: std_logic; attribute dont_touch of G8630: signal is true;
	signal G8631: std_logic; attribute dont_touch of G8631: signal is true;
	signal G8632: std_logic; attribute dont_touch of G8632: signal is true;
	signal G8635: std_logic; attribute dont_touch of G8635: signal is true;
	signal G8639: std_logic; attribute dont_touch of G8639: signal is true;
	signal G8643: std_logic; attribute dont_touch of G8643: signal is true;
	signal G8644: std_logic; attribute dont_touch of G8644: signal is true;
	signal G8647: std_logic; attribute dont_touch of G8647: signal is true;
	signal G8650: std_logic; attribute dont_touch of G8650: signal is true;
	signal G8651: std_logic; attribute dont_touch of G8651: signal is true;
	signal G8654: std_logic; attribute dont_touch of G8654: signal is true;
	signal G8655: std_logic; attribute dont_touch of G8655: signal is true;
	signal G8659: std_logic; attribute dont_touch of G8659: signal is true;
	signal G8663: std_logic; attribute dont_touch of G8663: signal is true;
	signal G8666: std_logic; attribute dont_touch of G8666: signal is true;
	signal G8669: std_logic; attribute dont_touch of G8669: signal is true;
	signal G8672: std_logic; attribute dont_touch of G8672: signal is true;
	signal G8673: std_logic; attribute dont_touch of G8673: signal is true;
	signal G8676: std_logic; attribute dont_touch of G8676: signal is true;
	signal G8677: std_logic; attribute dont_touch of G8677: signal is true;
	signal G8678: std_logic; attribute dont_touch of G8678: signal is true;
	signal G8679: std_logic; attribute dont_touch of G8679: signal is true;
	signal G8680: std_logic; attribute dont_touch of G8680: signal is true;
	signal G8681: std_logic; attribute dont_touch of G8681: signal is true;
	signal G8685: std_logic; attribute dont_touch of G8685: signal is true;
	signal G8686: std_logic; attribute dont_touch of G8686: signal is true;
	signal G8690: std_logic; attribute dont_touch of G8690: signal is true;
	signal G8691: std_logic; attribute dont_touch of G8691: signal is true;
	signal G8696: std_logic; attribute dont_touch of G8696: signal is true;
	signal G8697: std_logic; attribute dont_touch of G8697: signal is true;
	signal G8700: std_logic; attribute dont_touch of G8700: signal is true;
	signal G8703: std_logic; attribute dont_touch of G8703: signal is true;
	signal G8712: std_logic; attribute dont_touch of G8712: signal is true;
	signal G8713: std_logic; attribute dont_touch of G8713: signal is true;
	signal G8714: std_logic; attribute dont_touch of G8714: signal is true;
	signal G8715: std_logic; attribute dont_touch of G8715: signal is true;
	signal G8718: std_logic; attribute dont_touch of G8718: signal is true;
	signal G8720: std_logic; attribute dont_touch of G8720: signal is true;
	signal G8721: std_logic; attribute dont_touch of G8721: signal is true;
	signal G8725: std_logic; attribute dont_touch of G8725: signal is true;
	signal G8728: std_logic; attribute dont_touch of G8728: signal is true;
	signal G8733: std_logic; attribute dont_touch of G8733: signal is true;
	signal G8734: std_logic; attribute dont_touch of G8734: signal is true;
	signal G8737: std_logic; attribute dont_touch of G8737: signal is true;
	signal G8740: std_logic; attribute dont_touch of G8740: signal is true;
	signal G8741: std_logic; attribute dont_touch of G8741: signal is true;
	signal G8742: std_logic; attribute dont_touch of G8742: signal is true;
	signal G8743: std_logic; attribute dont_touch of G8743: signal is true;
	signal G8744: std_logic; attribute dont_touch of G8744: signal is true;
	signal G8745: std_logic; attribute dont_touch of G8745: signal is true;
	signal G8748: std_logic; attribute dont_touch of G8748: signal is true;
	signal G8751: std_logic; attribute dont_touch of G8751: signal is true;
	signal G8756: std_logic; attribute dont_touch of G8756: signal is true;
	signal G8757: std_logic; attribute dont_touch of G8757: signal is true;
	signal G8763: std_logic; attribute dont_touch of G8763: signal is true;
	signal G8764: std_logic; attribute dont_touch of G8764: signal is true;
	signal G8765: std_logic; attribute dont_touch of G8765: signal is true;
	signal G8766: std_logic; attribute dont_touch of G8766: signal is true;
	signal G8769: std_logic; attribute dont_touch of G8769: signal is true;
	signal G8770: std_logic; attribute dont_touch of G8770: signal is true;
	signal G8774: std_logic; attribute dont_touch of G8774: signal is true;
	signal G8778: std_logic; attribute dont_touch of G8778: signal is true;
	signal G8790: std_logic; attribute dont_touch of G8790: signal is true;
	signal G8791: std_logic; attribute dont_touch of G8791: signal is true;
	signal G8792: std_logic; attribute dont_touch of G8792: signal is true;
	signal G8795: std_logic; attribute dont_touch of G8795: signal is true;
	signal G8796: std_logic; attribute dont_touch of G8796: signal is true;
	signal G8803: std_logic; attribute dont_touch of G8803: signal is true;
	signal G8804: std_logic; attribute dont_touch of G8804: signal is true;
	signal G8805: std_logic; attribute dont_touch of G8805: signal is true;
	signal G8806: std_logic; attribute dont_touch of G8806: signal is true;
	signal G8807: std_logic; attribute dont_touch of G8807: signal is true;
	signal G8808: std_logic; attribute dont_touch of G8808: signal is true;
	signal G8812: std_logic; attribute dont_touch of G8812: signal is true;
	signal G8818: std_logic; attribute dont_touch of G8818: signal is true;
	signal G8821: std_logic; attribute dont_touch of G8821: signal is true;
	signal G8822: std_logic; attribute dont_touch of G8822: signal is true;
	signal G8829: std_logic; attribute dont_touch of G8829: signal is true;
	signal G8830: std_logic; attribute dont_touch of G8830: signal is true;
	signal G8833: std_logic; attribute dont_touch of G8833: signal is true;
	signal G8836: std_logic; attribute dont_touch of G8836: signal is true;
	signal G8840: std_logic; attribute dont_touch of G8840: signal is true;
	signal G8841: std_logic; attribute dont_touch of G8841: signal is true;
	signal G8844: std_logic; attribute dont_touch of G8844: signal is true;
	signal G8847: std_logic; attribute dont_touch of G8847: signal is true;
	signal G8848: std_logic; attribute dont_touch of G8848: signal is true;
	signal G8851: std_logic; attribute dont_touch of G8851: signal is true;
	signal G8854: std_logic; attribute dont_touch of G8854: signal is true;
	signal G8858: std_logic; attribute dont_touch of G8858: signal is true;
	signal G8859: std_logic; attribute dont_touch of G8859: signal is true;
	signal G8863: std_logic; attribute dont_touch of G8863: signal is true;
	signal G8864: std_logic; attribute dont_touch of G8864: signal is true;
	signal G8871: std_logic; attribute dont_touch of G8871: signal is true;
	signal G8872: std_logic; attribute dont_touch of G8872: signal is true;
	signal G8873: std_logic; attribute dont_touch of G8873: signal is true;
	signal G8876: std_logic; attribute dont_touch of G8876: signal is true;
	signal G8879: std_logic; attribute dont_touch of G8879: signal is true;
	signal G8880: std_logic; attribute dont_touch of G8880: signal is true;
	signal G8883: std_logic; attribute dont_touch of G8883: signal is true;
	signal G8889: std_logic; attribute dont_touch of G8889: signal is true;
	signal G8890: std_logic; attribute dont_touch of G8890: signal is true;
	signal G8891: std_logic; attribute dont_touch of G8891: signal is true;
	signal G8895: std_logic; attribute dont_touch of G8895: signal is true;
	signal G8898: std_logic; attribute dont_touch of G8898: signal is true;
	signal G8899: std_logic; attribute dont_touch of G8899: signal is true;
	signal G8903: std_logic; attribute dont_touch of G8903: signal is true;
	signal G8904: std_logic; attribute dont_touch of G8904: signal is true;
	signal G8905: std_logic; attribute dont_touch of G8905: signal is true;
	signal G8906: std_logic; attribute dont_touch of G8906: signal is true;
	signal G8912: std_logic; attribute dont_touch of G8912: signal is true;
	signal G8913: std_logic; attribute dont_touch of G8913: signal is true;
	signal G8914: std_logic; attribute dont_touch of G8914: signal is true;
	signal G8921: std_logic; attribute dont_touch of G8921: signal is true;
	signal G8922: std_logic; attribute dont_touch of G8922: signal is true;
	signal G8925: std_logic; attribute dont_touch of G8925: signal is true;
	signal G8928: std_logic; attribute dont_touch of G8928: signal is true;
	signal G8933: std_logic; attribute dont_touch of G8933: signal is true;
	signal G8938: std_logic; attribute dont_touch of G8938: signal is true;
	signal G8944: std_logic; attribute dont_touch of G8944: signal is true;
	signal G8945: std_logic; attribute dont_touch of G8945: signal is true;
	signal G8948: std_logic; attribute dont_touch of G8948: signal is true;
	signal G8951: std_logic; attribute dont_touch of G8951: signal is true;
	signal G8954: std_logic; attribute dont_touch of G8954: signal is true;
	signal G8955: std_logic; attribute dont_touch of G8955: signal is true;
	signal G8956: std_logic; attribute dont_touch of G8956: signal is true;
	signal G8957: std_logic; attribute dont_touch of G8957: signal is true;
	signal G8958: std_logic; attribute dont_touch of G8958: signal is true;
	signal G8964: std_logic; attribute dont_touch of G8964: signal is true;
	signal G8967: std_logic; attribute dont_touch of G8967: signal is true;
	signal G8971: std_logic; attribute dont_touch of G8971: signal is true;
	signal G8974: std_logic; attribute dont_touch of G8974: signal is true;
	signal G8977: std_logic; attribute dont_touch of G8977: signal is true;
	signal G8984: std_logic; attribute dont_touch of G8984: signal is true;
	signal G8989: std_logic; attribute dont_touch of G8989: signal is true;
	signal G8990: std_logic; attribute dont_touch of G8990: signal is true;
	signal G8993: std_logic; attribute dont_touch of G8993: signal is true;
	signal G8997: std_logic; attribute dont_touch of G8997: signal is true;
	signal G9000: std_logic; attribute dont_touch of G9000: signal is true;
	signal G9003: std_logic; attribute dont_touch of G9003: signal is true;
	signal G9007: std_logic; attribute dont_touch of G9007: signal is true;
	signal G9011: std_logic; attribute dont_touch of G9011: signal is true;
	signal G9012: std_logic; attribute dont_touch of G9012: signal is true;
	signal G9013: std_logic; attribute dont_touch of G9013: signal is true;
	signal G9014: std_logic; attribute dont_touch of G9014: signal is true;
	signal G9015: std_logic; attribute dont_touch of G9015: signal is true;
	signal G9018: std_logic; attribute dont_touch of G9018: signal is true;
	signal G9020: std_logic; attribute dont_touch of G9020: signal is true;
	signal G9021: std_logic; attribute dont_touch of G9021: signal is true;
	signal G9024: std_logic; attribute dont_touch of G9024: signal is true;
	signal G9030: std_logic; attribute dont_touch of G9030: signal is true;
	signal G9036: std_logic; attribute dont_touch of G9036: signal is true;
	signal G9037: std_logic; attribute dont_touch of G9037: signal is true;
	signal G9040: std_logic; attribute dont_touch of G9040: signal is true;
	signal G9044: std_logic; attribute dont_touch of G9044: signal is true;
	signal G9049: std_logic; attribute dont_touch of G9049: signal is true;
	signal G9050: std_logic; attribute dont_touch of G9050: signal is true;
	signal G9051: std_logic; attribute dont_touch of G9051: signal is true;
	signal G9055: std_logic; attribute dont_touch of G9055: signal is true;
	signal G9056: std_logic; attribute dont_touch of G9056: signal is true;
	signal G9060: std_logic; attribute dont_touch of G9060: signal is true;
	signal G9061: std_logic; attribute dont_touch of G9061: signal is true;
	signal G9064: std_logic; attribute dont_touch of G9064: signal is true;
	signal G9070: std_logic; attribute dont_touch of G9070: signal is true;
	signal G9071: std_logic; attribute dont_touch of G9071: signal is true;
	signal G9072: std_logic; attribute dont_touch of G9072: signal is true;
	signal G9073: std_logic; attribute dont_touch of G9073: signal is true;
	signal G9077: std_logic; attribute dont_touch of G9077: signal is true;
	signal G9083: std_logic; attribute dont_touch of G9083: signal is true;
	signal G9086: std_logic; attribute dont_touch of G9086: signal is true;
	signal G9091: std_logic; attribute dont_touch of G9091: signal is true;
	signal G9092: std_logic; attribute dont_touch of G9092: signal is true;
	signal G9095: std_logic; attribute dont_touch of G9095: signal is true;
	signal G9099: std_logic; attribute dont_touch of G9099: signal is true;
	signal G9100: std_logic; attribute dont_touch of G9100: signal is true;
	signal G9103: std_logic; attribute dont_touch of G9103: signal is true;
	signal G9104: std_logic; attribute dont_touch of G9104: signal is true;
	signal G9152: std_logic; attribute dont_touch of G9152: signal is true;
	signal G9153: std_logic; attribute dont_touch of G9153: signal is true;
	signal G9154: std_logic; attribute dont_touch of G9154: signal is true;
	signal G9155: std_logic; attribute dont_touch of G9155: signal is true;
	signal G9158: std_logic; attribute dont_touch of G9158: signal is true;
	signal G9162: std_logic; attribute dont_touch of G9162: signal is true;
	signal G9166: std_logic; attribute dont_touch of G9166: signal is true;
	signal G9174: std_logic; attribute dont_touch of G9174: signal is true;
	signal G9177: std_logic; attribute dont_touch of G9177: signal is true;
	signal G9180: std_logic; attribute dont_touch of G9180: signal is true;
	signal G9184: std_logic; attribute dont_touch of G9184: signal is true;
	signal G9185: std_logic; attribute dont_touch of G9185: signal is true;
	signal G9186: std_logic; attribute dont_touch of G9186: signal is true;
	signal G9187: std_logic; attribute dont_touch of G9187: signal is true;
	signal G9194: std_logic; attribute dont_touch of G9194: signal is true;
	signal G9197: std_logic; attribute dont_touch of G9197: signal is true;
	signal G9200: std_logic; attribute dont_touch of G9200: signal is true;
	signal G9203: std_logic; attribute dont_touch of G9203: signal is true;
	signal G9206: std_logic; attribute dont_touch of G9206: signal is true;
	signal G9212: std_logic; attribute dont_touch of G9212: signal is true;
	signal G9213: std_logic; attribute dont_touch of G9213: signal is true;
	signal G9214: std_logic; attribute dont_touch of G9214: signal is true;
	signal G9217: std_logic; attribute dont_touch of G9217: signal is true;
	signal G9220: std_logic; attribute dont_touch of G9220: signal is true;
	signal G9223: std_logic; attribute dont_touch of G9223: signal is true;
	signal G9226: std_logic; attribute dont_touch of G9226: signal is true;
	signal G9229: std_logic; attribute dont_touch of G9229: signal is true;
	signal G9234: std_logic; attribute dont_touch of G9234: signal is true;
	signal G9239: std_logic; attribute dont_touch of G9239: signal is true;
	signal G9245: std_logic; attribute dont_touch of G9245: signal is true;
	signal G9246: std_logic; attribute dont_touch of G9246: signal is true;
	signal G9247: std_logic; attribute dont_touch of G9247: signal is true;
	signal G9250: std_logic; attribute dont_touch of G9250: signal is true;
	signal G9252: std_logic; attribute dont_touch of G9252: signal is true;
	signal G9253: std_logic; attribute dont_touch of G9253: signal is true;
	signal G9257: std_logic; attribute dont_touch of G9257: signal is true;
	signal G9258: std_logic; attribute dont_touch of G9258: signal is true;
	signal G9259: std_logic; attribute dont_touch of G9259: signal is true;
	signal G9264: std_logic; attribute dont_touch of G9264: signal is true;
	signal G9269: std_logic; attribute dont_touch of G9269: signal is true;
	signal G9274: std_logic; attribute dont_touch of G9274: signal is true;
	signal G9280: std_logic; attribute dont_touch of G9280: signal is true;
	signal G9281: std_logic; attribute dont_touch of G9281: signal is true;
	signal G9282: std_logic; attribute dont_touch of G9282: signal is true;
	signal G9283: std_logic; attribute dont_touch of G9283: signal is true;
	signal G9284: std_logic; attribute dont_touch of G9284: signal is true;
	signal G9285: std_logic; attribute dont_touch of G9285: signal is true;
	signal G9291: std_logic; attribute dont_touch of G9291: signal is true;
	signal G9295: std_logic; attribute dont_touch of G9295: signal is true;
	signal G9298: std_logic; attribute dont_touch of G9298: signal is true;
	signal G9299: std_logic; attribute dont_touch of G9299: signal is true;
	signal G9300: std_logic; attribute dont_touch of G9300: signal is true;
	signal G9305: std_logic; attribute dont_touch of G9305: signal is true;
	signal G9309: std_logic; attribute dont_touch of G9309: signal is true;
	signal G9310: std_logic; attribute dont_touch of G9310: signal is true;
	signal G9311: std_logic; attribute dont_touch of G9311: signal is true;
	signal G9316: std_logic; attribute dont_touch of G9316: signal is true;
	signal G9321: std_logic; attribute dont_touch of G9321: signal is true;
	signal G9326: std_logic; attribute dont_touch of G9326: signal is true;
	signal G9332: std_logic; attribute dont_touch of G9332: signal is true;
	signal G9333: std_logic; attribute dont_touch of G9333: signal is true;
	signal G9334: std_logic; attribute dont_touch of G9334: signal is true;
	signal G9337: std_logic; attribute dont_touch of G9337: signal is true;
	signal G9338: std_logic; attribute dont_touch of G9338: signal is true;
	signal G9339: std_logic; attribute dont_touch of G9339: signal is true;
	signal G9340: std_logic; attribute dont_touch of G9340: signal is true;
	signal G9354: std_logic; attribute dont_touch of G9354: signal is true;
	signal G9360: std_logic; attribute dont_touch of G9360: signal is true;
	signal G9364: std_logic; attribute dont_touch of G9364: signal is true;
	signal G9369: std_logic; attribute dont_touch of G9369: signal is true;
	signal G9372: std_logic; attribute dont_touch of G9372: signal is true;
	signal G9373: std_logic; attribute dont_touch of G9373: signal is true;
	signal G9374: std_logic; attribute dont_touch of G9374: signal is true;
	signal G9379: std_logic; attribute dont_touch of G9379: signal is true;
	signal G9380: std_logic; attribute dont_touch of G9380: signal is true;
	signal G9381: std_logic; attribute dont_touch of G9381: signal is true;
	signal G9386: std_logic; attribute dont_touch of G9386: signal is true;
	signal G9390: std_logic; attribute dont_touch of G9390: signal is true;
	signal G9391: std_logic; attribute dont_touch of G9391: signal is true;
	signal G9392: std_logic; attribute dont_touch of G9392: signal is true;
	signal G9397: std_logic; attribute dont_touch of G9397: signal is true;
	signal G9402: std_logic; attribute dont_touch of G9402: signal is true;
	signal G9407: std_logic; attribute dont_touch of G9407: signal is true;
	signal G9413: std_logic; attribute dont_touch of G9413: signal is true;
	signal G9414: std_logic; attribute dont_touch of G9414: signal is true;
	signal G9415: std_logic; attribute dont_touch of G9415: signal is true;
	signal G9416: std_logic; attribute dont_touch of G9416: signal is true;
	signal G9417: std_logic; attribute dont_touch of G9417: signal is true;
	signal G9429: std_logic; attribute dont_touch of G9429: signal is true;
	signal G9433: std_logic; attribute dont_touch of G9433: signal is true;
	signal G9434: std_logic; attribute dont_touch of G9434: signal is true;
	signal G9439: std_logic; attribute dont_touch of G9439: signal is true;
	signal G9442: std_logic; attribute dont_touch of G9442: signal is true;
	signal G9443: std_logic; attribute dont_touch of G9443: signal is true;
	signal G9444: std_logic; attribute dont_touch of G9444: signal is true;
	signal G9449: std_logic; attribute dont_touch of G9449: signal is true;
	signal G9450: std_logic; attribute dont_touch of G9450: signal is true;
	signal G9451: std_logic; attribute dont_touch of G9451: signal is true;
	signal G9456: std_logic; attribute dont_touch of G9456: signal is true;
	signal G9460: std_logic; attribute dont_touch of G9460: signal is true;
	signal G9461: std_logic; attribute dont_touch of G9461: signal is true;
	signal G9462: std_logic; attribute dont_touch of G9462: signal is true;
	signal G9467: std_logic; attribute dont_touch of G9467: signal is true;
	signal G9472: std_logic; attribute dont_touch of G9472: signal is true;
	signal G9477: std_logic; attribute dont_touch of G9477: signal is true;
	signal G9478: std_logic; attribute dont_touch of G9478: signal is true;
	signal G9479: std_logic; attribute dont_touch of G9479: signal is true;
	signal G9480: std_logic; attribute dont_touch of G9480: signal is true;
	signal G9483: std_logic; attribute dont_touch of G9483: signal is true;
	signal G9484: std_logic; attribute dont_touch of G9484: signal is true;
	signal G9485: std_logic; attribute dont_touch of G9485: signal is true;
	signal G9488: std_logic; attribute dont_touch of G9488: signal is true;
	signal G9489: std_logic; attribute dont_touch of G9489: signal is true;
	signal G9490: std_logic; attribute dont_touch of G9490: signal is true;
	signal G9491: std_logic; attribute dont_touch of G9491: signal is true;
	signal G9492: std_logic; attribute dont_touch of G9492: signal is true;
	signal G9496: std_logic; attribute dont_touch of G9496: signal is true;
	signal G9498: std_logic; attribute dont_touch of G9498: signal is true;
	signal G9499: std_logic; attribute dont_touch of G9499: signal is true;
	signal G9500: std_logic; attribute dont_touch of G9500: signal is true;
	signal G9501: std_logic; attribute dont_touch of G9501: signal is true;
	signal G9506: std_logic; attribute dont_touch of G9506: signal is true;
	signal G9509: std_logic; attribute dont_touch of G9509: signal is true;
	signal G9510: std_logic; attribute dont_touch of G9510: signal is true;
	signal G9511: std_logic; attribute dont_touch of G9511: signal is true;
	signal G9516: std_logic; attribute dont_touch of G9516: signal is true;
	signal G9517: std_logic; attribute dont_touch of G9517: signal is true;
	signal G9518: std_logic; attribute dont_touch of G9518: signal is true;
	signal G9523: std_logic; attribute dont_touch of G9523: signal is true;
	signal G9527: std_logic; attribute dont_touch of G9527: signal is true;
	signal G9528: std_logic; attribute dont_touch of G9528: signal is true;
	signal G9529: std_logic; attribute dont_touch of G9529: signal is true;
	signal G9534: std_logic; attribute dont_touch of G9534: signal is true;
	signal G9535: std_logic; attribute dont_touch of G9535: signal is true;
	signal G9536: std_logic; attribute dont_touch of G9536: signal is true;
	signal G9537: std_logic; attribute dont_touch of G9537: signal is true;
	signal G9538: std_logic; attribute dont_touch of G9538: signal is true;
	signal G9541: std_logic; attribute dont_touch of G9541: signal is true;
	signal G9542: std_logic; attribute dont_touch of G9542: signal is true;
	signal G9543: std_logic; attribute dont_touch of G9543: signal is true;
	signal G9546: std_logic; attribute dont_touch of G9546: signal is true;
	signal G9547: std_logic; attribute dont_touch of G9547: signal is true;
	signal G9551: std_logic; attribute dont_touch of G9551: signal is true;
	signal G9552: std_logic; attribute dont_touch of G9552: signal is true;
	signal G9554: std_logic; attribute dont_touch of G9554: signal is true;
	signal G9556: std_logic; attribute dont_touch of G9556: signal is true;
	signal G9557: std_logic; attribute dont_touch of G9557: signal is true;
	signal G9558: std_logic; attribute dont_touch of G9558: signal is true;
	signal G9559: std_logic; attribute dont_touch of G9559: signal is true;
	signal G9564: std_logic; attribute dont_touch of G9564: signal is true;
	signal G9567: std_logic; attribute dont_touch of G9567: signal is true;
	signal G9568: std_logic; attribute dont_touch of G9568: signal is true;
	signal G9569: std_logic; attribute dont_touch of G9569: signal is true;
	signal G9574: std_logic; attribute dont_touch of G9574: signal is true;
	signal G9575: std_logic; attribute dont_touch of G9575: signal is true;
	signal G9576: std_logic; attribute dont_touch of G9576: signal is true;
	signal G9581: std_logic; attribute dont_touch of G9581: signal is true;
	signal G9582: std_logic; attribute dont_touch of G9582: signal is true;
	signal G9585: std_logic; attribute dont_touch of G9585: signal is true;
	signal G9586: std_logic; attribute dont_touch of G9586: signal is true;
	signal G9590: std_logic; attribute dont_touch of G9590: signal is true;
	signal G9591: std_logic; attribute dont_touch of G9591: signal is true;
	signal G9594: std_logic; attribute dont_touch of G9594: signal is true;
	signal G9595: std_logic; attribute dont_touch of G9595: signal is true;
	signal G9598: std_logic; attribute dont_touch of G9598: signal is true;
	signal G9599: std_logic; attribute dont_touch of G9599: signal is true;
	signal G9600: std_logic; attribute dont_touch of G9600: signal is true;
	signal G9601: std_logic; attribute dont_touch of G9601: signal is true;
	signal G9602: std_logic; attribute dont_touch of G9602: signal is true;
	signal G9607: std_logic; attribute dont_touch of G9607: signal is true;
	signal G9613: std_logic; attribute dont_touch of G9613: signal is true;
	signal G9614: std_logic; attribute dont_touch of G9614: signal is true;
	signal G9616: std_logic; attribute dont_touch of G9616: signal is true;
	signal G9618: std_logic; attribute dont_touch of G9618: signal is true;
	signal G9619: std_logic; attribute dont_touch of G9619: signal is true;
	signal G9620: std_logic; attribute dont_touch of G9620: signal is true;
	signal G9621: std_logic; attribute dont_touch of G9621: signal is true;
	signal G9626: std_logic; attribute dont_touch of G9626: signal is true;
	signal G9629: std_logic; attribute dont_touch of G9629: signal is true;
	signal G9630: std_logic; attribute dont_touch of G9630: signal is true;
	signal G9631: std_logic; attribute dont_touch of G9631: signal is true;
	signal G9636: std_logic; attribute dont_touch of G9636: signal is true;
	signal G9637: std_logic; attribute dont_touch of G9637: signal is true;
	signal G9638: std_logic; attribute dont_touch of G9638: signal is true;
	signal G9639: std_logic; attribute dont_touch of G9639: signal is true;
	signal G9640: std_logic; attribute dont_touch of G9640: signal is true;
	signal G9644: std_logic; attribute dont_touch of G9644: signal is true;
	signal G9645: std_logic; attribute dont_touch of G9645: signal is true;
	signal G9648: std_logic; attribute dont_touch of G9648: signal is true;
	signal G9649: std_logic; attribute dont_touch of G9649: signal is true;
	signal G9653: std_logic; attribute dont_touch of G9653: signal is true;
	signal G9654: std_logic; attribute dont_touch of G9654: signal is true;
	signal G9657: std_logic; attribute dont_touch of G9657: signal is true;
	signal G9660: std_logic; attribute dont_touch of G9660: signal is true;
	signal G9661: std_logic; attribute dont_touch of G9661: signal is true;
	signal G9662: std_logic; attribute dont_touch of G9662: signal is true;
	signal G9663: std_logic; attribute dont_touch of G9663: signal is true;
	signal G9664: std_logic; attribute dont_touch of G9664: signal is true;
	signal G9669: std_logic; attribute dont_touch of G9669: signal is true;
	signal G9670: std_logic; attribute dont_touch of G9670: signal is true;
	signal G9671: std_logic; attribute dont_touch of G9671: signal is true;
	signal G9672: std_logic; attribute dont_touch of G9672: signal is true;
	signal G9678: std_logic; attribute dont_touch of G9678: signal is true;
	signal G9679: std_logic; attribute dont_touch of G9679: signal is true;
	signal G9681: std_logic; attribute dont_touch of G9681: signal is true;
	signal G9683: std_logic; attribute dont_touch of G9683: signal is true;
	signal G9684: std_logic; attribute dont_touch of G9684: signal is true;
	signal G9685: std_logic; attribute dont_touch of G9685: signal is true;
	signal G9686: std_logic; attribute dont_touch of G9686: signal is true;
	signal G9687: std_logic; attribute dont_touch of G9687: signal is true;
	signal G9688: std_logic; attribute dont_touch of G9688: signal is true;
	signal G9689: std_logic; attribute dont_touch of G9689: signal is true;
	signal G9690: std_logic; attribute dont_touch of G9690: signal is true;
	signal G9691: std_logic; attribute dont_touch of G9691: signal is true;
	signal G9692: std_logic; attribute dont_touch of G9692: signal is true;
	signal G9693: std_logic; attribute dont_touch of G9693: signal is true;
	signal G9694: std_logic; attribute dont_touch of G9694: signal is true;
	signal G9698: std_logic; attribute dont_touch of G9698: signal is true;
	signal G9699: std_logic; attribute dont_touch of G9699: signal is true;
	signal G9700: std_logic; attribute dont_touch of G9700: signal is true;
	signal G9704: std_logic; attribute dont_touch of G9704: signal is true;
	signal G9705: std_logic; attribute dont_touch of G9705: signal is true;
	signal G9708: std_logic; attribute dont_touch of G9708: signal is true;
	signal G9713: std_logic; attribute dont_touch of G9713: signal is true;
	signal G9714: std_logic; attribute dont_touch of G9714: signal is true;
	signal G9715: std_logic; attribute dont_touch of G9715: signal is true;
	signal G9716: std_logic; attribute dont_touch of G9716: signal is true;
	signal G9721: std_logic; attribute dont_touch of G9721: signal is true;
	signal G9724: std_logic; attribute dont_touch of G9724: signal is true;
	signal G9728: std_logic; attribute dont_touch of G9728: signal is true;
	signal G9729: std_logic; attribute dont_touch of G9729: signal is true;
	signal G9730: std_logic; attribute dont_touch of G9730: signal is true;
	signal G9731: std_logic; attribute dont_touch of G9731: signal is true;
	signal G9732: std_logic; attribute dont_touch of G9732: signal is true;
	signal G9733: std_logic; attribute dont_touch of G9733: signal is true;
	signal G9739: std_logic; attribute dont_touch of G9739: signal is true;
	signal G9740: std_logic; attribute dont_touch of G9740: signal is true;
	signal G9742: std_logic; attribute dont_touch of G9742: signal is true;
	signal G9744: std_logic; attribute dont_touch of G9744: signal is true;
	signal G9745: std_logic; attribute dont_touch of G9745: signal is true;
	signal G9746: std_logic; attribute dont_touch of G9746: signal is true;
	signal G9747: std_logic; attribute dont_touch of G9747: signal is true;
	signal G9748: std_logic; attribute dont_touch of G9748: signal is true;
	signal G9749: std_logic; attribute dont_touch of G9749: signal is true;
	signal G9750: std_logic; attribute dont_touch of G9750: signal is true;
	signal G9751: std_logic; attribute dont_touch of G9751: signal is true;
	signal G9752: std_logic; attribute dont_touch of G9752: signal is true;
	signal G9753: std_logic; attribute dont_touch of G9753: signal is true;
	signal G9754: std_logic; attribute dont_touch of G9754: signal is true;
	signal G9755: std_logic; attribute dont_touch of G9755: signal is true;
	signal G9759: std_logic; attribute dont_touch of G9759: signal is true;
	signal G9760: std_logic; attribute dont_touch of G9760: signal is true;
	signal G9761: std_logic; attribute dont_touch of G9761: signal is true;
	signal G9762: std_logic; attribute dont_touch of G9762: signal is true;
	signal G9766: std_logic; attribute dont_touch of G9766: signal is true;
	signal G9771: std_logic; attribute dont_touch of G9771: signal is true;
	signal G9772: std_logic; attribute dont_touch of G9772: signal is true;
	signal G9775: std_logic; attribute dont_touch of G9775: signal is true;
	signal G9776: std_logic; attribute dont_touch of G9776: signal is true;
	signal G9777: std_logic; attribute dont_touch of G9777: signal is true;
	signal G9778: std_logic; attribute dont_touch of G9778: signal is true;
	signal G9779: std_logic; attribute dont_touch of G9779: signal is true;
	signal G9780: std_logic; attribute dont_touch of G9780: signal is true;
	signal G9792: std_logic; attribute dont_touch of G9792: signal is true;
	signal G9797: std_logic; attribute dont_touch of G9797: signal is true;
	signal G9800: std_logic; attribute dont_touch of G9800: signal is true;
	signal G9804: std_logic; attribute dont_touch of G9804: signal is true;
	signal G9805: std_logic; attribute dont_touch of G9805: signal is true;
	signal G9806: std_logic; attribute dont_touch of G9806: signal is true;
	signal G9807: std_logic; attribute dont_touch of G9807: signal is true;
	signal G9808: std_logic; attribute dont_touch of G9808: signal is true;
	signal G9809: std_logic; attribute dont_touch of G9809: signal is true;
	signal G9815: std_logic; attribute dont_touch of G9815: signal is true;
	signal G9816: std_logic; attribute dont_touch of G9816: signal is true;
	signal G9818: std_logic; attribute dont_touch of G9818: signal is true;
	signal G9819: std_logic; attribute dont_touch of G9819: signal is true;
	signal G9820: std_logic; attribute dont_touch of G9820: signal is true;
	signal G9821: std_logic; attribute dont_touch of G9821: signal is true;
	signal G9822: std_logic; attribute dont_touch of G9822: signal is true;
	signal G9823: std_logic; attribute dont_touch of G9823: signal is true;
	signal G9824: std_logic; attribute dont_touch of G9824: signal is true;
	signal G9825: std_logic; attribute dont_touch of G9825: signal is true;
	signal G9826: std_logic; attribute dont_touch of G9826: signal is true;
	signal G9827: std_logic; attribute dont_touch of G9827: signal is true;
	signal G9828: std_logic; attribute dont_touch of G9828: signal is true;
	signal G9829: std_logic; attribute dont_touch of G9829: signal is true;
	signal G9830: std_logic; attribute dont_touch of G9830: signal is true;
	signal G9831: std_logic; attribute dont_touch of G9831: signal is true;
	signal G9832: std_logic; attribute dont_touch of G9832: signal is true;
	signal G9833: std_logic; attribute dont_touch of G9833: signal is true;
	signal G9834: std_logic; attribute dont_touch of G9834: signal is true;
	signal G9835: std_logic; attribute dont_touch of G9835: signal is true;
	signal G9839: std_logic; attribute dont_touch of G9839: signal is true;
	signal G9842: std_logic; attribute dont_touch of G9842: signal is true;
	signal G9843: std_logic; attribute dont_touch of G9843: signal is true;
	signal G9848: std_logic; attribute dont_touch of G9848: signal is true;
	signal G9852: std_logic; attribute dont_touch of G9852: signal is true;
	signal G9853: std_logic; attribute dont_touch of G9853: signal is true;
	signal G9856: std_logic; attribute dont_touch of G9856: signal is true;
	signal G9860: std_logic; attribute dont_touch of G9860: signal is true;
	signal G9861: std_logic; attribute dont_touch of G9861: signal is true;
	signal G9862: std_logic; attribute dont_touch of G9862: signal is true;
	signal G9863: std_logic; attribute dont_touch of G9863: signal is true;
	signal G9864: std_logic; attribute dont_touch of G9864: signal is true;
	signal G9875: std_logic; attribute dont_touch of G9875: signal is true;
	signal G9880: std_logic; attribute dont_touch of G9880: signal is true;
	signal G9883: std_logic; attribute dont_touch of G9883: signal is true;
	signal G9887: std_logic; attribute dont_touch of G9887: signal is true;
	signal G9888: std_logic; attribute dont_touch of G9888: signal is true;
	signal G9889: std_logic; attribute dont_touch of G9889: signal is true;
	signal G9890: std_logic; attribute dont_touch of G9890: signal is true;
	signal G9891: std_logic; attribute dont_touch of G9891: signal is true;
	signal G9892: std_logic; attribute dont_touch of G9892: signal is true;
	signal G9898: std_logic; attribute dont_touch of G9898: signal is true;
	signal G9899: std_logic; attribute dont_touch of G9899: signal is true;
	signal G9900: std_logic; attribute dont_touch of G9900: signal is true;
	signal G9901: std_logic; attribute dont_touch of G9901: signal is true;
	signal G9902: std_logic; attribute dont_touch of G9902: signal is true;
	signal G9903: std_logic; attribute dont_touch of G9903: signal is true;
	signal G9904: std_logic; attribute dont_touch of G9904: signal is true;
	signal G9905: std_logic; attribute dont_touch of G9905: signal is true;
	signal G9906: std_logic; attribute dont_touch of G9906: signal is true;
	signal G9907: std_logic; attribute dont_touch of G9907: signal is true;
	signal G9908: std_logic; attribute dont_touch of G9908: signal is true;
	signal G9909: std_logic; attribute dont_touch of G9909: signal is true;
	signal G9910: std_logic; attribute dont_touch of G9910: signal is true;
	signal G9911: std_logic; attribute dont_touch of G9911: signal is true;
	signal G9912: std_logic; attribute dont_touch of G9912: signal is true;
	signal G9913: std_logic; attribute dont_touch of G9913: signal is true;
	signal G9914: std_logic; attribute dont_touch of G9914: signal is true;
	signal G9915: std_logic; attribute dont_touch of G9915: signal is true;
	signal G9916: std_logic; attribute dont_touch of G9916: signal is true;
	signal G9917: std_logic; attribute dont_touch of G9917: signal is true;
	signal G9920: std_logic; attribute dont_touch of G9920: signal is true;
	signal G9924: std_logic; attribute dont_touch of G9924: signal is true;
	signal G9927: std_logic; attribute dont_touch of G9927: signal is true;
	signal G9931: std_logic; attribute dont_touch of G9931: signal is true;
	signal G9932: std_logic; attribute dont_touch of G9932: signal is true;
	signal G9933: std_logic; attribute dont_touch of G9933: signal is true;
	signal G9934: std_logic; attribute dont_touch of G9934: signal is true;
	signal G9935: std_logic; attribute dont_touch of G9935: signal is true;
	signal G9946: std_logic; attribute dont_touch of G9946: signal is true;
	signal G9951: std_logic; attribute dont_touch of G9951: signal is true;
	signal G9954: std_logic; attribute dont_touch of G9954: signal is true;
	signal G9958: std_logic; attribute dont_touch of G9958: signal is true;
	signal G9959: std_logic; attribute dont_touch of G9959: signal is true;
	signal G9960: std_logic; attribute dont_touch of G9960: signal is true;
	signal G9961: std_logic; attribute dont_touch of G9961: signal is true;
	signal G9962: std_logic; attribute dont_touch of G9962: signal is true;
	signal G9963: std_logic; attribute dont_touch of G9963: signal is true;
	signal G9964: std_logic; attribute dont_touch of G9964: signal is true;
	signal G9965: std_logic; attribute dont_touch of G9965: signal is true;
	signal G9966: std_logic; attribute dont_touch of G9966: signal is true;
	signal G9967: std_logic; attribute dont_touch of G9967: signal is true;
	signal G9968: std_logic; attribute dont_touch of G9968: signal is true;
	signal G9969: std_logic; attribute dont_touch of G9969: signal is true;
	signal G9970: std_logic; attribute dont_touch of G9970: signal is true;
	signal G9971: std_logic; attribute dont_touch of G9971: signal is true;
	signal G9972: std_logic; attribute dont_touch of G9972: signal is true;
	signal G9973: std_logic; attribute dont_touch of G9973: signal is true;
	signal G9974: std_logic; attribute dont_touch of G9974: signal is true;
	signal G9975: std_logic; attribute dont_touch of G9975: signal is true;
	signal G9976: std_logic; attribute dont_touch of G9976: signal is true;
	signal G9977: std_logic; attribute dont_touch of G9977: signal is true;
	signal G9978: std_logic; attribute dont_touch of G9978: signal is true;
	signal G9982: std_logic; attribute dont_touch of G9982: signal is true;
	signal G9983: std_logic; attribute dont_touch of G9983: signal is true;
	signal G9984: std_logic; attribute dont_touch of G9984: signal is true;
	signal G9985: std_logic; attribute dont_touch of G9985: signal is true;
	signal G9989: std_logic; attribute dont_touch of G9989: signal is true;
	signal G9992: std_logic; attribute dont_touch of G9992: signal is true;
	signal G9995: std_logic; attribute dont_touch of G9995: signal is true;
	signal G9999: std_logic; attribute dont_touch of G9999: signal is true;
	signal G10000: std_logic; attribute dont_touch of G10000: signal is true;
	signal G10001: std_logic; attribute dont_touch of G10001: signal is true;
	signal G10002: std_logic; attribute dont_touch of G10002: signal is true;
	signal G10003: std_logic; attribute dont_touch of G10003: signal is true;
	signal G10014: std_logic; attribute dont_touch of G10014: signal is true;
	signal G10019: std_logic; attribute dont_touch of G10019: signal is true;
	signal G10022: std_logic; attribute dont_touch of G10022: signal is true;
	signal G10026: std_logic; attribute dont_touch of G10026: signal is true;
	signal G10027: std_logic; attribute dont_touch of G10027: signal is true;
	signal G10028: std_logic; attribute dont_touch of G10028: signal is true;
	signal G10029: std_logic; attribute dont_touch of G10029: signal is true;
	signal G10030: std_logic; attribute dont_touch of G10030: signal is true;
	signal G10031: std_logic; attribute dont_touch of G10031: signal is true;
	signal G10032: std_logic; attribute dont_touch of G10032: signal is true;
	signal G10033: std_logic; attribute dont_touch of G10033: signal is true;
	signal G10034: std_logic; attribute dont_touch of G10034: signal is true;
	signal G10035: std_logic; attribute dont_touch of G10035: signal is true;
	signal G10036: std_logic; attribute dont_touch of G10036: signal is true;
	signal G10037: std_logic; attribute dont_touch of G10037: signal is true;
	signal G10038: std_logic; attribute dont_touch of G10038: signal is true;
	signal G10039: std_logic; attribute dont_touch of G10039: signal is true;
	signal G10040: std_logic; attribute dont_touch of G10040: signal is true;
	signal G10041: std_logic; attribute dont_touch of G10041: signal is true;
	signal G10042: std_logic; attribute dont_touch of G10042: signal is true;
	signal G10043: std_logic; attribute dont_touch of G10043: signal is true;
	signal G10044: std_logic; attribute dont_touch of G10044: signal is true;
	signal G10047: std_logic; attribute dont_touch of G10047: signal is true;
	signal G10050: std_logic; attribute dont_touch of G10050: signal is true;
	signal G10053: std_logic; attribute dont_touch of G10053: signal is true;
	signal G10057: std_logic; attribute dont_touch of G10057: signal is true;
	signal G10058: std_logic; attribute dont_touch of G10058: signal is true;
	signal G10059: std_logic; attribute dont_touch of G10059: signal is true;
	signal G10060: std_logic; attribute dont_touch of G10060: signal is true;
	signal G10061: std_logic; attribute dont_touch of G10061: signal is true;
	signal G10072: std_logic; attribute dont_touch of G10072: signal is true;
	signal G10073: std_logic; attribute dont_touch of G10073: signal is true;
	signal G10074: std_logic; attribute dont_touch of G10074: signal is true;
	signal G10077: std_logic; attribute dont_touch of G10077: signal is true;
	signal G10078: std_logic; attribute dont_touch of G10078: signal is true;
	signal G10079: std_logic; attribute dont_touch of G10079: signal is true;
	signal G10080: std_logic; attribute dont_touch of G10080: signal is true;
	signal G10081: std_logic; attribute dont_touch of G10081: signal is true;
	signal G10082: std_logic; attribute dont_touch of G10082: signal is true;
	signal G10083: std_logic; attribute dont_touch of G10083: signal is true;
	signal G10084: std_logic; attribute dont_touch of G10084: signal is true;
	signal G10085: std_logic; attribute dont_touch of G10085: signal is true;
	signal G10086: std_logic; attribute dont_touch of G10086: signal is true;
	signal G10087: std_logic; attribute dont_touch of G10087: signal is true;
	signal G10090: std_logic; attribute dont_touch of G10090: signal is true;
	signal G10093: std_logic; attribute dont_touch of G10093: signal is true;
	signal G10096: std_logic; attribute dont_touch of G10096: signal is true;
	signal G10099: std_logic; attribute dont_touch of G10099: signal is true;
	signal G10102: std_logic; attribute dont_touch of G10102: signal is true;
	signal G10106: std_logic; attribute dont_touch of G10106: signal is true;
	signal G10107: std_logic; attribute dont_touch of G10107: signal is true;
	signal G10108: std_logic; attribute dont_touch of G10108: signal is true;
	signal G10109: std_logic; attribute dont_touch of G10109: signal is true;
	signal G10110: std_logic; attribute dont_touch of G10110: signal is true;
	signal G10111: std_logic; attribute dont_touch of G10111: signal is true;
	signal G10112: std_logic; attribute dont_touch of G10112: signal is true;
	signal G10113: std_logic; attribute dont_touch of G10113: signal is true;
	signal G10114: std_logic; attribute dont_touch of G10114: signal is true;
	signal G10115: std_logic; attribute dont_touch of G10115: signal is true;
	signal G10116: std_logic; attribute dont_touch of G10116: signal is true;
	signal G10117: std_logic; attribute dont_touch of G10117: signal is true;
	signal G10118: std_logic; attribute dont_touch of G10118: signal is true;
	signal G10119: std_logic; attribute dont_touch of G10119: signal is true;
	signal G10120: std_logic; attribute dont_touch of G10120: signal is true;
	signal G10121: std_logic; attribute dont_touch of G10121: signal is true;
	signal G10123: std_logic; attribute dont_touch of G10123: signal is true;
	signal G10124: std_logic; attribute dont_touch of G10124: signal is true;
	signal G10129: std_logic; attribute dont_touch of G10129: signal is true;
	signal G10130: std_logic; attribute dont_touch of G10130: signal is true;
	signal G10133: std_logic; attribute dont_touch of G10133: signal is true;
	signal G10136: std_logic; attribute dont_touch of G10136: signal is true;
	signal G10139: std_logic; attribute dont_touch of G10139: signal is true;
	signal G10140: std_logic; attribute dont_touch of G10140: signal is true;
	signal G10141: std_logic; attribute dont_touch of G10141: signal is true;
	signal G10142: std_logic; attribute dont_touch of G10142: signal is true;
	signal G10143: std_logic; attribute dont_touch of G10143: signal is true;
	signal G10147: std_logic; attribute dont_touch of G10147: signal is true;
	signal G10150: std_logic; attribute dont_touch of G10150: signal is true;
	signal G10151: std_logic; attribute dont_touch of G10151: signal is true;
	signal G10152: std_logic; attribute dont_touch of G10152: signal is true;
	signal G10153: std_logic; attribute dont_touch of G10153: signal is true;
	signal G10154: std_logic; attribute dont_touch of G10154: signal is true;
	signal G10155: std_logic; attribute dont_touch of G10155: signal is true;
	signal G10156: std_logic; attribute dont_touch of G10156: signal is true;
	signal G10157: std_logic; attribute dont_touch of G10157: signal is true;
	signal G10158: std_logic; attribute dont_touch of G10158: signal is true;
	signal G10159: std_logic; attribute dont_touch of G10159: signal is true;
	signal G10160: std_logic; attribute dont_touch of G10160: signal is true;
	signal G10165: std_logic; attribute dont_touch of G10165: signal is true;
	signal G10166: std_logic; attribute dont_touch of G10166: signal is true;
	signal G10169: std_logic; attribute dont_touch of G10169: signal is true;
	signal G10172: std_logic; attribute dont_touch of G10172: signal is true;
	signal G10175: std_logic; attribute dont_touch of G10175: signal is true;
	signal G10176: std_logic; attribute dont_touch of G10176: signal is true;
	signal G10177: std_logic; attribute dont_touch of G10177: signal is true;
	signal G10178: std_logic; attribute dont_touch of G10178: signal is true;
	signal G10179: std_logic; attribute dont_touch of G10179: signal is true;
	signal G10180: std_logic; attribute dont_touch of G10180: signal is true;
	signal G10181: std_logic; attribute dont_touch of G10181: signal is true;
	signal G10182: std_logic; attribute dont_touch of G10182: signal is true;
	signal G10183: std_logic; attribute dont_touch of G10183: signal is true;
	signal G10184: std_logic; attribute dont_touch of G10184: signal is true;
	signal G10185: std_logic; attribute dont_touch of G10185: signal is true;
	signal G10190: std_logic; attribute dont_touch of G10190: signal is true;
	signal G10191: std_logic; attribute dont_touch of G10191: signal is true;
	signal G10194: std_logic; attribute dont_touch of G10194: signal is true;
	signal G10197: std_logic; attribute dont_touch of G10197: signal is true;
	signal G10198: std_logic; attribute dont_touch of G10198: signal is true;
	signal G10199: std_logic; attribute dont_touch of G10199: signal is true;
	signal G10200: std_logic; attribute dont_touch of G10200: signal is true;
	signal G10203: std_logic; attribute dont_touch of G10203: signal is true;
	signal G10204: std_logic; attribute dont_touch of G10204: signal is true;
	signal G10205: std_logic; attribute dont_touch of G10205: signal is true;
	signal G10206: std_logic; attribute dont_touch of G10206: signal is true;
	signal G10207: std_logic; attribute dont_touch of G10207: signal is true;
	signal G10212: std_logic; attribute dont_touch of G10212: signal is true;
	signal G10213: std_logic; attribute dont_touch of G10213: signal is true;
	signal G10216: std_logic; attribute dont_touch of G10216: signal is true;
	signal G10217: std_logic; attribute dont_touch of G10217: signal is true;
	signal G10218: std_logic; attribute dont_touch of G10218: signal is true;
	signal G10219: std_logic; attribute dont_touch of G10219: signal is true;
	signal G10222: std_logic; attribute dont_touch of G10222: signal is true;
	signal G10223: std_logic; attribute dont_touch of G10223: signal is true;
	signal G10224: std_logic; attribute dont_touch of G10224: signal is true;
	signal G10229: std_logic; attribute dont_touch of G10229: signal is true;
	signal G10230: std_logic; attribute dont_touch of G10230: signal is true;
	signal G10231: std_logic; attribute dont_touch of G10231: signal is true;
	signal G10232: std_logic; attribute dont_touch of G10232: signal is true;
	signal G10233: std_logic; attribute dont_touch of G10233: signal is true;
	signal G10261: std_logic; attribute dont_touch of G10261: signal is true;
	signal G10262: std_logic; attribute dont_touch of G10262: signal is true;
	signal G10266: std_logic; attribute dont_touch of G10266: signal is true;
	signal G10272: std_logic; attribute dont_touch of G10272: signal is true;
	signal G10273: std_logic; attribute dont_touch of G10273: signal is true;
	signal G10274: std_logic; attribute dont_touch of G10274: signal is true;
	signal G10275: std_logic; attribute dont_touch of G10275: signal is true;
	signal G10278: std_logic; attribute dont_touch of G10278: signal is true;
	signal G10281: std_logic; attribute dont_touch of G10281: signal is true;
	signal G10287: std_logic; attribute dont_touch of G10287: signal is true;
	signal G10288: std_logic; attribute dont_touch of G10288: signal is true;
	signal G10289: std_logic; attribute dont_touch of G10289: signal is true;
	signal G10290: std_logic; attribute dont_touch of G10290: signal is true;
	signal G10295: std_logic; attribute dont_touch of G10295: signal is true;
	signal G10307: std_logic; attribute dont_touch of G10307: signal is true;
	signal G10308: std_logic; attribute dont_touch of G10308: signal is true;
	signal G10311: std_logic; attribute dont_touch of G10311: signal is true;
	signal G10312: std_logic; attribute dont_touch of G10312: signal is true;
	signal G10318: std_logic; attribute dont_touch of G10318: signal is true;
	signal G10319: std_logic; attribute dont_touch of G10319: signal is true;
	signal G10320: std_logic; attribute dont_touch of G10320: signal is true;
	signal G10323: std_logic; attribute dont_touch of G10323: signal is true;
	signal G10334: std_logic; attribute dont_touch of G10334: signal is true;
	signal G10335: std_logic; attribute dont_touch of G10335: signal is true;
	signal G10336: std_logic; attribute dont_touch of G10336: signal is true;
	signal G10337: std_logic; attribute dont_touch of G10337: signal is true;
	signal G10338: std_logic; attribute dont_touch of G10338: signal is true;
	signal G10341: std_logic; attribute dont_touch of G10341: signal is true;
	signal G10347: std_logic; attribute dont_touch of G10347: signal is true;
	signal G10348: std_logic; attribute dont_touch of G10348: signal is true;
	signal G10349: std_logic; attribute dont_touch of G10349: signal is true;
	signal G10350: std_logic; attribute dont_touch of G10350: signal is true;
	signal G10351: std_logic; attribute dont_touch of G10351: signal is true;
	signal G10352: std_logic; attribute dont_touch of G10352: signal is true;
	signal G10353: std_logic; attribute dont_touch of G10353: signal is true;
	signal G10354: std_logic; attribute dont_touch of G10354: signal is true;
	signal G10355: std_logic; attribute dont_touch of G10355: signal is true;
	signal G10356: std_logic; attribute dont_touch of G10356: signal is true;
	signal G10357: std_logic; attribute dont_touch of G10357: signal is true;
	signal G10358: std_logic; attribute dont_touch of G10358: signal is true;
	signal G10359: std_logic; attribute dont_touch of G10359: signal is true;
	signal G10360: std_logic; attribute dont_touch of G10360: signal is true;
	signal G10361: std_logic; attribute dont_touch of G10361: signal is true;
	signal G10362: std_logic; attribute dont_touch of G10362: signal is true;
	signal G10363: std_logic; attribute dont_touch of G10363: signal is true;
	signal G10364: std_logic; attribute dont_touch of G10364: signal is true;
	signal G10365: std_logic; attribute dont_touch of G10365: signal is true;
	signal G10366: std_logic; attribute dont_touch of G10366: signal is true;
	signal G10367: std_logic; attribute dont_touch of G10367: signal is true;
	signal G10368: std_logic; attribute dont_touch of G10368: signal is true;
	signal G10369: std_logic; attribute dont_touch of G10369: signal is true;
	signal G10370: std_logic; attribute dont_touch of G10370: signal is true;
	signal G10371: std_logic; attribute dont_touch of G10371: signal is true;
	signal G10372: std_logic; attribute dont_touch of G10372: signal is true;
	signal G10373: std_logic; attribute dont_touch of G10373: signal is true;
	signal G10374: std_logic; attribute dont_touch of G10374: signal is true;
	signal G10375: std_logic; attribute dont_touch of G10375: signal is true;
	signal G10376: std_logic; attribute dont_touch of G10376: signal is true;
	signal G10377: std_logic; attribute dont_touch of G10377: signal is true;
	signal G10378: std_logic; attribute dont_touch of G10378: signal is true;
	signal G10379: std_logic; attribute dont_touch of G10379: signal is true;
	signal G10380: std_logic; attribute dont_touch of G10380: signal is true;
	signal G10381: std_logic; attribute dont_touch of G10381: signal is true;
	signal G10382: std_logic; attribute dont_touch of G10382: signal is true;
	signal G10383: std_logic; attribute dont_touch of G10383: signal is true;
	signal G10384: std_logic; attribute dont_touch of G10384: signal is true;
	signal G10385: std_logic; attribute dont_touch of G10385: signal is true;
	signal G10386: std_logic; attribute dont_touch of G10386: signal is true;
	signal G10387: std_logic; attribute dont_touch of G10387: signal is true;
	signal G10388: std_logic; attribute dont_touch of G10388: signal is true;
	signal G10389: std_logic; attribute dont_touch of G10389: signal is true;
	signal G10390: std_logic; attribute dont_touch of G10390: signal is true;
	signal G10391: std_logic; attribute dont_touch of G10391: signal is true;
	signal G10392: std_logic; attribute dont_touch of G10392: signal is true;
	signal G10393: std_logic; attribute dont_touch of G10393: signal is true;
	signal G10394: std_logic; attribute dont_touch of G10394: signal is true;
	signal G10395: std_logic; attribute dont_touch of G10395: signal is true;
	signal G10396: std_logic; attribute dont_touch of G10396: signal is true;
	signal G10397: std_logic; attribute dont_touch of G10397: signal is true;
	signal G10398: std_logic; attribute dont_touch of G10398: signal is true;
	signal G10399: std_logic; attribute dont_touch of G10399: signal is true;
	signal G10400: std_logic; attribute dont_touch of G10400: signal is true;
	signal G10401: std_logic; attribute dont_touch of G10401: signal is true;
	signal G10402: std_logic; attribute dont_touch of G10402: signal is true;
	signal G10403: std_logic; attribute dont_touch of G10403: signal is true;
	signal G10404: std_logic; attribute dont_touch of G10404: signal is true;
	signal G10405: std_logic; attribute dont_touch of G10405: signal is true;
	signal G10406: std_logic; attribute dont_touch of G10406: signal is true;
	signal G10407: std_logic; attribute dont_touch of G10407: signal is true;
	signal G10408: std_logic; attribute dont_touch of G10408: signal is true;
	signal G10409: std_logic; attribute dont_touch of G10409: signal is true;
	signal G10410: std_logic; attribute dont_touch of G10410: signal is true;
	signal G10411: std_logic; attribute dont_touch of G10411: signal is true;
	signal G10412: std_logic; attribute dont_touch of G10412: signal is true;
	signal G10413: std_logic; attribute dont_touch of G10413: signal is true;
	signal G10414: std_logic; attribute dont_touch of G10414: signal is true;
	signal G10415: std_logic; attribute dont_touch of G10415: signal is true;
	signal G10416: std_logic; attribute dont_touch of G10416: signal is true;
	signal G10417: std_logic; attribute dont_touch of G10417: signal is true;
	signal G10418: std_logic; attribute dont_touch of G10418: signal is true;
	signal G10419: std_logic; attribute dont_touch of G10419: signal is true;
	signal G10420: std_logic; attribute dont_touch of G10420: signal is true;
	signal G10421: std_logic; attribute dont_touch of G10421: signal is true;
	signal G10427: std_logic; attribute dont_touch of G10427: signal is true;
	signal G10428: std_logic; attribute dont_touch of G10428: signal is true;
	signal G10429: std_logic; attribute dont_touch of G10429: signal is true;
	signal G10430: std_logic; attribute dont_touch of G10430: signal is true;
	signal G10472: std_logic; attribute dont_touch of G10472: signal is true;
	signal G10473: std_logic; attribute dont_touch of G10473: signal is true;
	signal G10474: std_logic; attribute dont_touch of G10474: signal is true;
	signal G10475: std_logic; attribute dont_touch of G10475: signal is true;
	signal G10476: std_logic; attribute dont_touch of G10476: signal is true;
	signal G10487: std_logic; attribute dont_touch of G10487: signal is true;
	signal G10488: std_logic; attribute dont_touch of G10488: signal is true;
	signal G10489: std_logic; attribute dont_touch of G10489: signal is true;
	signal G10490: std_logic; attribute dont_touch of G10490: signal is true;
	signal G10491: std_logic; attribute dont_touch of G10491: signal is true;
	signal G10497: std_logic; attribute dont_touch of G10497: signal is true;
	signal G10498: std_logic; attribute dont_touch of G10498: signal is true;
	signal G10499: std_logic; attribute dont_touch of G10499: signal is true;
	signal G10501: std_logic; attribute dont_touch of G10501: signal is true;
	signal G10502: std_logic; attribute dont_touch of G10502: signal is true;
	signal G10503: std_logic; attribute dont_touch of G10503: signal is true;
	signal G10504: std_logic; attribute dont_touch of G10504: signal is true;
	signal G10509: std_logic; attribute dont_touch of G10509: signal is true;
	signal G10510: std_logic; attribute dont_touch of G10510: signal is true;
	signal G10511: std_logic; attribute dont_touch of G10511: signal is true;
	signal G10515: std_logic; attribute dont_touch of G10515: signal is true;
	signal G10518: std_logic; attribute dont_touch of G10518: signal is true;
	signal G10519: std_logic; attribute dont_touch of G10519: signal is true;
	signal G10520: std_logic; attribute dont_touch of G10520: signal is true;
	signal G10521: std_logic; attribute dont_touch of G10521: signal is true;
	signal G10528: std_logic; attribute dont_touch of G10528: signal is true;
	signal G10529: std_logic; attribute dont_touch of G10529: signal is true;
	signal G10530: std_logic; attribute dont_touch of G10530: signal is true;
	signal G10531: std_logic; attribute dont_touch of G10531: signal is true;
	signal G10532: std_logic; attribute dont_touch of G10532: signal is true;
	signal G10533: std_logic; attribute dont_touch of G10533: signal is true;
	signal G10537: std_logic; attribute dont_touch of G10537: signal is true;
	signal G10540: std_logic; attribute dont_touch of G10540: signal is true;
	signal G10541: std_logic; attribute dont_touch of G10541: signal is true;
	signal G10542: std_logic; attribute dont_touch of G10542: signal is true;
	signal G10543: std_logic; attribute dont_touch of G10543: signal is true;
	signal G10544: std_logic; attribute dont_touch of G10544: signal is true;
	signal G10550: std_logic; attribute dont_touch of G10550: signal is true;
	signal G10551: std_logic; attribute dont_touch of G10551: signal is true;
	signal G10552: std_logic; attribute dont_touch of G10552: signal is true;
	signal G10553: std_logic; attribute dont_touch of G10553: signal is true;
	signal G10554: std_logic; attribute dont_touch of G10554: signal is true;
	signal G10555: std_logic; attribute dont_touch of G10555: signal is true;
	signal G10556: std_logic; attribute dont_touch of G10556: signal is true;
	signal G10561: std_logic; attribute dont_touch of G10561: signal is true;
	signal G10564: std_logic; attribute dont_touch of G10564: signal is true;
	signal G10565: std_logic; attribute dont_touch of G10565: signal is true;
	signal G10566: std_logic; attribute dont_touch of G10566: signal is true;
	signal G10567: std_logic; attribute dont_touch of G10567: signal is true;
	signal G10568: std_logic; attribute dont_touch of G10568: signal is true;
	signal G10569: std_logic; attribute dont_touch of G10569: signal is true;
	signal G10570: std_logic; attribute dont_touch of G10570: signal is true;
	signal G10571: std_logic; attribute dont_touch of G10571: signal is true;
	signal G10572: std_logic; attribute dont_touch of G10572: signal is true;
	signal G10573: std_logic; attribute dont_touch of G10573: signal is true;
	signal G10578: std_logic; attribute dont_touch of G10578: signal is true;
	signal G10581: std_logic; attribute dont_touch of G10581: signal is true;
	signal G10582: std_logic; attribute dont_touch of G10582: signal is true;
	signal G10583: std_logic; attribute dont_touch of G10583: signal is true;
	signal G10584: std_logic; attribute dont_touch of G10584: signal is true;
	signal G10585: std_logic; attribute dont_touch of G10585: signal is true;
	signal G10586: std_logic; attribute dont_touch of G10586: signal is true;
	signal G10587: std_logic; attribute dont_touch of G10587: signal is true;
	signal G10588: std_logic; attribute dont_touch of G10588: signal is true;
	signal G10589: std_logic; attribute dont_touch of G10589: signal is true;
	signal G10590: std_logic; attribute dont_touch of G10590: signal is true;
	signal G10597: std_logic; attribute dont_touch of G10597: signal is true;
	signal G10598: std_logic; attribute dont_touch of G10598: signal is true;
	signal G10601: std_logic; attribute dont_touch of G10601: signal is true;
	signal G10602: std_logic; attribute dont_touch of G10602: signal is true;
	signal G10603: std_logic; attribute dont_touch of G10603: signal is true;
	signal G10604: std_logic; attribute dont_touch of G10604: signal is true;
	signal G10605: std_logic; attribute dont_touch of G10605: signal is true;
	signal G10606: std_logic; attribute dont_touch of G10606: signal is true;
	signal G10607: std_logic; attribute dont_touch of G10607: signal is true;
	signal G10608: std_logic; attribute dont_touch of G10608: signal is true;
	signal G10609: std_logic; attribute dont_touch of G10609: signal is true;
	signal G10610: std_logic; attribute dont_touch of G10610: signal is true;
	signal G10611: std_logic; attribute dont_touch of G10611: signal is true;
	signal G10612: std_logic; attribute dont_touch of G10612: signal is true;
	signal G10613: std_logic; attribute dont_touch of G10613: signal is true;
	signal G10614: std_logic; attribute dont_touch of G10614: signal is true;
	signal G10615: std_logic; attribute dont_touch of G10615: signal is true;
	signal G10616: std_logic; attribute dont_touch of G10616: signal is true;
	signal G10617: std_logic; attribute dont_touch of G10617: signal is true;
	signal G10618: std_logic; attribute dont_touch of G10618: signal is true;
	signal G10619: std_logic; attribute dont_touch of G10619: signal is true;
	signal G10620: std_logic; attribute dont_touch of G10620: signal is true;
	signal G10621: std_logic; attribute dont_touch of G10621: signal is true;
	signal G10622: std_logic; attribute dont_touch of G10622: signal is true;
	signal G10623: std_logic; attribute dont_touch of G10623: signal is true;
	signal G10624: std_logic; attribute dont_touch of G10624: signal is true;
	signal G10625: std_logic; attribute dont_touch of G10625: signal is true;
	signal G10626: std_logic; attribute dont_touch of G10626: signal is true;
	signal G10627: std_logic; attribute dont_touch of G10627: signal is true;
	signal G10632: std_logic; attribute dont_touch of G10632: signal is true;
	signal G10649: std_logic; attribute dont_touch of G10649: signal is true;
	signal G10652: std_logic; attribute dont_touch of G10652: signal is true;
	signal G10653: std_logic; attribute dont_touch of G10653: signal is true;
	signal G10654: std_logic; attribute dont_touch of G10654: signal is true;
	signal G10655: std_logic; attribute dont_touch of G10655: signal is true;
	signal G10656: std_logic; attribute dont_touch of G10656: signal is true;
	signal G10657: std_logic; attribute dont_touch of G10657: signal is true;
	signal G10658: std_logic; attribute dont_touch of G10658: signal is true;
	signal G10664: std_logic; attribute dont_touch of G10664: signal is true;
	signal G10665: std_logic; attribute dont_touch of G10665: signal is true;
	signal G10666: std_logic; attribute dont_touch of G10666: signal is true;
	signal G10671: std_logic; attribute dont_touch of G10671: signal is true;
	signal G10674: std_logic; attribute dont_touch of G10674: signal is true;
	signal G10675: std_logic; attribute dont_touch of G10675: signal is true;
	signal G10676: std_logic; attribute dont_touch of G10676: signal is true;
	signal G10677: std_logic; attribute dont_touch of G10677: signal is true;
	signal G10678: std_logic; attribute dont_touch of G10678: signal is true;
	signal G10683: std_logic; attribute dont_touch of G10683: signal is true;
	signal G10684: std_logic; attribute dont_touch of G10684: signal is true;
	signal G10685: std_logic; attribute dont_touch of G10685: signal is true;
	signal G10695: std_logic; attribute dont_touch of G10695: signal is true;
	signal G10699: std_logic; attribute dont_touch of G10699: signal is true;
	signal G10704: std_logic; attribute dont_touch of G10704: signal is true;
	signal G10705: std_logic; attribute dont_touch of G10705: signal is true;
	signal G10706: std_logic; attribute dont_touch of G10706: signal is true;
	signal G10707: std_logic; attribute dont_touch of G10707: signal is true;
	signal G10708: std_logic; attribute dont_touch of G10708: signal is true;
	signal G10709: std_logic; attribute dont_touch of G10709: signal is true;
	signal G10710: std_logic; attribute dont_touch of G10710: signal is true;
	signal G10715: std_logic; attribute dont_touch of G10715: signal is true;
	signal G10719: std_logic; attribute dont_touch of G10719: signal is true;
	signal G10720: std_logic; attribute dont_touch of G10720: signal is true;
	signal G10721: std_logic; attribute dont_touch of G10721: signal is true;
	signal G10724: std_logic; attribute dont_touch of G10724: signal is true;
	signal G10725: std_logic; attribute dont_touch of G10725: signal is true;
	signal G10726: std_logic; attribute dont_touch of G10726: signal is true;
	signal G10727: std_logic; attribute dont_touch of G10727: signal is true;
	signal G10732: std_logic; attribute dont_touch of G10732: signal is true;
	signal G10733: std_logic; attribute dont_touch of G10733: signal is true;
	signal G10736: std_logic; attribute dont_touch of G10736: signal is true;
	signal G10737: std_logic; attribute dont_touch of G10737: signal is true;
	signal G10738: std_logic; attribute dont_touch of G10738: signal is true;
	signal G10741: std_logic; attribute dont_touch of G10741: signal is true;
	signal G10754: std_logic; attribute dont_touch of G10754: signal is true;
	signal G10755: std_logic; attribute dont_touch of G10755: signal is true;
	signal G10756: std_logic; attribute dont_touch of G10756: signal is true;
	signal G10759: std_logic; attribute dont_touch of G10759: signal is true;
	signal G10760: std_logic; attribute dont_touch of G10760: signal is true;
	signal G10761: std_logic; attribute dont_touch of G10761: signal is true;
	signal G10762: std_logic; attribute dont_touch of G10762: signal is true;
	signal G10775: std_logic; attribute dont_touch of G10775: signal is true;
	signal G10776: std_logic; attribute dont_touch of G10776: signal is true;
	signal G10793: std_logic; attribute dont_touch of G10793: signal is true;
	signal G10794: std_logic; attribute dont_touch of G10794: signal is true;
	signal G10795: std_logic; attribute dont_touch of G10795: signal is true;
	signal G10796: std_logic; attribute dont_touch of G10796: signal is true;
	signal G10799: std_logic; attribute dont_touch of G10799: signal is true;
	signal G10800: std_logic; attribute dont_touch of G10800: signal is true;
	signal G10801: std_logic; attribute dont_touch of G10801: signal is true;
	signal G10802: std_logic; attribute dont_touch of G10802: signal is true;
	signal G10803: std_logic; attribute dont_touch of G10803: signal is true;
	signal G10804: std_logic; attribute dont_touch of G10804: signal is true;
	signal G10805: std_logic; attribute dont_touch of G10805: signal is true;
	signal G10808: std_logic; attribute dont_touch of G10808: signal is true;
	signal G10812: std_logic; attribute dont_touch of G10812: signal is true;
	signal G10815: std_logic; attribute dont_touch of G10815: signal is true;
	signal G10816: std_logic; attribute dont_touch of G10816: signal is true;
	signal G10819: std_logic; attribute dont_touch of G10819: signal is true;
	signal G10820: std_logic; attribute dont_touch of G10820: signal is true;
	signal G10821: std_logic; attribute dont_touch of G10821: signal is true;
	signal G10822: std_logic; attribute dont_touch of G10822: signal is true;
	signal G10823: std_logic; attribute dont_touch of G10823: signal is true;
	signal G10827: std_logic; attribute dont_touch of G10827: signal is true;
	signal G10828: std_logic; attribute dont_touch of G10828: signal is true;
	signal G10829: std_logic; attribute dont_touch of G10829: signal is true;
	signal G10830: std_logic; attribute dont_touch of G10830: signal is true;
	signal G10831: std_logic; attribute dont_touch of G10831: signal is true;
	signal G10838: std_logic; attribute dont_touch of G10838: signal is true;
	signal G10841: std_logic; attribute dont_touch of G10841: signal is true;
	signal G10851: std_logic; attribute dont_touch of G10851: signal is true;
	signal G10856: std_logic; attribute dont_touch of G10856: signal is true;
	signal G10857: std_logic; attribute dont_touch of G10857: signal is true;
	signal G10862: std_logic; attribute dont_touch of G10862: signal is true;
	signal G10869: std_logic; attribute dont_touch of G10869: signal is true;
	signal G10872: std_logic; attribute dont_touch of G10872: signal is true;
	signal G10873: std_logic; attribute dont_touch of G10873: signal is true;
	signal G10874: std_logic; attribute dont_touch of G10874: signal is true;
	signal G10877: std_logic; attribute dont_touch of G10877: signal is true;
	signal G10878: std_logic; attribute dont_touch of G10878: signal is true;
	signal G10881: std_logic; attribute dont_touch of G10881: signal is true;
	signal G10882: std_logic; attribute dont_touch of G10882: signal is true;
	signal G10883: std_logic; attribute dont_touch of G10883: signal is true;
	signal G10884: std_logic; attribute dont_touch of G10884: signal is true;
	signal G10887: std_logic; attribute dont_touch of G10887: signal is true;
	signal G10890: std_logic; attribute dont_touch of G10890: signal is true;
	signal G10893: std_logic; attribute dont_touch of G10893: signal is true;
	signal G10896: std_logic; attribute dont_touch of G10896: signal is true;
	signal G10897: std_logic; attribute dont_touch of G10897: signal is true;
	signal G10898: std_logic; attribute dont_touch of G10898: signal is true;
	signal G10899: std_logic; attribute dont_touch of G10899: signal is true;
	signal G10902: std_logic; attribute dont_touch of G10902: signal is true;
	signal G10905: std_logic; attribute dont_touch of G10905: signal is true;
	signal G10909: std_logic; attribute dont_touch of G10909: signal is true;
	signal G10916: std_logic; attribute dont_touch of G10916: signal is true;
	signal G10917: std_logic; attribute dont_touch of G10917: signal is true;
	signal G10918: std_logic; attribute dont_touch of G10918: signal is true;
	signal G10921: std_logic; attribute dont_touch of G10921: signal is true;
	signal G10922: std_logic; attribute dont_touch of G10922: signal is true;
	signal G10925: std_logic; attribute dont_touch of G10925: signal is true;
	signal G10928: std_logic; attribute dont_touch of G10928: signal is true;
	signal G10929: std_logic; attribute dont_touch of G10929: signal is true;
	signal G10934: std_logic; attribute dont_touch of G10934: signal is true;
	signal G10935: std_logic; attribute dont_touch of G10935: signal is true;
	signal G10939: std_logic; attribute dont_touch of G10939: signal is true;
	signal G10946: std_logic; attribute dont_touch of G10946: signal is true;
	signal G10947: std_logic; attribute dont_touch of G10947: signal is true;
	signal G10948: std_logic; attribute dont_touch of G10948: signal is true;
	signal G10951: std_logic; attribute dont_touch of G10951: signal is true;
	signal G10960: std_logic; attribute dont_touch of G10960: signal is true;
	signal G10961: std_logic; attribute dont_touch of G10961: signal is true;
	signal G10966: std_logic; attribute dont_touch of G10966: signal is true;
	signal G10967: std_logic; attribute dont_touch of G10967: signal is true;
	signal G10970: std_logic; attribute dont_touch of G10970: signal is true;
	signal G10971: std_logic; attribute dont_touch of G10971: signal is true;
	signal G10980: std_logic; attribute dont_touch of G10980: signal is true;
	signal G10981: std_logic; attribute dont_touch of G10981: signal is true;
	signal G10998: std_logic; attribute dont_touch of G10998: signal is true;
	signal G10999: std_logic; attribute dont_touch of G10999: signal is true;
	signal G11002: std_logic; attribute dont_touch of G11002: signal is true;
	signal G11003: std_logic; attribute dont_touch of G11003: signal is true;
	signal G11006: std_logic; attribute dont_touch of G11006: signal is true;
	signal G11010: std_logic; attribute dont_touch of G11010: signal is true;
	signal G11011: std_logic; attribute dont_touch of G11011: signal is true;
	signal G11012: std_logic; attribute dont_touch of G11012: signal is true;
	signal G11016: std_logic; attribute dont_touch of G11016: signal is true;
	signal G11017: std_logic; attribute dont_touch of G11017: signal is true;
	signal G11018: std_logic; attribute dont_touch of G11018: signal is true;
	signal G11019: std_logic; attribute dont_touch of G11019: signal is true;
	signal G11020: std_logic; attribute dont_touch of G11020: signal is true;
	signal G11023: std_logic; attribute dont_touch of G11023: signal is true;
	signal G11024: std_logic; attribute dont_touch of G11024: signal is true;
	signal G11025: std_logic; attribute dont_touch of G11025: signal is true;
	signal G11026: std_logic; attribute dont_touch of G11026: signal is true;
	signal G11027: std_logic; attribute dont_touch of G11027: signal is true;
	signal G11028: std_logic; attribute dont_touch of G11028: signal is true;
	signal G11029: std_logic; attribute dont_touch of G11029: signal is true;
	signal G11030: std_logic; attribute dont_touch of G11030: signal is true;
	signal G11031: std_logic; attribute dont_touch of G11031: signal is true;
	signal G11032: std_logic; attribute dont_touch of G11032: signal is true;
	signal G11033: std_logic; attribute dont_touch of G11033: signal is true;
	signal G11034: std_logic; attribute dont_touch of G11034: signal is true;
	signal G11035: std_logic; attribute dont_touch of G11035: signal is true;
	signal G11036: std_logic; attribute dont_touch of G11036: signal is true;
	signal G11037: std_logic; attribute dont_touch of G11037: signal is true;
	signal G11038: std_logic; attribute dont_touch of G11038: signal is true;
	signal G11039: std_logic; attribute dont_touch of G11039: signal is true;
	signal G11042: std_logic; attribute dont_touch of G11042: signal is true;
	signal G11043: std_logic; attribute dont_touch of G11043: signal is true;
	signal G11044: std_logic; attribute dont_touch of G11044: signal is true;
	signal G11045: std_logic; attribute dont_touch of G11045: signal is true;
	signal G11046: std_logic; attribute dont_touch of G11046: signal is true;
	signal G11047: std_logic; attribute dont_touch of G11047: signal is true;
	signal G11048: std_logic; attribute dont_touch of G11048: signal is true;
	signal G11083: std_logic; attribute dont_touch of G11083: signal is true;
	signal G11107: std_logic; attribute dont_touch of G11107: signal is true;
	signal G11110: std_logic; attribute dont_touch of G11110: signal is true;
	signal G11111: std_logic; attribute dont_touch of G11111: signal is true;
	signal G11114: std_logic; attribute dont_touch of G11114: signal is true;
	signal G11115: std_logic; attribute dont_touch of G11115: signal is true;
	signal G11116: std_logic; attribute dont_touch of G11116: signal is true;
	signal G11117: std_logic; attribute dont_touch of G11117: signal is true;
	signal G11118: std_logic; attribute dont_touch of G11118: signal is true;
	signal G11119: std_logic; attribute dont_touch of G11119: signal is true;
	signal G11122: std_logic; attribute dont_touch of G11122: signal is true;
	signal G11123: std_logic; attribute dont_touch of G11123: signal is true;
	signal G11126: std_logic; attribute dont_touch of G11126: signal is true;
	signal G11127: std_logic; attribute dont_touch of G11127: signal is true;
	signal G11128: std_logic; attribute dont_touch of G11128: signal is true;
	signal G11129: std_logic; attribute dont_touch of G11129: signal is true;
	signal G11130: std_logic; attribute dont_touch of G11130: signal is true;
	signal G11134: std_logic; attribute dont_touch of G11134: signal is true;
	signal G11135: std_logic; attribute dont_touch of G11135: signal is true;
	signal G11136: std_logic; attribute dont_touch of G11136: signal is true;
	signal G11139: std_logic; attribute dont_touch of G11139: signal is true;
	signal G11142: std_logic; attribute dont_touch of G11142: signal is true;
	signal G11143: std_logic; attribute dont_touch of G11143: signal is true;
	signal G11144: std_logic; attribute dont_touch of G11144: signal is true;
	signal G11147: std_logic; attribute dont_touch of G11147: signal is true;
	signal G11148: std_logic; attribute dont_touch of G11148: signal is true;
	signal G11149: std_logic; attribute dont_touch of G11149: signal is true;
	signal G11153: std_logic; attribute dont_touch of G11153: signal is true;
	signal G11154: std_logic; attribute dont_touch of G11154: signal is true;
	signal G11155: std_logic; attribute dont_touch of G11155: signal is true;
	signal G11160: std_logic; attribute dont_touch of G11160: signal is true;
	signal G11163: std_logic; attribute dont_touch of G11163: signal is true;
	signal G11164: std_logic; attribute dont_touch of G11164: signal is true;
	signal G11165: std_logic; attribute dont_touch of G11165: signal is true;
	signal G11166: std_logic; attribute dont_touch of G11166: signal is true;
	signal G11169: std_logic; attribute dont_touch of G11169: signal is true;
	signal G11170: std_logic; attribute dont_touch of G11170: signal is true;
	signal G11171: std_logic; attribute dont_touch of G11171: signal is true;
	signal G11172: std_logic; attribute dont_touch of G11172: signal is true;
	signal G11173: std_logic; attribute dont_touch of G11173: signal is true;
	signal G11178: std_logic; attribute dont_touch of G11178: signal is true;
	signal G11181: std_logic; attribute dont_touch of G11181: signal is true;
	signal G11182: std_logic; attribute dont_touch of G11182: signal is true;
	signal G11183: std_logic; attribute dont_touch of G11183: signal is true;
	signal G11184: std_logic; attribute dont_touch of G11184: signal is true;
	signal G11185: std_logic; attribute dont_touch of G11185: signal is true;
	signal G11189: std_logic; attribute dont_touch of G11189: signal is true;
	signal G11190: std_logic; attribute dont_touch of G11190: signal is true;
	signal G11191: std_logic; attribute dont_touch of G11191: signal is true;
	signal G11192: std_logic; attribute dont_touch of G11192: signal is true;
	signal G11193: std_logic; attribute dont_touch of G11193: signal is true;
	signal G11194: std_logic; attribute dont_touch of G11194: signal is true;
	signal G11200: std_logic; attribute dont_touch of G11200: signal is true;
	signal G11201: std_logic; attribute dont_touch of G11201: signal is true;
	signal G11202: std_logic; attribute dont_touch of G11202: signal is true;
	signal G11203: std_logic; attribute dont_touch of G11203: signal is true;
	signal G11204: std_logic; attribute dont_touch of G11204: signal is true;
	signal G11205: std_logic; attribute dont_touch of G11205: signal is true;
	signal G11206: std_logic; attribute dont_touch of G11206: signal is true;
	signal G11207: std_logic; attribute dont_touch of G11207: signal is true;
	signal G11213: std_logic; attribute dont_touch of G11213: signal is true;
	signal G11214: std_logic; attribute dont_touch of G11214: signal is true;
	signal G11215: std_logic; attribute dont_touch of G11215: signal is true;
	signal G11216: std_logic; attribute dont_touch of G11216: signal is true;
	signal G11217: std_logic; attribute dont_touch of G11217: signal is true;
	signal G11223: std_logic; attribute dont_touch of G11223: signal is true;
	signal G11224: std_logic; attribute dont_touch of G11224: signal is true;
	signal G11225: std_logic; attribute dont_touch of G11225: signal is true;
	signal G11231: std_logic; attribute dont_touch of G11231: signal is true;
	signal G11232: std_logic; attribute dont_touch of G11232: signal is true;
	signal G11233: std_logic; attribute dont_touch of G11233: signal is true;
	signal G11234: std_logic; attribute dont_touch of G11234: signal is true;
	signal G11235: std_logic; attribute dont_touch of G11235: signal is true;
	signal G11236: std_logic; attribute dont_touch of G11236: signal is true;
	signal G11237: std_logic; attribute dont_touch of G11237: signal is true;
	signal G11238: std_logic; attribute dont_touch of G11238: signal is true;
	signal G11244: std_logic; attribute dont_touch of G11244: signal is true;
	signal G11245: std_logic; attribute dont_touch of G11245: signal is true;
	signal G11248: std_logic; attribute dont_touch of G11248: signal is true;
	signal G11249: std_logic; attribute dont_touch of G11249: signal is true;
	signal G11250: std_logic; attribute dont_touch of G11250: signal is true;
	signal G11251: std_logic; attribute dont_touch of G11251: signal is true;
	signal G11252: std_logic; attribute dont_touch of G11252: signal is true;
	signal G11255: std_logic; attribute dont_touch of G11255: signal is true;
	signal G11261: std_logic; attribute dont_touch of G11261: signal is true;
	signal G11268: std_logic; attribute dont_touch of G11268: signal is true;
	signal G11269: std_logic; attribute dont_touch of G11269: signal is true;
	signal G11270: std_logic; attribute dont_touch of G11270: signal is true;
	signal G11273: std_logic; attribute dont_touch of G11273: signal is true;
	signal G11276: std_logic; attribute dont_touch of G11276: signal is true;
	signal G11279: std_logic; attribute dont_touch of G11279: signal is true;
	signal G11280: std_logic; attribute dont_touch of G11280: signal is true;
	signal G11283: std_logic; attribute dont_touch of G11283: signal is true;
	signal G11290: std_logic; attribute dont_touch of G11290: signal is true;
	signal G11291: std_logic; attribute dont_touch of G11291: signal is true;
	signal G11292: std_logic; attribute dont_touch of G11292: signal is true;
	signal G11293: std_logic; attribute dont_touch of G11293: signal is true;
	signal G11294: std_logic; attribute dont_touch of G11294: signal is true;
	signal G11302: std_logic; attribute dont_touch of G11302: signal is true;
	signal G11303: std_logic; attribute dont_touch of G11303: signal is true;
	signal G11306: std_logic; attribute dont_touch of G11306: signal is true;
	signal G11309: std_logic; attribute dont_touch of G11309: signal is true;
	signal G11312: std_logic; attribute dont_touch of G11312: signal is true;
	signal G11313: std_logic; attribute dont_touch of G11313: signal is true;
	signal G11316: std_logic; attribute dont_touch of G11316: signal is true;
	signal G11317: std_logic; attribute dont_touch of G11317: signal is true;
	signal G11320: std_logic; attribute dont_touch of G11320: signal is true;
	signal G11323: std_logic; attribute dont_touch of G11323: signal is true;
	signal G11324: std_logic; attribute dont_touch of G11324: signal is true;
	signal G11325: std_logic; attribute dont_touch of G11325: signal is true;
	signal G11326: std_logic; attribute dont_touch of G11326: signal is true;
	signal G11330: std_logic; attribute dont_touch of G11330: signal is true;
	signal G11336: std_logic; attribute dont_touch of G11336: signal is true;
	signal G11344: std_logic; attribute dont_touch of G11344: signal is true;
	signal G11345: std_logic; attribute dont_touch of G11345: signal is true;
	signal G11346: std_logic; attribute dont_touch of G11346: signal is true;
	signal G11350: std_logic; attribute dont_touch of G11350: signal is true;
	signal G11355: std_logic; attribute dont_touch of G11355: signal is true;
	signal G11356: std_logic; attribute dont_touch of G11356: signal is true;
	signal G11357: std_logic; attribute dont_touch of G11357: signal is true;
	signal G11360: std_logic; attribute dont_touch of G11360: signal is true;
	signal G11363: std_logic; attribute dont_touch of G11363: signal is true;
	signal G11366: std_logic; attribute dont_touch of G11366: signal is true;
	signal G11367: std_logic; attribute dont_touch of G11367: signal is true;
	signal G11370: std_logic; attribute dont_touch of G11370: signal is true;
	signal G11371: std_logic; attribute dont_touch of G11371: signal is true;
	signal G11372: std_logic; attribute dont_touch of G11372: signal is true;
	signal G11373: std_logic; attribute dont_touch of G11373: signal is true;
	signal G11374: std_logic; attribute dont_touch of G11374: signal is true;
	signal G11380: std_logic; attribute dont_touch of G11380: signal is true;
	signal G11381: std_logic; attribute dont_touch of G11381: signal is true;
	signal G11382: std_logic; attribute dont_touch of G11382: signal is true;
	signal G11383: std_logic; attribute dont_touch of G11383: signal is true;
	signal G11384: std_logic; attribute dont_touch of G11384: signal is true;
	signal G11385: std_logic; attribute dont_touch of G11385: signal is true;
	signal G11389: std_logic; attribute dont_touch of G11389: signal is true;
	signal G11394: std_logic; attribute dont_touch of G11394: signal is true;
	signal G11395: std_logic; attribute dont_touch of G11395: signal is true;
	signal G11396: std_logic; attribute dont_touch of G11396: signal is true;
	signal G11397: std_logic; attribute dont_touch of G11397: signal is true;
	signal G11398: std_logic; attribute dont_touch of G11398: signal is true;
	signal G11401: std_logic; attribute dont_touch of G11401: signal is true;
	signal G11402: std_logic; attribute dont_touch of G11402: signal is true;
	signal G11403: std_logic; attribute dont_touch of G11403: signal is true;
	signal G11404: std_logic; attribute dont_touch of G11404: signal is true;
	signal G11405: std_logic; attribute dont_touch of G11405: signal is true;
	signal G11409: std_logic; attribute dont_touch of G11409: signal is true;
	signal G11410: std_logic; attribute dont_touch of G11410: signal is true;
	signal G11411: std_logic; attribute dont_touch of G11411: signal is true;
	signal G11412: std_logic; attribute dont_touch of G11412: signal is true;
	signal G11413: std_logic; attribute dont_touch of G11413: signal is true;
	signal G11414: std_logic; attribute dont_touch of G11414: signal is true;
	signal G11415: std_logic; attribute dont_touch of G11415: signal is true;
	signal G11419: std_logic; attribute dont_touch of G11419: signal is true;
	signal G11424: std_logic; attribute dont_touch of G11424: signal is true;
	signal G11425: std_logic; attribute dont_touch of G11425: signal is true;
	signal G11426: std_logic; attribute dont_touch of G11426: signal is true;
	signal G11427: std_logic; attribute dont_touch of G11427: signal is true;
	signal G11428: std_logic; attribute dont_touch of G11428: signal is true;
	signal G11429: std_logic; attribute dont_touch of G11429: signal is true;
	signal G11430: std_logic; attribute dont_touch of G11430: signal is true;
	signal G11431: std_logic; attribute dont_touch of G11431: signal is true;
	signal G11432: std_logic; attribute dont_touch of G11432: signal is true;
	signal G11435: std_logic; attribute dont_touch of G11435: signal is true;
	signal G11441: std_logic; attribute dont_touch of G11441: signal is true;
	signal G11442: std_logic; attribute dont_touch of G11442: signal is true;
	signal G11443: std_logic; attribute dont_touch of G11443: signal is true;
	signal G11444: std_logic; attribute dont_touch of G11444: signal is true;
	signal G11445: std_logic; attribute dont_touch of G11445: signal is true;
	signal G11446: std_logic; attribute dont_touch of G11446: signal is true;
	signal G11448: std_logic; attribute dont_touch of G11448: signal is true;
	signal G11449: std_logic; attribute dont_touch of G11449: signal is true;
	signal G11450: std_logic; attribute dont_touch of G11450: signal is true;
	signal G11467: std_logic; attribute dont_touch of G11467: signal is true;
	signal G11468: std_logic; attribute dont_touch of G11468: signal is true;
	signal G11469: std_logic; attribute dont_touch of G11469: signal is true;
	signal G11470: std_logic; attribute dont_touch of G11470: signal is true;
	signal G11471: std_logic; attribute dont_touch of G11471: signal is true;
	signal G11472: std_logic; attribute dont_touch of G11472: signal is true;
	signal G11473: std_logic; attribute dont_touch of G11473: signal is true;
	signal G11479: std_logic; attribute dont_touch of G11479: signal is true;
	signal G11480: std_logic; attribute dont_touch of G11480: signal is true;
	signal G11483: std_logic; attribute dont_touch of G11483: signal is true;
	signal G11489: std_logic; attribute dont_touch of G11489: signal is true;
	signal G11490: std_logic; attribute dont_touch of G11490: signal is true;
	signal G11491: std_logic; attribute dont_touch of G11491: signal is true;
	signal G11492: std_logic; attribute dont_touch of G11492: signal is true;
	signal G11493: std_logic; attribute dont_touch of G11493: signal is true;
	signal G11496: std_logic; attribute dont_touch of G11496: signal is true;
	signal G11497: std_logic; attribute dont_touch of G11497: signal is true;
	signal G11498: std_logic; attribute dont_touch of G11498: signal is true;
	signal G11509: std_logic; attribute dont_touch of G11509: signal is true;
	signal G11510: std_logic; attribute dont_touch of G11510: signal is true;
	signal G11511: std_logic; attribute dont_touch of G11511: signal is true;
	signal G11512: std_logic; attribute dont_touch of G11512: signal is true;
	signal G11513: std_logic; attribute dont_touch of G11513: signal is true;
	signal G11514: std_logic; attribute dont_touch of G11514: signal is true;
	signal G11519: std_logic; attribute dont_touch of G11519: signal is true;
	signal G11527: std_logic; attribute dont_touch of G11527: signal is true;
	signal G11533: std_logic; attribute dont_touch of G11533: signal is true;
	signal G11534: std_logic; attribute dont_touch of G11534: signal is true;
	signal G11537: std_logic; attribute dont_touch of G11537: signal is true;
	signal G11543: std_logic; attribute dont_touch of G11543: signal is true;
	signal G11544: std_logic; attribute dont_touch of G11544: signal is true;
	signal G11545: std_logic; attribute dont_touch of G11545: signal is true;
	signal G11546: std_logic; attribute dont_touch of G11546: signal is true;
	signal G11547: std_logic; attribute dont_touch of G11547: signal is true;
	signal G11559: std_logic; attribute dont_touch of G11559: signal is true;
	signal G11560: std_logic; attribute dont_touch of G11560: signal is true;
	signal G11561: std_logic; attribute dont_touch of G11561: signal is true;
	signal G11562: std_logic; attribute dont_touch of G11562: signal is true;
	signal G11563: std_logic; attribute dont_touch of G11563: signal is true;
	signal G11566: std_logic; attribute dont_touch of G11566: signal is true;
	signal G11571: std_logic; attribute dont_touch of G11571: signal is true;
	signal G11576: std_logic; attribute dont_touch of G11576: signal is true;
	signal G11584: std_logic; attribute dont_touch of G11584: signal is true;
	signal G11590: std_logic; attribute dont_touch of G11590: signal is true;
	signal G11591: std_logic; attribute dont_touch of G11591: signal is true;
	signal G11592: std_logic; attribute dont_touch of G11592: signal is true;
	signal G11607: std_logic; attribute dont_touch of G11607: signal is true;
	signal G11608: std_logic; attribute dont_touch of G11608: signal is true;
	signal G11609: std_logic; attribute dont_touch of G11609: signal is true;
	signal G11610: std_logic; attribute dont_touch of G11610: signal is true;
	signal G11615: std_logic; attribute dont_touch of G11615: signal is true;
	signal G11618: std_logic; attribute dont_touch of G11618: signal is true;
	signal G11621: std_logic; attribute dont_touch of G11621: signal is true;
	signal G11626: std_logic; attribute dont_touch of G11626: signal is true;
	signal G11631: std_logic; attribute dont_touch of G11631: signal is true;
	signal G11639: std_logic; attribute dont_touch of G11639: signal is true;
	signal G11640: std_logic; attribute dont_touch of G11640: signal is true;
	signal G11652: std_logic; attribute dont_touch of G11652: signal is true;
	signal G11653: std_logic; attribute dont_touch of G11653: signal is true;
	signal G11658: std_logic; attribute dont_touch of G11658: signal is true;
	signal G11663: std_logic; attribute dont_touch of G11663: signal is true;
	signal G11666: std_logic; attribute dont_touch of G11666: signal is true;
	signal G11669: std_logic; attribute dont_touch of G11669: signal is true;
	signal G11674: std_logic; attribute dont_touch of G11674: signal is true;
	signal G11675: std_logic; attribute dont_touch of G11675: signal is true;
	signal G11676: std_logic; attribute dont_touch of G11676: signal is true;
	signal G11677: std_logic; attribute dont_touch of G11677: signal is true;
	signal G11679: std_logic; attribute dont_touch of G11679: signal is true;
	signal G11686: std_logic; attribute dont_touch of G11686: signal is true;
	signal G11691: std_logic; attribute dont_touch of G11691: signal is true;
	signal G11692: std_logic; attribute dont_touch of G11692: signal is true;
	signal G11697: std_logic; attribute dont_touch of G11697: signal is true;
	signal G11702: std_logic; attribute dont_touch of G11702: signal is true;
	signal G11705: std_logic; attribute dont_touch of G11705: signal is true;
	signal G11706: std_logic; attribute dont_touch of G11706: signal is true;
	signal G11707: std_logic; attribute dont_touch of G11707: signal is true;
	signal G11708: std_logic; attribute dont_touch of G11708: signal is true;
	signal G11709: std_logic; attribute dont_touch of G11709: signal is true;
	signal G11714: std_logic; attribute dont_touch of G11714: signal is true;
	signal G11715: std_logic; attribute dont_touch of G11715: signal is true;
	signal G11720: std_logic; attribute dont_touch of G11720: signal is true;
	signal G11721: std_logic; attribute dont_touch of G11721: signal is true;
	signal G11724: std_logic; attribute dont_touch of G11724: signal is true;
	signal G11729: std_logic; attribute dont_touch of G11729: signal is true;
	signal G11735: std_logic; attribute dont_touch of G11735: signal is true;
	signal G11736: std_logic; attribute dont_touch of G11736: signal is true;
	signal G11737: std_logic; attribute dont_touch of G11737: signal is true;
	signal G11740: std_logic; attribute dont_touch of G11740: signal is true;
	signal G11741: std_logic; attribute dont_touch of G11741: signal is true;
	signal G11744: std_logic; attribute dont_touch of G11744: signal is true;
	signal G11747: std_logic; attribute dont_touch of G11747: signal is true;
	signal G11753: std_logic; attribute dont_touch of G11753: signal is true;
	signal G11754: std_logic; attribute dont_touch of G11754: signal is true;
	signal G11755: std_logic; attribute dont_touch of G11755: signal is true;
	signal G11761: std_logic; attribute dont_touch of G11761: signal is true;
	signal G11762: std_logic; attribute dont_touch of G11762: signal is true;
	signal G11763: std_logic; attribute dont_touch of G11763: signal is true;
	signal G11769: std_logic; attribute dont_touch of G11769: signal is true;
	signal G11771: std_logic; attribute dont_touch of G11771: signal is true;
	signal G11772: std_logic; attribute dont_touch of G11772: signal is true;
	signal G11773: std_logic; attribute dont_touch of G11773: signal is true;
	signal G11779: std_logic; attribute dont_touch of G11779: signal is true;
	signal G11780: std_logic; attribute dont_touch of G11780: signal is true;
	signal G11786: std_logic; attribute dont_touch of G11786: signal is true;
	signal G11790: std_logic; attribute dont_touch of G11790: signal is true;
	signal G11793: std_logic; attribute dont_touch of G11793: signal is true;
	signal G11796: std_logic; attribute dont_touch of G11796: signal is true;
	signal G11797: std_logic; attribute dont_touch of G11797: signal is true;
	signal G11804: std_logic; attribute dont_touch of G11804: signal is true;
	signal G11810: std_logic; attribute dont_touch of G11810: signal is true;
	signal G11811: std_logic; attribute dont_touch of G11811: signal is true;
	signal G11812: std_logic; attribute dont_touch of G11812: signal is true;
	signal G11815: std_logic; attribute dont_touch of G11815: signal is true;
	signal G11819: std_logic; attribute dont_touch of G11819: signal is true;
	signal G11820: std_logic; attribute dont_touch of G11820: signal is true;
	signal G11823: std_logic; attribute dont_touch of G11823: signal is true;
	signal G11826: std_logic; attribute dont_touch of G11826: signal is true;
	signal G11829: std_logic; attribute dont_touch of G11829: signal is true;
	signal G11832: std_logic; attribute dont_touch of G11832: signal is true;
	signal G11833: std_logic; attribute dont_touch of G11833: signal is true;
	signal G11834: std_logic; attribute dont_touch of G11834: signal is true;
	signal G11841: std_logic; attribute dont_touch of G11841: signal is true;
	signal G11842: std_logic; attribute dont_touch of G11842: signal is true;
	signal G11845: std_logic; attribute dont_touch of G11845: signal is true;
	signal G11846: std_logic; attribute dont_touch of G11846: signal is true;
	signal G11849: std_logic; attribute dont_touch of G11849: signal is true;
	signal G11852: std_logic; attribute dont_touch of G11852: signal is true;
	signal G11855: std_logic; attribute dont_touch of G11855: signal is true;
	signal G11858: std_logic; attribute dont_touch of G11858: signal is true;
	signal G11861: std_logic; attribute dont_touch of G11861: signal is true;
	signal G11862: std_logic; attribute dont_touch of G11862: signal is true;
	signal G11865: std_logic; attribute dont_touch of G11865: signal is true;
	signal G11866: std_logic; attribute dont_touch of G11866: signal is true;
	signal G11867: std_logic; attribute dont_touch of G11867: signal is true;
	signal G11868: std_logic; attribute dont_touch of G11868: signal is true;
	signal G11869: std_logic; attribute dont_touch of G11869: signal is true;
	signal G11872: std_logic; attribute dont_touch of G11872: signal is true;
	signal G11875: std_logic; attribute dont_touch of G11875: signal is true;
	signal G11878: std_logic; attribute dont_touch of G11878: signal is true;
	signal G11881: std_logic; attribute dont_touch of G11881: signal is true;
	signal G11884: std_logic; attribute dont_touch of G11884: signal is true;
	signal G11885: std_logic; attribute dont_touch of G11885: signal is true;
	signal G11888: std_logic; attribute dont_touch of G11888: signal is true;
	signal G11889: std_logic; attribute dont_touch of G11889: signal is true;
	signal G11890: std_logic; attribute dont_touch of G11890: signal is true;
	signal G11891: std_logic; attribute dont_touch of G11891: signal is true;
	signal G11892: std_logic; attribute dont_touch of G11892: signal is true;
	signal G11893: std_logic; attribute dont_touch of G11893: signal is true;
	signal G11894: std_logic; attribute dont_touch of G11894: signal is true;
	signal G11897: std_logic; attribute dont_touch of G11897: signal is true;
	signal G11900: std_logic; attribute dont_touch of G11900: signal is true;
	signal G11903: std_logic; attribute dont_touch of G11903: signal is true;
	signal G11906: std_logic; attribute dont_touch of G11906: signal is true;
	signal G11907: std_logic; attribute dont_touch of G11907: signal is true;
	signal G11910: std_logic; attribute dont_touch of G11910: signal is true;
	signal G11911: std_logic; attribute dont_touch of G11911: signal is true;
	signal G11912: std_logic; attribute dont_touch of G11912: signal is true;
	signal G11913: std_logic; attribute dont_touch of G11913: signal is true;
	signal G11914: std_logic; attribute dont_touch of G11914: signal is true;
	signal G11915: std_logic; attribute dont_touch of G11915: signal is true;
	signal G11916: std_logic; attribute dont_touch of G11916: signal is true;
	signal G11917: std_logic; attribute dont_touch of G11917: signal is true;
	signal G11920: std_logic; attribute dont_touch of G11920: signal is true;
	signal G11923: std_logic; attribute dont_touch of G11923: signal is true;
	signal G11924: std_logic; attribute dont_touch of G11924: signal is true;
	signal G11927: std_logic; attribute dont_touch of G11927: signal is true;
	signal G11928: std_logic; attribute dont_touch of G11928: signal is true;
	signal G11929: std_logic; attribute dont_touch of G11929: signal is true;
	signal G11930: std_logic; attribute dont_touch of G11930: signal is true;
	signal G11931: std_logic; attribute dont_touch of G11931: signal is true;
	signal G11932: std_logic; attribute dont_touch of G11932: signal is true;
	signal G11933: std_logic; attribute dont_touch of G11933: signal is true;
	signal G11934: std_logic; attribute dont_touch of G11934: signal is true;
	signal G11935: std_logic; attribute dont_touch of G11935: signal is true;
	signal G11936: std_logic; attribute dont_touch of G11936: signal is true;
	signal G11937: std_logic; attribute dont_touch of G11937: signal is true;
	signal G11938: std_logic; attribute dont_touch of G11938: signal is true;
	signal G11939: std_logic; attribute dont_touch of G11939: signal is true;
	signal G11940: std_logic; attribute dont_touch of G11940: signal is true;
	signal G11941: std_logic; attribute dont_touch of G11941: signal is true;
	signal G11944: std_logic; attribute dont_touch of G11944: signal is true;
	signal G11945: std_logic; attribute dont_touch of G11945: signal is true;
	signal G11948: std_logic; attribute dont_touch of G11948: signal is true;
	signal G11949: std_logic; attribute dont_touch of G11949: signal is true;
	signal G11950: std_logic; attribute dont_touch of G11950: signal is true;
	signal G11951: std_logic; attribute dont_touch of G11951: signal is true;
	signal G11952: std_logic; attribute dont_touch of G11952: signal is true;
	signal G11953: std_logic; attribute dont_touch of G11953: signal is true;
	signal G11954: std_logic; attribute dont_touch of G11954: signal is true;
	signal G11955: std_logic; attribute dont_touch of G11955: signal is true;
	signal G11956: std_logic; attribute dont_touch of G11956: signal is true;
	signal G11957: std_logic; attribute dont_touch of G11957: signal is true;
	signal G11958: std_logic; attribute dont_touch of G11958: signal is true;
	signal G11959: std_logic; attribute dont_touch of G11959: signal is true;
	signal G11960: std_logic; attribute dont_touch of G11960: signal is true;
	signal G11961: std_logic; attribute dont_touch of G11961: signal is true;
	signal G11962: std_logic; attribute dont_touch of G11962: signal is true;
	signal G11963: std_logic; attribute dont_touch of G11963: signal is true;
	signal G11964: std_logic; attribute dont_touch of G11964: signal is true;
	signal G11965: std_logic; attribute dont_touch of G11965: signal is true;
	signal G11966: std_logic; attribute dont_touch of G11966: signal is true;
	signal G11967: std_logic; attribute dont_touch of G11967: signal is true;
	signal G11968: std_logic; attribute dont_touch of G11968: signal is true;
	signal G11969: std_logic; attribute dont_touch of G11969: signal is true;
	signal G11970: std_logic; attribute dont_touch of G11970: signal is true;
	signal G11971: std_logic; attribute dont_touch of G11971: signal is true;
	signal G11972: std_logic; attribute dont_touch of G11972: signal is true;
	signal G11973: std_logic; attribute dont_touch of G11973: signal is true;
	signal G11974: std_logic; attribute dont_touch of G11974: signal is true;
	signal G11975: std_logic; attribute dont_touch of G11975: signal is true;
	signal G11976: std_logic; attribute dont_touch of G11976: signal is true;
	signal G11977: std_logic; attribute dont_touch of G11977: signal is true;
	signal G11978: std_logic; attribute dont_touch of G11978: signal is true;
	signal G11979: std_logic; attribute dont_touch of G11979: signal is true;
	signal G11980: std_logic; attribute dont_touch of G11980: signal is true;
	signal G11981: std_logic; attribute dont_touch of G11981: signal is true;
	signal G11984: std_logic; attribute dont_touch of G11984: signal is true;
	signal G11985: std_logic; attribute dont_touch of G11985: signal is true;
	signal G11986: std_logic; attribute dont_touch of G11986: signal is true;
	signal G11987: std_logic; attribute dont_touch of G11987: signal is true;
	signal G11988: std_logic; attribute dont_touch of G11988: signal is true;
	signal G11989: std_logic; attribute dont_touch of G11989: signal is true;
	signal G11990: std_logic; attribute dont_touch of G11990: signal is true;
	signal G11991: std_logic; attribute dont_touch of G11991: signal is true;
	signal G11992: std_logic; attribute dont_touch of G11992: signal is true;
	signal G11993: std_logic; attribute dont_touch of G11993: signal is true;
	signal G11994: std_logic; attribute dont_touch of G11994: signal is true;
	signal G11995: std_logic; attribute dont_touch of G11995: signal is true;
	signal G11996: std_logic; attribute dont_touch of G11996: signal is true;
	signal G11997: std_logic; attribute dont_touch of G11997: signal is true;
	signal G11998: std_logic; attribute dont_touch of G11998: signal is true;
	signal G11999: std_logic; attribute dont_touch of G11999: signal is true;
	signal G12000: std_logic; attribute dont_touch of G12000: signal is true;
	signal G12001: std_logic; attribute dont_touch of G12001: signal is true;
	signal G12002: std_logic; attribute dont_touch of G12002: signal is true;
	signal G12008: std_logic; attribute dont_touch of G12008: signal is true;
	signal G12009: std_logic; attribute dont_touch of G12009: signal is true;
	signal G12012: std_logic; attribute dont_touch of G12012: signal is true;
	signal G12013: std_logic; attribute dont_touch of G12013: signal is true;
	signal G12014: std_logic; attribute dont_touch of G12014: signal is true;
	signal G12015: std_logic; attribute dont_touch of G12015: signal is true;
	signal G12016: std_logic; attribute dont_touch of G12016: signal is true;
	signal G12017: std_logic; attribute dont_touch of G12017: signal is true;
	signal G12018: std_logic; attribute dont_touch of G12018: signal is true;
	signal G12019: std_logic; attribute dont_touch of G12019: signal is true;
	signal G12020: std_logic; attribute dont_touch of G12020: signal is true;
	signal G12021: std_logic; attribute dont_touch of G12021: signal is true;
	signal G12022: std_logic; attribute dont_touch of G12022: signal is true;
	signal G12023: std_logic; attribute dont_touch of G12023: signal is true;
	signal G12024: std_logic; attribute dont_touch of G12024: signal is true;
	signal G12025: std_logic; attribute dont_touch of G12025: signal is true;
	signal G12026: std_logic; attribute dont_touch of G12026: signal is true;
	signal G12027: std_logic; attribute dont_touch of G12027: signal is true;
	signal G12028: std_logic; attribute dont_touch of G12028: signal is true;
	signal G12029: std_logic; attribute dont_touch of G12029: signal is true;
	signal G12035: std_logic; attribute dont_touch of G12035: signal is true;
	signal G12036: std_logic; attribute dont_touch of G12036: signal is true;
	signal G12037: std_logic; attribute dont_touch of G12037: signal is true;
	signal G12038: std_logic; attribute dont_touch of G12038: signal is true;
	signal G12039: std_logic; attribute dont_touch of G12039: signal is true;
	signal G12040: std_logic; attribute dont_touch of G12040: signal is true;
	signal G12041: std_logic; attribute dont_touch of G12041: signal is true;
	signal G12042: std_logic; attribute dont_touch of G12042: signal is true;
	signal G12043: std_logic; attribute dont_touch of G12043: signal is true;
	signal G12044: std_logic; attribute dont_touch of G12044: signal is true;
	signal G12045: std_logic; attribute dont_touch of G12045: signal is true;
	signal G12046: std_logic; attribute dont_touch of G12046: signal is true;
	signal G12047: std_logic; attribute dont_touch of G12047: signal is true;
	signal G12048: std_logic; attribute dont_touch of G12048: signal is true;
	signal G12049: std_logic; attribute dont_touch of G12049: signal is true;
	signal G12050: std_logic; attribute dont_touch of G12050: signal is true;
	signal G12051: std_logic; attribute dont_touch of G12051: signal is true;
	signal G12052: std_logic; attribute dont_touch of G12052: signal is true;
	signal G12053: std_logic; attribute dont_touch of G12053: signal is true;
	signal G12054: std_logic; attribute dont_touch of G12054: signal is true;
	signal G12059: std_logic; attribute dont_touch of G12059: signal is true;
	signal G12065: std_logic; attribute dont_touch of G12065: signal is true;
	signal G12066: std_logic; attribute dont_touch of G12066: signal is true;
	signal G12067: std_logic; attribute dont_touch of G12067: signal is true;
	signal G12073: std_logic; attribute dont_touch of G12073: signal is true;
	signal G12074: std_logic; attribute dont_touch of G12074: signal is true;
	signal G12075: std_logic; attribute dont_touch of G12075: signal is true;
	signal G12076: std_logic; attribute dont_touch of G12076: signal is true;
	signal G12077: std_logic; attribute dont_touch of G12077: signal is true;
	signal G12078: std_logic; attribute dont_touch of G12078: signal is true;
	signal G12079: std_logic; attribute dont_touch of G12079: signal is true;
	signal G12080: std_logic; attribute dont_touch of G12080: signal is true;
	signal G12081: std_logic; attribute dont_touch of G12081: signal is true;
	signal G12082: std_logic; attribute dont_touch of G12082: signal is true;
	signal G12083: std_logic; attribute dont_touch of G12083: signal is true;
	signal G12084: std_logic; attribute dont_touch of G12084: signal is true;
	signal G12085: std_logic; attribute dont_touch of G12085: signal is true;
	signal G12086: std_logic; attribute dont_touch of G12086: signal is true;
	signal G12087: std_logic; attribute dont_touch of G12087: signal is true;
	signal G12088: std_logic; attribute dont_touch of G12088: signal is true;
	signal G12093: std_logic; attribute dont_touch of G12093: signal is true;
	signal G12099: std_logic; attribute dont_touch of G12099: signal is true;
	signal G12100: std_logic; attribute dont_touch of G12100: signal is true;
	signal G12101: std_logic; attribute dont_touch of G12101: signal is true;
	signal G12107: std_logic; attribute dont_touch of G12107: signal is true;
	signal G12108: std_logic; attribute dont_touch of G12108: signal is true;
	signal G12109: std_logic; attribute dont_touch of G12109: signal is true;
	signal G12110: std_logic; attribute dont_touch of G12110: signal is true;
	signal G12111: std_logic; attribute dont_touch of G12111: signal is true;
	signal G12112: std_logic; attribute dont_touch of G12112: signal is true;
	signal G12113: std_logic; attribute dont_touch of G12113: signal is true;
	signal G12114: std_logic; attribute dont_touch of G12114: signal is true;
	signal G12115: std_logic; attribute dont_touch of G12115: signal is true;
	signal G12116: std_logic; attribute dont_touch of G12116: signal is true;
	signal G12117: std_logic; attribute dont_touch of G12117: signal is true;
	signal G12118: std_logic; attribute dont_touch of G12118: signal is true;
	signal G12119: std_logic; attribute dont_touch of G12119: signal is true;
	signal G12120: std_logic; attribute dont_touch of G12120: signal is true;
	signal G12121: std_logic; attribute dont_touch of G12121: signal is true;
	signal G12122: std_logic; attribute dont_touch of G12122: signal is true;
	signal G12123: std_logic; attribute dont_touch of G12123: signal is true;
	signal G12124: std_logic; attribute dont_touch of G12124: signal is true;
	signal G12125: std_logic; attribute dont_touch of G12125: signal is true;
	signal G12126: std_logic; attribute dont_touch of G12126: signal is true;
	signal G12129: std_logic; attribute dont_touch of G12129: signal is true;
	signal G12135: std_logic; attribute dont_touch of G12135: signal is true;
	signal G12136: std_logic; attribute dont_touch of G12136: signal is true;
	signal G12137: std_logic; attribute dont_touch of G12137: signal is true;
	signal G12143: std_logic; attribute dont_touch of G12143: signal is true;
	signal G12144: std_logic; attribute dont_touch of G12144: signal is true;
	signal G12145: std_logic; attribute dont_touch of G12145: signal is true;
	signal G12146: std_logic; attribute dont_touch of G12146: signal is true;
	signal G12147: std_logic; attribute dont_touch of G12147: signal is true;
	signal G12148: std_logic; attribute dont_touch of G12148: signal is true;
	signal G12149: std_logic; attribute dont_touch of G12149: signal is true;
	signal G12150: std_logic; attribute dont_touch of G12150: signal is true;
	signal G12151: std_logic; attribute dont_touch of G12151: signal is true;
	signal G12152: std_logic; attribute dont_touch of G12152: signal is true;
	signal G12153: std_logic; attribute dont_touch of G12153: signal is true;
	signal G12154: std_logic; attribute dont_touch of G12154: signal is true;
	signal G12155: std_logic; attribute dont_touch of G12155: signal is true;
	signal G12159: std_logic; attribute dont_touch of G12159: signal is true;
	signal G12160: std_logic; attribute dont_touch of G12160: signal is true;
	signal G12163: std_logic; attribute dont_touch of G12163: signal is true;
	signal G12166: std_logic; attribute dont_touch of G12166: signal is true;
	signal G12169: std_logic; attribute dont_touch of G12169: signal is true;
	signal G12170: std_logic; attribute dont_touch of G12170: signal is true;
	signal G12173: std_logic; attribute dont_touch of G12173: signal is true;
	signal G12179: std_logic; attribute dont_touch of G12179: signal is true;
	signal G12180: std_logic; attribute dont_touch of G12180: signal is true;
	signal G12181: std_logic; attribute dont_touch of G12181: signal is true;
	signal G12182: std_logic; attribute dont_touch of G12182: signal is true;
	signal G12183: std_logic; attribute dont_touch of G12183: signal is true;
	signal G12185: std_logic; attribute dont_touch of G12185: signal is true;
	signal G12186: std_logic; attribute dont_touch of G12186: signal is true;
	signal G12187: std_logic; attribute dont_touch of G12187: signal is true;
	signal G12188: std_logic; attribute dont_touch of G12188: signal is true;
	signal G12189: std_logic; attribute dont_touch of G12189: signal is true;
	signal G12190: std_logic; attribute dont_touch of G12190: signal is true;
	signal G12191: std_logic; attribute dont_touch of G12191: signal is true;
	signal G12192: std_logic; attribute dont_touch of G12192: signal is true;
	signal G12193: std_logic; attribute dont_touch of G12193: signal is true;
	signal G12194: std_logic; attribute dont_touch of G12194: signal is true;
	signal G12195: std_logic; attribute dont_touch of G12195: signal is true;
	signal G12196: std_logic; attribute dont_touch of G12196: signal is true;
	signal G12197: std_logic; attribute dont_touch of G12197: signal is true;
	signal G12198: std_logic; attribute dont_touch of G12198: signal is true;
	signal G12201: std_logic; attribute dont_touch of G12201: signal is true;
	signal G12204: std_logic; attribute dont_touch of G12204: signal is true;
	signal G12207: std_logic; attribute dont_touch of G12207: signal is true;
	signal G12208: std_logic; attribute dont_touch of G12208: signal is true;
	signal G12211: std_logic; attribute dont_touch of G12211: signal is true;
	signal G12217: std_logic; attribute dont_touch of G12217: signal is true;
	signal G12218: std_logic; attribute dont_touch of G12218: signal is true;
	signal G12219: std_logic; attribute dont_touch of G12219: signal is true;
	signal G12220: std_logic; attribute dont_touch of G12220: signal is true;
	signal G12221: std_logic; attribute dont_touch of G12221: signal is true;
	signal G12222: std_logic; attribute dont_touch of G12222: signal is true;
	signal G12223: std_logic; attribute dont_touch of G12223: signal is true;
	signal G12224: std_logic; attribute dont_touch of G12224: signal is true;
	signal G12225: std_logic; attribute dont_touch of G12225: signal is true;
	signal G12226: std_logic; attribute dont_touch of G12226: signal is true;
	signal G12227: std_logic; attribute dont_touch of G12227: signal is true;
	signal G12228: std_logic; attribute dont_touch of G12228: signal is true;
	signal G12232: std_logic; attribute dont_touch of G12232: signal is true;
	signal G12233: std_logic; attribute dont_touch of G12233: signal is true;
	signal G12234: std_logic; attribute dont_touch of G12234: signal is true;
	signal G12235: std_logic; attribute dont_touch of G12235: signal is true;
	signal G12239: std_logic; attribute dont_touch of G12239: signal is true;
	signal G12244: std_logic; attribute dont_touch of G12244: signal is true;
	signal G12245: std_logic; attribute dont_touch of G12245: signal is true;
	signal G12246: std_logic; attribute dont_touch of G12246: signal is true;
	signal G12249: std_logic; attribute dont_touch of G12249: signal is true;
	signal G12252: std_logic; attribute dont_touch of G12252: signal is true;
	signal G12255: std_logic; attribute dont_touch of G12255: signal is true;
	signal G12256: std_logic; attribute dont_touch of G12256: signal is true;
	signal G12259: std_logic; attribute dont_touch of G12259: signal is true;
	signal G12284: std_logic; attribute dont_touch of G12284: signal is true;
	signal G12285: std_logic; attribute dont_touch of G12285: signal is true;
	signal G12286: std_logic; attribute dont_touch of G12286: signal is true;
	signal G12287: std_logic; attribute dont_touch of G12287: signal is true;
	signal G12288: std_logic; attribute dont_touch of G12288: signal is true;
	signal G12289: std_logic; attribute dont_touch of G12289: signal is true;
	signal G12292: std_logic; attribute dont_touch of G12292: signal is true;
	signal G12293: std_logic; attribute dont_touch of G12293: signal is true;
	signal G12294: std_logic; attribute dont_touch of G12294: signal is true;
	signal G12295: std_logic; attribute dont_touch of G12295: signal is true;
	signal G12296: std_logic; attribute dont_touch of G12296: signal is true;
	signal G12297: std_logic; attribute dont_touch of G12297: signal is true;
	signal G12301: std_logic; attribute dont_touch of G12301: signal is true;
	signal G12306: std_logic; attribute dont_touch of G12306: signal is true;
	signal G12307: std_logic; attribute dont_touch of G12307: signal is true;
	signal G12308: std_logic; attribute dont_touch of G12308: signal is true;
	signal G12311: std_logic; attribute dont_touch of G12311: signal is true;
	signal G12314: std_logic; attribute dont_touch of G12314: signal is true;
	signal G12317: std_logic; attribute dont_touch of G12317: signal is true;
	signal G12318: std_logic; attribute dont_touch of G12318: signal is true;
	signal G12321: std_logic; attribute dont_touch of G12321: signal is true;
	signal G12322: std_logic; attribute dont_touch of G12322: signal is true;
	signal G12323: std_logic; attribute dont_touch of G12323: signal is true;
	signal G12332: std_logic; attribute dont_touch of G12332: signal is true;
	signal G12333: std_logic; attribute dont_touch of G12333: signal is true;
	signal G12336: std_logic; attribute dont_touch of G12336: signal is true;
	signal G12337: std_logic; attribute dont_touch of G12337: signal is true;
	signal G12340: std_logic; attribute dont_touch of G12340: signal is true;
	signal G12341: std_logic; attribute dont_touch of G12341: signal is true;
	signal G12342: std_logic; attribute dont_touch of G12342: signal is true;
	signal G12343: std_logic; attribute dont_touch of G12343: signal is true;
	signal G12344: std_logic; attribute dont_touch of G12344: signal is true;
	signal G12345: std_logic; attribute dont_touch of G12345: signal is true;
	signal G12346: std_logic; attribute dont_touch of G12346: signal is true;
	signal G12347: std_logic; attribute dont_touch of G12347: signal is true;
	signal G12351: std_logic; attribute dont_touch of G12351: signal is true;
	signal G12356: std_logic; attribute dont_touch of G12356: signal is true;
	signal G12357: std_logic; attribute dont_touch of G12357: signal is true;
	signal G12358: std_logic; attribute dont_touch of G12358: signal is true;
	signal G12361: std_logic; attribute dont_touch of G12361: signal is true;
	signal G12364: std_logic; attribute dont_touch of G12364: signal is true;
	signal G12367: std_logic; attribute dont_touch of G12367: signal is true;
	signal G12369: std_logic; attribute dont_touch of G12369: signal is true;
	signal G12370: std_logic; attribute dont_touch of G12370: signal is true;
	signal G12371: std_logic; attribute dont_touch of G12371: signal is true;
	signal G12374: std_logic; attribute dont_touch of G12374: signal is true;
	signal G12377: std_logic; attribute dont_touch of G12377: signal is true;
	signal G12378: std_logic; attribute dont_touch of G12378: signal is true;
	signal G12381: std_logic; attribute dont_touch of G12381: signal is true;
	signal G12399: std_logic; attribute dont_touch of G12399: signal is true;
	signal G12402: std_logic; attribute dont_touch of G12402: signal is true;
	signal G12405: std_logic; attribute dont_touch of G12405: signal is true;
	signal G12411: std_logic; attribute dont_touch of G12411: signal is true;
	signal G12412: std_logic; attribute dont_touch of G12412: signal is true;
	signal G12413: std_logic; attribute dont_touch of G12413: signal is true;
	signal G12414: std_logic; attribute dont_touch of G12414: signal is true;
	signal G12415: std_logic; attribute dont_touch of G12415: signal is true;
	signal G12416: std_logic; attribute dont_touch of G12416: signal is true;
	signal G12417: std_logic; attribute dont_touch of G12417: signal is true;
	signal G12418: std_logic; attribute dont_touch of G12418: signal is true;
	signal G12419: std_logic; attribute dont_touch of G12419: signal is true;
	signal G12423: std_logic; attribute dont_touch of G12423: signal is true;
	signal G12428: std_logic; attribute dont_touch of G12428: signal is true;
	signal G12429: std_logic; attribute dont_touch of G12429: signal is true;
	signal G12430: std_logic; attribute dont_touch of G12430: signal is true;
	signal G12431: std_logic; attribute dont_touch of G12431: signal is true;
	signal G12432: std_logic; attribute dont_touch of G12432: signal is true;
	signal G12435: std_logic; attribute dont_touch of G12435: signal is true;
	signal G12436: std_logic; attribute dont_touch of G12436: signal is true;
	signal G12437: std_logic; attribute dont_touch of G12437: signal is true;
	signal G12440: std_logic; attribute dont_touch of G12440: signal is true;
	signal G12443: std_logic; attribute dont_touch of G12443: signal is true;
	signal G12449: std_logic; attribute dont_touch of G12449: signal is true;
	signal G12450: std_logic; attribute dont_touch of G12450: signal is true;
	signal G12453: std_logic; attribute dont_touch of G12453: signal is true;
	signal G12459: std_logic; attribute dont_touch of G12459: signal is true;
	signal G12460: std_logic; attribute dont_touch of G12460: signal is true;
	signal G12461: std_logic; attribute dont_touch of G12461: signal is true;
	signal G12462: std_logic; attribute dont_touch of G12462: signal is true;
	signal G12463: std_logic; attribute dont_touch of G12463: signal is true;
	signal G12464: std_logic; attribute dont_touch of G12464: signal is true;
	signal G12465: std_logic; attribute dont_touch of G12465: signal is true;
	signal G12466: std_logic; attribute dont_touch of G12466: signal is true;
	signal G12467: std_logic; attribute dont_touch of G12467: signal is true;
	signal G12471: std_logic; attribute dont_touch of G12471: signal is true;
	signal G12476: std_logic; attribute dont_touch of G12476: signal is true;
	signal G12477: std_logic; attribute dont_touch of G12477: signal is true;
	signal G12478: std_logic; attribute dont_touch of G12478: signal is true;
	signal G12479: std_logic; attribute dont_touch of G12479: signal is true;
	signal G12482: std_logic; attribute dont_touch of G12482: signal is true;
	signal G12483: std_logic; attribute dont_touch of G12483: signal is true;
	signal G12486: std_logic; attribute dont_touch of G12486: signal is true;
	signal G12487: std_logic; attribute dont_touch of G12487: signal is true;
	signal G12490: std_logic; attribute dont_touch of G12490: signal is true;
	signal G12491: std_logic; attribute dont_touch of G12491: signal is true;
	signal G12492: std_logic; attribute dont_touch of G12492: signal is true;
	signal G12497: std_logic; attribute dont_touch of G12497: signal is true;
	signal G12505: std_logic; attribute dont_touch of G12505: signal is true;
	signal G12511: std_logic; attribute dont_touch of G12511: signal is true;
	signal G12512: std_logic; attribute dont_touch of G12512: signal is true;
	signal G12515: std_logic; attribute dont_touch of G12515: signal is true;
	signal G12521: std_logic; attribute dont_touch of G12521: signal is true;
	signal G12522: std_logic; attribute dont_touch of G12522: signal is true;
	signal G12523: std_logic; attribute dont_touch of G12523: signal is true;
	signal G12524: std_logic; attribute dont_touch of G12524: signal is true;
	signal G12525: std_logic; attribute dont_touch of G12525: signal is true;
	signal G12526: std_logic; attribute dont_touch of G12526: signal is true;
	signal G12527: std_logic; attribute dont_touch of G12527: signal is true;
	signal G12538: std_logic; attribute dont_touch of G12538: signal is true;
	signal G12539: std_logic; attribute dont_touch of G12539: signal is true;
	signal G12540: std_logic; attribute dont_touch of G12540: signal is true;
	signal G12543: std_logic; attribute dont_touch of G12543: signal is true;
	signal G12546: std_logic; attribute dont_touch of G12546: signal is true;
	signal G12550: std_logic; attribute dont_touch of G12550: signal is true;
	signal G12553: std_logic; attribute dont_touch of G12553: signal is true;
	signal G12558: std_logic; attribute dont_touch of G12558: signal is true;
	signal G12563: std_logic; attribute dont_touch of G12563: signal is true;
	signal G12571: std_logic; attribute dont_touch of G12571: signal is true;
	signal G12577: std_logic; attribute dont_touch of G12577: signal is true;
	signal G12578: std_logic; attribute dont_touch of G12578: signal is true;
	signal G12581: std_logic; attribute dont_touch of G12581: signal is true;
	signal G12587: std_logic; attribute dont_touch of G12587: signal is true;
	signal G12588: std_logic; attribute dont_touch of G12588: signal is true;
	signal G12589: std_logic; attribute dont_touch of G12589: signal is true;
	signal G12590: std_logic; attribute dont_touch of G12590: signal is true;
	signal G12591: std_logic; attribute dont_touch of G12591: signal is true;
	signal G12592: std_logic; attribute dont_touch of G12592: signal is true;
	signal G12593: std_logic; attribute dont_touch of G12593: signal is true;
	signal G12598: std_logic; attribute dont_touch of G12598: signal is true;
	signal G12601: std_logic; attribute dont_touch of G12601: signal is true;
	signal G12604: std_logic; attribute dont_touch of G12604: signal is true;
	signal G12609: std_logic; attribute dont_touch of G12609: signal is true;
	signal G12614: std_logic; attribute dont_touch of G12614: signal is true;
	signal G12622: std_logic; attribute dont_touch of G12622: signal is true;
	signal G12628: std_logic; attribute dont_touch of G12628: signal is true;
	signal G12629: std_logic; attribute dont_touch of G12629: signal is true;
	signal G12632: std_logic; attribute dont_touch of G12632: signal is true;
	signal G12638: std_logic; attribute dont_touch of G12638: signal is true;
	signal G12639: std_logic; attribute dont_touch of G12639: signal is true;
	signal G12640: std_logic; attribute dont_touch of G12640: signal is true;
	signal G12641: std_logic; attribute dont_touch of G12641: signal is true;
	signal G12644: std_logic; attribute dont_touch of G12644: signal is true;
	signal G12645: std_logic; attribute dont_touch of G12645: signal is true;
	signal G12646: std_logic; attribute dont_touch of G12646: signal is true;
	signal G12651: std_logic; attribute dont_touch of G12651: signal is true;
	signal G12656: std_logic; attribute dont_touch of G12656: signal is true;
	signal G12659: std_logic; attribute dont_touch of G12659: signal is true;
	signal G12662: std_logic; attribute dont_touch of G12662: signal is true;
	signal G12667: std_logic; attribute dont_touch of G12667: signal is true;
	signal G12672: std_logic; attribute dont_touch of G12672: signal is true;
	signal G12680: std_logic; attribute dont_touch of G12680: signal is true;
	signal G12686: std_logic; attribute dont_touch of G12686: signal is true;
	signal G12687: std_logic; attribute dont_touch of G12687: signal is true;
	signal G12692: std_logic; attribute dont_touch of G12692: signal is true;
	signal G12695: std_logic; attribute dont_touch of G12695: signal is true;
	signal G12700: std_logic; attribute dont_touch of G12700: signal is true;
	signal G12705: std_logic; attribute dont_touch of G12705: signal is true;
	signal G12708: std_logic; attribute dont_touch of G12708: signal is true;
	signal G12711: std_logic; attribute dont_touch of G12711: signal is true;
	signal G12716: std_logic; attribute dont_touch of G12716: signal is true;
	signal G12721: std_logic; attribute dont_touch of G12721: signal is true;
	signal G12729: std_logic; attribute dont_touch of G12729: signal is true;
	signal G12730: std_logic; attribute dont_touch of G12730: signal is true;
	signal G12735: std_logic; attribute dont_touch of G12735: signal is true;
	signal G12738: std_logic; attribute dont_touch of G12738: signal is true;
	signal G12739: std_logic; attribute dont_touch of G12739: signal is true;
	signal G12744: std_logic; attribute dont_touch of G12744: signal is true;
	signal G12749: std_logic; attribute dont_touch of G12749: signal is true;
	signal G12752: std_logic; attribute dont_touch of G12752: signal is true;
	signal G12755: std_logic; attribute dont_touch of G12755: signal is true;
	signal G12760: std_logic; attribute dont_touch of G12760: signal is true;
	signal G12761: std_logic; attribute dont_touch of G12761: signal is true;
	signal G12762: std_logic; attribute dont_touch of G12762: signal is true;
	signal G12767: std_logic; attribute dont_touch of G12767: signal is true;
	signal G12768: std_logic; attribute dont_touch of G12768: signal is true;
	signal G12772: std_logic; attribute dont_touch of G12772: signal is true;
	signal G12778: std_logic; attribute dont_touch of G12778: signal is true;
	signal G12779: std_logic; attribute dont_touch of G12779: signal is true;
	signal G12780: std_logic; attribute dont_touch of G12780: signal is true;
	signal G12785: std_logic; attribute dont_touch of G12785: signal is true;
	signal G12790: std_logic; attribute dont_touch of G12790: signal is true;
	signal G12793: std_logic; attribute dont_touch of G12793: signal is true;
	signal G12794: std_logic; attribute dont_touch of G12794: signal is true;
	signal G12795: std_logic; attribute dont_touch of G12795: signal is true;
	signal G12796: std_logic; attribute dont_touch of G12796: signal is true;
	signal G12797: std_logic; attribute dont_touch of G12797: signal is true;
	signal G12798: std_logic; attribute dont_touch of G12798: signal is true;
	signal G12804: std_logic; attribute dont_touch of G12804: signal is true;
	signal G12805: std_logic; attribute dont_touch of G12805: signal is true;
	signal G12806: std_logic; attribute dont_touch of G12806: signal is true;
	signal G12811: std_logic; attribute dont_touch of G12811: signal is true;
	signal G12812: std_logic; attribute dont_touch of G12812: signal is true;
	signal G12817: std_logic; attribute dont_touch of G12817: signal is true;
	signal G12818: std_logic; attribute dont_touch of G12818: signal is true;
	signal G12819: std_logic; attribute dont_touch of G12819: signal is true;
	signal G12820: std_logic; attribute dont_touch of G12820: signal is true;
	signal G12821: std_logic; attribute dont_touch of G12821: signal is true;
	signal G12822: std_logic; attribute dont_touch of G12822: signal is true;
	signal G12823: std_logic; attribute dont_touch of G12823: signal is true;
	signal G12824: std_logic; attribute dont_touch of G12824: signal is true;
	signal G12830: std_logic; attribute dont_touch of G12830: signal is true;
	signal G12831: std_logic; attribute dont_touch of G12831: signal is true;
	signal G12834: std_logic; attribute dont_touch of G12834: signal is true;
	signal G12835: std_logic; attribute dont_touch of G12835: signal is true;
	signal G12836: std_logic; attribute dont_touch of G12836: signal is true;
	signal G12837: std_logic; attribute dont_touch of G12837: signal is true;
	signal G12838: std_logic; attribute dont_touch of G12838: signal is true;
	signal G12839: std_logic; attribute dont_touch of G12839: signal is true;
	signal G12840: std_logic; attribute dont_touch of G12840: signal is true;
	signal G12841: std_logic; attribute dont_touch of G12841: signal is true;
	signal G12842: std_logic; attribute dont_touch of G12842: signal is true;
	signal G12843: std_logic; attribute dont_touch of G12843: signal is true;
	signal G12844: std_logic; attribute dont_touch of G12844: signal is true;
	signal G12845: std_logic; attribute dont_touch of G12845: signal is true;
	signal G12846: std_logic; attribute dont_touch of G12846: signal is true;
	signal G12847: std_logic; attribute dont_touch of G12847: signal is true;
	signal G12848: std_logic; attribute dont_touch of G12848: signal is true;
	signal G12849: std_logic; attribute dont_touch of G12849: signal is true;
	signal G12850: std_logic; attribute dont_touch of G12850: signal is true;
	signal G12851: std_logic; attribute dont_touch of G12851: signal is true;
	signal G12852: std_logic; attribute dont_touch of G12852: signal is true;
	signal G12853: std_logic; attribute dont_touch of G12853: signal is true;
	signal G12854: std_logic; attribute dont_touch of G12854: signal is true;
	signal G12855: std_logic; attribute dont_touch of G12855: signal is true;
	signal G12856: std_logic; attribute dont_touch of G12856: signal is true;
	signal G12857: std_logic; attribute dont_touch of G12857: signal is true;
	signal G12858: std_logic; attribute dont_touch of G12858: signal is true;
	signal G12859: std_logic; attribute dont_touch of G12859: signal is true;
	signal G12860: std_logic; attribute dont_touch of G12860: signal is true;
	signal G12861: std_logic; attribute dont_touch of G12861: signal is true;
	signal G12862: std_logic; attribute dont_touch of G12862: signal is true;
	signal G12863: std_logic; attribute dont_touch of G12863: signal is true;
	signal G12864: std_logic; attribute dont_touch of G12864: signal is true;
	signal G12865: std_logic; attribute dont_touch of G12865: signal is true;
	signal G12866: std_logic; attribute dont_touch of G12866: signal is true;
	signal G12867: std_logic; attribute dont_touch of G12867: signal is true;
	signal G12868: std_logic; attribute dont_touch of G12868: signal is true;
	signal G12869: std_logic; attribute dont_touch of G12869: signal is true;
	signal G12870: std_logic; attribute dont_touch of G12870: signal is true;
	signal G12871: std_logic; attribute dont_touch of G12871: signal is true;
	signal G12872: std_logic; attribute dont_touch of G12872: signal is true;
	signal G12873: std_logic; attribute dont_touch of G12873: signal is true;
	signal G12874: std_logic; attribute dont_touch of G12874: signal is true;
	signal G12875: std_logic; attribute dont_touch of G12875: signal is true;
	signal G12878: std_logic; attribute dont_touch of G12878: signal is true;
	signal G12879: std_logic; attribute dont_touch of G12879: signal is true;
	signal G12880: std_logic; attribute dont_touch of G12880: signal is true;
	signal G12881: std_logic; attribute dont_touch of G12881: signal is true;
	signal G12882: std_logic; attribute dont_touch of G12882: signal is true;
	signal G12883: std_logic; attribute dont_touch of G12883: signal is true;
	signal G12884: std_logic; attribute dont_touch of G12884: signal is true;
	signal G12885: std_logic; attribute dont_touch of G12885: signal is true;
	signal G12886: std_logic; attribute dont_touch of G12886: signal is true;
	signal G12887: std_logic; attribute dont_touch of G12887: signal is true;
	signal G12888: std_logic; attribute dont_touch of G12888: signal is true;
	signal G12889: std_logic; attribute dont_touch of G12889: signal is true;
	signal G12890: std_logic; attribute dont_touch of G12890: signal is true;
	signal G12891: std_logic; attribute dont_touch of G12891: signal is true;
	signal G12892: std_logic; attribute dont_touch of G12892: signal is true;
	signal G12893: std_logic; attribute dont_touch of G12893: signal is true;
	signal G12894: std_logic; attribute dont_touch of G12894: signal is true;
	signal G12895: std_logic; attribute dont_touch of G12895: signal is true;
	signal G12896: std_logic; attribute dont_touch of G12896: signal is true;
	signal G12897: std_logic; attribute dont_touch of G12897: signal is true;
	signal G12898: std_logic; attribute dont_touch of G12898: signal is true;
	signal G12899: std_logic; attribute dont_touch of G12899: signal is true;
	signal G12900: std_logic; attribute dont_touch of G12900: signal is true;
	signal G12901: std_logic; attribute dont_touch of G12901: signal is true;
	signal G12902: std_logic; attribute dont_touch of G12902: signal is true;
	signal G12903: std_logic; attribute dont_touch of G12903: signal is true;
	signal G12904: std_logic; attribute dont_touch of G12904: signal is true;
	signal G12905: std_logic; attribute dont_touch of G12905: signal is true;
	signal G12906: std_logic; attribute dont_touch of G12906: signal is true;
	signal G12907: std_logic; attribute dont_touch of G12907: signal is true;
	signal G12908: std_logic; attribute dont_touch of G12908: signal is true;
	signal G12909: std_logic; attribute dont_touch of G12909: signal is true;
	signal G12910: std_logic; attribute dont_touch of G12910: signal is true;
	signal G12911: std_logic; attribute dont_touch of G12911: signal is true;
	signal G12914: std_logic; attribute dont_touch of G12914: signal is true;
	signal G12915: std_logic; attribute dont_touch of G12915: signal is true;
	signal G12918: std_logic; attribute dont_touch of G12918: signal is true;
	signal G12920: std_logic; attribute dont_touch of G12920: signal is true;
	signal G12921: std_logic; attribute dont_touch of G12921: signal is true;
	signal G12922: std_logic; attribute dont_touch of G12922: signal is true;
	signal G12924: std_logic; attribute dont_touch of G12924: signal is true;
	signal G12925: std_logic; attribute dont_touch of G12925: signal is true;
	signal G12929: std_logic; attribute dont_touch of G12929: signal is true;
	signal G12930: std_logic; attribute dont_touch of G12930: signal is true;
	signal G12931: std_logic; attribute dont_touch of G12931: signal is true;
	signal G12932: std_logic; attribute dont_touch of G12932: signal is true;
	signal G12933: std_logic; attribute dont_touch of G12933: signal is true;
	signal G12936: std_logic; attribute dont_touch of G12936: signal is true;
	signal G12937: std_logic; attribute dont_touch of G12937: signal is true;
	signal G12938: std_logic; attribute dont_touch of G12938: signal is true;
	signal G12939: std_logic; attribute dont_touch of G12939: signal is true;
	signal G12940: std_logic; attribute dont_touch of G12940: signal is true;
	signal G12941: std_logic; attribute dont_touch of G12941: signal is true;
	signal G12944: std_logic; attribute dont_touch of G12944: signal is true;
	signal G12945: std_logic; attribute dont_touch of G12945: signal is true;
	signal G12946: std_logic; attribute dont_touch of G12946: signal is true;
	signal G12947: std_logic; attribute dont_touch of G12947: signal is true;
	signal G12950: std_logic; attribute dont_touch of G12950: signal is true;
	signal G12951: std_logic; attribute dont_touch of G12951: signal is true;
	signal G12952: std_logic; attribute dont_touch of G12952: signal is true;
	signal G12953: std_logic; attribute dont_touch of G12953: signal is true;
	signal G12954: std_logic; attribute dont_touch of G12954: signal is true;
	signal G12955: std_logic; attribute dont_touch of G12955: signal is true;
	signal G12967: std_logic; attribute dont_touch of G12967: signal is true;
	signal G12968: std_logic; attribute dont_touch of G12968: signal is true;
	signal G12969: std_logic; attribute dont_touch of G12969: signal is true;
	signal G12970: std_logic; attribute dont_touch of G12970: signal is true;
	signal G12971: std_logic; attribute dont_touch of G12971: signal is true;
	signal G12972: std_logic; attribute dont_touch of G12972: signal is true;
	signal G12975: std_logic; attribute dont_touch of G12975: signal is true;
	signal G12976: std_logic; attribute dont_touch of G12976: signal is true;
	signal G12977: std_logic; attribute dont_touch of G12977: signal is true;
	signal G12978: std_logic; attribute dont_touch of G12978: signal is true;
	signal G12979: std_logic; attribute dont_touch of G12979: signal is true;
	signal G12980: std_logic; attribute dont_touch of G12980: signal is true;
	signal G12981: std_logic; attribute dont_touch of G12981: signal is true;
	signal G12982: std_logic; attribute dont_touch of G12982: signal is true;
	signal G12983: std_logic; attribute dont_touch of G12983: signal is true;
	signal G12995: std_logic; attribute dont_touch of G12995: signal is true;
	signal G12996: std_logic; attribute dont_touch of G12996: signal is true;
	signal G12997: std_logic; attribute dont_touch of G12997: signal is true;
	signal G12998: std_logic; attribute dont_touch of G12998: signal is true;
	signal G12999: std_logic; attribute dont_touch of G12999: signal is true;
	signal G13000: std_logic; attribute dont_touch of G13000: signal is true;
	signal G13003: std_logic; attribute dont_touch of G13003: signal is true;
	signal G13004: std_logic; attribute dont_touch of G13004: signal is true;
	signal G13005: std_logic; attribute dont_touch of G13005: signal is true;
	signal G13006: std_logic; attribute dont_touch of G13006: signal is true;
	signal G13007: std_logic; attribute dont_touch of G13007: signal is true;
	signal G13008: std_logic; attribute dont_touch of G13008: signal is true;
	signal G13009: std_logic; attribute dont_touch of G13009: signal is true;
	signal G13010: std_logic; attribute dont_touch of G13010: signal is true;
	signal G13011: std_logic; attribute dont_touch of G13011: signal is true;
	signal G13012: std_logic; attribute dont_touch of G13012: signal is true;
	signal G13013: std_logic; attribute dont_touch of G13013: signal is true;
	signal G13014: std_logic; attribute dont_touch of G13014: signal is true;
	signal G13015: std_logic; attribute dont_touch of G13015: signal is true;
	signal G13016: std_logic; attribute dont_touch of G13016: signal is true;
	signal G13017: std_logic; attribute dont_touch of G13017: signal is true;
	signal G13018: std_logic; attribute dont_touch of G13018: signal is true;
	signal G13019: std_logic; attribute dont_touch of G13019: signal is true;
	signal G13020: std_logic; attribute dont_touch of G13020: signal is true;
	signal G13021: std_logic; attribute dont_touch of G13021: signal is true;
	signal G13022: std_logic; attribute dont_touch of G13022: signal is true;
	signal G13023: std_logic; attribute dont_touch of G13023: signal is true;
	signal G13024: std_logic; attribute dont_touch of G13024: signal is true;
	signal G13025: std_logic; attribute dont_touch of G13025: signal is true;
	signal G13026: std_logic; attribute dont_touch of G13026: signal is true;
	signal G13027: std_logic; attribute dont_touch of G13027: signal is true;
	signal G13028: std_logic; attribute dont_touch of G13028: signal is true;
	signal G13029: std_logic; attribute dont_touch of G13029: signal is true;
	signal G13030: std_logic; attribute dont_touch of G13030: signal is true;
	signal G13031: std_logic; attribute dont_touch of G13031: signal is true;
	signal G13032: std_logic; attribute dont_touch of G13032: signal is true;
	signal G13033: std_logic; attribute dont_touch of G13033: signal is true;
	signal G13034: std_logic; attribute dont_touch of G13034: signal is true;
	signal G13035: std_logic; attribute dont_touch of G13035: signal is true;
	signal G13036: std_logic; attribute dont_touch of G13036: signal is true;
	signal G13037: std_logic; attribute dont_touch of G13037: signal is true;
	signal G13038: std_logic; attribute dont_touch of G13038: signal is true;
	signal G13040: std_logic; attribute dont_touch of G13040: signal is true;
	signal G13041: std_logic; attribute dont_touch of G13041: signal is true;
	signal G13042: std_logic; attribute dont_touch of G13042: signal is true;
	signal G13043: std_logic; attribute dont_touch of G13043: signal is true;
	signal G13044: std_logic; attribute dont_touch of G13044: signal is true;
	signal G13045: std_logic; attribute dont_touch of G13045: signal is true;
	signal G13046: std_logic; attribute dont_touch of G13046: signal is true;
	signal G13047: std_logic; attribute dont_touch of G13047: signal is true;
	signal G13048: std_logic; attribute dont_touch of G13048: signal is true;
	signal G13050: std_logic; attribute dont_touch of G13050: signal is true;
	signal G13051: std_logic; attribute dont_touch of G13051: signal is true;
	signal G13055: std_logic; attribute dont_touch of G13055: signal is true;
	signal G13056: std_logic; attribute dont_touch of G13056: signal is true;
	signal G13057: std_logic; attribute dont_touch of G13057: signal is true;
	signal G13058: std_logic; attribute dont_touch of G13058: signal is true;
	signal G13059: std_logic; attribute dont_touch of G13059: signal is true;
	signal G13060: std_logic; attribute dont_touch of G13060: signal is true;
	signal G13061: std_logic; attribute dont_touch of G13061: signal is true;
	signal G13062: std_logic; attribute dont_touch of G13062: signal is true;
	signal G13063: std_logic; attribute dont_touch of G13063: signal is true;
	signal G13064: std_logic; attribute dont_touch of G13064: signal is true;
	signal G13065: std_logic; attribute dont_touch of G13065: signal is true;
	signal G13066: std_logic; attribute dont_touch of G13066: signal is true;
	signal G13067: std_logic; attribute dont_touch of G13067: signal is true;
	signal G13069: std_logic; attribute dont_touch of G13069: signal is true;
	signal G13070: std_logic; attribute dont_touch of G13070: signal is true;
	signal G13074: std_logic; attribute dont_touch of G13074: signal is true;
	signal G13075: std_logic; attribute dont_touch of G13075: signal is true;
	signal G13076: std_logic; attribute dont_touch of G13076: signal is true;
	signal G13077: std_logic; attribute dont_touch of G13077: signal is true;
	signal G13078: std_logic; attribute dont_touch of G13078: signal is true;
	signal G13079: std_logic; attribute dont_touch of G13079: signal is true;
	signal G13080: std_logic; attribute dont_touch of G13080: signal is true;
	signal G13081: std_logic; attribute dont_touch of G13081: signal is true;
	signal G13082: std_logic; attribute dont_touch of G13082: signal is true;
	signal G13083: std_logic; attribute dont_touch of G13083: signal is true;
	signal G13084: std_logic; attribute dont_touch of G13084: signal is true;
	signal G13086: std_logic; attribute dont_touch of G13086: signal is true;
	signal G13087: std_logic; attribute dont_touch of G13087: signal is true;
	signal G13091: std_logic; attribute dont_touch of G13091: signal is true;
	signal G13092: std_logic; attribute dont_touch of G13092: signal is true;
	signal G13093: std_logic; attribute dont_touch of G13093: signal is true;
	signal G13094: std_logic; attribute dont_touch of G13094: signal is true;
	signal G13095: std_logic; attribute dont_touch of G13095: signal is true;
	signal G13096: std_logic; attribute dont_touch of G13096: signal is true;
	signal G13097: std_logic; attribute dont_touch of G13097: signal is true;
	signal G13098: std_logic; attribute dont_touch of G13098: signal is true;
	signal G13100: std_logic; attribute dont_touch of G13100: signal is true;
	signal G13101: std_logic; attribute dont_touch of G13101: signal is true;
	signal G13102: std_logic; attribute dont_touch of G13102: signal is true;
	signal G13103: std_logic; attribute dont_touch of G13103: signal is true;
	signal G13104: std_logic; attribute dont_touch of G13104: signal is true;
	signal G13105: std_logic; attribute dont_touch of G13105: signal is true;
	signal G13106: std_logic; attribute dont_touch of G13106: signal is true;
	signal G13107: std_logic; attribute dont_touch of G13107: signal is true;
	signal G13108: std_logic; attribute dont_touch of G13108: signal is true;
	signal G13109: std_logic; attribute dont_touch of G13109: signal is true;
	signal G13110: std_logic; attribute dont_touch of G13110: signal is true;
	signal G13114: std_logic; attribute dont_touch of G13114: signal is true;
	signal G13115: std_logic; attribute dont_touch of G13115: signal is true;
	signal G13116: std_logic; attribute dont_touch of G13116: signal is true;
	signal G13117: std_logic; attribute dont_touch of G13117: signal is true;
	signal G13118: std_logic; attribute dont_touch of G13118: signal is true;
	signal G13119: std_logic; attribute dont_touch of G13119: signal is true;
	signal G13120: std_logic; attribute dont_touch of G13120: signal is true;
	signal G13121: std_logic; attribute dont_touch of G13121: signal is true;
	signal G13124: std_logic; attribute dont_touch of G13124: signal is true;
	signal G13125: std_logic; attribute dont_touch of G13125: signal is true;
	signal G13129: std_logic; attribute dont_touch of G13129: signal is true;
	signal G13130: std_logic; attribute dont_touch of G13130: signal is true;
	signal G13131: std_logic; attribute dont_touch of G13131: signal is true;
	signal G13132: std_logic; attribute dont_touch of G13132: signal is true;
	signal G13133: std_logic; attribute dont_touch of G13133: signal is true;
	signal G13134: std_logic; attribute dont_touch of G13134: signal is true;
	signal G13137: std_logic; attribute dont_touch of G13137: signal is true;
	signal G13138: std_logic; attribute dont_touch of G13138: signal is true;
	signal G13139: std_logic; attribute dont_touch of G13139: signal is true;
	signal G13140: std_logic; attribute dont_touch of G13140: signal is true;
	signal G13141: std_logic; attribute dont_touch of G13141: signal is true;
	signal G13142: std_logic; attribute dont_touch of G13142: signal is true;
	signal G13143: std_logic; attribute dont_touch of G13143: signal is true;
	signal G13144: std_logic; attribute dont_touch of G13144: signal is true;
	signal G13155: std_logic; attribute dont_touch of G13155: signal is true;
	signal G13156: std_logic; attribute dont_touch of G13156: signal is true;
	signal G13173: std_logic; attribute dont_touch of G13173: signal is true;
	signal G13174: std_logic; attribute dont_touch of G13174: signal is true;
	signal G13175: std_logic; attribute dont_touch of G13175: signal is true;
	signal G13176: std_logic; attribute dont_touch of G13176: signal is true;
	signal G13177: std_logic; attribute dont_touch of G13177: signal is true;
	signal G13188: std_logic; attribute dont_touch of G13188: signal is true;
	signal G13189: std_logic; attribute dont_touch of G13189: signal is true;
	signal G13190: std_logic; attribute dont_touch of G13190: signal is true;
	signal G13191: std_logic; attribute dont_touch of G13191: signal is true;
	signal G13202: std_logic; attribute dont_touch of G13202: signal is true;
	signal G13209: std_logic; attribute dont_touch of G13209: signal is true;
	signal G13210: std_logic; attribute dont_touch of G13210: signal is true;
	signal G13211: std_logic; attribute dont_touch of G13211: signal is true;
	signal G13215: std_logic; attribute dont_touch of G13215: signal is true;
	signal G13216: std_logic; attribute dont_touch of G13216: signal is true;
	signal G13217: std_logic; attribute dont_touch of G13217: signal is true;
	signal G13221: std_logic; attribute dont_touch of G13221: signal is true;
	signal G13222: std_logic; attribute dont_touch of G13222: signal is true;
	signal G13223: std_logic; attribute dont_touch of G13223: signal is true;
	signal G13239: std_logic; attribute dont_touch of G13239: signal is true;
	signal G13240: std_logic; attribute dont_touch of G13240: signal is true;
	signal G13241: std_logic; attribute dont_touch of G13241: signal is true;
	signal G13242: std_logic; attribute dont_touch of G13242: signal is true;
	signal G13246: std_logic; attribute dont_touch of G13246: signal is true;
	signal G13247: std_logic; attribute dont_touch of G13247: signal is true;
	signal G13248: std_logic; attribute dont_touch of G13248: signal is true;
	signal G13249: std_logic; attribute dont_touch of G13249: signal is true;
	signal G13250: std_logic; attribute dont_touch of G13250: signal is true;
	signal G13251: std_logic; attribute dont_touch of G13251: signal is true;
	signal G13252: std_logic; attribute dont_touch of G13252: signal is true;
	signal G13255: std_logic; attribute dont_touch of G13255: signal is true;
	signal G13256: std_logic; attribute dont_touch of G13256: signal is true;
	signal G13257: std_logic; attribute dont_touch of G13257: signal is true;
	signal G13258: std_logic; attribute dont_touch of G13258: signal is true;
	signal G13260: std_logic; attribute dont_touch of G13260: signal is true;
	signal G13264: std_logic; attribute dont_touch of G13264: signal is true;
	signal G13265: std_logic; attribute dont_touch of G13265: signal is true;
	signal G13266: std_logic; attribute dont_touch of G13266: signal is true;
	signal G13267: std_logic; attribute dont_touch of G13267: signal is true;
	signal G13271: std_logic; attribute dont_touch of G13271: signal is true;
	signal G13273: std_logic; attribute dont_touch of G13273: signal is true;
	signal G13277: std_logic; attribute dont_touch of G13277: signal is true;
	signal G13278: std_logic; attribute dont_touch of G13278: signal is true;
	signal G13279: std_logic; attribute dont_touch of G13279: signal is true;
	signal G13280: std_logic; attribute dont_touch of G13280: signal is true;
	signal G13281: std_logic; attribute dont_touch of G13281: signal is true;
	signal G13282: std_logic; attribute dont_touch of G13282: signal is true;
	signal G13283: std_logic; attribute dont_touch of G13283: signal is true;
	signal G13284: std_logic; attribute dont_touch of G13284: signal is true;
	signal G13287: std_logic; attribute dont_touch of G13287: signal is true;
	signal G13288: std_logic; attribute dont_touch of G13288: signal is true;
	signal G13289: std_logic; attribute dont_touch of G13289: signal is true;
	signal G13290: std_logic; attribute dont_touch of G13290: signal is true;
	signal G13291: std_logic; attribute dont_touch of G13291: signal is true;
	signal G13294: std_logic; attribute dont_touch of G13294: signal is true;
	signal G13295: std_logic; attribute dont_touch of G13295: signal is true;
	signal G13296: std_logic; attribute dont_touch of G13296: signal is true;
	signal G13297: std_logic; attribute dont_touch of G13297: signal is true;
	signal G13298: std_logic; attribute dont_touch of G13298: signal is true;
	signal G13299: std_logic; attribute dont_touch of G13299: signal is true;
	signal G13300: std_logic; attribute dont_touch of G13300: signal is true;
	signal G13301: std_logic; attribute dont_touch of G13301: signal is true;
	signal G13302: std_logic; attribute dont_touch of G13302: signal is true;
	signal G13303: std_logic; attribute dont_touch of G13303: signal is true;
	signal G13304: std_logic; attribute dont_touch of G13304: signal is true;
	signal G13305: std_logic; attribute dont_touch of G13305: signal is true;
	signal G13306: std_logic; attribute dont_touch of G13306: signal is true;
	signal G13307: std_logic; attribute dont_touch of G13307: signal is true;
	signal G13311: std_logic; attribute dont_touch of G13311: signal is true;
	signal G13312: std_logic; attribute dont_touch of G13312: signal is true;
	signal G13313: std_logic; attribute dont_touch of G13313: signal is true;
	signal G13314: std_logic; attribute dont_touch of G13314: signal is true;
	signal G13315: std_logic; attribute dont_touch of G13315: signal is true;
	signal G13319: std_logic; attribute dont_touch of G13319: signal is true;
	signal G13320: std_logic; attribute dont_touch of G13320: signal is true;
	signal G13321: std_logic; attribute dont_touch of G13321: signal is true;
	signal G13322: std_logic; attribute dont_touch of G13322: signal is true;
	signal G13323: std_logic; attribute dont_touch of G13323: signal is true;
	signal G13324: std_logic; attribute dont_touch of G13324: signal is true;
	signal G13325: std_logic; attribute dont_touch of G13325: signal is true;
	signal G13326: std_logic; attribute dont_touch of G13326: signal is true;
	signal G13329: std_logic; attribute dont_touch of G13329: signal is true;
	signal G13330: std_logic; attribute dont_touch of G13330: signal is true;
	signal G13333: std_logic; attribute dont_touch of G13333: signal is true;
	signal G13334: std_logic; attribute dont_touch of G13334: signal is true;
	signal G13335: std_logic; attribute dont_touch of G13335: signal is true;
	signal G13336: std_logic; attribute dont_touch of G13336: signal is true;
	signal G13341: std_logic; attribute dont_touch of G13341: signal is true;
	signal G13342: std_logic; attribute dont_touch of G13342: signal is true;
	signal G13345: std_logic; attribute dont_touch of G13345: signal is true;
	signal G13346: std_logic; attribute dont_touch of G13346: signal is true;
	signal G13349: std_logic; attribute dont_touch of G13349: signal is true;
	signal G13350: std_logic; attribute dont_touch of G13350: signal is true;
	signal G13377: std_logic; attribute dont_touch of G13377: signal is true;
	signal G13378: std_logic; attribute dont_touch of G13378: signal is true;
	signal G13383: std_logic; attribute dont_touch of G13383: signal is true;
	signal G13384: std_logic; attribute dont_touch of G13384: signal is true;
	signal G13385: std_logic; attribute dont_touch of G13385: signal is true;
	signal G13393: std_logic; attribute dont_touch of G13393: signal is true;
	signal G13394: std_logic; attribute dont_touch of G13394: signal is true;
	signal G13409: std_logic; attribute dont_touch of G13409: signal is true;
	signal G13410: std_logic; attribute dont_touch of G13410: signal is true;
	signal G13411: std_logic; attribute dont_touch of G13411: signal is true;
	signal G13412: std_logic; attribute dont_touch of G13412: signal is true;
	signal G13413: std_logic; attribute dont_touch of G13413: signal is true;
	signal G13414: std_logic; attribute dont_touch of G13414: signal is true;
	signal G13415: std_logic; attribute dont_touch of G13415: signal is true;
	signal G13416: std_logic; attribute dont_touch of G13416: signal is true;
	signal G13431: std_logic; attribute dont_touch of G13431: signal is true;
	signal G13432: std_logic; attribute dont_touch of G13432: signal is true;
	signal G13436: std_logic; attribute dont_touch of G13436: signal is true;
	signal G13437: std_logic; attribute dont_touch of G13437: signal is true;
	signal G13458: std_logic; attribute dont_touch of G13458: signal is true;
	signal G13459: std_logic; attribute dont_touch of G13459: signal is true;
	signal G13460: std_logic; attribute dont_touch of G13460: signal is true;
	signal G13461: std_logic; attribute dont_touch of G13461: signal is true;
	signal G13462: std_logic; attribute dont_touch of G13462: signal is true;
	signal G13463: std_logic; attribute dont_touch of G13463: signal is true;
	signal G13464: std_logic; attribute dont_touch of G13464: signal is true;
	signal G13469: std_logic; attribute dont_touch of G13469: signal is true;
	signal G13473: std_logic; attribute dont_touch of G13473: signal is true;
	signal G13474: std_logic; attribute dont_touch of G13474: signal is true;
	signal G13475: std_logic; attribute dont_touch of G13475: signal is true;
	signal G13476: std_logic; attribute dont_touch of G13476: signal is true;
	signal G13477: std_logic; attribute dont_touch of G13477: signal is true;
	signal G13478: std_logic; attribute dont_touch of G13478: signal is true;
	signal G13479: std_logic; attribute dont_touch of G13479: signal is true;
	signal G13480: std_logic; attribute dont_touch of G13480: signal is true;
	signal G13483: std_logic; attribute dont_touch of G13483: signal is true;
	signal G13484: std_logic; attribute dont_touch of G13484: signal is true;
	signal G13485: std_logic; attribute dont_touch of G13485: signal is true;
	signal G13486: std_logic; attribute dont_touch of G13486: signal is true;
	signal G13491: std_logic; attribute dont_touch of G13491: signal is true;
	signal G13492: std_logic; attribute dont_touch of G13492: signal is true;
	signal G13493: std_logic; attribute dont_touch of G13493: signal is true;
	signal G13494: std_logic; attribute dont_touch of G13494: signal is true;
	signal G13495: std_logic; attribute dont_touch of G13495: signal is true;
	signal G13496: std_logic; attribute dont_touch of G13496: signal is true;
	signal G13497: std_logic; attribute dont_touch of G13497: signal is true;
	signal G13498: std_logic; attribute dont_touch of G13498: signal is true;
	signal G13499: std_logic; attribute dont_touch of G13499: signal is true;
	signal G13500: std_logic; attribute dont_touch of G13500: signal is true;
	signal G13501: std_logic; attribute dont_touch of G13501: signal is true;
	signal G13504: std_logic; attribute dont_touch of G13504: signal is true;
	signal G13505: std_logic; attribute dont_touch of G13505: signal is true;
	signal G13506: std_logic; attribute dont_touch of G13506: signal is true;
	signal G13507: std_logic; attribute dont_touch of G13507: signal is true;
	signal G13508: std_logic; attribute dont_touch of G13508: signal is true;
	signal G13509: std_logic; attribute dont_touch of G13509: signal is true;
	signal G13510: std_logic; attribute dont_touch of G13510: signal is true;
	signal G13511: std_logic; attribute dont_touch of G13511: signal is true;
	signal G13512: std_logic; attribute dont_touch of G13512: signal is true;
	signal G13513: std_logic; attribute dont_touch of G13513: signal is true;
	signal G13514: std_logic; attribute dont_touch of G13514: signal is true;
	signal G13515: std_logic; attribute dont_touch of G13515: signal is true;
	signal G13516: std_logic; attribute dont_touch of G13516: signal is true;
	signal G13517: std_logic; attribute dont_touch of G13517: signal is true;
	signal G13518: std_logic; attribute dont_touch of G13518: signal is true;
	signal G13521: std_logic; attribute dont_touch of G13521: signal is true;
	signal G13522: std_logic; attribute dont_touch of G13522: signal is true;
	signal G13523: std_logic; attribute dont_touch of G13523: signal is true;
	signal G13524: std_logic; attribute dont_touch of G13524: signal is true;
	signal G13525: std_logic; attribute dont_touch of G13525: signal is true;
	signal G13526: std_logic; attribute dont_touch of G13526: signal is true;
	signal G13527: std_logic; attribute dont_touch of G13527: signal is true;
	signal G13528: std_logic; attribute dont_touch of G13528: signal is true;
	signal G13529: std_logic; attribute dont_touch of G13529: signal is true;
	signal G13530: std_logic; attribute dont_touch of G13530: signal is true;
	signal G13539: std_logic; attribute dont_touch of G13539: signal is true;
	signal G13540: std_logic; attribute dont_touch of G13540: signal is true;
	signal G13541: std_logic; attribute dont_touch of G13541: signal is true;
	signal G13542: std_logic; attribute dont_touch of G13542: signal is true;
	signal G13543: std_logic; attribute dont_touch of G13543: signal is true;
	signal G13544: std_logic; attribute dont_touch of G13544: signal is true;
	signal G13545: std_logic; attribute dont_touch of G13545: signal is true;
	signal G13551: std_logic; attribute dont_touch of G13551: signal is true;
	signal G13554: std_logic; attribute dont_touch of G13554: signal is true;
	signal G13555: std_logic; attribute dont_touch of G13555: signal is true;
	signal G13564: std_logic; attribute dont_touch of G13564: signal is true;
	signal G13565: std_logic; attribute dont_touch of G13565: signal is true;
	signal G13566: std_logic; attribute dont_touch of G13566: signal is true;
	signal G13567: std_logic; attribute dont_touch of G13567: signal is true;
	signal G13568: std_logic; attribute dont_touch of G13568: signal is true;
	signal G13569: std_logic; attribute dont_touch of G13569: signal is true;
	signal G13570: std_logic; attribute dont_touch of G13570: signal is true;
	signal G13573: std_logic; attribute dont_touch of G13573: signal is true;
	signal G13574: std_logic; attribute dont_touch of G13574: signal is true;
	signal G13580: std_logic; attribute dont_touch of G13580: signal is true;
	signal G13583: std_logic; attribute dont_touch of G13583: signal is true;
	signal G13584: std_logic; attribute dont_touch of G13584: signal is true;
	signal G13593: std_logic; attribute dont_touch of G13593: signal is true;
	signal G13594: std_logic; attribute dont_touch of G13594: signal is true;
	signal G13595: std_logic; attribute dont_touch of G13595: signal is true;
	signal G13596: std_logic; attribute dont_touch of G13596: signal is true;
	signal G13597: std_logic; attribute dont_touch of G13597: signal is true;
	signal G13600: std_logic; attribute dont_touch of G13600: signal is true;
	signal G13603: std_logic; attribute dont_touch of G13603: signal is true;
	signal G13604: std_logic; attribute dont_touch of G13604: signal is true;
	signal G13605: std_logic; attribute dont_touch of G13605: signal is true;
	signal G13620: std_logic; attribute dont_touch of G13620: signal is true;
	signal G13621: std_logic; attribute dont_touch of G13621: signal is true;
	signal G13622: std_logic; attribute dont_touch of G13622: signal is true;
	signal G13623: std_logic; attribute dont_touch of G13623: signal is true;
	signal G13624: std_logic; attribute dont_touch of G13624: signal is true;
	signal G13625: std_logic; attribute dont_touch of G13625: signal is true;
	signal G13626: std_logic; attribute dont_touch of G13626: signal is true;
	signal G13627: std_logic; attribute dont_touch of G13627: signal is true;
	signal G13628: std_logic; attribute dont_touch of G13628: signal is true;
	signal G13631: std_logic; attribute dont_touch of G13631: signal is true;
	signal G13632: std_logic; attribute dont_touch of G13632: signal is true;
	signal G13633: std_logic; attribute dont_touch of G13633: signal is true;
	signal G13634: std_logic; attribute dont_touch of G13634: signal is true;
	signal G13637: std_logic; attribute dont_touch of G13637: signal is true;
	signal G13638: std_logic; attribute dont_touch of G13638: signal is true;
	signal G13655: std_logic; attribute dont_touch of G13655: signal is true;
	signal G13656: std_logic; attribute dont_touch of G13656: signal is true;
	signal G13657: std_logic; attribute dont_touch of G13657: signal is true;
	signal G13660: std_logic; attribute dont_touch of G13660: signal is true;
	signal G13661: std_logic; attribute dont_touch of G13661: signal is true;
	signal G13662: std_logic; attribute dont_touch of G13662: signal is true;
	signal G13663: std_logic; attribute dont_touch of G13663: signal is true;
	signal G13664: std_logic; attribute dont_touch of G13664: signal is true;
	signal G13665: std_logic; attribute dont_touch of G13665: signal is true;
	signal G13666: std_logic; attribute dont_touch of G13666: signal is true;
	signal G13667: std_logic; attribute dont_touch of G13667: signal is true;
	signal G13670: std_logic; attribute dont_touch of G13670: signal is true;
	signal G13671: std_logic; attribute dont_touch of G13671: signal is true;
	signal G13672: std_logic; attribute dont_touch of G13672: signal is true;
	signal G13675: std_logic; attribute dont_touch of G13675: signal is true;
	signal G13676: std_logic; attribute dont_touch of G13676: signal is true;
	signal G13679: std_logic; attribute dont_touch of G13679: signal is true;
	signal G13680: std_logic; attribute dont_touch of G13680: signal is true;
	signal G13697: std_logic; attribute dont_touch of G13697: signal is true;
	signal G13698: std_logic; attribute dont_touch of G13698: signal is true;
	signal G13699: std_logic; attribute dont_touch of G13699: signal is true;
	signal G13700: std_logic; attribute dont_touch of G13700: signal is true;
	signal G13706: std_logic; attribute dont_touch of G13706: signal is true;
	signal G13707: std_logic; attribute dont_touch of G13707: signal is true;
	signal G13708: std_logic; attribute dont_touch of G13708: signal is true;
	signal G13709: std_logic; attribute dont_touch of G13709: signal is true;
	signal G13712: std_logic; attribute dont_touch of G13712: signal is true;
	signal G13715: std_logic; attribute dont_touch of G13715: signal is true;
	signal G13716: std_logic; attribute dont_touch of G13716: signal is true;
	signal G13727: std_logic; attribute dont_touch of G13727: signal is true;
	signal G13728: std_logic; attribute dont_touch of G13728: signal is true;
	signal G13729: std_logic; attribute dont_touch of G13729: signal is true;
	signal G13730: std_logic; attribute dont_touch of G13730: signal is true;
	signal G13736: std_logic; attribute dont_touch of G13736: signal is true;
	signal G13737: std_logic; attribute dont_touch of G13737: signal is true;
	signal G13738: std_logic; attribute dont_touch of G13738: signal is true;
	signal G13739: std_logic; attribute dont_touch of G13739: signal is true;
	signal G13742: std_logic; attribute dont_touch of G13742: signal is true;
	signal G13745: std_logic; attribute dont_touch of G13745: signal is true;
	signal G13756: std_logic; attribute dont_touch of G13756: signal is true;
	signal G13761: std_logic; attribute dont_touch of G13761: signal is true;
	signal G13762: std_logic; attribute dont_touch of G13762: signal is true;
	signal G13763: std_logic; attribute dont_touch of G13763: signal is true;
	signal G13764: std_logic; attribute dont_touch of G13764: signal is true;
	signal G13765: std_logic; attribute dont_touch of G13765: signal is true;
	signal G13771: std_logic; attribute dont_touch of G13771: signal is true;
	signal G13772: std_logic; attribute dont_touch of G13772: signal is true;
	signal G13778: std_logic; attribute dont_touch of G13778: signal is true;
	signal G13779: std_logic; attribute dont_touch of G13779: signal is true;
	signal G13782: std_logic; attribute dont_touch of G13782: signal is true;
	signal G13793: std_logic; attribute dont_touch of G13793: signal is true;
	signal G13794: std_logic; attribute dont_touch of G13794: signal is true;
	signal G13795: std_logic; attribute dont_touch of G13795: signal is true;
	signal G13796: std_logic; attribute dont_touch of G13796: signal is true;
	signal G13797: std_logic; attribute dont_touch of G13797: signal is true;
	signal G13798: std_logic; attribute dont_touch of G13798: signal is true;
	signal G13799: std_logic; attribute dont_touch of G13799: signal is true;
	signal G13805: std_logic; attribute dont_touch of G13805: signal is true;
	signal G13806: std_logic; attribute dont_touch of G13806: signal is true;
	signal G13807: std_logic; attribute dont_touch of G13807: signal is true;
	signal G13808: std_logic; attribute dont_touch of G13808: signal is true;
	signal G13809: std_logic; attribute dont_touch of G13809: signal is true;
	signal G13820: std_logic; attribute dont_touch of G13820: signal is true;
	signal G13821: std_logic; attribute dont_touch of G13821: signal is true;
	signal G13822: std_logic; attribute dont_touch of G13822: signal is true;
	signal G13823: std_logic; attribute dont_touch of G13823: signal is true;
	signal G13824: std_logic; attribute dont_touch of G13824: signal is true;
	signal G13830: std_logic; attribute dont_touch of G13830: signal is true;
	signal G13831: std_logic; attribute dont_touch of G13831: signal is true;
	signal G13832: std_logic; attribute dont_touch of G13832: signal is true;
	signal G13833: std_logic; attribute dont_touch of G13833: signal is true;
	signal G13834: std_logic; attribute dont_touch of G13834: signal is true;
	signal G13835: std_logic; attribute dont_touch of G13835: signal is true;
	signal G13846: std_logic; attribute dont_touch of G13846: signal is true;
	signal G13850: std_logic; attribute dont_touch of G13850: signal is true;
	signal G13851: std_logic; attribute dont_touch of G13851: signal is true;
	signal G13852: std_logic; attribute dont_touch of G13852: signal is true;
	signal G13853: std_logic; attribute dont_touch of G13853: signal is true;
	signal G13854: std_logic; attribute dont_touch of G13854: signal is true;
	signal G13855: std_logic; attribute dont_touch of G13855: signal is true;
	signal G13856: std_logic; attribute dont_touch of G13856: signal is true;
	signal G13857: std_logic; attribute dont_touch of G13857: signal is true;
	signal G13858: std_logic; attribute dont_touch of G13858: signal is true;
	signal G13861: std_logic; attribute dont_touch of G13861: signal is true;
	signal G13866: std_logic; attribute dont_touch of G13866: signal is true;
	signal G13867: std_logic; attribute dont_touch of G13867: signal is true;
	signal G13868: std_logic; attribute dont_touch of G13868: signal is true;
	signal G13869: std_logic; attribute dont_touch of G13869: signal is true;
	signal G13870: std_logic; attribute dont_touch of G13870: signal is true;
	signal G13871: std_logic; attribute dont_touch of G13871: signal is true;
	signal G13872: std_logic; attribute dont_touch of G13872: signal is true;
	signal G13873: std_logic; attribute dont_touch of G13873: signal is true;
	signal G13876: std_logic; attribute dont_touch of G13876: signal is true;
	signal G13877: std_logic; attribute dont_touch of G13877: signal is true;
	signal G13882: std_logic; attribute dont_touch of G13882: signal is true;
	signal G13883: std_logic; attribute dont_touch of G13883: signal is true;
	signal G13884: std_logic; attribute dont_touch of G13884: signal is true;
	signal G13885: std_logic; attribute dont_touch of G13885: signal is true;
	signal G13886: std_logic; attribute dont_touch of G13886: signal is true;
	signal G13887: std_logic; attribute dont_touch of G13887: signal is true;
	signal G13888: std_logic; attribute dont_touch of G13888: signal is true;
	signal G13889: std_logic; attribute dont_touch of G13889: signal is true;
	signal G13892: std_logic; attribute dont_touch of G13892: signal is true;
	signal G13896: std_logic; attribute dont_touch of G13896: signal is true;
	signal G13897: std_logic; attribute dont_touch of G13897: signal is true;
	signal G13898: std_logic; attribute dont_touch of G13898: signal is true;
	signal G13901: std_logic; attribute dont_touch of G13901: signal is true;
	signal G13902: std_logic; attribute dont_touch of G13902: signal is true;
	signal G13907: std_logic; attribute dont_touch of G13907: signal is true;
	signal G13908: std_logic; attribute dont_touch of G13908: signal is true;
	signal G13909: std_logic; attribute dont_touch of G13909: signal is true;
	signal G13910: std_logic; attribute dont_touch of G13910: signal is true;
	signal G13911: std_logic; attribute dont_touch of G13911: signal is true;
	signal G13912: std_logic; attribute dont_touch of G13912: signal is true;
	signal G13913: std_logic; attribute dont_touch of G13913: signal is true;
	signal G13914: std_logic; attribute dont_touch of G13914: signal is true;
	signal G13915: std_logic; attribute dont_touch of G13915: signal is true;
	signal G13918: std_logic; attribute dont_touch of G13918: signal is true;
	signal G13919: std_logic; attribute dont_touch of G13919: signal is true;
	signal G13920: std_logic; attribute dont_touch of G13920: signal is true;
	signal G13923: std_logic; attribute dont_touch of G13923: signal is true;
	signal G13927: std_logic; attribute dont_touch of G13927: signal is true;
	signal G13928: std_logic; attribute dont_touch of G13928: signal is true;
	signal G13929: std_logic; attribute dont_touch of G13929: signal is true;
	signal G13932: std_logic; attribute dont_touch of G13932: signal is true;
	signal G13933: std_logic; attribute dont_touch of G13933: signal is true;
	signal G13937: std_logic; attribute dont_touch of G13937: signal is true;
	signal G13938: std_logic; attribute dont_touch of G13938: signal is true;
	signal G13939: std_logic; attribute dont_touch of G13939: signal is true;
	signal G13940: std_logic; attribute dont_touch of G13940: signal is true;
	signal G13941: std_logic; attribute dont_touch of G13941: signal is true;
	signal G13942: std_logic; attribute dont_touch of G13942: signal is true;
	signal G13943: std_logic; attribute dont_touch of G13943: signal is true;
	signal G13944: std_logic; attribute dont_touch of G13944: signal is true;
	signal G13945: std_logic; attribute dont_touch of G13945: signal is true;
	signal G13946: std_logic; attribute dont_touch of G13946: signal is true;
	signal G13947: std_logic; attribute dont_touch of G13947: signal is true;
	signal G13948: std_logic; attribute dont_touch of G13948: signal is true;
	signal G13951: std_logic; attribute dont_touch of G13951: signal is true;
	signal G13954: std_logic; attribute dont_touch of G13954: signal is true;
	signal G13955: std_logic; attribute dont_touch of G13955: signal is true;
	signal G13958: std_logic; attribute dont_touch of G13958: signal is true;
	signal G13959: std_logic; attribute dont_touch of G13959: signal is true;
	signal G13960: std_logic; attribute dont_touch of G13960: signal is true;
	signal G13963: std_logic; attribute dont_touch of G13963: signal is true;
	signal G13967: std_logic; attribute dont_touch of G13967: signal is true;
	signal G13968: std_logic; attribute dont_touch of G13968: signal is true;
	signal G13969: std_logic; attribute dont_touch of G13969: signal is true;
	signal G13970: std_logic; attribute dont_touch of G13970: signal is true;
	signal G13971: std_logic; attribute dont_touch of G13971: signal is true;
	signal G13972: std_logic; attribute dont_touch of G13972: signal is true;
	signal G13973: std_logic; attribute dont_touch of G13973: signal is true;
	signal G13974: std_logic; attribute dont_touch of G13974: signal is true;
	signal G13975: std_logic; attribute dont_touch of G13975: signal is true;
	signal G13976: std_logic; attribute dont_touch of G13976: signal is true;
	signal G13977: std_logic; attribute dont_touch of G13977: signal is true;
	signal G13980: std_logic; attribute dont_touch of G13980: signal is true;
	signal G13983: std_logic; attribute dont_touch of G13983: signal is true;
	signal G13986: std_logic; attribute dont_touch of G13986: signal is true;
	signal G13989: std_logic; attribute dont_touch of G13989: signal is true;
	signal G13990: std_logic; attribute dont_touch of G13990: signal is true;
	signal G13993: std_logic; attribute dont_touch of G13993: signal is true;
	signal G13994: std_logic; attribute dont_touch of G13994: signal is true;
	signal G13995: std_logic; attribute dont_touch of G13995: signal is true;
	signal G13996: std_logic; attribute dont_touch of G13996: signal is true;
	signal G13997: std_logic; attribute dont_touch of G13997: signal is true;
	signal G13998: std_logic; attribute dont_touch of G13998: signal is true;
	signal G13999: std_logic; attribute dont_touch of G13999: signal is true;
	signal G14000: std_logic; attribute dont_touch of G14000: signal is true;
	signal G14001: std_logic; attribute dont_touch of G14001: signal is true;
	signal G14002: std_logic; attribute dont_touch of G14002: signal is true;
	signal G14003: std_logic; attribute dont_touch of G14003: signal is true;
	signal G14004: std_logic; attribute dont_touch of G14004: signal is true;
	signal G14005: std_logic; attribute dont_touch of G14005: signal is true;
	signal G14008: std_logic; attribute dont_touch of G14008: signal is true;
	signal G14011: std_logic; attribute dont_touch of G14011: signal is true;
	signal G14014: std_logic; attribute dont_touch of G14014: signal is true;
	signal G14015: std_logic; attribute dont_touch of G14015: signal is true;
	signal G14018: std_logic; attribute dont_touch of G14018: signal is true;
	signal G14021: std_logic; attribute dont_touch of G14021: signal is true;
	signal G14024: std_logic; attribute dont_touch of G14024: signal is true;
	signal G14027: std_logic; attribute dont_touch of G14027: signal is true;
	signal G14028: std_logic; attribute dont_touch of G14028: signal is true;
	signal G14029: std_logic; attribute dont_touch of G14029: signal is true;
	signal G14030: std_logic; attribute dont_touch of G14030: signal is true;
	signal G14031: std_logic; attribute dont_touch of G14031: signal is true;
	signal G14032: std_logic; attribute dont_touch of G14032: signal is true;
	signal G14033: std_logic; attribute dont_touch of G14033: signal is true;
	signal G14034: std_logic; attribute dont_touch of G14034: signal is true;
	signal G14035: std_logic; attribute dont_touch of G14035: signal is true;
	signal G14036: std_logic; attribute dont_touch of G14036: signal is true;
	signal G14037: std_logic; attribute dont_touch of G14037: signal is true;
	signal G14038: std_logic; attribute dont_touch of G14038: signal is true;
	signal G14041: std_logic; attribute dont_touch of G14041: signal is true;
	signal G14044: std_logic; attribute dont_touch of G14044: signal is true;
	signal G14045: std_logic; attribute dont_touch of G14045: signal is true;
	signal G14048: std_logic; attribute dont_touch of G14048: signal is true;
	signal G14051: std_logic; attribute dont_touch of G14051: signal is true;
	signal G14054: std_logic; attribute dont_touch of G14054: signal is true;
	signal G14055: std_logic; attribute dont_touch of G14055: signal is true;
	signal G14058: std_logic; attribute dont_touch of G14058: signal is true;
	signal G14061: std_logic; attribute dont_touch of G14061: signal is true;
	signal G14062: std_logic; attribute dont_touch of G14062: signal is true;
	signal G14063: std_logic; attribute dont_touch of G14063: signal is true;
	signal G14064: std_logic; attribute dont_touch of G14064: signal is true;
	signal G14065: std_logic; attribute dont_touch of G14065: signal is true;
	signal G14066: std_logic; attribute dont_touch of G14066: signal is true;
	signal G14069: std_logic; attribute dont_touch of G14069: signal is true;
	signal G14072: std_logic; attribute dont_touch of G14072: signal is true;
	signal G14075: std_logic; attribute dont_touch of G14075: signal is true;
	signal G14078: std_logic; attribute dont_touch of G14078: signal is true;
	signal G14079: std_logic; attribute dont_touch of G14079: signal is true;
	signal G14082: std_logic; attribute dont_touch of G14082: signal is true;
	signal G14085: std_logic; attribute dont_touch of G14085: signal is true;
	signal G14088: std_logic; attribute dont_touch of G14088: signal is true;
	signal G14089: std_logic; attribute dont_touch of G14089: signal is true;
	signal G14090: std_logic; attribute dont_touch of G14090: signal is true;
	signal G14091: std_logic; attribute dont_touch of G14091: signal is true;
	signal G14092: std_logic; attribute dont_touch of G14092: signal is true;
	signal G14093: std_logic; attribute dont_touch of G14093: signal is true;
	signal G14094: std_logic; attribute dont_touch of G14094: signal is true;
	signal G14095: std_logic; attribute dont_touch of G14095: signal is true;
	signal G14097: std_logic; attribute dont_touch of G14097: signal is true;
	signal G14098: std_logic; attribute dont_touch of G14098: signal is true;
	signal G14101: std_logic; attribute dont_touch of G14101: signal is true;
	signal G14104: std_logic; attribute dont_touch of G14104: signal is true;
	signal G14107: std_logic; attribute dont_touch of G14107: signal is true;
	signal G14110: std_logic; attribute dont_touch of G14110: signal is true;
	signal G14113: std_logic; attribute dont_touch of G14113: signal is true;
	signal G14116: std_logic; attribute dont_touch of G14116: signal is true;
	signal G14119: std_logic; attribute dont_touch of G14119: signal is true;
	signal G14120: std_logic; attribute dont_touch of G14120: signal is true;
	signal G14121: std_logic; attribute dont_touch of G14121: signal is true;
	signal G14122: std_logic; attribute dont_touch of G14122: signal is true;
	signal G14123: std_logic; attribute dont_touch of G14123: signal is true;
	signal G14124: std_logic; attribute dont_touch of G14124: signal is true;
	signal G14126: std_logic; attribute dont_touch of G14126: signal is true;
	signal G14127: std_logic; attribute dont_touch of G14127: signal is true;
	signal G14130: std_logic; attribute dont_touch of G14130: signal is true;
	signal G14133: std_logic; attribute dont_touch of G14133: signal is true;
	signal G14136: std_logic; attribute dont_touch of G14136: signal is true;
	signal G14139: std_logic; attribute dont_touch of G14139: signal is true;
	signal G14142: std_logic; attribute dont_touch of G14142: signal is true;
	signal G14145: std_logic; attribute dont_touch of G14145: signal is true;
	signal G14146: std_logic; attribute dont_touch of G14146: signal is true;
	signal G14148: std_logic; attribute dont_touch of G14148: signal is true;
	signal G14149: std_logic; attribute dont_touch of G14149: signal is true;
	signal G14150: std_logic; attribute dont_touch of G14150: signal is true;
	signal G14151: std_logic; attribute dont_touch of G14151: signal is true;
	signal G14154: std_logic; attribute dont_touch of G14154: signal is true;
	signal G14157: std_logic; attribute dont_touch of G14157: signal is true;
	signal G14160: std_logic; attribute dont_touch of G14160: signal is true;
	signal G14163: std_logic; attribute dont_touch of G14163: signal is true;
	signal G14164: std_logic; attribute dont_touch of G14164: signal is true;
	signal G14165: std_logic; attribute dont_touch of G14165: signal is true;
	signal G14166: std_logic; attribute dont_touch of G14166: signal is true;
	signal G14168: std_logic; attribute dont_touch of G14168: signal is true;
	signal G14169: std_logic; attribute dont_touch of G14169: signal is true;
	signal G14170: std_logic; attribute dont_touch of G14170: signal is true;
	signal G14173: std_logic; attribute dont_touch of G14173: signal is true;
	signal G14176: std_logic; attribute dont_touch of G14176: signal is true;
	signal G14177: std_logic; attribute dont_touch of G14177: signal is true;
	signal G14178: std_logic; attribute dont_touch of G14178: signal is true;
	signal G14179: std_logic; attribute dont_touch of G14179: signal is true;
	signal G14180: std_logic; attribute dont_touch of G14180: signal is true;
	signal G14181: std_logic; attribute dont_touch of G14181: signal is true;
	signal G14182: std_logic; attribute dont_touch of G14182: signal is true;
	signal G14183: std_logic; attribute dont_touch of G14183: signal is true;
	signal G14184: std_logic; attribute dont_touch of G14184: signal is true;
	signal G14185: std_logic; attribute dont_touch of G14185: signal is true;
	signal G14186: std_logic; attribute dont_touch of G14186: signal is true;
	signal G14187: std_logic; attribute dont_touch of G14187: signal is true;
	signal G14188: std_logic; attribute dont_touch of G14188: signal is true;
	signal G14190: std_logic; attribute dont_touch of G14190: signal is true;
	signal G14191: std_logic; attribute dont_touch of G14191: signal is true;
	signal G14192: std_logic; attribute dont_touch of G14192: signal is true;
	signal G14193: std_logic; attribute dont_touch of G14193: signal is true;
	signal G14194: std_logic; attribute dont_touch of G14194: signal is true;
	signal G14197: std_logic; attribute dont_touch of G14197: signal is true;
	signal G14198: std_logic; attribute dont_touch of G14198: signal is true;
	signal G14202: std_logic; attribute dont_touch of G14202: signal is true;
	signal G14203: std_logic; attribute dont_touch of G14203: signal is true;
	signal G14204: std_logic; attribute dont_touch of G14204: signal is true;
	signal G14205: std_logic; attribute dont_touch of G14205: signal is true;
	signal G14206: std_logic; attribute dont_touch of G14206: signal is true;
	signal G14207: std_logic; attribute dont_touch of G14207: signal is true;
	signal G14208: std_logic; attribute dont_touch of G14208: signal is true;
	signal G14209: std_logic; attribute dont_touch of G14209: signal is true;
	signal G14210: std_logic; attribute dont_touch of G14210: signal is true;
	signal G14211: std_logic; attribute dont_touch of G14211: signal is true;
	signal G14212: std_logic; attribute dont_touch of G14212: signal is true;
	signal G14215: std_logic; attribute dont_touch of G14215: signal is true;
	signal G14216: std_logic; attribute dont_touch of G14216: signal is true;
	signal G14218: std_logic; attribute dont_touch of G14218: signal is true;
	signal G14219: std_logic; attribute dont_touch of G14219: signal is true;
	signal G14220: std_logic; attribute dont_touch of G14220: signal is true;
	signal G14221: std_logic; attribute dont_touch of G14221: signal is true;
	signal G14222: std_logic; attribute dont_touch of G14222: signal is true;
	signal G14223: std_logic; attribute dont_touch of G14223: signal is true;
	signal G14226: std_logic; attribute dont_touch of G14226: signal is true;
	signal G14227: std_logic; attribute dont_touch of G14227: signal is true;
	signal G14228: std_logic; attribute dont_touch of G14228: signal is true;
	signal G14231: std_logic; attribute dont_touch of G14231: signal is true;
	signal G14232: std_logic; attribute dont_touch of G14232: signal is true;
	signal G14233: std_logic; attribute dont_touch of G14233: signal is true;
	signal G14234: std_logic; attribute dont_touch of G14234: signal is true;
	signal G14237: std_logic; attribute dont_touch of G14237: signal is true;
	signal G14238: std_logic; attribute dont_touch of G14238: signal is true;
	signal G14247: std_logic; attribute dont_touch of G14247: signal is true;
	signal G14248: std_logic; attribute dont_touch of G14248: signal is true;
	signal G14251: std_logic; attribute dont_touch of G14251: signal is true;
	signal G14252: std_logic; attribute dont_touch of G14252: signal is true;
	signal G14253: std_logic; attribute dont_touch of G14253: signal is true;
	signal G14254: std_logic; attribute dont_touch of G14254: signal is true;
	signal G14255: std_logic; attribute dont_touch of G14255: signal is true;
	signal G14256: std_logic; attribute dont_touch of G14256: signal is true;
	signal G14257: std_logic; attribute dont_touch of G14257: signal is true;
	signal G14258: std_logic; attribute dont_touch of G14258: signal is true;
	signal G14261: std_logic; attribute dont_touch of G14261: signal is true;
	signal G14262: std_logic; attribute dont_touch of G14262: signal is true;
	signal G14271: std_logic; attribute dont_touch of G14271: signal is true;
	signal G14272: std_logic; attribute dont_touch of G14272: signal is true;
	signal G14275: std_logic; attribute dont_touch of G14275: signal is true;
	signal G14276: std_logic; attribute dont_touch of G14276: signal is true;
	signal G14277: std_logic; attribute dont_touch of G14277: signal is true;
	signal G14278: std_logic; attribute dont_touch of G14278: signal is true;
	signal G14279: std_logic; attribute dont_touch of G14279: signal is true;
	signal G14290: std_logic; attribute dont_touch of G14290: signal is true;
	signal G14291: std_logic; attribute dont_touch of G14291: signal is true;
	signal G14295: std_logic; attribute dont_touch of G14295: signal is true;
	signal G14296: std_logic; attribute dont_touch of G14296: signal is true;
	signal G14297: std_logic; attribute dont_touch of G14297: signal is true;
	signal G14306: std_logic; attribute dont_touch of G14306: signal is true;
	signal G14307: std_logic; attribute dont_touch of G14307: signal is true;
	signal G14308: std_logic; attribute dont_touch of G14308: signal is true;
	signal G14309: std_logic; attribute dont_touch of G14309: signal is true;
	signal G14313: std_logic; attribute dont_touch of G14313: signal is true;
	signal G14314: std_logic; attribute dont_touch of G14314: signal is true;
	signal G14315: std_logic; attribute dont_touch of G14315: signal is true;
	signal G14316: std_logic; attribute dont_touch of G14316: signal is true;
	signal G14317: std_logic; attribute dont_touch of G14317: signal is true;
	signal G14320: std_logic; attribute dont_touch of G14320: signal is true;
	signal G14321: std_logic; attribute dont_touch of G14321: signal is true;
	signal G14330: std_logic; attribute dont_touch of G14330: signal is true;
	signal G14331: std_logic; attribute dont_touch of G14331: signal is true;
	signal G14332: std_logic; attribute dont_touch of G14332: signal is true;
	signal G14333: std_logic; attribute dont_touch of G14333: signal is true;
	signal G14334: std_logic; attribute dont_touch of G14334: signal is true;
	signal G14335: std_logic; attribute dont_touch of G14335: signal is true;
	signal G14336: std_logic; attribute dont_touch of G14336: signal is true;
	signal G14337: std_logic; attribute dont_touch of G14337: signal is true;
	signal G14338: std_logic; attribute dont_touch of G14338: signal is true;
	signal G14339: std_logic; attribute dont_touch of G14339: signal is true;
	signal G14342: std_logic; attribute dont_touch of G14342: signal is true;
	signal G14343: std_logic; attribute dont_touch of G14343: signal is true;
	signal G14344: std_logic; attribute dont_touch of G14344: signal is true;
	signal G14347: std_logic; attribute dont_touch of G14347: signal is true;
	signal G14348: std_logic; attribute dont_touch of G14348: signal is true;
	signal G14357: std_logic; attribute dont_touch of G14357: signal is true;
	signal G14358: std_logic; attribute dont_touch of G14358: signal is true;
	signal G14359: std_logic; attribute dont_touch of G14359: signal is true;
	signal G14360: std_logic; attribute dont_touch of G14360: signal is true;
	signal G14361: std_logic; attribute dont_touch of G14361: signal is true;
	signal G14362: std_logic; attribute dont_touch of G14362: signal is true;
	signal G14363: std_logic; attribute dont_touch of G14363: signal is true;
	signal G14364: std_logic; attribute dont_touch of G14364: signal is true;
	signal G14365: std_logic; attribute dont_touch of G14365: signal is true;
	signal G14366: std_logic; attribute dont_touch of G14366: signal is true;
	signal G14367: std_logic; attribute dont_touch of G14367: signal is true;
	signal G14376: std_logic; attribute dont_touch of G14376: signal is true;
	signal G14377: std_logic; attribute dont_touch of G14377: signal is true;
	signal G14378: std_logic; attribute dont_touch of G14378: signal is true;
	signal G14379: std_logic; attribute dont_touch of G14379: signal is true;
	signal G14382: std_logic; attribute dont_touch of G14382: signal is true;
	signal G14383: std_logic; attribute dont_touch of G14383: signal is true;
	signal G14384: std_logic; attribute dont_touch of G14384: signal is true;
	signal G14385: std_logic; attribute dont_touch of G14385: signal is true;
	signal G14386: std_logic; attribute dont_touch of G14386: signal is true;
	signal G14387: std_logic; attribute dont_touch of G14387: signal is true;
	signal G14391: std_logic; attribute dont_touch of G14391: signal is true;
	signal G14392: std_logic; attribute dont_touch of G14392: signal is true;
	signal G14393: std_logic; attribute dont_touch of G14393: signal is true;
	signal G14394: std_logic; attribute dont_touch of G14394: signal is true;
	signal G14395: std_logic; attribute dont_touch of G14395: signal is true;
	signal G14396: std_logic; attribute dont_touch of G14396: signal is true;
	signal G14397: std_logic; attribute dont_touch of G14397: signal is true;
	signal G14398: std_logic; attribute dont_touch of G14398: signal is true;
	signal G14399: std_logic; attribute dont_touch of G14399: signal is true;
	signal G14405: std_logic; attribute dont_touch of G14405: signal is true;
	signal G14406: std_logic; attribute dont_touch of G14406: signal is true;
	signal G14407: std_logic; attribute dont_touch of G14407: signal is true;
	signal G14408: std_logic; attribute dont_touch of G14408: signal is true;
	signal G14411: std_logic; attribute dont_touch of G14411: signal is true;
	signal G14412: std_logic; attribute dont_touch of G14412: signal is true;
	signal G14413: std_logic; attribute dont_touch of G14413: signal is true;
	signal G14414: std_logic; attribute dont_touch of G14414: signal is true;
	signal G14415: std_logic; attribute dont_touch of G14415: signal is true;
	signal G14416: std_logic; attribute dont_touch of G14416: signal is true;
	signal G14417: std_logic; attribute dont_touch of G14417: signal is true;
	signal G14418: std_logic; attribute dont_touch of G14418: signal is true;
	signal G14419: std_logic; attribute dont_touch of G14419: signal is true;
	signal G14420: std_logic; attribute dont_touch of G14420: signal is true;
	signal G14422: std_logic; attribute dont_touch of G14422: signal is true;
	signal G14423: std_logic; attribute dont_touch of G14423: signal is true;
	signal G14424: std_logic; attribute dont_touch of G14424: signal is true;
	signal G14425: std_logic; attribute dont_touch of G14425: signal is true;
	signal G14431: std_logic; attribute dont_touch of G14431: signal is true;
	signal G14432: std_logic; attribute dont_touch of G14432: signal is true;
	signal G14433: std_logic; attribute dont_touch of G14433: signal is true;
	signal G14434: std_logic; attribute dont_touch of G14434: signal is true;
	signal G14437: std_logic; attribute dont_touch of G14437: signal is true;
	signal G14438: std_logic; attribute dont_touch of G14438: signal is true;
	signal G14441: std_logic; attribute dont_touch of G14441: signal is true;
	signal G14442: std_logic; attribute dont_touch of G14442: signal is true;
	signal G14443: std_logic; attribute dont_touch of G14443: signal is true;
	signal G14444: std_logic; attribute dont_touch of G14444: signal is true;
	signal G14445: std_logic; attribute dont_touch of G14445: signal is true;
	signal G14446: std_logic; attribute dont_touch of G14446: signal is true;
	signal G14447: std_logic; attribute dont_touch of G14447: signal is true;
	signal G14448: std_logic; attribute dont_touch of G14448: signal is true;
	signal G14449: std_logic; attribute dont_touch of G14449: signal is true;
	signal G14450: std_logic; attribute dont_touch of G14450: signal is true;
	signal G14452: std_logic; attribute dont_touch of G14452: signal is true;
	signal G14453: std_logic; attribute dont_touch of G14453: signal is true;
	signal G14454: std_logic; attribute dont_touch of G14454: signal is true;
	signal G14489: std_logic; attribute dont_touch of G14489: signal is true;
	signal G14490: std_logic; attribute dont_touch of G14490: signal is true;
	signal G14496: std_logic; attribute dont_touch of G14496: signal is true;
	signal G14497: std_logic; attribute dont_touch of G14497: signal is true;
	signal G14503: std_logic; attribute dont_touch of G14503: signal is true;
	signal G14504: std_logic; attribute dont_touch of G14504: signal is true;
	signal G14505: std_logic; attribute dont_touch of G14505: signal is true;
	signal G14506: std_logic; attribute dont_touch of G14506: signal is true;
	signal G14509: std_logic; attribute dont_touch of G14509: signal is true;
	signal G14510: std_logic; attribute dont_touch of G14510: signal is true;
	signal G14511: std_logic; attribute dont_touch of G14511: signal is true;
	signal G14512: std_logic; attribute dont_touch of G14512: signal is true;
	signal G14513: std_logic; attribute dont_touch of G14513: signal is true;
	signal G14514: std_logic; attribute dont_touch of G14514: signal is true;
	signal G14515: std_logic; attribute dont_touch of G14515: signal is true;
	signal G14516: std_logic; attribute dont_touch of G14516: signal is true;
	signal G14517: std_logic; attribute dont_touch of G14517: signal is true;
	signal G14519: std_logic; attribute dont_touch of G14519: signal is true;
	signal G14520: std_logic; attribute dont_touch of G14520: signal is true;
	signal G14521: std_logic; attribute dont_touch of G14521: signal is true;
	signal G14522: std_logic; attribute dont_touch of G14522: signal is true;
	signal G14528: std_logic; attribute dont_touch of G14528: signal is true;
	signal G14529: std_logic; attribute dont_touch of G14529: signal is true;
	signal G14535: std_logic; attribute dont_touch of G14535: signal is true;
	signal G14536: std_logic; attribute dont_touch of G14536: signal is true;
	signal G14537: std_logic; attribute dont_touch of G14537: signal is true;
	signal G14538: std_logic; attribute dont_touch of G14538: signal is true;
	signal G14539: std_logic; attribute dont_touch of G14539: signal is true;
	signal G14540: std_logic; attribute dont_touch of G14540: signal is true;
	signal G14541: std_logic; attribute dont_touch of G14541: signal is true;
	signal G14542: std_logic; attribute dont_touch of G14542: signal is true;
	signal G14543: std_logic; attribute dont_touch of G14543: signal is true;
	signal G14544: std_logic; attribute dont_touch of G14544: signal is true;
	signal G14545: std_logic; attribute dont_touch of G14545: signal is true;
	signal G14546: std_logic; attribute dont_touch of G14546: signal is true;
	signal G14547: std_logic; attribute dont_touch of G14547: signal is true;
	signal G14548: std_logic; attribute dont_touch of G14548: signal is true;
	signal G14549: std_logic; attribute dont_touch of G14549: signal is true;
	signal G14555: std_logic; attribute dont_touch of G14555: signal is true;
	signal G14556: std_logic; attribute dont_touch of G14556: signal is true;
	signal G14562: std_logic; attribute dont_touch of G14562: signal is true;
	signal G14563: std_logic; attribute dont_touch of G14563: signal is true;
	signal G14564: std_logic; attribute dont_touch of G14564: signal is true;
	signal G14565: std_logic; attribute dont_touch of G14565: signal is true;
	signal G14566: std_logic; attribute dont_touch of G14566: signal is true;
	signal G14567: std_logic; attribute dont_touch of G14567: signal is true;
	signal G14568: std_logic; attribute dont_touch of G14568: signal is true;
	signal G14569: std_logic; attribute dont_touch of G14569: signal is true;
	signal G14570: std_logic; attribute dont_touch of G14570: signal is true;
	signal G14571: std_logic; attribute dont_touch of G14571: signal is true;
	signal G14572: std_logic; attribute dont_touch of G14572: signal is true;
	signal G14573: std_logic; attribute dont_touch of G14573: signal is true;
	signal G14574: std_logic; attribute dont_touch of G14574: signal is true;
	signal G14575: std_logic; attribute dont_touch of G14575: signal is true;
	signal G14581: std_logic; attribute dont_touch of G14581: signal is true;
	signal G14582: std_logic; attribute dont_touch of G14582: signal is true;
	signal G14583: std_logic; attribute dont_touch of G14583: signal is true;
	signal G14584: std_logic; attribute dont_touch of G14584: signal is true;
	signal G14585: std_logic; attribute dont_touch of G14585: signal is true;
	signal G14586: std_logic; attribute dont_touch of G14586: signal is true;
	signal G14587: std_logic; attribute dont_touch of G14587: signal is true;
	signal G14588: std_logic; attribute dont_touch of G14588: signal is true;
	signal G14589: std_logic; attribute dont_touch of G14589: signal is true;
	signal G14590: std_logic; attribute dont_touch of G14590: signal is true;
	signal G14591: std_logic; attribute dont_touch of G14591: signal is true;
	signal G14596: std_logic; attribute dont_touch of G14596: signal is true;
	signal G14598: std_logic; attribute dont_touch of G14598: signal is true;
	signal G14599: std_logic; attribute dont_touch of G14599: signal is true;
	signal G14600: std_logic; attribute dont_touch of G14600: signal is true;
	signal G14601: std_logic; attribute dont_touch of G14601: signal is true;
	signal G14602: std_logic; attribute dont_touch of G14602: signal is true;
	signal G14608: std_logic; attribute dont_touch of G14608: signal is true;
	signal G14609: std_logic; attribute dont_touch of G14609: signal is true;
	signal G14610: std_logic; attribute dont_touch of G14610: signal is true;
	signal G14611: std_logic; attribute dont_touch of G14611: signal is true;
	signal G14612: std_logic; attribute dont_touch of G14612: signal is true;
	signal G14613: std_logic; attribute dont_touch of G14613: signal is true;
	signal G14614: std_logic; attribute dont_touch of G14614: signal is true;
	signal G14615: std_logic; attribute dont_touch of G14615: signal is true;
	signal G14616: std_logic; attribute dont_touch of G14616: signal is true;
	signal G14625: std_logic; attribute dont_touch of G14625: signal is true;
	signal G14626: std_logic; attribute dont_touch of G14626: signal is true;
	signal G14627: std_logic; attribute dont_touch of G14627: signal is true;
	signal G14630: std_logic; attribute dont_touch of G14630: signal is true;
	signal G14631: std_logic; attribute dont_touch of G14631: signal is true;
	signal G14636: std_logic; attribute dont_touch of G14636: signal is true;
	signal G14637: std_logic; attribute dont_touch of G14637: signal is true;
	signal G14638: std_logic; attribute dont_touch of G14638: signal is true;
	signal G14639: std_logic; attribute dont_touch of G14639: signal is true;
	signal G14640: std_logic; attribute dont_touch of G14640: signal is true;
	signal G14641: std_logic; attribute dont_touch of G14641: signal is true;
	signal G14642: std_logic; attribute dont_touch of G14642: signal is true;
	signal G14643: std_logic; attribute dont_touch of G14643: signal is true;
	signal G14644: std_logic; attribute dont_touch of G14644: signal is true;
	signal G14645: std_logic; attribute dont_touch of G14645: signal is true;
	signal G14654: std_logic; attribute dont_touch of G14654: signal is true;
	signal G14655: std_logic; attribute dont_touch of G14655: signal is true;
	signal G14656: std_logic; attribute dont_touch of G14656: signal is true;
	signal G14659: std_logic; attribute dont_touch of G14659: signal is true;
	signal G14663: std_logic; attribute dont_touch of G14663: signal is true;
	signal G14664: std_logic; attribute dont_touch of G14664: signal is true;
	signal G14665: std_logic; attribute dont_touch of G14665: signal is true;
	signal G14668: std_logic; attribute dont_touch of G14668: signal is true;
	signal G14669: std_logic; attribute dont_touch of G14669: signal is true;
	signal G14674: std_logic; attribute dont_touch of G14674: signal is true;
	signal G14675: std_logic; attribute dont_touch of G14675: signal is true;
	signal G14676: std_logic; attribute dont_touch of G14676: signal is true;
	signal G14677: std_logic; attribute dont_touch of G14677: signal is true;
	signal G14678: std_logic; attribute dont_touch of G14678: signal is true;
	signal G14679: std_logic; attribute dont_touch of G14679: signal is true;
	signal G14680: std_logic; attribute dont_touch of G14680: signal is true;
	signal G14681: std_logic; attribute dont_touch of G14681: signal is true;
	signal G14682: std_logic; attribute dont_touch of G14682: signal is true;
	signal G14683: std_logic; attribute dont_touch of G14683: signal is true;
	signal G14686: std_logic; attribute dont_touch of G14686: signal is true;
	signal G14687: std_logic; attribute dont_touch of G14687: signal is true;
	signal G14688: std_logic; attribute dont_touch of G14688: signal is true;
	signal G14691: std_logic; attribute dont_touch of G14691: signal is true;
	signal G14695: std_logic; attribute dont_touch of G14695: signal is true;
	signal G14696: std_logic; attribute dont_touch of G14696: signal is true;
	signal G14697: std_logic; attribute dont_touch of G14697: signal is true;
	signal G14700: std_logic; attribute dont_touch of G14700: signal is true;
	signal G14701: std_logic; attribute dont_touch of G14701: signal is true;
	signal G14706: std_logic; attribute dont_touch of G14706: signal is true;
	signal G14707: std_logic; attribute dont_touch of G14707: signal is true;
	signal G14708: std_logic; attribute dont_touch of G14708: signal is true;
	signal G14712: std_logic; attribute dont_touch of G14712: signal is true;
	signal G14713: std_logic; attribute dont_touch of G14713: signal is true;
	signal G14714: std_logic; attribute dont_touch of G14714: signal is true;
	signal G14719: std_logic; attribute dont_touch of G14719: signal is true;
	signal G14720: std_logic; attribute dont_touch of G14720: signal is true;
	signal G14723: std_logic; attribute dont_touch of G14723: signal is true;
	signal G14726: std_logic; attribute dont_touch of G14726: signal is true;
	signal G14727: std_logic; attribute dont_touch of G14727: signal is true;
	signal G14730: std_logic; attribute dont_touch of G14730: signal is true;
	signal G14731: std_logic; attribute dont_touch of G14731: signal is true;
	signal G14732: std_logic; attribute dont_touch of G14732: signal is true;
	signal G14735: std_logic; attribute dont_touch of G14735: signal is true;
	signal G14739: std_logic; attribute dont_touch of G14739: signal is true;
	signal G14740: std_logic; attribute dont_touch of G14740: signal is true;
	signal G14741: std_logic; attribute dont_touch of G14741: signal is true;
	signal G14744: std_logic; attribute dont_touch of G14744: signal is true;
	signal G14745: std_logic; attribute dont_touch of G14745: signal is true;
	signal G14750: std_logic; attribute dont_touch of G14750: signal is true;
	signal G14751: std_logic; attribute dont_touch of G14751: signal is true;
	signal G14752: std_logic; attribute dont_touch of G14752: signal is true;
	signal G14753: std_logic; attribute dont_touch of G14753: signal is true;
	signal G14754: std_logic; attribute dont_touch of G14754: signal is true;
	signal G14755: std_logic; attribute dont_touch of G14755: signal is true;
	signal G14758: std_logic; attribute dont_touch of G14758: signal is true;
	signal G14761: std_logic; attribute dont_touch of G14761: signal is true;
	signal G14764: std_logic; attribute dont_touch of G14764: signal is true;
	signal G14767: std_logic; attribute dont_touch of G14767: signal is true;
	signal G14768: std_logic; attribute dont_touch of G14768: signal is true;
	signal G14771: std_logic; attribute dont_touch of G14771: signal is true;
	signal G14772: std_logic; attribute dont_touch of G14772: signal is true;
	signal G14773: std_logic; attribute dont_touch of G14773: signal is true;
	signal G14776: std_logic; attribute dont_touch of G14776: signal is true;
	signal G14780: std_logic; attribute dont_touch of G14780: signal is true;
	signal G14781: std_logic; attribute dont_touch of G14781: signal is true;
	signal G14782: std_logic; attribute dont_touch of G14782: signal is true;
	signal G14785: std_logic; attribute dont_touch of G14785: signal is true;
	signal G14786: std_logic; attribute dont_touch of G14786: signal is true;
	signal G14790: std_logic; attribute dont_touch of G14790: signal is true;
	signal G14791: std_logic; attribute dont_touch of G14791: signal is true;
	signal G14792: std_logic; attribute dont_touch of G14792: signal is true;
	signal G14793: std_logic; attribute dont_touch of G14793: signal is true;
	signal G14794: std_logic; attribute dont_touch of G14794: signal is true;
	signal G14797: std_logic; attribute dont_touch of G14797: signal is true;
	signal G14800: std_logic; attribute dont_touch of G14800: signal is true;
	signal G14803: std_logic; attribute dont_touch of G14803: signal is true;
	signal G14804: std_logic; attribute dont_touch of G14804: signal is true;
	signal G14807: std_logic; attribute dont_touch of G14807: signal is true;
	signal G14810: std_logic; attribute dont_touch of G14810: signal is true;
	signal G14813: std_logic; attribute dont_touch of G14813: signal is true;
	signal G14816: std_logic; attribute dont_touch of G14816: signal is true;
	signal G14817: std_logic; attribute dont_touch of G14817: signal is true;
	signal G14820: std_logic; attribute dont_touch of G14820: signal is true;
	signal G14821: std_logic; attribute dont_touch of G14821: signal is true;
	signal G14822: std_logic; attribute dont_touch of G14822: signal is true;
	signal G14825: std_logic; attribute dont_touch of G14825: signal is true;
	signal G14829: std_logic; attribute dont_touch of G14829: signal is true;
	signal G14830: std_logic; attribute dont_touch of G14830: signal is true;
	signal G14831: std_logic; attribute dont_touch of G14831: signal is true;
	signal G14832: std_logic; attribute dont_touch of G14832: signal is true;
	signal G14833: std_logic; attribute dont_touch of G14833: signal is true;
	signal G14838: std_logic; attribute dont_touch of G14838: signal is true;
	signal G14841: std_logic; attribute dont_touch of G14841: signal is true;
	signal G14844: std_logic; attribute dont_touch of G14844: signal is true;
	signal G14845: std_logic; attribute dont_touch of G14845: signal is true;
	signal G14848: std_logic; attribute dont_touch of G14848: signal is true;
	signal G14851: std_logic; attribute dont_touch of G14851: signal is true;
	signal G14854: std_logic; attribute dont_touch of G14854: signal is true;
	signal G14855: std_logic; attribute dont_touch of G14855: signal is true;
	signal G14858: std_logic; attribute dont_touch of G14858: signal is true;
	signal G14861: std_logic; attribute dont_touch of G14861: signal is true;
	signal G14864: std_logic; attribute dont_touch of G14864: signal is true;
	signal G14867: std_logic; attribute dont_touch of G14867: signal is true;
	signal G14868: std_logic; attribute dont_touch of G14868: signal is true;
	signal G14871: std_logic; attribute dont_touch of G14871: signal is true;
	signal G14872: std_logic; attribute dont_touch of G14872: signal is true;
	signal G14873: std_logic; attribute dont_touch of G14873: signal is true;
	signal G14874: std_logic; attribute dont_touch of G14874: signal is true;
	signal G14875: std_logic; attribute dont_touch of G14875: signal is true;
	signal G14876: std_logic; attribute dont_touch of G14876: signal is true;
	signal G14879: std_logic; attribute dont_touch of G14879: signal is true;
	signal G14882: std_logic; attribute dont_touch of G14882: signal is true;
	signal G14885: std_logic; attribute dont_touch of G14885: signal is true;
	signal G14888: std_logic; attribute dont_touch of G14888: signal is true;
	signal G14889: std_logic; attribute dont_touch of G14889: signal is true;
	signal G14892: std_logic; attribute dont_touch of G14892: signal is true;
	signal G14895: std_logic; attribute dont_touch of G14895: signal is true;
	signal G14898: std_logic; attribute dont_touch of G14898: signal is true;
	signal G14899: std_logic; attribute dont_touch of G14899: signal is true;
	signal G14902: std_logic; attribute dont_touch of G14902: signal is true;
	signal G14905: std_logic; attribute dont_touch of G14905: signal is true;
	signal G14908: std_logic; attribute dont_touch of G14908: signal is true;
	signal G14911: std_logic; attribute dont_touch of G14911: signal is true;
	signal G14912: std_logic; attribute dont_touch of G14912: signal is true;
	signal G14913: std_logic; attribute dont_touch of G14913: signal is true;
	signal G14914: std_logic; attribute dont_touch of G14914: signal is true;
	signal G14915: std_logic; attribute dont_touch of G14915: signal is true;
	signal G14918: std_logic; attribute dont_touch of G14918: signal is true;
	signal G14921: std_logic; attribute dont_touch of G14921: signal is true;
	signal G14924: std_logic; attribute dont_touch of G14924: signal is true;
	signal G14927: std_logic; attribute dont_touch of G14927: signal is true;
	signal G14930: std_logic; attribute dont_touch of G14930: signal is true;
	signal G14933: std_logic; attribute dont_touch of G14933: signal is true;
	signal G14936: std_logic; attribute dont_touch of G14936: signal is true;
	signal G14937: std_logic; attribute dont_touch of G14937: signal is true;
	signal G14940: std_logic; attribute dont_touch of G14940: signal is true;
	signal G14943: std_logic; attribute dont_touch of G14943: signal is true;
	signal G14946: std_logic; attribute dont_touch of G14946: signal is true;
	signal G14947: std_logic; attribute dont_touch of G14947: signal is true;
	signal G14950: std_logic; attribute dont_touch of G14950: signal is true;
	signal G14953: std_logic; attribute dont_touch of G14953: signal is true;
	signal G14956: std_logic; attribute dont_touch of G14956: signal is true;
	signal G14959: std_logic; attribute dont_touch of G14959: signal is true;
	signal G14962: std_logic; attribute dont_touch of G14962: signal is true;
	signal G14965: std_logic; attribute dont_touch of G14965: signal is true;
	signal G14968: std_logic; attribute dont_touch of G14968: signal is true;
	signal G14971: std_logic; attribute dont_touch of G14971: signal is true;
	signal G14974: std_logic; attribute dont_touch of G14974: signal is true;
	signal G14977: std_logic; attribute dont_touch of G14977: signal is true;
	signal G14978: std_logic; attribute dont_touch of G14978: signal is true;
	signal G14981: std_logic; attribute dont_touch of G14981: signal is true;
	signal G14984: std_logic; attribute dont_touch of G14984: signal is true;
	signal G14987: std_logic; attribute dont_touch of G14987: signal is true;
	signal G14988: std_logic; attribute dont_touch of G14988: signal is true;
	signal G14993: std_logic; attribute dont_touch of G14993: signal is true;
	signal G14996: std_logic; attribute dont_touch of G14996: signal is true;
	signal G14999: std_logic; attribute dont_touch of G14999: signal is true;
	signal G15002: std_logic; attribute dont_touch of G15002: signal is true;
	signal G15005: std_logic; attribute dont_touch of G15005: signal is true;
	signal G15008: std_logic; attribute dont_touch of G15008: signal is true;
	signal G15011: std_logic; attribute dont_touch of G15011: signal is true;
	signal G15014: std_logic; attribute dont_touch of G15014: signal is true;
	signal G15017: std_logic; attribute dont_touch of G15017: signal is true;
	signal G15018: std_logic; attribute dont_touch of G15018: signal is true;
	signal G15021: std_logic; attribute dont_touch of G15021: signal is true;
	signal G15024: std_logic; attribute dont_touch of G15024: signal is true;
	signal G15027: std_logic; attribute dont_touch of G15027: signal is true;
	signal G15030: std_logic; attribute dont_touch of G15030: signal is true;
	signal G15033: std_logic; attribute dont_touch of G15033: signal is true;
	signal G15036: std_logic; attribute dont_touch of G15036: signal is true;
	signal G15039: std_logic; attribute dont_touch of G15039: signal is true;
	signal G15042: std_logic; attribute dont_touch of G15042: signal is true;
	signal G15045: std_logic; attribute dont_touch of G15045: signal is true;
	signal G15048: std_logic; attribute dont_touch of G15048: signal is true;
	signal G15049: std_logic; attribute dont_touch of G15049: signal is true;
	signal G15050: std_logic; attribute dont_touch of G15050: signal is true;
	signal G15051: std_logic; attribute dont_touch of G15051: signal is true;
	signal G15052: std_logic; attribute dont_touch of G15052: signal is true;
	signal G15053: std_logic; attribute dont_touch of G15053: signal is true;
	signal G15054: std_logic; attribute dont_touch of G15054: signal is true;
	signal G15055: std_logic; attribute dont_touch of G15055: signal is true;
	signal G15056: std_logic; attribute dont_touch of G15056: signal is true;
	signal G15057: std_logic; attribute dont_touch of G15057: signal is true;
	signal G15058: std_logic; attribute dont_touch of G15058: signal is true;
	signal G15059: std_logic; attribute dont_touch of G15059: signal is true;
	signal G15060: std_logic; attribute dont_touch of G15060: signal is true;
	signal G15061: std_logic; attribute dont_touch of G15061: signal is true;
	signal G15062: std_logic; attribute dont_touch of G15062: signal is true;
	signal G15063: std_logic; attribute dont_touch of G15063: signal is true;
	signal G15064: std_logic; attribute dont_touch of G15064: signal is true;
	signal G15065: std_logic; attribute dont_touch of G15065: signal is true;
	signal G15066: std_logic; attribute dont_touch of G15066: signal is true;
	signal G15067: std_logic; attribute dont_touch of G15067: signal is true;
	signal G15068: std_logic; attribute dont_touch of G15068: signal is true;
	signal G15069: std_logic; attribute dont_touch of G15069: signal is true;
	signal G15070: std_logic; attribute dont_touch of G15070: signal is true;
	signal G15071: std_logic; attribute dont_touch of G15071: signal is true;
	signal G15072: std_logic; attribute dont_touch of G15072: signal is true;
	signal G15073: std_logic; attribute dont_touch of G15073: signal is true;
	signal G15074: std_logic; attribute dont_touch of G15074: signal is true;
	signal G15075: std_logic; attribute dont_touch of G15075: signal is true;
	signal G15076: std_logic; attribute dont_touch of G15076: signal is true;
	signal G15077: std_logic; attribute dont_touch of G15077: signal is true;
	signal G15078: std_logic; attribute dont_touch of G15078: signal is true;
	signal G15079: std_logic; attribute dont_touch of G15079: signal is true;
	signal G15080: std_logic; attribute dont_touch of G15080: signal is true;
	signal G15081: std_logic; attribute dont_touch of G15081: signal is true;
	signal G15082: std_logic; attribute dont_touch of G15082: signal is true;
	signal G15083: std_logic; attribute dont_touch of G15083: signal is true;
	signal G15084: std_logic; attribute dont_touch of G15084: signal is true;
	signal G15085: std_logic; attribute dont_touch of G15085: signal is true;
	signal G15086: std_logic; attribute dont_touch of G15086: signal is true;
	signal G15087: std_logic; attribute dont_touch of G15087: signal is true;
	signal G15088: std_logic; attribute dont_touch of G15088: signal is true;
	signal G15089: std_logic; attribute dont_touch of G15089: signal is true;
	signal G15090: std_logic; attribute dont_touch of G15090: signal is true;
	signal G15091: std_logic; attribute dont_touch of G15091: signal is true;
	signal G15092: std_logic; attribute dont_touch of G15092: signal is true;
	signal G15093: std_logic; attribute dont_touch of G15093: signal is true;
	signal G15094: std_logic; attribute dont_touch of G15094: signal is true;
	signal G15095: std_logic; attribute dont_touch of G15095: signal is true;
	signal G15096: std_logic; attribute dont_touch of G15096: signal is true;
	signal G15097: std_logic; attribute dont_touch of G15097: signal is true;
	signal G15098: std_logic; attribute dont_touch of G15098: signal is true;
	signal G15099: std_logic; attribute dont_touch of G15099: signal is true;
	signal G15100: std_logic; attribute dont_touch of G15100: signal is true;
	signal G15101: std_logic; attribute dont_touch of G15101: signal is true;
	signal G15102: std_logic; attribute dont_touch of G15102: signal is true;
	signal G15103: std_logic; attribute dont_touch of G15103: signal is true;
	signal G15104: std_logic; attribute dont_touch of G15104: signal is true;
	signal G15105: std_logic; attribute dont_touch of G15105: signal is true;
	signal G15106: std_logic; attribute dont_touch of G15106: signal is true;
	signal G15107: std_logic; attribute dont_touch of G15107: signal is true;
	signal G15108: std_logic; attribute dont_touch of G15108: signal is true;
	signal G15109: std_logic; attribute dont_touch of G15109: signal is true;
	signal G15110: std_logic; attribute dont_touch of G15110: signal is true;
	signal G15111: std_logic; attribute dont_touch of G15111: signal is true;
	signal G15112: std_logic; attribute dont_touch of G15112: signal is true;
	signal G15113: std_logic; attribute dont_touch of G15113: signal is true;
	signal G15114: std_logic; attribute dont_touch of G15114: signal is true;
	signal G15115: std_logic; attribute dont_touch of G15115: signal is true;
	signal G15116: std_logic; attribute dont_touch of G15116: signal is true;
	signal G15117: std_logic; attribute dont_touch of G15117: signal is true;
	signal G15118: std_logic; attribute dont_touch of G15118: signal is true;
	signal G15119: std_logic; attribute dont_touch of G15119: signal is true;
	signal G15120: std_logic; attribute dont_touch of G15120: signal is true;
	signal G15121: std_logic; attribute dont_touch of G15121: signal is true;
	signal G15122: std_logic; attribute dont_touch of G15122: signal is true;
	signal G15123: std_logic; attribute dont_touch of G15123: signal is true;
	signal G15124: std_logic; attribute dont_touch of G15124: signal is true;
	signal G15125: std_logic; attribute dont_touch of G15125: signal is true;
	signal G15126: std_logic; attribute dont_touch of G15126: signal is true;
	signal G15127: std_logic; attribute dont_touch of G15127: signal is true;
	signal G15128: std_logic; attribute dont_touch of G15128: signal is true;
	signal G15129: std_logic; attribute dont_touch of G15129: signal is true;
	signal G15130: std_logic; attribute dont_touch of G15130: signal is true;
	signal G15131: std_logic; attribute dont_touch of G15131: signal is true;
	signal G15132: std_logic; attribute dont_touch of G15132: signal is true;
	signal G15133: std_logic; attribute dont_touch of G15133: signal is true;
	signal G15134: std_logic; attribute dont_touch of G15134: signal is true;
	signal G15135: std_logic; attribute dont_touch of G15135: signal is true;
	signal G15136: std_logic; attribute dont_touch of G15136: signal is true;
	signal G15137: std_logic; attribute dont_touch of G15137: signal is true;
	signal G15138: std_logic; attribute dont_touch of G15138: signal is true;
	signal G15139: std_logic; attribute dont_touch of G15139: signal is true;
	signal G15140: std_logic; attribute dont_touch of G15140: signal is true;
	signal G15141: std_logic; attribute dont_touch of G15141: signal is true;
	signal G15142: std_logic; attribute dont_touch of G15142: signal is true;
	signal G15143: std_logic; attribute dont_touch of G15143: signal is true;
	signal G15144: std_logic; attribute dont_touch of G15144: signal is true;
	signal G15145: std_logic; attribute dont_touch of G15145: signal is true;
	signal G15146: std_logic; attribute dont_touch of G15146: signal is true;
	signal G15147: std_logic; attribute dont_touch of G15147: signal is true;
	signal G15148: std_logic; attribute dont_touch of G15148: signal is true;
	signal G15149: std_logic; attribute dont_touch of G15149: signal is true;
	signal G15150: std_logic; attribute dont_touch of G15150: signal is true;
	signal G15151: std_logic; attribute dont_touch of G15151: signal is true;
	signal G15152: std_logic; attribute dont_touch of G15152: signal is true;
	signal G15153: std_logic; attribute dont_touch of G15153: signal is true;
	signal G15154: std_logic; attribute dont_touch of G15154: signal is true;
	signal G15155: std_logic; attribute dont_touch of G15155: signal is true;
	signal G15156: std_logic; attribute dont_touch of G15156: signal is true;
	signal G15157: std_logic; attribute dont_touch of G15157: signal is true;
	signal G15158: std_logic; attribute dont_touch of G15158: signal is true;
	signal G15159: std_logic; attribute dont_touch of G15159: signal is true;
	signal G15160: std_logic; attribute dont_touch of G15160: signal is true;
	signal G15161: std_logic; attribute dont_touch of G15161: signal is true;
	signal G15162: std_logic; attribute dont_touch of G15162: signal is true;
	signal G15163: std_logic; attribute dont_touch of G15163: signal is true;
	signal G15164: std_logic; attribute dont_touch of G15164: signal is true;
	signal G15165: std_logic; attribute dont_touch of G15165: signal is true;
	signal G15166: std_logic; attribute dont_touch of G15166: signal is true;
	signal G15167: std_logic; attribute dont_touch of G15167: signal is true;
	signal G15168: std_logic; attribute dont_touch of G15168: signal is true;
	signal G15169: std_logic; attribute dont_touch of G15169: signal is true;
	signal G15170: std_logic; attribute dont_touch of G15170: signal is true;
	signal G15171: std_logic; attribute dont_touch of G15171: signal is true;
	signal G15224: std_logic; attribute dont_touch of G15224: signal is true;
	signal G15277: std_logic; attribute dont_touch of G15277: signal is true;
	signal G15344: std_logic; attribute dont_touch of G15344: signal is true;
	signal G15345: std_logic; attribute dont_touch of G15345: signal is true;
	signal G15348: std_logic; attribute dont_touch of G15348: signal is true;
	signal G15371: std_logic; attribute dont_touch of G15371: signal is true;
	signal G15372: std_logic; attribute dont_touch of G15372: signal is true;
	signal G15373: std_logic; attribute dont_touch of G15373: signal is true;
	signal G15426: std_logic; attribute dont_touch of G15426: signal is true;
	signal G15479: std_logic; attribute dont_touch of G15479: signal is true;
	signal G15480: std_logic; attribute dont_touch of G15480: signal is true;
	signal G15483: std_logic; attribute dont_touch of G15483: signal is true;
	signal G15506: std_logic; attribute dont_touch of G15506: signal is true;
	signal G15507: std_logic; attribute dont_touch of G15507: signal is true;
	signal G15508: std_logic; attribute dont_touch of G15508: signal is true;
	signal G15509: std_logic; attribute dont_touch of G15509: signal is true;
	signal G15562: std_logic; attribute dont_touch of G15562: signal is true;
	signal G15563: std_logic; attribute dont_touch of G15563: signal is true;
	signal G15566: std_logic; attribute dont_touch of G15566: signal is true;
	signal G15567: std_logic; attribute dont_touch of G15567: signal is true;
	signal G15568: std_logic; attribute dont_touch of G15568: signal is true;
	signal G15569: std_logic; attribute dont_touch of G15569: signal is true;
	signal G15570: std_logic; attribute dont_touch of G15570: signal is true;
	signal G15571: std_logic; attribute dont_touch of G15571: signal is true;
	signal G15572: std_logic; attribute dont_touch of G15572: signal is true;
	signal G15573: std_logic; attribute dont_touch of G15573: signal is true;
	signal G15574: std_logic; attribute dont_touch of G15574: signal is true;
	signal G15578: std_logic; attribute dont_touch of G15578: signal is true;
	signal G15579: std_logic; attribute dont_touch of G15579: signal is true;
	signal G15580: std_logic; attribute dont_touch of G15580: signal is true;
	signal G15581: std_logic; attribute dont_touch of G15581: signal is true;
	signal G15582: std_logic; attribute dont_touch of G15582: signal is true;
	signal G15585: std_logic; attribute dont_touch of G15585: signal is true;
	signal G15588: std_logic; attribute dont_touch of G15588: signal is true;
	signal G15589: std_logic; attribute dont_touch of G15589: signal is true;
	signal G15590: std_logic; attribute dont_touch of G15590: signal is true;
	signal G15591: std_logic; attribute dont_touch of G15591: signal is true;
	signal G15594: std_logic; attribute dont_touch of G15594: signal is true;
	signal G15595: std_logic; attribute dont_touch of G15595: signal is true;
	signal G15608: std_logic; attribute dont_touch of G15608: signal is true;
	signal G15611: std_logic; attribute dont_touch of G15611: signal is true;
	signal G15612: std_logic; attribute dont_touch of G15612: signal is true;
	signal G15613: std_logic; attribute dont_touch of G15613: signal is true;
	signal G15614: std_logic; attribute dont_touch of G15614: signal is true;
	signal G15615: std_logic; attribute dont_touch of G15615: signal is true;
	signal G15628: std_logic; attribute dont_touch of G15628: signal is true;
	signal G15631: std_logic; attribute dont_touch of G15631: signal is true;
	signal G15632: std_logic; attribute dont_touch of G15632: signal is true;
	signal G15633: std_logic; attribute dont_touch of G15633: signal is true;
	signal G15634: std_logic; attribute dont_touch of G15634: signal is true;
	signal G15647: std_logic; attribute dont_touch of G15647: signal is true;
	signal G15650: std_logic; attribute dont_touch of G15650: signal is true;
	signal G15651: std_logic; attribute dont_touch of G15651: signal is true;
	signal G15652: std_logic; attribute dont_touch of G15652: signal is true;
	signal G15653: std_logic; attribute dont_touch of G15653: signal is true;
	signal G15654: std_logic; attribute dont_touch of G15654: signal is true;
	signal G15655: std_logic; attribute dont_touch of G15655: signal is true;
	signal G15656: std_logic; attribute dont_touch of G15656: signal is true;
	signal G15669: std_logic; attribute dont_touch of G15669: signal is true;
	signal G15672: std_logic; attribute dont_touch of G15672: signal is true;
	signal G15673: std_logic; attribute dont_touch of G15673: signal is true;
	signal G15674: std_logic; attribute dont_touch of G15674: signal is true;
	signal G15678: std_logic; attribute dont_touch of G15678: signal is true;
	signal G15679: std_logic; attribute dont_touch of G15679: signal is true;
	signal G15680: std_logic; attribute dont_touch of G15680: signal is true;
	signal G15693: std_logic; attribute dont_touch of G15693: signal is true;
	signal G15694: std_logic; attribute dont_touch of G15694: signal is true;
	signal G15695: std_logic; attribute dont_touch of G15695: signal is true;
	signal G15699: std_logic; attribute dont_touch of G15699: signal is true;
	signal G15700: std_logic; attribute dont_touch of G15700: signal is true;
	signal G15701: std_logic; attribute dont_touch of G15701: signal is true;
	signal G15702: std_logic; attribute dont_touch of G15702: signal is true;
	signal G15703: std_logic; attribute dont_touch of G15703: signal is true;
	signal G15704: std_logic; attribute dont_touch of G15704: signal is true;
	signal G15705: std_logic; attribute dont_touch of G15705: signal is true;
	signal G15706: std_logic; attribute dont_touch of G15706: signal is true;
	signal G15707: std_logic; attribute dont_touch of G15707: signal is true;
	signal G15708: std_logic; attribute dont_touch of G15708: signal is true;
	signal G15709: std_logic; attribute dont_touch of G15709: signal is true;
	signal G15710: std_logic; attribute dont_touch of G15710: signal is true;
	signal G15711: std_logic; attribute dont_touch of G15711: signal is true;
	signal G15712: std_logic; attribute dont_touch of G15712: signal is true;
	signal G15713: std_logic; attribute dont_touch of G15713: signal is true;
	signal G15714: std_logic; attribute dont_touch of G15714: signal is true;
	signal G15715: std_logic; attribute dont_touch of G15715: signal is true;
	signal G15716: std_logic; attribute dont_touch of G15716: signal is true;
	signal G15717: std_logic; attribute dont_touch of G15717: signal is true;
	signal G15718: std_logic; attribute dont_touch of G15718: signal is true;
	signal G15719: std_logic; attribute dont_touch of G15719: signal is true;
	signal G15720: std_logic; attribute dont_touch of G15720: signal is true;
	signal G15721: std_logic; attribute dont_touch of G15721: signal is true;
	signal G15722: std_logic; attribute dont_touch of G15722: signal is true;
	signal G15723: std_logic; attribute dont_touch of G15723: signal is true;
	signal G15724: std_logic; attribute dont_touch of G15724: signal is true;
	signal G15725: std_logic; attribute dont_touch of G15725: signal is true;
	signal G15726: std_logic; attribute dont_touch of G15726: signal is true;
	signal G15727: std_logic; attribute dont_touch of G15727: signal is true;
	signal G15728: std_logic; attribute dont_touch of G15728: signal is true;
	signal G15729: std_logic; attribute dont_touch of G15729: signal is true;
	signal G15730: std_logic; attribute dont_touch of G15730: signal is true;
	signal G15731: std_logic; attribute dont_touch of G15731: signal is true;
	signal G15732: std_logic; attribute dont_touch of G15732: signal is true;
	signal G15733: std_logic; attribute dont_touch of G15733: signal is true;
	signal G15734: std_logic; attribute dont_touch of G15734: signal is true;
	signal G15735: std_logic; attribute dont_touch of G15735: signal is true;
	signal G15736: std_logic; attribute dont_touch of G15736: signal is true;
	signal G15737: std_logic; attribute dont_touch of G15737: signal is true;
	signal G15738: std_logic; attribute dont_touch of G15738: signal is true;
	signal G15739: std_logic; attribute dont_touch of G15739: signal is true;
	signal G15740: std_logic; attribute dont_touch of G15740: signal is true;
	signal G15741: std_logic; attribute dont_touch of G15741: signal is true;
	signal G15742: std_logic; attribute dont_touch of G15742: signal is true;
	signal G15743: std_logic; attribute dont_touch of G15743: signal is true;
	signal G15744: std_logic; attribute dont_touch of G15744: signal is true;
	signal G15745: std_logic; attribute dont_touch of G15745: signal is true;
	signal G15746: std_logic; attribute dont_touch of G15746: signal is true;
	signal G15747: std_logic; attribute dont_touch of G15747: signal is true;
	signal G15748: std_logic; attribute dont_touch of G15748: signal is true;
	signal G15749: std_logic; attribute dont_touch of G15749: signal is true;
	signal G15750: std_logic; attribute dont_touch of G15750: signal is true;
	signal G15751: std_logic; attribute dont_touch of G15751: signal is true;
	signal G15752: std_logic; attribute dont_touch of G15752: signal is true;
	signal G15753: std_logic; attribute dont_touch of G15753: signal is true;
	signal G15754: std_logic; attribute dont_touch of G15754: signal is true;
	signal G15755: std_logic; attribute dont_touch of G15755: signal is true;
	signal G15756: std_logic; attribute dont_touch of G15756: signal is true;
	signal G15757: std_logic; attribute dont_touch of G15757: signal is true;
	signal G15758: std_logic; attribute dont_touch of G15758: signal is true;
	signal G15779: std_logic; attribute dont_touch of G15779: signal is true;
	signal G15780: std_logic; attribute dont_touch of G15780: signal is true;
	signal G15781: std_logic; attribute dont_touch of G15781: signal is true;
	signal G15782: std_logic; attribute dont_touch of G15782: signal is true;
	signal G15783: std_logic; attribute dont_touch of G15783: signal is true;
	signal G15784: std_logic; attribute dont_touch of G15784: signal is true;
	signal G15785: std_logic; attribute dont_touch of G15785: signal is true;
	signal G15786: std_logic; attribute dont_touch of G15786: signal is true;
	signal G15787: std_logic; attribute dont_touch of G15787: signal is true;
	signal G15788: std_logic; attribute dont_touch of G15788: signal is true;
	signal G15789: std_logic; attribute dont_touch of G15789: signal is true;
	signal G15792: std_logic; attribute dont_touch of G15792: signal is true;
	signal G15793: std_logic; attribute dont_touch of G15793: signal is true;
	signal G15794: std_logic; attribute dont_touch of G15794: signal is true;
	signal G15795: std_logic; attribute dont_touch of G15795: signal is true;
	signal G15796: std_logic; attribute dont_touch of G15796: signal is true;
	signal G15797: std_logic; attribute dont_touch of G15797: signal is true;
	signal G15798: std_logic; attribute dont_touch of G15798: signal is true;
	signal G15799: std_logic; attribute dont_touch of G15799: signal is true;
	signal G15800: std_logic; attribute dont_touch of G15800: signal is true;
	signal G15803: std_logic; attribute dont_touch of G15803: signal is true;
	signal G15804: std_logic; attribute dont_touch of G15804: signal is true;
	signal G15805: std_logic; attribute dont_touch of G15805: signal is true;
	signal G15806: std_logic; attribute dont_touch of G15806: signal is true;
	signal G15807: std_logic; attribute dont_touch of G15807: signal is true;
	signal G15808: std_logic; attribute dont_touch of G15808: signal is true;
	signal G15809: std_logic; attribute dont_touch of G15809: signal is true;
	signal G15810: std_logic; attribute dont_touch of G15810: signal is true;
	signal G15811: std_logic; attribute dont_touch of G15811: signal is true;
	signal G15812: std_logic; attribute dont_touch of G15812: signal is true;
	signal G15813: std_logic; attribute dont_touch of G15813: signal is true;
	signal G15814: std_logic; attribute dont_touch of G15814: signal is true;
	signal G15815: std_logic; attribute dont_touch of G15815: signal is true;
	signal G15816: std_logic; attribute dont_touch of G15816: signal is true;
	signal G15817: std_logic; attribute dont_touch of G15817: signal is true;
	signal G15818: std_logic; attribute dont_touch of G15818: signal is true;
	signal G15819: std_logic; attribute dont_touch of G15819: signal is true;
	signal G15820: std_logic; attribute dont_touch of G15820: signal is true;
	signal G15821: std_logic; attribute dont_touch of G15821: signal is true;
	signal G15822: std_logic; attribute dont_touch of G15822: signal is true;
	signal G15823: std_logic; attribute dont_touch of G15823: signal is true;
	signal G15824: std_logic; attribute dont_touch of G15824: signal is true;
	signal G15825: std_logic; attribute dont_touch of G15825: signal is true;
	signal G15829: std_logic; attribute dont_touch of G15829: signal is true;
	signal G15830: std_logic; attribute dont_touch of G15830: signal is true;
	signal G15831: std_logic; attribute dont_touch of G15831: signal is true;
	signal G15832: std_logic; attribute dont_touch of G15832: signal is true;
	signal G15833: std_logic; attribute dont_touch of G15833: signal is true;
	signal G15836: std_logic; attribute dont_touch of G15836: signal is true;
	signal G15837: std_logic; attribute dont_touch of G15837: signal is true;
	signal G15838: std_logic; attribute dont_touch of G15838: signal is true;
	signal G15839: std_logic; attribute dont_touch of G15839: signal is true;
	signal G15840: std_logic; attribute dont_touch of G15840: signal is true;
	signal G15841: std_logic; attribute dont_touch of G15841: signal is true;
	signal G15842: std_logic; attribute dont_touch of G15842: signal is true;
	signal G15843: std_logic; attribute dont_touch of G15843: signal is true;
	signal G15844: std_logic; attribute dont_touch of G15844: signal is true;
	signal G15847: std_logic; attribute dont_touch of G15847: signal is true;
	signal G15848: std_logic; attribute dont_touch of G15848: signal is true;
	signal G15849: std_logic; attribute dont_touch of G15849: signal is true;
	signal G15850: std_logic; attribute dont_touch of G15850: signal is true;
	signal G15851: std_logic; attribute dont_touch of G15851: signal is true;
	signal G15852: std_logic; attribute dont_touch of G15852: signal is true;
	signal G15853: std_logic; attribute dont_touch of G15853: signal is true;
	signal G15856: std_logic; attribute dont_touch of G15856: signal is true;
	signal G15857: std_logic; attribute dont_touch of G15857: signal is true;
	signal G15858: std_logic; attribute dont_touch of G15858: signal is true;
	signal G15859: std_logic; attribute dont_touch of G15859: signal is true;
	signal G15860: std_logic; attribute dont_touch of G15860: signal is true;
	signal G15861: std_logic; attribute dont_touch of G15861: signal is true;
	signal G15862: std_logic; attribute dont_touch of G15862: signal is true;
	signal G15863: std_logic; attribute dont_touch of G15863: signal is true;
	signal G15864: std_logic; attribute dont_touch of G15864: signal is true;
	signal G15867: std_logic; attribute dont_touch of G15867: signal is true;
	signal G15870: std_logic; attribute dont_touch of G15870: signal is true;
	signal G15871: std_logic; attribute dont_touch of G15871: signal is true;
	signal G15872: std_logic; attribute dont_touch of G15872: signal is true;
	signal G15873: std_logic; attribute dont_touch of G15873: signal is true;
	signal G15874: std_logic; attribute dont_touch of G15874: signal is true;
	signal G15875: std_logic; attribute dont_touch of G15875: signal is true;
	signal G15876: std_logic; attribute dont_touch of G15876: signal is true;
	signal G15877: std_logic; attribute dont_touch of G15877: signal is true;
	signal G15880: std_logic; attribute dont_touch of G15880: signal is true;
	signal G15881: std_logic; attribute dont_touch of G15881: signal is true;
	signal G15882: std_logic; attribute dont_touch of G15882: signal is true;
	signal G15883: std_logic; attribute dont_touch of G15883: signal is true;
	signal G15884: std_logic; attribute dont_touch of G15884: signal is true;
	signal G15885: std_logic; attribute dont_touch of G15885: signal is true;
	signal G15902: std_logic; attribute dont_touch of G15902: signal is true;
	signal G15903: std_logic; attribute dont_touch of G15903: signal is true;
	signal G15904: std_logic; attribute dont_touch of G15904: signal is true;
	signal G15907: std_logic; attribute dont_touch of G15907: signal is true;
	signal G15910: std_logic; attribute dont_touch of G15910: signal is true;
	signal G15911: std_logic; attribute dont_touch of G15911: signal is true;
	signal G15912: std_logic; attribute dont_touch of G15912: signal is true;
	signal G15913: std_logic; attribute dont_touch of G15913: signal is true;
	signal G15914: std_logic; attribute dont_touch of G15914: signal is true;
	signal G15915: std_logic; attribute dont_touch of G15915: signal is true;
	signal G15932: std_logic; attribute dont_touch of G15932: signal is true;
	signal G15935: std_logic; attribute dont_touch of G15935: signal is true;
	signal G15936: std_logic; attribute dont_touch of G15936: signal is true;
	signal G15937: std_logic; attribute dont_touch of G15937: signal is true;
	signal G15938: std_logic; attribute dont_touch of G15938: signal is true;
	signal G15959: std_logic; attribute dont_touch of G15959: signal is true;
	signal G15962: std_logic; attribute dont_touch of G15962: signal is true;
	signal G15965: std_logic; attribute dont_touch of G15965: signal is true;
	signal G15966: std_logic; attribute dont_touch of G15966: signal is true;
	signal G15967: std_logic; attribute dont_touch of G15967: signal is true;
	signal G15968: std_logic; attribute dont_touch of G15968: signal is true;
	signal G15969: std_logic; attribute dont_touch of G15969: signal is true;
	signal G15978: std_logic; attribute dont_touch of G15978: signal is true;
	signal G15979: std_logic; attribute dont_touch of G15979: signal is true;
	signal G15992: std_logic; attribute dont_touch of G15992: signal is true;
	signal G15995: std_logic; attribute dont_touch of G15995: signal is true;
	signal G16000: std_logic; attribute dont_touch of G16000: signal is true;
	signal G16021: std_logic; attribute dont_touch of G16021: signal is true;
	signal G16022: std_logic; attribute dont_touch of G16022: signal is true;
	signal G16023: std_logic; attribute dont_touch of G16023: signal is true;
	signal G16024: std_logic; attribute dont_touch of G16024: signal is true;
	signal G16025: std_logic; attribute dont_touch of G16025: signal is true;
	signal G16026: std_logic; attribute dont_touch of G16026: signal is true;
	signal G16027: std_logic; attribute dont_touch of G16027: signal is true;
	signal G16030: std_logic; attribute dont_touch of G16030: signal is true;
	signal G16031: std_logic; attribute dont_touch of G16031: signal is true;
	signal G16044: std_logic; attribute dont_touch of G16044: signal is true;
	signal G16047: std_logic; attribute dont_touch of G16047: signal is true;
	signal G16052: std_logic; attribute dont_touch of G16052: signal is true;
	signal G16053: std_logic; attribute dont_touch of G16053: signal is true;
	signal G16066: std_logic; attribute dont_touch of G16066: signal is true;
	signal G16069: std_logic; attribute dont_touch of G16069: signal is true;
	signal G16072: std_logic; attribute dont_touch of G16072: signal is true;
	signal G16075: std_logic; attribute dont_touch of G16075: signal is true;
	signal G16076: std_logic; attribute dont_touch of G16076: signal is true;
	signal G16077: std_logic; attribute dont_touch of G16077: signal is true;
	signal G16090: std_logic; attribute dont_touch of G16090: signal is true;
	signal G16093: std_logic; attribute dont_touch of G16093: signal is true;
	signal G16096: std_logic; attribute dont_touch of G16096: signal is true;
	signal G16097: std_logic; attribute dont_touch of G16097: signal is true;
	signal G16098: std_logic; attribute dont_touch of G16098: signal is true;
	signal G16099: std_logic; attribute dont_touch of G16099: signal is true;
	signal G16100: std_logic; attribute dont_touch of G16100: signal is true;
	signal G16119: std_logic; attribute dont_touch of G16119: signal is true;
	signal G16122: std_logic; attribute dont_touch of G16122: signal is true;
	signal G16123: std_logic; attribute dont_touch of G16123: signal is true;
	signal G16124: std_logic; attribute dont_touch of G16124: signal is true;
	signal G16125: std_logic; attribute dont_touch of G16125: signal is true;
	signal G16126: std_logic; attribute dont_touch of G16126: signal is true;
	signal G16127: std_logic; attribute dont_touch of G16127: signal is true;
	signal G16128: std_logic; attribute dont_touch of G16128: signal is true;
	signal G16129: std_logic; attribute dont_touch of G16129: signal is true;
	signal G16136: std_logic; attribute dont_touch of G16136: signal is true;
	signal G16155: std_logic; attribute dont_touch of G16155: signal is true;
	signal G16158: std_logic; attribute dont_touch of G16158: signal is true;
	signal G16159: std_logic; attribute dont_touch of G16159: signal is true;
	signal G16160: std_logic; attribute dont_touch of G16160: signal is true;
	signal G16161: std_logic; attribute dont_touch of G16161: signal is true;
	signal G16162: std_logic; attribute dont_touch of G16162: signal is true;
	signal G16163: std_logic; attribute dont_touch of G16163: signal is true;
	signal G16164: std_logic; attribute dont_touch of G16164: signal is true;
	signal G16171: std_logic; attribute dont_touch of G16171: signal is true;
	signal G16172: std_logic; attribute dont_touch of G16172: signal is true;
	signal G16173: std_logic; attribute dont_touch of G16173: signal is true;
	signal G16176: std_logic; attribute dont_touch of G16176: signal is true;
	signal G16177: std_logic; attribute dont_touch of G16177: signal is true;
	signal G16178: std_logic; attribute dont_touch of G16178: signal is true;
	signal G16179: std_logic; attribute dont_touch of G16179: signal is true;
	signal G16180: std_logic; attribute dont_touch of G16180: signal is true;
	signal G16181: std_logic; attribute dont_touch of G16181: signal is true;
	signal G16182: std_logic; attribute dont_touch of G16182: signal is true;
	signal G16183: std_logic; attribute dont_touch of G16183: signal is true;
	signal G16184: std_logic; attribute dont_touch of G16184: signal is true;
	signal G16185: std_logic; attribute dont_touch of G16185: signal is true;
	signal G16186: std_logic; attribute dont_touch of G16186: signal is true;
	signal G16187: std_logic; attribute dont_touch of G16187: signal is true;
	signal G16190: std_logic; attribute dont_touch of G16190: signal is true;
	signal G16191: std_logic; attribute dont_touch of G16191: signal is true;
	signal G16192: std_logic; attribute dont_touch of G16192: signal is true;
	signal G16193: std_logic; attribute dont_touch of G16193: signal is true;
	signal G16194: std_logic; attribute dont_touch of G16194: signal is true;
	signal G16195: std_logic; attribute dont_touch of G16195: signal is true;
	signal G16196: std_logic; attribute dont_touch of G16196: signal is true;
	signal G16197: std_logic; attribute dont_touch of G16197: signal is true;
	signal G16198: std_logic; attribute dont_touch of G16198: signal is true;
	signal G16199: std_logic; attribute dont_touch of G16199: signal is true;
	signal G16200: std_logic; attribute dont_touch of G16200: signal is true;
	signal G16201: std_logic; attribute dont_touch of G16201: signal is true;
	signal G16202: std_logic; attribute dont_touch of G16202: signal is true;
	signal G16203: std_logic; attribute dont_touch of G16203: signal is true;
	signal G16204: std_logic; attribute dont_touch of G16204: signal is true;
	signal G16205: std_logic; attribute dont_touch of G16205: signal is true;
	signal G16206: std_logic; attribute dont_touch of G16206: signal is true;
	signal G16207: std_logic; attribute dont_touch of G16207: signal is true;
	signal G16208: std_logic; attribute dont_touch of G16208: signal is true;
	signal G16209: std_logic; attribute dont_touch of G16209: signal is true;
	signal G16210: std_logic; attribute dont_touch of G16210: signal is true;
	signal G16211: std_logic; attribute dont_touch of G16211: signal is true;
	signal G16212: std_logic; attribute dont_touch of G16212: signal is true;
	signal G16213: std_logic; attribute dont_touch of G16213: signal is true;
	signal G16214: std_logic; attribute dont_touch of G16214: signal is true;
	signal G16215: std_logic; attribute dont_touch of G16215: signal is true;
	signal G16216: std_logic; attribute dont_touch of G16216: signal is true;
	signal G16219: std_logic; attribute dont_touch of G16219: signal is true;
	signal G16220: std_logic; attribute dont_touch of G16220: signal is true;
	signal G16221: std_logic; attribute dont_touch of G16221: signal is true;
	signal G16222: std_logic; attribute dont_touch of G16222: signal is true;
	signal G16223: std_logic; attribute dont_touch of G16223: signal is true;
	signal G16224: std_logic; attribute dont_touch of G16224: signal is true;
	signal G16225: std_logic; attribute dont_touch of G16225: signal is true;
	signal G16226: std_logic; attribute dont_touch of G16226: signal is true;
	signal G16227: std_logic; attribute dont_touch of G16227: signal is true;
	signal G16228: std_logic; attribute dont_touch of G16228: signal is true;
	signal G16231: std_logic; attribute dont_touch of G16231: signal is true;
	signal G16232: std_logic; attribute dont_touch of G16232: signal is true;
	signal G16233: std_logic; attribute dont_touch of G16233: signal is true;
	signal G16234: std_logic; attribute dont_touch of G16234: signal is true;
	signal G16235: std_logic; attribute dont_touch of G16235: signal is true;
	signal G16236: std_logic; attribute dont_touch of G16236: signal is true;
	signal G16237: std_logic; attribute dont_touch of G16237: signal is true;
	signal G16238: std_logic; attribute dont_touch of G16238: signal is true;
	signal G16239: std_logic; attribute dont_touch of G16239: signal is true;
	signal G16242: std_logic; attribute dont_touch of G16242: signal is true;
	signal G16243: std_logic; attribute dont_touch of G16243: signal is true;
	signal G16244: std_logic; attribute dont_touch of G16244: signal is true;
	signal G16245: std_logic; attribute dont_touch of G16245: signal is true;
	signal G16246: std_logic; attribute dont_touch of G16246: signal is true;
	signal G16249: std_logic; attribute dont_touch of G16249: signal is true;
	signal G16258: std_logic; attribute dont_touch of G16258: signal is true;
	signal G16259: std_logic; attribute dont_touch of G16259: signal is true;
	signal G16260: std_logic; attribute dont_touch of G16260: signal is true;
	signal G16261: std_logic; attribute dont_touch of G16261: signal is true;
	signal G16264: std_logic; attribute dont_touch of G16264: signal is true;
	signal G16268: std_logic; attribute dont_touch of G16268: signal is true;
	signal G16272: std_logic; attribute dont_touch of G16272: signal is true;
	signal G16275: std_logic; attribute dont_touch of G16275: signal is true;
	signal G16278: std_logic; attribute dont_touch of G16278: signal is true;
	signal G16279: std_logic; attribute dont_touch of G16279: signal is true;
	signal G16280: std_logic; attribute dont_touch of G16280: signal is true;
	signal G16281: std_logic; attribute dont_touch of G16281: signal is true;
	signal G16282: std_logic; attribute dont_touch of G16282: signal is true;
	signal G16283: std_logic; attribute dont_touch of G16283: signal is true;
	signal G16284: std_logic; attribute dont_touch of G16284: signal is true;
	signal G16285: std_logic; attribute dont_touch of G16285: signal is true;
	signal G16286: std_logic; attribute dont_touch of G16286: signal is true;
	signal G16287: std_logic; attribute dont_touch of G16287: signal is true;
	signal G16288: std_logic; attribute dont_touch of G16288: signal is true;
	signal G16289: std_logic; attribute dont_touch of G16289: signal is true;
	signal G16290: std_logic; attribute dont_touch of G16290: signal is true;
	signal G16291: std_logic; attribute dont_touch of G16291: signal is true;
	signal G16292: std_logic; attribute dont_touch of G16292: signal is true;
	signal G16296: std_logic; attribute dont_touch of G16296: signal is true;
	signal G16299: std_logic; attribute dont_touch of G16299: signal is true;
	signal G16300: std_logic; attribute dont_touch of G16300: signal is true;
	signal G16303: std_logic; attribute dont_touch of G16303: signal is true;
	signal G16304: std_logic; attribute dont_touch of G16304: signal is true;
	signal G16305: std_logic; attribute dont_touch of G16305: signal is true;
	signal G16306: std_logic; attribute dont_touch of G16306: signal is true;
	signal G16307: std_logic; attribute dont_touch of G16307: signal is true;
	signal G16308: std_logic; attribute dont_touch of G16308: signal is true;
	signal G16309: std_logic; attribute dont_touch of G16309: signal is true;
	signal G16310: std_logic; attribute dont_touch of G16310: signal is true;
	signal G16311: std_logic; attribute dont_touch of G16311: signal is true;
	signal G16312: std_logic; attribute dont_touch of G16312: signal is true;
	signal G16313: std_logic; attribute dont_touch of G16313: signal is true;
	signal G16316: std_logic; attribute dont_touch of G16316: signal is true;
	signal G16319: std_logic; attribute dont_touch of G16319: signal is true;
	signal G16320: std_logic; attribute dont_touch of G16320: signal is true;
	signal G16321: std_logic; attribute dont_touch of G16321: signal is true;
	signal G16322: std_logic; attribute dont_touch of G16322: signal is true;
	signal G16323: std_logic; attribute dont_touch of G16323: signal is true;
	signal G16324: std_logic; attribute dont_touch of G16324: signal is true;
	signal G16325: std_logic; attribute dont_touch of G16325: signal is true;
	signal G16326: std_logic; attribute dont_touch of G16326: signal is true;
	signal G16349: std_logic; attribute dont_touch of G16349: signal is true;
	signal G16422: std_logic; attribute dont_touch of G16422: signal is true;
	signal G16423: std_logic; attribute dont_touch of G16423: signal is true;
	signal G16424: std_logic; attribute dont_touch of G16424: signal is true;
	signal G16427: std_logic; attribute dont_touch of G16427: signal is true;
	signal G16428: std_logic; attribute dont_touch of G16428: signal is true;
	signal G16429: std_logic; attribute dont_touch of G16429: signal is true;
	signal G16430: std_logic; attribute dont_touch of G16430: signal is true;
	signal G16431: std_logic; attribute dont_touch of G16431: signal is true;
	signal G16448: std_logic; attribute dont_touch of G16448: signal is true;
	signal G16449: std_logic; attribute dont_touch of G16449: signal is true;
	signal G16472: std_logic; attribute dont_touch of G16472: signal is true;
	signal G16473: std_logic; attribute dont_touch of G16473: signal is true;
	signal G16474: std_logic; attribute dont_touch of G16474: signal is true;
	signal G16475: std_logic; attribute dont_touch of G16475: signal is true;
	signal G16476: std_logic; attribute dont_touch of G16476: signal is true;
	signal G16479: std_logic; attribute dont_touch of G16479: signal is true;
	signal G16482: std_logic; attribute dont_touch of G16482: signal is true;
	signal G16483: std_logic; attribute dont_touch of G16483: signal is true;
	signal G16484: std_logic; attribute dont_touch of G16484: signal is true;
	signal G16485: std_logic; attribute dont_touch of G16485: signal is true;
	signal G16486: std_logic; attribute dont_touch of G16486: signal is true;
	signal G16487: std_logic; attribute dont_touch of G16487: signal is true;
	signal G16488: std_logic; attribute dont_touch of G16488: signal is true;
	signal G16489: std_logic; attribute dont_touch of G16489: signal is true;
	signal G16506: std_logic; attribute dont_touch of G16506: signal is true;
	signal G16507: std_logic; attribute dont_touch of G16507: signal is true;
	signal G16508: std_logic; attribute dont_touch of G16508: signal is true;
	signal G16509: std_logic; attribute dont_touch of G16509: signal is true;
	signal G16510: std_logic; attribute dont_touch of G16510: signal is true;
	signal G16511: std_logic; attribute dont_touch of G16511: signal is true;
	signal G16512: std_logic; attribute dont_touch of G16512: signal is true;
	signal G16513: std_logic; attribute dont_touch of G16513: signal is true;
	signal G16514: std_logic; attribute dont_touch of G16514: signal is true;
	signal G16515: std_logic; attribute dont_touch of G16515: signal is true;
	signal G16516: std_logic; attribute dont_touch of G16516: signal is true;
	signal G16517: std_logic; attribute dont_touch of G16517: signal is true;
	signal G16518: std_logic; attribute dont_touch of G16518: signal is true;
	signal G16519: std_logic; attribute dont_touch of G16519: signal is true;
	signal G16520: std_logic; attribute dont_touch of G16520: signal is true;
	signal G16521: std_logic; attribute dont_touch of G16521: signal is true;
	signal G16522: std_logic; attribute dont_touch of G16522: signal is true;
	signal G16523: std_logic; attribute dont_touch of G16523: signal is true;
	signal G16524: std_logic; attribute dont_touch of G16524: signal is true;
	signal G16525: std_logic; attribute dont_touch of G16525: signal is true;
	signal G16526: std_logic; attribute dont_touch of G16526: signal is true;
	signal G16527: std_logic; attribute dont_touch of G16527: signal is true;
	signal G16528: std_logic; attribute dont_touch of G16528: signal is true;
	signal G16529: std_logic; attribute dont_touch of G16529: signal is true;
	signal G16530: std_logic; attribute dont_touch of G16530: signal is true;
	signal G16531: std_logic; attribute dont_touch of G16531: signal is true;
	signal G16532: std_logic; attribute dont_touch of G16532: signal is true;
	signal G16533: std_logic; attribute dont_touch of G16533: signal is true;
	signal G16534: std_logic; attribute dont_touch of G16534: signal is true;
	signal G16535: std_logic; attribute dont_touch of G16535: signal is true;
	signal G16536: std_logic; attribute dont_touch of G16536: signal is true;
	signal G16537: std_logic; attribute dont_touch of G16537: signal is true;
	signal G16538: std_logic; attribute dont_touch of G16538: signal is true;
	signal G16539: std_logic; attribute dont_touch of G16539: signal is true;
	signal G16540: std_logic; attribute dont_touch of G16540: signal is true;
	signal G16577: std_logic; attribute dont_touch of G16577: signal is true;
	signal G16578: std_logic; attribute dont_touch of G16578: signal is true;
	signal G16579: std_logic; attribute dont_touch of G16579: signal is true;
	signal G16580: std_logic; attribute dont_touch of G16580: signal is true;
	signal G16581: std_logic; attribute dont_touch of G16581: signal is true;
	signal G16582: std_logic; attribute dont_touch of G16582: signal is true;
	signal G16583: std_logic; attribute dont_touch of G16583: signal is true;
	signal G16584: std_logic; attribute dont_touch of G16584: signal is true;
	signal G16585: std_logic; attribute dont_touch of G16585: signal is true;
	signal G16586: std_logic; attribute dont_touch of G16586: signal is true;
	signal G16587: std_logic; attribute dont_touch of G16587: signal is true;
	signal G16588: std_logic; attribute dont_touch of G16588: signal is true;
	signal G16589: std_logic; attribute dont_touch of G16589: signal is true;
	signal G16590: std_logic; attribute dont_touch of G16590: signal is true;
	signal G16591: std_logic; attribute dont_touch of G16591: signal is true;
	signal G16592: std_logic; attribute dont_touch of G16592: signal is true;
	signal G16593: std_logic; attribute dont_touch of G16593: signal is true;
	signal G16594: std_logic; attribute dont_touch of G16594: signal is true;
	signal G16595: std_logic; attribute dont_touch of G16595: signal is true;
	signal G16596: std_logic; attribute dont_touch of G16596: signal is true;
	signal G16597: std_logic; attribute dont_touch of G16597: signal is true;
	signal G16598: std_logic; attribute dont_touch of G16598: signal is true;
	signal G16599: std_logic; attribute dont_touch of G16599: signal is true;
	signal G16600: std_logic; attribute dont_touch of G16600: signal is true;
	signal G16601: std_logic; attribute dont_touch of G16601: signal is true;
	signal G16602: std_logic; attribute dont_touch of G16602: signal is true;
	signal G16604: std_logic; attribute dont_touch of G16604: signal is true;
	signal G16605: std_logic; attribute dont_touch of G16605: signal is true;
	signal G16606: std_logic; attribute dont_touch of G16606: signal is true;
	signal G16607: std_logic; attribute dont_touch of G16607: signal is true;
	signal G16608: std_logic; attribute dont_touch of G16608: signal is true;
	signal G16609: std_logic; attribute dont_touch of G16609: signal is true;
	signal G16610: std_logic; attribute dont_touch of G16610: signal is true;
	signal G16611: std_logic; attribute dont_touch of G16611: signal is true;
	signal G16612: std_logic; attribute dont_touch of G16612: signal is true;
	signal G16613: std_logic; attribute dont_touch of G16613: signal is true;
	signal G16614: std_logic; attribute dont_touch of G16614: signal is true;
	signal G16615: std_logic; attribute dont_touch of G16615: signal is true;
	signal G16616: std_logic; attribute dont_touch of G16616: signal is true;
	signal G16617: std_logic; attribute dont_touch of G16617: signal is true;
	signal G16618: std_logic; attribute dont_touch of G16618: signal is true;
	signal G16619: std_logic; attribute dont_touch of G16619: signal is true;
	signal G16620: std_logic; attribute dont_touch of G16620: signal is true;
	signal G16621: std_logic; attribute dont_touch of G16621: signal is true;
	signal G16622: std_logic; attribute dont_touch of G16622: signal is true;
	signal G16623: std_logic; attribute dont_touch of G16623: signal is true;
	signal G16625: std_logic; attribute dont_touch of G16625: signal is true;
	signal G16626: std_logic; attribute dont_touch of G16626: signal is true;
	signal G16628: std_logic; attribute dont_touch of G16628: signal is true;
	signal G16629: std_logic; attribute dont_touch of G16629: signal is true;
	signal G16630: std_logic; attribute dont_touch of G16630: signal is true;
	signal G16631: std_logic; attribute dont_touch of G16631: signal is true;
	signal G16632: std_logic; attribute dont_touch of G16632: signal is true;
	signal G16633: std_logic; attribute dont_touch of G16633: signal is true;
	signal G16634: std_logic; attribute dont_touch of G16634: signal is true;
	signal G16635: std_logic; attribute dont_touch of G16635: signal is true;
	signal G16636: std_logic; attribute dont_touch of G16636: signal is true;
	signal G16637: std_logic; attribute dont_touch of G16637: signal is true;
	signal G16638: std_logic; attribute dont_touch of G16638: signal is true;
	signal G16639: std_logic; attribute dont_touch of G16639: signal is true;
	signal G16640: std_logic; attribute dont_touch of G16640: signal is true;
	signal G16641: std_logic; attribute dont_touch of G16641: signal is true;
	signal G16642: std_logic; attribute dont_touch of G16642: signal is true;
	signal G16643: std_logic; attribute dont_touch of G16643: signal is true;
	signal G16644: std_logic; attribute dont_touch of G16644: signal is true;
	signal G16645: std_logic; attribute dont_touch of G16645: signal is true;
	signal G16646: std_logic; attribute dont_touch of G16646: signal is true;
	signal G16651: std_logic; attribute dont_touch of G16651: signal is true;
	signal G16652: std_logic; attribute dont_touch of G16652: signal is true;
	signal G16653: std_logic; attribute dont_touch of G16653: signal is true;
	signal G16654: std_logic; attribute dont_touch of G16654: signal is true;
	signal G16655: std_logic; attribute dont_touch of G16655: signal is true;
	signal G16657: std_logic; attribute dont_touch of G16657: signal is true;
	signal G16658: std_logic; attribute dont_touch of G16658: signal is true;
	signal G16660: std_logic; attribute dont_touch of G16660: signal is true;
	signal G16661: std_logic; attribute dont_touch of G16661: signal is true;
	signal G16662: std_logic; attribute dont_touch of G16662: signal is true;
	signal G16663: std_logic; attribute dont_touch of G16663: signal is true;
	signal G16666: std_logic; attribute dont_touch of G16666: signal is true;
	signal G16667: std_logic; attribute dont_touch of G16667: signal is true;
	signal G16668: std_logic; attribute dont_touch of G16668: signal is true;
	signal G16669: std_logic; attribute dont_touch of G16669: signal is true;
	signal G16670: std_logic; attribute dont_touch of G16670: signal is true;
	signal G16671: std_logic; attribute dont_touch of G16671: signal is true;
	signal G16672: std_logic; attribute dont_touch of G16672: signal is true;
	signal G16673: std_logic; attribute dont_touch of G16673: signal is true;
	signal G16674: std_logic; attribute dont_touch of G16674: signal is true;
	signal G16675: std_logic; attribute dont_touch of G16675: signal is true;
	signal G16676: std_logic; attribute dont_touch of G16676: signal is true;
	signal G16677: std_logic; attribute dont_touch of G16677: signal is true;
	signal G16680: std_logic; attribute dont_touch of G16680: signal is true;
	signal G16681: std_logic; attribute dont_touch of G16681: signal is true;
	signal G16684: std_logic; attribute dont_touch of G16684: signal is true;
	signal G16685: std_logic; attribute dont_touch of G16685: signal is true;
	signal G16687: std_logic; attribute dont_touch of G16687: signal is true;
	signal G16688: std_logic; attribute dont_touch of G16688: signal is true;
	signal G16689: std_logic; attribute dont_touch of G16689: signal is true;
	signal G16690: std_logic; attribute dont_touch of G16690: signal is true;
	signal G16691: std_logic; attribute dont_touch of G16691: signal is true;
	signal G16692: std_logic; attribute dont_touch of G16692: signal is true;
	signal G16694: std_logic; attribute dont_touch of G16694: signal is true;
	signal G16695: std_logic; attribute dont_touch of G16695: signal is true;
	signal G16696: std_logic; attribute dont_touch of G16696: signal is true;
	signal G16699: std_logic; attribute dont_touch of G16699: signal is true;
	signal G16700: std_logic; attribute dont_touch of G16700: signal is true;
	signal G16701: std_logic; attribute dont_touch of G16701: signal is true;
	signal G16702: std_logic; attribute dont_touch of G16702: signal is true;
	signal G16703: std_logic; attribute dont_touch of G16703: signal is true;
	signal G16704: std_logic; attribute dont_touch of G16704: signal is true;
	signal G16705: std_logic; attribute dont_touch of G16705: signal is true;
	signal G16706: std_logic; attribute dont_touch of G16706: signal is true;
	signal G16707: std_logic; attribute dont_touch of G16707: signal is true;
	signal G16708: std_logic; attribute dont_touch of G16708: signal is true;
	signal G16709: std_logic; attribute dont_touch of G16709: signal is true;
	signal G16712: std_logic; attribute dont_touch of G16712: signal is true;
	signal G16713: std_logic; attribute dont_touch of G16713: signal is true;
	signal G16716: std_logic; attribute dont_touch of G16716: signal is true;
	signal G16717: std_logic; attribute dont_touch of G16717: signal is true;
	signal G16719: std_logic; attribute dont_touch of G16719: signal is true;
	signal G16720: std_logic; attribute dont_touch of G16720: signal is true;
	signal G16721: std_logic; attribute dont_touch of G16721: signal is true;
	signal G16723: std_logic; attribute dont_touch of G16723: signal is true;
	signal G16724: std_logic; attribute dont_touch of G16724: signal is true;
	signal G16725: std_logic; attribute dont_touch of G16725: signal is true;
	signal G16726: std_logic; attribute dont_touch of G16726: signal is true;
	signal G16727: std_logic; attribute dont_touch of G16727: signal is true;
	signal G16728: std_logic; attribute dont_touch of G16728: signal is true;
	signal G16729: std_logic; attribute dont_touch of G16729: signal is true;
	signal G16730: std_logic; attribute dont_touch of G16730: signal is true;
	signal G16731: std_logic; attribute dont_touch of G16731: signal is true;
	signal G16732: std_logic; attribute dont_touch of G16732: signal is true;
	signal G16733: std_logic; attribute dont_touch of G16733: signal is true;
	signal G16734: std_logic; attribute dont_touch of G16734: signal is true;
	signal G16735: std_logic; attribute dont_touch of G16735: signal is true;
	signal G16736: std_logic; attribute dont_touch of G16736: signal is true;
	signal G16737: std_logic; attribute dont_touch of G16737: signal is true;
	signal G16738: std_logic; attribute dont_touch of G16738: signal is true;
	signal G16739: std_logic; attribute dont_touch of G16739: signal is true;
	signal G16740: std_logic; attribute dont_touch of G16740: signal is true;
	signal G16741: std_logic; attribute dont_touch of G16741: signal is true;
	signal G16742: std_logic; attribute dont_touch of G16742: signal is true;
	signal G16743: std_logic; attribute dont_touch of G16743: signal is true;
	signal G16745: std_logic; attribute dont_touch of G16745: signal is true;
	signal G16746: std_logic; attribute dont_touch of G16746: signal is true;
	signal G16747: std_logic; attribute dont_touch of G16747: signal is true;
	signal G16749: std_logic; attribute dont_touch of G16749: signal is true;
	signal G16750: std_logic; attribute dont_touch of G16750: signal is true;
	signal G16751: std_logic; attribute dont_touch of G16751: signal is true;
	signal G16752: std_logic; attribute dont_touch of G16752: signal is true;
	signal G16757: std_logic; attribute dont_touch of G16757: signal is true;
	signal G16758: std_logic; attribute dont_touch of G16758: signal is true;
	signal G16759: std_logic; attribute dont_touch of G16759: signal is true;
	signal G16760: std_logic; attribute dont_touch of G16760: signal is true;
	signal G16761: std_logic; attribute dont_touch of G16761: signal is true;
	signal G16762: std_logic; attribute dont_touch of G16762: signal is true;
	signal G16763: std_logic; attribute dont_touch of G16763: signal is true;
	signal G16764: std_logic; attribute dont_touch of G16764: signal is true;
	signal G16765: std_logic; attribute dont_touch of G16765: signal is true;
	signal G16766: std_logic; attribute dont_touch of G16766: signal is true;
	signal G16767: std_logic; attribute dont_touch of G16767: signal is true;
	signal G16768: std_logic; attribute dont_touch of G16768: signal is true;
	signal G16769: std_logic; attribute dont_touch of G16769: signal is true;
	signal G16770: std_logic; attribute dont_touch of G16770: signal is true;
	signal G16771: std_logic; attribute dont_touch of G16771: signal is true;
	signal G16772: std_logic; attribute dont_touch of G16772: signal is true;
	signal G16773: std_logic; attribute dont_touch of G16773: signal is true;
	signal G16774: std_logic; attribute dont_touch of G16774: signal is true;
	signal G16776: std_logic; attribute dont_touch of G16776: signal is true;
	signal G16777: std_logic; attribute dont_touch of G16777: signal is true;
	signal G16782: std_logic; attribute dont_touch of G16782: signal is true;
	signal G16795: std_logic; attribute dont_touch of G16795: signal is true;
	signal G16800: std_logic; attribute dont_touch of G16800: signal is true;
	signal G16801: std_logic; attribute dont_touch of G16801: signal is true;
	signal G16802: std_logic; attribute dont_touch of G16802: signal is true;
	signal G16803: std_logic; attribute dont_touch of G16803: signal is true;
	signal G16804: std_logic; attribute dont_touch of G16804: signal is true;
	signal G16805: std_logic; attribute dont_touch of G16805: signal is true;
	signal G16806: std_logic; attribute dont_touch of G16806: signal is true;
	signal G16807: std_logic; attribute dont_touch of G16807: signal is true;
	signal G16808: std_logic; attribute dont_touch of G16808: signal is true;
	signal G16809: std_logic; attribute dont_touch of G16809: signal is true;
	signal G16810: std_logic; attribute dont_touch of G16810: signal is true;
	signal G16811: std_logic; attribute dont_touch of G16811: signal is true;
	signal G16812: std_logic; attribute dont_touch of G16812: signal is true;
	signal G16813: std_logic; attribute dont_touch of G16813: signal is true;
	signal G16814: std_logic; attribute dont_touch of G16814: signal is true;
	signal G16815: std_logic; attribute dont_touch of G16815: signal is true;
	signal G16816: std_logic; attribute dont_touch of G16816: signal is true;
	signal G16821: std_logic; attribute dont_touch of G16821: signal is true;
	signal G16826: std_logic; attribute dont_touch of G16826: signal is true;
	signal G16839: std_logic; attribute dont_touch of G16839: signal is true;
	signal G16840: std_logic; attribute dont_touch of G16840: signal is true;
	signal G16841: std_logic; attribute dont_touch of G16841: signal is true;
	signal G16842: std_logic; attribute dont_touch of G16842: signal is true;
	signal G16843: std_logic; attribute dont_touch of G16843: signal is true;
	signal G16844: std_logic; attribute dont_touch of G16844: signal is true;
	signal G16845: std_logic; attribute dont_touch of G16845: signal is true;
	signal G16846: std_logic; attribute dont_touch of G16846: signal is true;
	signal G16853: std_logic; attribute dont_touch of G16853: signal is true;
	signal G16854: std_logic; attribute dont_touch of G16854: signal is true;
	signal G16855: std_logic; attribute dont_touch of G16855: signal is true;
	signal G16856: std_logic; attribute dont_touch of G16856: signal is true;
	signal G16861: std_logic; attribute dont_touch of G16861: signal is true;
	signal G16866: std_logic; attribute dont_touch of G16866: signal is true;
	signal G16867: std_logic; attribute dont_touch of G16867: signal is true;
	signal G16868: std_logic; attribute dont_touch of G16868: signal is true;
	signal G16869: std_logic; attribute dont_touch of G16869: signal is true;
	signal G16870: std_logic; attribute dont_touch of G16870: signal is true;
	signal G16871: std_logic; attribute dont_touch of G16871: signal is true;
	signal G16872: std_logic; attribute dont_touch of G16872: signal is true;
	signal G16873: std_logic; attribute dont_touch of G16873: signal is true;
	signal G16875: std_logic; attribute dont_touch of G16875: signal is true;
	signal G16876: std_logic; attribute dont_touch of G16876: signal is true;
	signal G16877: std_logic; attribute dont_touch of G16877: signal is true;
	signal G16882: std_logic; attribute dont_touch of G16882: signal is true;
	signal G16883: std_logic; attribute dont_touch of G16883: signal is true;
	signal G16884: std_logic; attribute dont_touch of G16884: signal is true;
	signal G16885: std_logic; attribute dont_touch of G16885: signal is true;
	signal G16886: std_logic; attribute dont_touch of G16886: signal is true;
	signal G16893: std_logic; attribute dont_touch of G16893: signal is true;
	signal G16896: std_logic; attribute dont_touch of G16896: signal is true;
	signal G16897: std_logic; attribute dont_touch of G16897: signal is true;
	signal G16920: std_logic; attribute dont_touch of G16920: signal is true;
	signal G16923: std_logic; attribute dont_touch of G16923: signal is true;
	signal G16925: std_logic; attribute dont_touch of G16925: signal is true;
	signal G16926: std_logic; attribute dont_touch of G16926: signal is true;
	signal G16927: std_logic; attribute dont_touch of G16927: signal is true;
	signal G16928: std_logic; attribute dont_touch of G16928: signal is true;
	signal G16929: std_logic; attribute dont_touch of G16929: signal is true;
	signal G16930: std_logic; attribute dont_touch of G16930: signal is true;
	signal G16931: std_logic; attribute dont_touch of G16931: signal is true;
	signal G16954: std_logic; attribute dont_touch of G16954: signal is true;
	signal G16956: std_logic; attribute dont_touch of G16956: signal is true;
	signal G16957: std_logic; attribute dont_touch of G16957: signal is true;
	signal G16958: std_logic; attribute dont_touch of G16958: signal is true;
	signal G16959: std_logic; attribute dont_touch of G16959: signal is true;
	signal G16960: std_logic; attribute dont_touch of G16960: signal is true;
	signal G16963: std_logic; attribute dont_touch of G16963: signal is true;
	signal G16964: std_logic; attribute dont_touch of G16964: signal is true;
	signal G16965: std_logic; attribute dont_touch of G16965: signal is true;
	signal G16966: std_logic; attribute dont_touch of G16966: signal is true;
	signal G16967: std_logic; attribute dont_touch of G16967: signal is true;
	signal G16968: std_logic; attribute dont_touch of G16968: signal is true;
	signal G16969: std_logic; attribute dont_touch of G16969: signal is true;
	signal G16970: std_logic; attribute dont_touch of G16970: signal is true;
	signal G16971: std_logic; attribute dont_touch of G16971: signal is true;
	signal G16986: std_logic; attribute dont_touch of G16986: signal is true;
	signal G16987: std_logic; attribute dont_touch of G16987: signal is true;
	signal G17010: std_logic; attribute dont_touch of G17010: signal is true;
	signal G17013: std_logic; attribute dont_touch of G17013: signal is true;
	signal G17014: std_logic; attribute dont_touch of G17014: signal is true;
	signal G17015: std_logic; attribute dont_touch of G17015: signal is true;
	signal G17056: std_logic; attribute dont_touch of G17056: signal is true;
	signal G17057: std_logic; attribute dont_touch of G17057: signal is true;
	signal G17058: std_logic; attribute dont_touch of G17058: signal is true;
	signal G17059: std_logic; attribute dont_touch of G17059: signal is true;
	signal G17062: std_logic; attribute dont_touch of G17062: signal is true;
	signal G17085: std_logic; attribute dont_touch of G17085: signal is true;
	signal G17086: std_logic; attribute dont_touch of G17086: signal is true;
	signal G17087: std_logic; attribute dont_touch of G17087: signal is true;
	signal G17088: std_logic; attribute dont_touch of G17088: signal is true;
	signal G17091: std_logic; attribute dont_touch of G17091: signal is true;
	signal G17092: std_logic; attribute dont_touch of G17092: signal is true;
	signal G17093: std_logic; attribute dont_touch of G17093: signal is true;
	signal G17096: std_logic; attribute dont_touch of G17096: signal is true;
	signal G17119: std_logic; attribute dont_touch of G17119: signal is true;
	signal G17120: std_logic; attribute dont_touch of G17120: signal is true;
	signal G17121: std_logic; attribute dont_touch of G17121: signal is true;
	signal G17122: std_logic; attribute dont_touch of G17122: signal is true;
	signal G17123: std_logic; attribute dont_touch of G17123: signal is true;
	signal G17124: std_logic; attribute dont_touch of G17124: signal is true;
	signal G17125: std_logic; attribute dont_touch of G17125: signal is true;
	signal G17128: std_logic; attribute dont_touch of G17128: signal is true;
	signal G17133: std_logic; attribute dont_touch of G17133: signal is true;
	signal G17134: std_logic; attribute dont_touch of G17134: signal is true;
	signal G17135: std_logic; attribute dont_touch of G17135: signal is true;
	signal G17136: std_logic; attribute dont_touch of G17136: signal is true;
	signal G17137: std_logic; attribute dont_touch of G17137: signal is true;
	signal G17138: std_logic; attribute dont_touch of G17138: signal is true;
	signal G17139: std_logic; attribute dont_touch of G17139: signal is true;
	signal G17140: std_logic; attribute dont_touch of G17140: signal is true;
	signal G17141: std_logic; attribute dont_touch of G17141: signal is true;
	signal G17144: std_logic; attribute dont_touch of G17144: signal is true;
	signal G17145: std_logic; attribute dont_touch of G17145: signal is true;
	signal G17146: std_logic; attribute dont_touch of G17146: signal is true;
	signal G17147: std_logic; attribute dont_touch of G17147: signal is true;
	signal G17148: std_logic; attribute dont_touch of G17148: signal is true;
	signal G17149: std_logic; attribute dont_touch of G17149: signal is true;
	signal G17150: std_logic; attribute dont_touch of G17150: signal is true;
	signal G17151: std_logic; attribute dont_touch of G17151: signal is true;
	signal G17152: std_logic; attribute dont_touch of G17152: signal is true;
	signal G17153: std_logic; attribute dont_touch of G17153: signal is true;
	signal G17154: std_logic; attribute dont_touch of G17154: signal is true;
	signal G17155: std_logic; attribute dont_touch of G17155: signal is true;
	signal G17156: std_logic; attribute dont_touch of G17156: signal is true;
	signal G17157: std_logic; attribute dont_touch of G17157: signal is true;
	signal G17174: std_logic; attribute dont_touch of G17174: signal is true;
	signal G17175: std_logic; attribute dont_touch of G17175: signal is true;
	signal G17176: std_logic; attribute dont_touch of G17176: signal is true;
	signal G17177: std_logic; attribute dont_touch of G17177: signal is true;
	signal G17178: std_logic; attribute dont_touch of G17178: signal is true;
	signal G17179: std_logic; attribute dont_touch of G17179: signal is true;
	signal G17180: std_logic; attribute dont_touch of G17180: signal is true;
	signal G17181: std_logic; attribute dont_touch of G17181: signal is true;
	signal G17182: std_logic; attribute dont_touch of G17182: signal is true;
	signal G17183: std_logic; attribute dont_touch of G17183: signal is true;
	signal G17188: std_logic; attribute dont_touch of G17188: signal is true;
	signal G17189: std_logic; attribute dont_touch of G17189: signal is true;
	signal G17190: std_logic; attribute dont_touch of G17190: signal is true;
	signal G17191: std_logic; attribute dont_touch of G17191: signal is true;
	signal G17192: std_logic; attribute dont_touch of G17192: signal is true;
	signal G17193: std_logic; attribute dont_touch of G17193: signal is true;
	signal G17194: std_logic; attribute dont_touch of G17194: signal is true;
	signal G17197: std_logic; attribute dont_touch of G17197: signal is true;
	signal G17198: std_logic; attribute dont_touch of G17198: signal is true;
	signal G17199: std_logic; attribute dont_touch of G17199: signal is true;
	signal G17200: std_logic; attribute dont_touch of G17200: signal is true;
	signal G17213: std_logic; attribute dont_touch of G17213: signal is true;
	signal G17216: std_logic; attribute dont_touch of G17216: signal is true;
	signal G17217: std_logic; attribute dont_touch of G17217: signal is true;
	signal G17220: std_logic; attribute dont_touch of G17220: signal is true;
	signal G17221: std_logic; attribute dont_touch of G17221: signal is true;
	signal G17224: std_logic; attribute dont_touch of G17224: signal is true;
	signal G17225: std_logic; attribute dont_touch of G17225: signal is true;
	signal G17226: std_logic; attribute dont_touch of G17226: signal is true;
	signal G17239: std_logic; attribute dont_touch of G17239: signal is true;
	signal G17242: std_logic; attribute dont_touch of G17242: signal is true;
	signal G17243: std_logic; attribute dont_touch of G17243: signal is true;
	signal G17246: std_logic; attribute dont_touch of G17246: signal is true;
	signal G17247: std_logic; attribute dont_touch of G17247: signal is true;
	signal G17248: std_logic; attribute dont_touch of G17248: signal is true;
	signal G17249: std_logic; attribute dont_touch of G17249: signal is true;
	signal G17264: std_logic; attribute dont_touch of G17264: signal is true;
	signal G17268: std_logic; attribute dont_touch of G17268: signal is true;
	signal G17271: std_logic; attribute dont_touch of G17271: signal is true;
	signal G17284: std_logic; attribute dont_touch of G17284: signal is true;
	signal G17287: std_logic; attribute dont_touch of G17287: signal is true;
	signal G17290: std_logic; attribute dont_touch of G17290: signal is true;
	signal G17292: std_logic; attribute dont_touch of G17292: signal is true;
	signal G17296: std_logic; attribute dont_touch of G17296: signal is true;
	signal G17297: std_logic; attribute dont_touch of G17297: signal is true;
	signal G17301: std_logic; attribute dont_touch of G17301: signal is true;
	signal G17302: std_logic; attribute dont_touch of G17302: signal is true;
	signal G17307: std_logic; attribute dont_touch of G17307: signal is true;
	signal G17308: std_logic; attribute dont_touch of G17308: signal is true;
	signal G17309: std_logic; attribute dont_touch of G17309: signal is true;
	signal G17312: std_logic; attribute dont_touch of G17312: signal is true;
	signal G17315: std_logic; attribute dont_touch of G17315: signal is true;
	signal G17317: std_logic; attribute dont_touch of G17317: signal is true;
	signal G17321: std_logic; attribute dont_touch of G17321: signal is true;
	signal G17324: std_logic; attribute dont_touch of G17324: signal is true;
	signal G17325: std_logic; attribute dont_touch of G17325: signal is true;
	signal G17326: std_logic; attribute dont_touch of G17326: signal is true;
	signal G17327: std_logic; attribute dont_touch of G17327: signal is true;
	signal G17328: std_logic; attribute dont_touch of G17328: signal is true;
	signal G17363: std_logic; attribute dont_touch of G17363: signal is true;
	signal G17364: std_logic; attribute dont_touch of G17364: signal is true;
	signal G17365: std_logic; attribute dont_touch of G17365: signal is true;
	signal G17366: std_logic; attribute dont_touch of G17366: signal is true;
	signal G17367: std_logic; attribute dont_touch of G17367: signal is true;
	signal G17384: std_logic; attribute dont_touch of G17384: signal is true;
	signal G17389: std_logic; attribute dont_touch of G17389: signal is true;
	signal G17390: std_logic; attribute dont_touch of G17390: signal is true;
	signal G17391: std_logic; attribute dont_touch of G17391: signal is true;
	signal G17392: std_logic; attribute dont_touch of G17392: signal is true;
	signal G17393: std_logic; attribute dont_touch of G17393: signal is true;
	signal G17396: std_logic; attribute dont_touch of G17396: signal is true;
	signal G17399: std_logic; attribute dont_touch of G17399: signal is true;
	signal G17401: std_logic; attribute dont_touch of G17401: signal is true;
	signal G17405: std_logic; attribute dont_touch of G17405: signal is true;
	signal G17408: std_logic; attribute dont_touch of G17408: signal is true;
	signal G17409: std_logic; attribute dont_touch of G17409: signal is true;
	signal G17410: std_logic; attribute dont_touch of G17410: signal is true;
	signal G17411: std_logic; attribute dont_touch of G17411: signal is true;
	signal G17412: std_logic; attribute dont_touch of G17412: signal is true;
	signal G17413: std_logic; attribute dont_touch of G17413: signal is true;
	signal G17414: std_logic; attribute dont_touch of G17414: signal is true;
	signal G17415: std_logic; attribute dont_touch of G17415: signal is true;
	signal G17416: std_logic; attribute dont_touch of G17416: signal is true;
	signal G17417: std_logic; attribute dont_touch of G17417: signal is true;
	signal G17418: std_logic; attribute dont_touch of G17418: signal is true;
	signal G17419: std_logic; attribute dont_touch of G17419: signal is true;
	signal G17420: std_logic; attribute dont_touch of G17420: signal is true;
	signal G17424: std_logic; attribute dont_touch of G17424: signal is true;
	signal G17427: std_logic; attribute dont_touch of G17427: signal is true;
	signal G17428: std_logic; attribute dont_touch of G17428: signal is true;
	signal G17429: std_logic; attribute dont_touch of G17429: signal is true;
	signal G17430: std_logic; attribute dont_touch of G17430: signal is true;
	signal G17431: std_logic; attribute dont_touch of G17431: signal is true;
	signal G17432: std_logic; attribute dont_touch of G17432: signal is true;
	signal G17433: std_logic; attribute dont_touch of G17433: signal is true;
	signal G17464: std_logic; attribute dont_touch of G17464: signal is true;
	signal G17465: std_logic; attribute dont_touch of G17465: signal is true;
	signal G17466: std_logic; attribute dont_touch of G17466: signal is true;
	signal G17467: std_logic; attribute dont_touch of G17467: signal is true;
	signal G17468: std_logic; attribute dont_touch of G17468: signal is true;
	signal G17469: std_logic; attribute dont_touch of G17469: signal is true;
	signal G17470: std_logic; attribute dont_touch of G17470: signal is true;
	signal G17471: std_logic; attribute dont_touch of G17471: signal is true;
	signal G17472: std_logic; attribute dont_touch of G17472: signal is true;
	signal G17473: std_logic; attribute dont_touch of G17473: signal is true;
	signal G17474: std_logic; attribute dont_touch of G17474: signal is true;
	signal G17475: std_logic; attribute dont_touch of G17475: signal is true;
	signal G17476: std_logic; attribute dont_touch of G17476: signal is true;
	signal G17477: std_logic; attribute dont_touch of G17477: signal is true;
	signal G17478: std_logic; attribute dont_touch of G17478: signal is true;
	signal G17479: std_logic; attribute dont_touch of G17479: signal is true;
	signal G17480: std_logic; attribute dont_touch of G17480: signal is true;
	signal G17481: std_logic; attribute dont_touch of G17481: signal is true;
	signal G17482: std_logic; attribute dont_touch of G17482: signal is true;
	signal G17485: std_logic; attribute dont_touch of G17485: signal is true;
	signal G17486: std_logic; attribute dont_touch of G17486: signal is true;
	signal G17487: std_logic; attribute dont_touch of G17487: signal is true;
	signal G17488: std_logic; attribute dont_touch of G17488: signal is true;
	signal G17489: std_logic; attribute dont_touch of G17489: signal is true;
	signal G17490: std_logic; attribute dont_touch of G17490: signal is true;
	signal G17491: std_logic; attribute dont_touch of G17491: signal is true;
	signal G17492: std_logic; attribute dont_touch of G17492: signal is true;
	signal G17493: std_logic; attribute dont_touch of G17493: signal is true;
	signal G17494: std_logic; attribute dont_touch of G17494: signal is true;
	signal G17495: std_logic; attribute dont_touch of G17495: signal is true;
	signal G17496: std_logic; attribute dont_touch of G17496: signal is true;
	signal G17497: std_logic; attribute dont_touch of G17497: signal is true;
	signal G17498: std_logic; attribute dont_touch of G17498: signal is true;
	signal G17499: std_logic; attribute dont_touch of G17499: signal is true;
	signal G17500: std_logic; attribute dont_touch of G17500: signal is true;
	signal G17501: std_logic; attribute dont_touch of G17501: signal is true;
	signal G17502: std_logic; attribute dont_touch of G17502: signal is true;
	signal G17503: std_logic; attribute dont_touch of G17503: signal is true;
	signal G17504: std_logic; attribute dont_touch of G17504: signal is true;
	signal G17505: std_logic; attribute dont_touch of G17505: signal is true;
	signal G17506: std_logic; attribute dont_touch of G17506: signal is true;
	signal G17507: std_logic; attribute dont_touch of G17507: signal is true;
	signal G17508: std_logic; attribute dont_touch of G17508: signal is true;
	signal G17509: std_logic; attribute dont_touch of G17509: signal is true;
	signal G17510: std_logic; attribute dont_touch of G17510: signal is true;
	signal G17511: std_logic; attribute dont_touch of G17511: signal is true;
	signal G17512: std_logic; attribute dont_touch of G17512: signal is true;
	signal G17513: std_logic; attribute dont_touch of G17513: signal is true;
	signal G17514: std_logic; attribute dont_touch of G17514: signal is true;
	signal G17515: std_logic; attribute dont_touch of G17515: signal is true;
	signal G17518: std_logic; attribute dont_touch of G17518: signal is true;
	signal G17520: std_logic; attribute dont_touch of G17520: signal is true;
	signal G17521: std_logic; attribute dont_touch of G17521: signal is true;
	signal G17522: std_logic; attribute dont_touch of G17522: signal is true;
	signal G17523: std_logic; attribute dont_touch of G17523: signal is true;
	signal G17524: std_logic; attribute dont_touch of G17524: signal is true;
	signal G17525: std_logic; attribute dont_touch of G17525: signal is true;
	signal G17526: std_logic; attribute dont_touch of G17526: signal is true;
	signal G17527: std_logic; attribute dont_touch of G17527: signal is true;
	signal G17528: std_logic; attribute dont_touch of G17528: signal is true;
	signal G17529: std_logic; attribute dont_touch of G17529: signal is true;
	signal G17530: std_logic; attribute dont_touch of G17530: signal is true;
	signal G17531: std_logic; attribute dont_touch of G17531: signal is true;
	signal G17532: std_logic; attribute dont_touch of G17532: signal is true;
	signal G17533: std_logic; attribute dont_touch of G17533: signal is true;
	signal G17568: std_logic; attribute dont_touch of G17568: signal is true;
	signal G17569: std_logic; attribute dont_touch of G17569: signal is true;
	signal G17570: std_logic; attribute dont_touch of G17570: signal is true;
	signal G17571: std_logic; attribute dont_touch of G17571: signal is true;
	signal G17572: std_logic; attribute dont_touch of G17572: signal is true;
	signal G17573: std_logic; attribute dont_touch of G17573: signal is true;
	signal G17574: std_logic; attribute dont_touch of G17574: signal is true;
	signal G17575: std_logic; attribute dont_touch of G17575: signal is true;
	signal G17576: std_logic; attribute dont_touch of G17576: signal is true;
	signal G17578: std_logic; attribute dont_touch of G17578: signal is true;
	signal G17579: std_logic; attribute dont_touch of G17579: signal is true;
	signal G17581: std_logic; attribute dont_touch of G17581: signal is true;
	signal G17582: std_logic; attribute dont_touch of G17582: signal is true;
	signal G17583: std_logic; attribute dont_touch of G17583: signal is true;
	signal G17584: std_logic; attribute dont_touch of G17584: signal is true;
	signal G17585: std_logic; attribute dont_touch of G17585: signal is true;
	signal G17586: std_logic; attribute dont_touch of G17586: signal is true;
	signal G17587: std_logic; attribute dont_touch of G17587: signal is true;
	signal G17588: std_logic; attribute dont_touch of G17588: signal is true;
	signal G17589: std_logic; attribute dont_touch of G17589: signal is true;
	signal G17590: std_logic; attribute dont_touch of G17590: signal is true;
	signal G17591: std_logic; attribute dont_touch of G17591: signal is true;
	signal G17592: std_logic; attribute dont_touch of G17592: signal is true;
	signal G17593: std_logic; attribute dont_touch of G17593: signal is true;
	signal G17594: std_logic; attribute dont_touch of G17594: signal is true;
	signal G17595: std_logic; attribute dont_touch of G17595: signal is true;
	signal G17596: std_logic; attribute dont_touch of G17596: signal is true;
	signal G17597: std_logic; attribute dont_touch of G17597: signal is true;
	signal G17598: std_logic; attribute dont_touch of G17598: signal is true;
	signal G17599: std_logic; attribute dont_touch of G17599: signal is true;
	signal G17600: std_logic; attribute dont_touch of G17600: signal is true;
	signal G17601: std_logic; attribute dont_touch of G17601: signal is true;
	signal G17602: std_logic; attribute dont_touch of G17602: signal is true;
	signal G17603: std_logic; attribute dont_touch of G17603: signal is true;
	signal G17605: std_logic; attribute dont_touch of G17605: signal is true;
	signal G17606: std_logic; attribute dont_touch of G17606: signal is true;
	signal G17608: std_logic; attribute dont_touch of G17608: signal is true;
	signal G17609: std_logic; attribute dont_touch of G17609: signal is true;
	signal G17610: std_logic; attribute dont_touch of G17610: signal is true;
	signal G17611: std_logic; attribute dont_touch of G17611: signal is true;
	signal G17612: std_logic; attribute dont_touch of G17612: signal is true;
	signal G17613: std_logic; attribute dont_touch of G17613: signal is true;
	signal G17614: std_logic; attribute dont_touch of G17614: signal is true;
	signal G17615: std_logic; attribute dont_touch of G17615: signal is true;
	signal G17616: std_logic; attribute dont_touch of G17616: signal is true;
	signal G17617: std_logic; attribute dont_touch of G17617: signal is true;
	signal G17618: std_logic; attribute dont_touch of G17618: signal is true;
	signal G17619: std_logic; attribute dont_touch of G17619: signal is true;
	signal G17624: std_logic; attribute dont_touch of G17624: signal is true;
	signal G17625: std_logic; attribute dont_touch of G17625: signal is true;
	signal G17634: std_logic; attribute dont_touch of G17634: signal is true;
	signal G17635: std_logic; attribute dont_touch of G17635: signal is true;
	signal G17636: std_logic; attribute dont_touch of G17636: signal is true;
	signal G17637: std_logic; attribute dont_touch of G17637: signal is true;
	signal G17638: std_logic; attribute dont_touch of G17638: signal is true;
	signal G17640: std_logic; attribute dont_touch of G17640: signal is true;
	signal G17641: std_logic; attribute dont_touch of G17641: signal is true;
	signal G17642: std_logic; attribute dont_touch of G17642: signal is true;
	signal G17643: std_logic; attribute dont_touch of G17643: signal is true;
	signal G17644: std_logic; attribute dont_touch of G17644: signal is true;
	signal G17645: std_logic; attribute dont_touch of G17645: signal is true;
	signal G17647: std_logic; attribute dont_touch of G17647: signal is true;
	signal G17648: std_logic; attribute dont_touch of G17648: signal is true;
	signal G17650: std_logic; attribute dont_touch of G17650: signal is true;
	signal G17651: std_logic; attribute dont_touch of G17651: signal is true;
	signal G17652: std_logic; attribute dont_touch of G17652: signal is true;
	signal G17653: std_logic; attribute dont_touch of G17653: signal is true;
	signal G17654: std_logic; attribute dont_touch of G17654: signal is true;
	signal G17655: std_logic; attribute dont_touch of G17655: signal is true;
	signal G17656: std_logic; attribute dont_touch of G17656: signal is true;
	signal G17657: std_logic; attribute dont_touch of G17657: signal is true;
	signal G17662: std_logic; attribute dont_touch of G17662: signal is true;
	signal G17663: std_logic; attribute dont_touch of G17663: signal is true;
	signal G17668: std_logic; attribute dont_touch of G17668: signal is true;
	signal G17669: std_logic; attribute dont_touch of G17669: signal is true;
	signal G17670: std_logic; attribute dont_touch of G17670: signal is true;
	signal G17671: std_logic; attribute dont_touch of G17671: signal is true;
	signal G17672: std_logic; attribute dont_touch of G17672: signal is true;
	signal G17673: std_logic; attribute dont_touch of G17673: signal is true;
	signal G17675: std_logic; attribute dont_touch of G17675: signal is true;
	signal G17676: std_logic; attribute dont_touch of G17676: signal is true;
	signal G17677: std_logic; attribute dont_touch of G17677: signal is true;
	signal G17679: std_logic; attribute dont_touch of G17679: signal is true;
	signal G17680: std_logic; attribute dont_touch of G17680: signal is true;
	signal G17681: std_logic; attribute dont_touch of G17681: signal is true;
	signal G17682: std_logic; attribute dont_touch of G17682: signal is true;
	signal G17683: std_logic; attribute dont_touch of G17683: signal is true;
	signal G17684: std_logic; attribute dont_touch of G17684: signal is true;
	signal G17686: std_logic; attribute dont_touch of G17686: signal is true;
	signal G17687: std_logic; attribute dont_touch of G17687: signal is true;
	signal G17689: std_logic; attribute dont_touch of G17689: signal is true;
	signal G17690: std_logic; attribute dont_touch of G17690: signal is true;
	signal G17691: std_logic; attribute dont_touch of G17691: signal is true;
	signal G17692: std_logic; attribute dont_touch of G17692: signal is true;
	signal G17693: std_logic; attribute dont_touch of G17693: signal is true;
	signal G17694: std_logic; attribute dont_touch of G17694: signal is true;
	signal G17699: std_logic; attribute dont_touch of G17699: signal is true;
	signal G17700: std_logic; attribute dont_touch of G17700: signal is true;
	signal G17705: std_logic; attribute dont_touch of G17705: signal is true;
	signal G17706: std_logic; attribute dont_touch of G17706: signal is true;
	signal G17707: std_logic; attribute dont_touch of G17707: signal is true;
	signal G17708: std_logic; attribute dont_touch of G17708: signal is true;
	signal G17709: std_logic; attribute dont_touch of G17709: signal is true;
	signal G17710: std_logic; attribute dont_touch of G17710: signal is true;
	signal G17712: std_logic; attribute dont_touch of G17712: signal is true;
	signal G17713: std_logic; attribute dont_touch of G17713: signal is true;
	signal G17714: std_logic; attribute dont_touch of G17714: signal is true;
	signal G17716: std_logic; attribute dont_touch of G17716: signal is true;
	signal G17717: std_logic; attribute dont_touch of G17717: signal is true;
	signal G17718: std_logic; attribute dont_touch of G17718: signal is true;
	signal G17719: std_logic; attribute dont_touch of G17719: signal is true;
	signal G17720: std_logic; attribute dont_touch of G17720: signal is true;
	signal G17721: std_logic; attribute dont_touch of G17721: signal is true;
	signal G17723: std_logic; attribute dont_touch of G17723: signal is true;
	signal G17724: std_logic; attribute dont_touch of G17724: signal is true;
	signal G17725: std_logic; attribute dont_touch of G17725: signal is true;
	signal G17726: std_logic; attribute dont_touch of G17726: signal is true;
	signal G17727: std_logic; attribute dont_touch of G17727: signal is true;
	signal G17732: std_logic; attribute dont_touch of G17732: signal is true;
	signal G17733: std_logic; attribute dont_touch of G17733: signal is true;
	signal G17734: std_logic; attribute dont_touch of G17734: signal is true;
	signal G17735: std_logic; attribute dont_touch of G17735: signal is true;
	signal G17736: std_logic; attribute dont_touch of G17736: signal is true;
	signal G17737: std_logic; attribute dont_touch of G17737: signal is true;
	signal G17738: std_logic; attribute dont_touch of G17738: signal is true;
	signal G17740: std_logic; attribute dont_touch of G17740: signal is true;
	signal G17741: std_logic; attribute dont_touch of G17741: signal is true;
	signal G17742: std_logic; attribute dont_touch of G17742: signal is true;
	signal G17744: std_logic; attribute dont_touch of G17744: signal is true;
	signal G17745: std_logic; attribute dont_touch of G17745: signal is true;
	signal G17746: std_logic; attribute dont_touch of G17746: signal is true;
	signal G17747: std_logic; attribute dont_touch of G17747: signal is true;
	signal G17748: std_logic; attribute dont_touch of G17748: signal is true;
	signal G17752: std_logic; attribute dont_touch of G17752: signal is true;
	signal G17753: std_logic; attribute dont_touch of G17753: signal is true;
	signal G17754: std_logic; attribute dont_touch of G17754: signal is true;
	signal G17755: std_logic; attribute dont_touch of G17755: signal is true;
	signal G17756: std_logic; attribute dont_touch of G17756: signal is true;
	signal G17757: std_logic; attribute dont_touch of G17757: signal is true;
	signal G17758: std_logic; attribute dont_touch of G17758: signal is true;
	signal G17759: std_logic; attribute dont_touch of G17759: signal is true;
	signal G17761: std_logic; attribute dont_touch of G17761: signal is true;
	signal G17762: std_logic; attribute dont_touch of G17762: signal is true;
	signal G17763: std_logic; attribute dont_touch of G17763: signal is true;
	signal G17765: std_logic; attribute dont_touch of G17765: signal is true;
	signal G17766: std_logic; attribute dont_touch of G17766: signal is true;
	signal G17767: std_logic; attribute dont_touch of G17767: signal is true;
	signal G17768: std_logic; attribute dont_touch of G17768: signal is true;
	signal G17769: std_logic; attribute dont_touch of G17769: signal is true;
	signal G17770: std_logic; attribute dont_touch of G17770: signal is true;
	signal G17771: std_logic; attribute dont_touch of G17771: signal is true;
	signal G17772: std_logic; attribute dont_touch of G17772: signal is true;
	signal G17773: std_logic; attribute dont_touch of G17773: signal is true;
	signal G17774: std_logic; attribute dont_touch of G17774: signal is true;
	signal G17775: std_logic; attribute dont_touch of G17775: signal is true;
	signal G17776: std_logic; attribute dont_touch of G17776: signal is true;
	signal G17777: std_logic; attribute dont_touch of G17777: signal is true;
	signal G17779: std_logic; attribute dont_touch of G17779: signal is true;
	signal G17780: std_logic; attribute dont_touch of G17780: signal is true;
	signal G17781: std_logic; attribute dont_touch of G17781: signal is true;
	signal G17782: std_logic; attribute dont_touch of G17782: signal is true;
	signal G17783: std_logic; attribute dont_touch of G17783: signal is true;
	signal G17784: std_logic; attribute dont_touch of G17784: signal is true;
	signal G17785: std_logic; attribute dont_touch of G17785: signal is true;
	signal G17786: std_logic; attribute dont_touch of G17786: signal is true;
	signal G17788: std_logic; attribute dont_touch of G17788: signal is true;
	signal G17789: std_logic; attribute dont_touch of G17789: signal is true;
	signal G17790: std_logic; attribute dont_touch of G17790: signal is true;
	signal G17791: std_logic; attribute dont_touch of G17791: signal is true;
	signal G17792: std_logic; attribute dont_touch of G17792: signal is true;
	signal G17793: std_logic; attribute dont_touch of G17793: signal is true;
	signal G17794: std_logic; attribute dont_touch of G17794: signal is true;
	signal G17809: std_logic; attribute dont_touch of G17809: signal is true;
	signal G17810: std_logic; attribute dont_touch of G17810: signal is true;
	signal G17811: std_logic; attribute dont_touch of G17811: signal is true;
	signal G17812: std_logic; attribute dont_touch of G17812: signal is true;
	signal G17814: std_logic; attribute dont_touch of G17814: signal is true;
	signal G17815: std_logic; attribute dont_touch of G17815: signal is true;
	signal G17816: std_logic; attribute dont_touch of G17816: signal is true;
	signal G17817: std_logic; attribute dont_touch of G17817: signal is true;
	signal G17818: std_logic; attribute dont_touch of G17818: signal is true;
	signal G17820: std_logic; attribute dont_touch of G17820: signal is true;
	signal G17821: std_logic; attribute dont_touch of G17821: signal is true;
	signal G17844: std_logic; attribute dont_touch of G17844: signal is true;
	signal G17846: std_logic; attribute dont_touch of G17846: signal is true;
	signal G17847: std_logic; attribute dont_touch of G17847: signal is true;
	signal G17870: std_logic; attribute dont_touch of G17870: signal is true;
	signal G17872: std_logic; attribute dont_touch of G17872: signal is true;
	signal G17873: std_logic; attribute dont_touch of G17873: signal is true;
	signal G17926: std_logic; attribute dont_touch of G17926: signal is true;
	signal G17929: std_logic; attribute dont_touch of G17929: signal is true;
	signal G17952: std_logic; attribute dont_touch of G17952: signal is true;
	signal G17953: std_logic; attribute dont_touch of G17953: signal is true;
	signal G17954: std_logic; attribute dont_touch of G17954: signal is true;
	signal G17955: std_logic; attribute dont_touch of G17955: signal is true;
	signal G18008: std_logic; attribute dont_touch of G18008: signal is true;
	signal G18061: std_logic; attribute dont_touch of G18061: signal is true;
	signal G18062: std_logic; attribute dont_touch of G18062: signal is true;
	signal G18065: std_logic; attribute dont_touch of G18065: signal is true;
	signal G18088: std_logic; attribute dont_touch of G18088: signal is true;
	signal G18091: std_logic; attribute dont_touch of G18091: signal is true;
	signal G18093: std_logic; attribute dont_touch of G18093: signal is true;
	signal G18102: std_logic; attribute dont_touch of G18102: signal is true;
	signal G18103: std_logic; attribute dont_touch of G18103: signal is true;
	signal G18104: std_logic; attribute dont_touch of G18104: signal is true;
	signal G18105: std_logic; attribute dont_touch of G18105: signal is true;
	signal G18106: std_logic; attribute dont_touch of G18106: signal is true;
	signal G18107: std_logic; attribute dont_touch of G18107: signal is true;
	signal G18108: std_logic; attribute dont_touch of G18108: signal is true;
	signal G18109: std_logic; attribute dont_touch of G18109: signal is true;
	signal G18110: std_logic; attribute dont_touch of G18110: signal is true;
	signal G18111: std_logic; attribute dont_touch of G18111: signal is true;
	signal G18112: std_logic; attribute dont_touch of G18112: signal is true;
	signal G18113: std_logic; attribute dont_touch of G18113: signal is true;
	signal G18114: std_logic; attribute dont_touch of G18114: signal is true;
	signal G18115: std_logic; attribute dont_touch of G18115: signal is true;
	signal G18116: std_logic; attribute dont_touch of G18116: signal is true;
	signal G18117: std_logic; attribute dont_touch of G18117: signal is true;
	signal G18118: std_logic; attribute dont_touch of G18118: signal is true;
	signal G18119: std_logic; attribute dont_touch of G18119: signal is true;
	signal G18120: std_logic; attribute dont_touch of G18120: signal is true;
	signal G18121: std_logic; attribute dont_touch of G18121: signal is true;
	signal G18122: std_logic; attribute dont_touch of G18122: signal is true;
	signal G18123: std_logic; attribute dont_touch of G18123: signal is true;
	signal G18124: std_logic; attribute dont_touch of G18124: signal is true;
	signal G18125: std_logic; attribute dont_touch of G18125: signal is true;
	signal G18126: std_logic; attribute dont_touch of G18126: signal is true;
	signal G18127: std_logic; attribute dont_touch of G18127: signal is true;
	signal G18128: std_logic; attribute dont_touch of G18128: signal is true;
	signal G18129: std_logic; attribute dont_touch of G18129: signal is true;
	signal G18130: std_logic; attribute dont_touch of G18130: signal is true;
	signal G18131: std_logic; attribute dont_touch of G18131: signal is true;
	signal G18132: std_logic; attribute dont_touch of G18132: signal is true;
	signal G18133: std_logic; attribute dont_touch of G18133: signal is true;
	signal G18134: std_logic; attribute dont_touch of G18134: signal is true;
	signal G18135: std_logic; attribute dont_touch of G18135: signal is true;
	signal G18136: std_logic; attribute dont_touch of G18136: signal is true;
	signal G18137: std_logic; attribute dont_touch of G18137: signal is true;
	signal G18138: std_logic; attribute dont_touch of G18138: signal is true;
	signal G18139: std_logic; attribute dont_touch of G18139: signal is true;
	signal G18140: std_logic; attribute dont_touch of G18140: signal is true;
	signal G18141: std_logic; attribute dont_touch of G18141: signal is true;
	signal G18142: std_logic; attribute dont_touch of G18142: signal is true;
	signal G18143: std_logic; attribute dont_touch of G18143: signal is true;
	signal G18144: std_logic; attribute dont_touch of G18144: signal is true;
	signal G18145: std_logic; attribute dont_touch of G18145: signal is true;
	signal G18146: std_logic; attribute dont_touch of G18146: signal is true;
	signal G18147: std_logic; attribute dont_touch of G18147: signal is true;
	signal G18148: std_logic; attribute dont_touch of G18148: signal is true;
	signal G18149: std_logic; attribute dont_touch of G18149: signal is true;
	signal G18150: std_logic; attribute dont_touch of G18150: signal is true;
	signal G18151: std_logic; attribute dont_touch of G18151: signal is true;
	signal G18152: std_logic; attribute dont_touch of G18152: signal is true;
	signal G18153: std_logic; attribute dont_touch of G18153: signal is true;
	signal G18154: std_logic; attribute dont_touch of G18154: signal is true;
	signal G18155: std_logic; attribute dont_touch of G18155: signal is true;
	signal G18156: std_logic; attribute dont_touch of G18156: signal is true;
	signal G18157: std_logic; attribute dont_touch of G18157: signal is true;
	signal G18158: std_logic; attribute dont_touch of G18158: signal is true;
	signal G18159: std_logic; attribute dont_touch of G18159: signal is true;
	signal G18160: std_logic; attribute dont_touch of G18160: signal is true;
	signal G18161: std_logic; attribute dont_touch of G18161: signal is true;
	signal G18162: std_logic; attribute dont_touch of G18162: signal is true;
	signal G18163: std_logic; attribute dont_touch of G18163: signal is true;
	signal G18164: std_logic; attribute dont_touch of G18164: signal is true;
	signal G18165: std_logic; attribute dont_touch of G18165: signal is true;
	signal G18166: std_logic; attribute dont_touch of G18166: signal is true;
	signal G18167: std_logic; attribute dont_touch of G18167: signal is true;
	signal G18168: std_logic; attribute dont_touch of G18168: signal is true;
	signal G18169: std_logic; attribute dont_touch of G18169: signal is true;
	signal G18170: std_logic; attribute dont_touch of G18170: signal is true;
	signal G18171: std_logic; attribute dont_touch of G18171: signal is true;
	signal G18172: std_logic; attribute dont_touch of G18172: signal is true;
	signal G18173: std_logic; attribute dont_touch of G18173: signal is true;
	signal G18174: std_logic; attribute dont_touch of G18174: signal is true;
	signal G18175: std_logic; attribute dont_touch of G18175: signal is true;
	signal G18176: std_logic; attribute dont_touch of G18176: signal is true;
	signal G18177: std_logic; attribute dont_touch of G18177: signal is true;
	signal G18178: std_logic; attribute dont_touch of G18178: signal is true;
	signal G18179: std_logic; attribute dont_touch of G18179: signal is true;
	signal G18180: std_logic; attribute dont_touch of G18180: signal is true;
	signal G18181: std_logic; attribute dont_touch of G18181: signal is true;
	signal G18182: std_logic; attribute dont_touch of G18182: signal is true;
	signal G18183: std_logic; attribute dont_touch of G18183: signal is true;
	signal G18184: std_logic; attribute dont_touch of G18184: signal is true;
	signal G18185: std_logic; attribute dont_touch of G18185: signal is true;
	signal G18186: std_logic; attribute dont_touch of G18186: signal is true;
	signal G18187: std_logic; attribute dont_touch of G18187: signal is true;
	signal G18188: std_logic; attribute dont_touch of G18188: signal is true;
	signal G18189: std_logic; attribute dont_touch of G18189: signal is true;
	signal G18190: std_logic; attribute dont_touch of G18190: signal is true;
	signal G18191: std_logic; attribute dont_touch of G18191: signal is true;
	signal G18192: std_logic; attribute dont_touch of G18192: signal is true;
	signal G18193: std_logic; attribute dont_touch of G18193: signal is true;
	signal G18194: std_logic; attribute dont_touch of G18194: signal is true;
	signal G18195: std_logic; attribute dont_touch of G18195: signal is true;
	signal G18196: std_logic; attribute dont_touch of G18196: signal is true;
	signal G18197: std_logic; attribute dont_touch of G18197: signal is true;
	signal G18198: std_logic; attribute dont_touch of G18198: signal is true;
	signal G18199: std_logic; attribute dont_touch of G18199: signal is true;
	signal G18200: std_logic; attribute dont_touch of G18200: signal is true;
	signal G18201: std_logic; attribute dont_touch of G18201: signal is true;
	signal G18202: std_logic; attribute dont_touch of G18202: signal is true;
	signal G18203: std_logic; attribute dont_touch of G18203: signal is true;
	signal G18204: std_logic; attribute dont_touch of G18204: signal is true;
	signal G18205: std_logic; attribute dont_touch of G18205: signal is true;
	signal G18206: std_logic; attribute dont_touch of G18206: signal is true;
	signal G18207: std_logic; attribute dont_touch of G18207: signal is true;
	signal G18208: std_logic; attribute dont_touch of G18208: signal is true;
	signal G18209: std_logic; attribute dont_touch of G18209: signal is true;
	signal G18210: std_logic; attribute dont_touch of G18210: signal is true;
	signal G18211: std_logic; attribute dont_touch of G18211: signal is true;
	signal G18212: std_logic; attribute dont_touch of G18212: signal is true;
	signal G18213: std_logic; attribute dont_touch of G18213: signal is true;
	signal G18214: std_logic; attribute dont_touch of G18214: signal is true;
	signal G18215: std_logic; attribute dont_touch of G18215: signal is true;
	signal G18216: std_logic; attribute dont_touch of G18216: signal is true;
	signal G18217: std_logic; attribute dont_touch of G18217: signal is true;
	signal G18218: std_logic; attribute dont_touch of G18218: signal is true;
	signal G18219: std_logic; attribute dont_touch of G18219: signal is true;
	signal G18220: std_logic; attribute dont_touch of G18220: signal is true;
	signal G18221: std_logic; attribute dont_touch of G18221: signal is true;
	signal G18222: std_logic; attribute dont_touch of G18222: signal is true;
	signal G18223: std_logic; attribute dont_touch of G18223: signal is true;
	signal G18224: std_logic; attribute dont_touch of G18224: signal is true;
	signal G18225: std_logic; attribute dont_touch of G18225: signal is true;
	signal G18226: std_logic; attribute dont_touch of G18226: signal is true;
	signal G18227: std_logic; attribute dont_touch of G18227: signal is true;
	signal G18228: std_logic; attribute dont_touch of G18228: signal is true;
	signal G18229: std_logic; attribute dont_touch of G18229: signal is true;
	signal G18230: std_logic; attribute dont_touch of G18230: signal is true;
	signal G18231: std_logic; attribute dont_touch of G18231: signal is true;
	signal G18232: std_logic; attribute dont_touch of G18232: signal is true;
	signal G18233: std_logic; attribute dont_touch of G18233: signal is true;
	signal G18234: std_logic; attribute dont_touch of G18234: signal is true;
	signal G18235: std_logic; attribute dont_touch of G18235: signal is true;
	signal G18236: std_logic; attribute dont_touch of G18236: signal is true;
	signal G18237: std_logic; attribute dont_touch of G18237: signal is true;
	signal G18238: std_logic; attribute dont_touch of G18238: signal is true;
	signal G18239: std_logic; attribute dont_touch of G18239: signal is true;
	signal G18240: std_logic; attribute dont_touch of G18240: signal is true;
	signal G18241: std_logic; attribute dont_touch of G18241: signal is true;
	signal G18242: std_logic; attribute dont_touch of G18242: signal is true;
	signal G18243: std_logic; attribute dont_touch of G18243: signal is true;
	signal G18244: std_logic; attribute dont_touch of G18244: signal is true;
	signal G18245: std_logic; attribute dont_touch of G18245: signal is true;
	signal G18246: std_logic; attribute dont_touch of G18246: signal is true;
	signal G18247: std_logic; attribute dont_touch of G18247: signal is true;
	signal G18248: std_logic; attribute dont_touch of G18248: signal is true;
	signal G18249: std_logic; attribute dont_touch of G18249: signal is true;
	signal G18250: std_logic; attribute dont_touch of G18250: signal is true;
	signal G18251: std_logic; attribute dont_touch of G18251: signal is true;
	signal G18252: std_logic; attribute dont_touch of G18252: signal is true;
	signal G18253: std_logic; attribute dont_touch of G18253: signal is true;
	signal G18254: std_logic; attribute dont_touch of G18254: signal is true;
	signal G18255: std_logic; attribute dont_touch of G18255: signal is true;
	signal G18256: std_logic; attribute dont_touch of G18256: signal is true;
	signal G18257: std_logic; attribute dont_touch of G18257: signal is true;
	signal G18258: std_logic; attribute dont_touch of G18258: signal is true;
	signal G18259: std_logic; attribute dont_touch of G18259: signal is true;
	signal G18260: std_logic; attribute dont_touch of G18260: signal is true;
	signal G18261: std_logic; attribute dont_touch of G18261: signal is true;
	signal G18262: std_logic; attribute dont_touch of G18262: signal is true;
	signal G18263: std_logic; attribute dont_touch of G18263: signal is true;
	signal G18264: std_logic; attribute dont_touch of G18264: signal is true;
	signal G18265: std_logic; attribute dont_touch of G18265: signal is true;
	signal G18266: std_logic; attribute dont_touch of G18266: signal is true;
	signal G18267: std_logic; attribute dont_touch of G18267: signal is true;
	signal G18268: std_logic; attribute dont_touch of G18268: signal is true;
	signal G18269: std_logic; attribute dont_touch of G18269: signal is true;
	signal G18270: std_logic; attribute dont_touch of G18270: signal is true;
	signal G18271: std_logic; attribute dont_touch of G18271: signal is true;
	signal G18272: std_logic; attribute dont_touch of G18272: signal is true;
	signal G18273: std_logic; attribute dont_touch of G18273: signal is true;
	signal G18274: std_logic; attribute dont_touch of G18274: signal is true;
	signal G18275: std_logic; attribute dont_touch of G18275: signal is true;
	signal G18276: std_logic; attribute dont_touch of G18276: signal is true;
	signal G18277: std_logic; attribute dont_touch of G18277: signal is true;
	signal G18278: std_logic; attribute dont_touch of G18278: signal is true;
	signal G18279: std_logic; attribute dont_touch of G18279: signal is true;
	signal G18280: std_logic; attribute dont_touch of G18280: signal is true;
	signal G18281: std_logic; attribute dont_touch of G18281: signal is true;
	signal G18282: std_logic; attribute dont_touch of G18282: signal is true;
	signal G18283: std_logic; attribute dont_touch of G18283: signal is true;
	signal G18284: std_logic; attribute dont_touch of G18284: signal is true;
	signal G18285: std_logic; attribute dont_touch of G18285: signal is true;
	signal G18286: std_logic; attribute dont_touch of G18286: signal is true;
	signal G18287: std_logic; attribute dont_touch of G18287: signal is true;
	signal G18288: std_logic; attribute dont_touch of G18288: signal is true;
	signal G18289: std_logic; attribute dont_touch of G18289: signal is true;
	signal G18290: std_logic; attribute dont_touch of G18290: signal is true;
	signal G18291: std_logic; attribute dont_touch of G18291: signal is true;
	signal G18292: std_logic; attribute dont_touch of G18292: signal is true;
	signal G18293: std_logic; attribute dont_touch of G18293: signal is true;
	signal G18294: std_logic; attribute dont_touch of G18294: signal is true;
	signal G18295: std_logic; attribute dont_touch of G18295: signal is true;
	signal G18296: std_logic; attribute dont_touch of G18296: signal is true;
	signal G18297: std_logic; attribute dont_touch of G18297: signal is true;
	signal G18298: std_logic; attribute dont_touch of G18298: signal is true;
	signal G18299: std_logic; attribute dont_touch of G18299: signal is true;
	signal G18300: std_logic; attribute dont_touch of G18300: signal is true;
	signal G18301: std_logic; attribute dont_touch of G18301: signal is true;
	signal G18302: std_logic; attribute dont_touch of G18302: signal is true;
	signal G18303: std_logic; attribute dont_touch of G18303: signal is true;
	signal G18304: std_logic; attribute dont_touch of G18304: signal is true;
	signal G18305: std_logic; attribute dont_touch of G18305: signal is true;
	signal G18306: std_logic; attribute dont_touch of G18306: signal is true;
	signal G18307: std_logic; attribute dont_touch of G18307: signal is true;
	signal G18308: std_logic; attribute dont_touch of G18308: signal is true;
	signal G18309: std_logic; attribute dont_touch of G18309: signal is true;
	signal G18310: std_logic; attribute dont_touch of G18310: signal is true;
	signal G18311: std_logic; attribute dont_touch of G18311: signal is true;
	signal G18312: std_logic; attribute dont_touch of G18312: signal is true;
	signal G18313: std_logic; attribute dont_touch of G18313: signal is true;
	signal G18314: std_logic; attribute dont_touch of G18314: signal is true;
	signal G18315: std_logic; attribute dont_touch of G18315: signal is true;
	signal G18316: std_logic; attribute dont_touch of G18316: signal is true;
	signal G18317: std_logic; attribute dont_touch of G18317: signal is true;
	signal G18318: std_logic; attribute dont_touch of G18318: signal is true;
	signal G18319: std_logic; attribute dont_touch of G18319: signal is true;
	signal G18320: std_logic; attribute dont_touch of G18320: signal is true;
	signal G18321: std_logic; attribute dont_touch of G18321: signal is true;
	signal G18322: std_logic; attribute dont_touch of G18322: signal is true;
	signal G18323: std_logic; attribute dont_touch of G18323: signal is true;
	signal G18324: std_logic; attribute dont_touch of G18324: signal is true;
	signal G18325: std_logic; attribute dont_touch of G18325: signal is true;
	signal G18326: std_logic; attribute dont_touch of G18326: signal is true;
	signal G18327: std_logic; attribute dont_touch of G18327: signal is true;
	signal G18328: std_logic; attribute dont_touch of G18328: signal is true;
	signal G18329: std_logic; attribute dont_touch of G18329: signal is true;
	signal G18330: std_logic; attribute dont_touch of G18330: signal is true;
	signal G18331: std_logic; attribute dont_touch of G18331: signal is true;
	signal G18332: std_logic; attribute dont_touch of G18332: signal is true;
	signal G18333: std_logic; attribute dont_touch of G18333: signal is true;
	signal G18334: std_logic; attribute dont_touch of G18334: signal is true;
	signal G18335: std_logic; attribute dont_touch of G18335: signal is true;
	signal G18336: std_logic; attribute dont_touch of G18336: signal is true;
	signal G18337: std_logic; attribute dont_touch of G18337: signal is true;
	signal G18338: std_logic; attribute dont_touch of G18338: signal is true;
	signal G18339: std_logic; attribute dont_touch of G18339: signal is true;
	signal G18340: std_logic; attribute dont_touch of G18340: signal is true;
	signal G18341: std_logic; attribute dont_touch of G18341: signal is true;
	signal G18342: std_logic; attribute dont_touch of G18342: signal is true;
	signal G18343: std_logic; attribute dont_touch of G18343: signal is true;
	signal G18344: std_logic; attribute dont_touch of G18344: signal is true;
	signal G18345: std_logic; attribute dont_touch of G18345: signal is true;
	signal G18346: std_logic; attribute dont_touch of G18346: signal is true;
	signal G18347: std_logic; attribute dont_touch of G18347: signal is true;
	signal G18348: std_logic; attribute dont_touch of G18348: signal is true;
	signal G18349: std_logic; attribute dont_touch of G18349: signal is true;
	signal G18350: std_logic; attribute dont_touch of G18350: signal is true;
	signal G18351: std_logic; attribute dont_touch of G18351: signal is true;
	signal G18352: std_logic; attribute dont_touch of G18352: signal is true;
	signal G18353: std_logic; attribute dont_touch of G18353: signal is true;
	signal G18354: std_logic; attribute dont_touch of G18354: signal is true;
	signal G18355: std_logic; attribute dont_touch of G18355: signal is true;
	signal G18356: std_logic; attribute dont_touch of G18356: signal is true;
	signal G18357: std_logic; attribute dont_touch of G18357: signal is true;
	signal G18358: std_logic; attribute dont_touch of G18358: signal is true;
	signal G18359: std_logic; attribute dont_touch of G18359: signal is true;
	signal G18360: std_logic; attribute dont_touch of G18360: signal is true;
	signal G18361: std_logic; attribute dont_touch of G18361: signal is true;
	signal G18362: std_logic; attribute dont_touch of G18362: signal is true;
	signal G18363: std_logic; attribute dont_touch of G18363: signal is true;
	signal G18364: std_logic; attribute dont_touch of G18364: signal is true;
	signal G18365: std_logic; attribute dont_touch of G18365: signal is true;
	signal G18366: std_logic; attribute dont_touch of G18366: signal is true;
	signal G18367: std_logic; attribute dont_touch of G18367: signal is true;
	signal G18368: std_logic; attribute dont_touch of G18368: signal is true;
	signal G18369: std_logic; attribute dont_touch of G18369: signal is true;
	signal G18370: std_logic; attribute dont_touch of G18370: signal is true;
	signal G18371: std_logic; attribute dont_touch of G18371: signal is true;
	signal G18372: std_logic; attribute dont_touch of G18372: signal is true;
	signal G18373: std_logic; attribute dont_touch of G18373: signal is true;
	signal G18374: std_logic; attribute dont_touch of G18374: signal is true;
	signal G18375: std_logic; attribute dont_touch of G18375: signal is true;
	signal G18376: std_logic; attribute dont_touch of G18376: signal is true;
	signal G18377: std_logic; attribute dont_touch of G18377: signal is true;
	signal G18378: std_logic; attribute dont_touch of G18378: signal is true;
	signal G18379: std_logic; attribute dont_touch of G18379: signal is true;
	signal G18380: std_logic; attribute dont_touch of G18380: signal is true;
	signal G18381: std_logic; attribute dont_touch of G18381: signal is true;
	signal G18382: std_logic; attribute dont_touch of G18382: signal is true;
	signal G18383: std_logic; attribute dont_touch of G18383: signal is true;
	signal G18384: std_logic; attribute dont_touch of G18384: signal is true;
	signal G18385: std_logic; attribute dont_touch of G18385: signal is true;
	signal G18386: std_logic; attribute dont_touch of G18386: signal is true;
	signal G18387: std_logic; attribute dont_touch of G18387: signal is true;
	signal G18388: std_logic; attribute dont_touch of G18388: signal is true;
	signal G18389: std_logic; attribute dont_touch of G18389: signal is true;
	signal G18390: std_logic; attribute dont_touch of G18390: signal is true;
	signal G18391: std_logic; attribute dont_touch of G18391: signal is true;
	signal G18392: std_logic; attribute dont_touch of G18392: signal is true;
	signal G18393: std_logic; attribute dont_touch of G18393: signal is true;
	signal G18394: std_logic; attribute dont_touch of G18394: signal is true;
	signal G18395: std_logic; attribute dont_touch of G18395: signal is true;
	signal G18396: std_logic; attribute dont_touch of G18396: signal is true;
	signal G18397: std_logic; attribute dont_touch of G18397: signal is true;
	signal G18398: std_logic; attribute dont_touch of G18398: signal is true;
	signal G18399: std_logic; attribute dont_touch of G18399: signal is true;
	signal G18400: std_logic; attribute dont_touch of G18400: signal is true;
	signal G18401: std_logic; attribute dont_touch of G18401: signal is true;
	signal G18402: std_logic; attribute dont_touch of G18402: signal is true;
	signal G18403: std_logic; attribute dont_touch of G18403: signal is true;
	signal G18404: std_logic; attribute dont_touch of G18404: signal is true;
	signal G18405: std_logic; attribute dont_touch of G18405: signal is true;
	signal G18406: std_logic; attribute dont_touch of G18406: signal is true;
	signal G18407: std_logic; attribute dont_touch of G18407: signal is true;
	signal G18408: std_logic; attribute dont_touch of G18408: signal is true;
	signal G18409: std_logic; attribute dont_touch of G18409: signal is true;
	signal G18410: std_logic; attribute dont_touch of G18410: signal is true;
	signal G18411: std_logic; attribute dont_touch of G18411: signal is true;
	signal G18412: std_logic; attribute dont_touch of G18412: signal is true;
	signal G18413: std_logic; attribute dont_touch of G18413: signal is true;
	signal G18414: std_logic; attribute dont_touch of G18414: signal is true;
	signal G18415: std_logic; attribute dont_touch of G18415: signal is true;
	signal G18416: std_logic; attribute dont_touch of G18416: signal is true;
	signal G18417: std_logic; attribute dont_touch of G18417: signal is true;
	signal G18418: std_logic; attribute dont_touch of G18418: signal is true;
	signal G18419: std_logic; attribute dont_touch of G18419: signal is true;
	signal G18420: std_logic; attribute dont_touch of G18420: signal is true;
	signal G18421: std_logic; attribute dont_touch of G18421: signal is true;
	signal G18422: std_logic; attribute dont_touch of G18422: signal is true;
	signal G18423: std_logic; attribute dont_touch of G18423: signal is true;
	signal G18424: std_logic; attribute dont_touch of G18424: signal is true;
	signal G18425: std_logic; attribute dont_touch of G18425: signal is true;
	signal G18426: std_logic; attribute dont_touch of G18426: signal is true;
	signal G18427: std_logic; attribute dont_touch of G18427: signal is true;
	signal G18428: std_logic; attribute dont_touch of G18428: signal is true;
	signal G18429: std_logic; attribute dont_touch of G18429: signal is true;
	signal G18430: std_logic; attribute dont_touch of G18430: signal is true;
	signal G18431: std_logic; attribute dont_touch of G18431: signal is true;
	signal G18432: std_logic; attribute dont_touch of G18432: signal is true;
	signal G18433: std_logic; attribute dont_touch of G18433: signal is true;
	signal G18434: std_logic; attribute dont_touch of G18434: signal is true;
	signal G18435: std_logic; attribute dont_touch of G18435: signal is true;
	signal G18436: std_logic; attribute dont_touch of G18436: signal is true;
	signal G18437: std_logic; attribute dont_touch of G18437: signal is true;
	signal G18438: std_logic; attribute dont_touch of G18438: signal is true;
	signal G18439: std_logic; attribute dont_touch of G18439: signal is true;
	signal G18440: std_logic; attribute dont_touch of G18440: signal is true;
	signal G18441: std_logic; attribute dont_touch of G18441: signal is true;
	signal G18442: std_logic; attribute dont_touch of G18442: signal is true;
	signal G18443: std_logic; attribute dont_touch of G18443: signal is true;
	signal G18444: std_logic; attribute dont_touch of G18444: signal is true;
	signal G18445: std_logic; attribute dont_touch of G18445: signal is true;
	signal G18446: std_logic; attribute dont_touch of G18446: signal is true;
	signal G18447: std_logic; attribute dont_touch of G18447: signal is true;
	signal G18448: std_logic; attribute dont_touch of G18448: signal is true;
	signal G18449: std_logic; attribute dont_touch of G18449: signal is true;
	signal G18450: std_logic; attribute dont_touch of G18450: signal is true;
	signal G18451: std_logic; attribute dont_touch of G18451: signal is true;
	signal G18452: std_logic; attribute dont_touch of G18452: signal is true;
	signal G18453: std_logic; attribute dont_touch of G18453: signal is true;
	signal G18454: std_logic; attribute dont_touch of G18454: signal is true;
	signal G18455: std_logic; attribute dont_touch of G18455: signal is true;
	signal G18456: std_logic; attribute dont_touch of G18456: signal is true;
	signal G18457: std_logic; attribute dont_touch of G18457: signal is true;
	signal G18458: std_logic; attribute dont_touch of G18458: signal is true;
	signal G18459: std_logic; attribute dont_touch of G18459: signal is true;
	signal G18460: std_logic; attribute dont_touch of G18460: signal is true;
	signal G18461: std_logic; attribute dont_touch of G18461: signal is true;
	signal G18462: std_logic; attribute dont_touch of G18462: signal is true;
	signal G18463: std_logic; attribute dont_touch of G18463: signal is true;
	signal G18464: std_logic; attribute dont_touch of G18464: signal is true;
	signal G18465: std_logic; attribute dont_touch of G18465: signal is true;
	signal G18466: std_logic; attribute dont_touch of G18466: signal is true;
	signal G18467: std_logic; attribute dont_touch of G18467: signal is true;
	signal G18468: std_logic; attribute dont_touch of G18468: signal is true;
	signal G18469: std_logic; attribute dont_touch of G18469: signal is true;
	signal G18470: std_logic; attribute dont_touch of G18470: signal is true;
	signal G18471: std_logic; attribute dont_touch of G18471: signal is true;
	signal G18472: std_logic; attribute dont_touch of G18472: signal is true;
	signal G18473: std_logic; attribute dont_touch of G18473: signal is true;
	signal G18474: std_logic; attribute dont_touch of G18474: signal is true;
	signal G18475: std_logic; attribute dont_touch of G18475: signal is true;
	signal G18476: std_logic; attribute dont_touch of G18476: signal is true;
	signal G18477: std_logic; attribute dont_touch of G18477: signal is true;
	signal G18478: std_logic; attribute dont_touch of G18478: signal is true;
	signal G18479: std_logic; attribute dont_touch of G18479: signal is true;
	signal G18480: std_logic; attribute dont_touch of G18480: signal is true;
	signal G18481: std_logic; attribute dont_touch of G18481: signal is true;
	signal G18482: std_logic; attribute dont_touch of G18482: signal is true;
	signal G18483: std_logic; attribute dont_touch of G18483: signal is true;
	signal G18484: std_logic; attribute dont_touch of G18484: signal is true;
	signal G18485: std_logic; attribute dont_touch of G18485: signal is true;
	signal G18486: std_logic; attribute dont_touch of G18486: signal is true;
	signal G18487: std_logic; attribute dont_touch of G18487: signal is true;
	signal G18488: std_logic; attribute dont_touch of G18488: signal is true;
	signal G18489: std_logic; attribute dont_touch of G18489: signal is true;
	signal G18490: std_logic; attribute dont_touch of G18490: signal is true;
	signal G18491: std_logic; attribute dont_touch of G18491: signal is true;
	signal G18492: std_logic; attribute dont_touch of G18492: signal is true;
	signal G18493: std_logic; attribute dont_touch of G18493: signal is true;
	signal G18494: std_logic; attribute dont_touch of G18494: signal is true;
	signal G18495: std_logic; attribute dont_touch of G18495: signal is true;
	signal G18496: std_logic; attribute dont_touch of G18496: signal is true;
	signal G18497: std_logic; attribute dont_touch of G18497: signal is true;
	signal G18498: std_logic; attribute dont_touch of G18498: signal is true;
	signal G18499: std_logic; attribute dont_touch of G18499: signal is true;
	signal G18500: std_logic; attribute dont_touch of G18500: signal is true;
	signal G18501: std_logic; attribute dont_touch of G18501: signal is true;
	signal G18502: std_logic; attribute dont_touch of G18502: signal is true;
	signal G18503: std_logic; attribute dont_touch of G18503: signal is true;
	signal G18504: std_logic; attribute dont_touch of G18504: signal is true;
	signal G18505: std_logic; attribute dont_touch of G18505: signal is true;
	signal G18506: std_logic; attribute dont_touch of G18506: signal is true;
	signal G18507: std_logic; attribute dont_touch of G18507: signal is true;
	signal G18508: std_logic; attribute dont_touch of G18508: signal is true;
	signal G18509: std_logic; attribute dont_touch of G18509: signal is true;
	signal G18510: std_logic; attribute dont_touch of G18510: signal is true;
	signal G18511: std_logic; attribute dont_touch of G18511: signal is true;
	signal G18512: std_logic; attribute dont_touch of G18512: signal is true;
	signal G18513: std_logic; attribute dont_touch of G18513: signal is true;
	signal G18514: std_logic; attribute dont_touch of G18514: signal is true;
	signal G18515: std_logic; attribute dont_touch of G18515: signal is true;
	signal G18516: std_logic; attribute dont_touch of G18516: signal is true;
	signal G18517: std_logic; attribute dont_touch of G18517: signal is true;
	signal G18518: std_logic; attribute dont_touch of G18518: signal is true;
	signal G18519: std_logic; attribute dont_touch of G18519: signal is true;
	signal G18520: std_logic; attribute dont_touch of G18520: signal is true;
	signal G18521: std_logic; attribute dont_touch of G18521: signal is true;
	signal G18522: std_logic; attribute dont_touch of G18522: signal is true;
	signal G18523: std_logic; attribute dont_touch of G18523: signal is true;
	signal G18524: std_logic; attribute dont_touch of G18524: signal is true;
	signal G18525: std_logic; attribute dont_touch of G18525: signal is true;
	signal G18526: std_logic; attribute dont_touch of G18526: signal is true;
	signal G18527: std_logic; attribute dont_touch of G18527: signal is true;
	signal G18528: std_logic; attribute dont_touch of G18528: signal is true;
	signal G18529: std_logic; attribute dont_touch of G18529: signal is true;
	signal G18530: std_logic; attribute dont_touch of G18530: signal is true;
	signal G18531: std_logic; attribute dont_touch of G18531: signal is true;
	signal G18532: std_logic; attribute dont_touch of G18532: signal is true;
	signal G18533: std_logic; attribute dont_touch of G18533: signal is true;
	signal G18534: std_logic; attribute dont_touch of G18534: signal is true;
	signal G18535: std_logic; attribute dont_touch of G18535: signal is true;
	signal G18536: std_logic; attribute dont_touch of G18536: signal is true;
	signal G18537: std_logic; attribute dont_touch of G18537: signal is true;
	signal G18538: std_logic; attribute dont_touch of G18538: signal is true;
	signal G18539: std_logic; attribute dont_touch of G18539: signal is true;
	signal G18540: std_logic; attribute dont_touch of G18540: signal is true;
	signal G18541: std_logic; attribute dont_touch of G18541: signal is true;
	signal G18542: std_logic; attribute dont_touch of G18542: signal is true;
	signal G18543: std_logic; attribute dont_touch of G18543: signal is true;
	signal G18544: std_logic; attribute dont_touch of G18544: signal is true;
	signal G18545: std_logic; attribute dont_touch of G18545: signal is true;
	signal G18546: std_logic; attribute dont_touch of G18546: signal is true;
	signal G18547: std_logic; attribute dont_touch of G18547: signal is true;
	signal G18548: std_logic; attribute dont_touch of G18548: signal is true;
	signal G18549: std_logic; attribute dont_touch of G18549: signal is true;
	signal G18550: std_logic; attribute dont_touch of G18550: signal is true;
	signal G18551: std_logic; attribute dont_touch of G18551: signal is true;
	signal G18552: std_logic; attribute dont_touch of G18552: signal is true;
	signal G18553: std_logic; attribute dont_touch of G18553: signal is true;
	signal G18554: std_logic; attribute dont_touch of G18554: signal is true;
	signal G18555: std_logic; attribute dont_touch of G18555: signal is true;
	signal G18556: std_logic; attribute dont_touch of G18556: signal is true;
	signal G18557: std_logic; attribute dont_touch of G18557: signal is true;
	signal G18558: std_logic; attribute dont_touch of G18558: signal is true;
	signal G18559: std_logic; attribute dont_touch of G18559: signal is true;
	signal G18560: std_logic; attribute dont_touch of G18560: signal is true;
	signal G18561: std_logic; attribute dont_touch of G18561: signal is true;
	signal G18562: std_logic; attribute dont_touch of G18562: signal is true;
	signal G18563: std_logic; attribute dont_touch of G18563: signal is true;
	signal G18564: std_logic; attribute dont_touch of G18564: signal is true;
	signal G18565: std_logic; attribute dont_touch of G18565: signal is true;
	signal G18566: std_logic; attribute dont_touch of G18566: signal is true;
	signal G18567: std_logic; attribute dont_touch of G18567: signal is true;
	signal G18568: std_logic; attribute dont_touch of G18568: signal is true;
	signal G18569: std_logic; attribute dont_touch of G18569: signal is true;
	signal G18570: std_logic; attribute dont_touch of G18570: signal is true;
	signal G18571: std_logic; attribute dont_touch of G18571: signal is true;
	signal G18572: std_logic; attribute dont_touch of G18572: signal is true;
	signal G18573: std_logic; attribute dont_touch of G18573: signal is true;
	signal G18574: std_logic; attribute dont_touch of G18574: signal is true;
	signal G18575: std_logic; attribute dont_touch of G18575: signal is true;
	signal G18576: std_logic; attribute dont_touch of G18576: signal is true;
	signal G18577: std_logic; attribute dont_touch of G18577: signal is true;
	signal G18578: std_logic; attribute dont_touch of G18578: signal is true;
	signal G18579: std_logic; attribute dont_touch of G18579: signal is true;
	signal G18580: std_logic; attribute dont_touch of G18580: signal is true;
	signal G18581: std_logic; attribute dont_touch of G18581: signal is true;
	signal G18582: std_logic; attribute dont_touch of G18582: signal is true;
	signal G18583: std_logic; attribute dont_touch of G18583: signal is true;
	signal G18584: std_logic; attribute dont_touch of G18584: signal is true;
	signal G18585: std_logic; attribute dont_touch of G18585: signal is true;
	signal G18586: std_logic; attribute dont_touch of G18586: signal is true;
	signal G18587: std_logic; attribute dont_touch of G18587: signal is true;
	signal G18588: std_logic; attribute dont_touch of G18588: signal is true;
	signal G18589: std_logic; attribute dont_touch of G18589: signal is true;
	signal G18590: std_logic; attribute dont_touch of G18590: signal is true;
	signal G18591: std_logic; attribute dont_touch of G18591: signal is true;
	signal G18592: std_logic; attribute dont_touch of G18592: signal is true;
	signal G18593: std_logic; attribute dont_touch of G18593: signal is true;
	signal G18594: std_logic; attribute dont_touch of G18594: signal is true;
	signal G18595: std_logic; attribute dont_touch of G18595: signal is true;
	signal G18596: std_logic; attribute dont_touch of G18596: signal is true;
	signal G18597: std_logic; attribute dont_touch of G18597: signal is true;
	signal G18598: std_logic; attribute dont_touch of G18598: signal is true;
	signal G18599: std_logic; attribute dont_touch of G18599: signal is true;
	signal G18600: std_logic; attribute dont_touch of G18600: signal is true;
	signal G18601: std_logic; attribute dont_touch of G18601: signal is true;
	signal G18602: std_logic; attribute dont_touch of G18602: signal is true;
	signal G18603: std_logic; attribute dont_touch of G18603: signal is true;
	signal G18604: std_logic; attribute dont_touch of G18604: signal is true;
	signal G18605: std_logic; attribute dont_touch of G18605: signal is true;
	signal G18606: std_logic; attribute dont_touch of G18606: signal is true;
	signal G18607: std_logic; attribute dont_touch of G18607: signal is true;
	signal G18608: std_logic; attribute dont_touch of G18608: signal is true;
	signal G18609: std_logic; attribute dont_touch of G18609: signal is true;
	signal G18610: std_logic; attribute dont_touch of G18610: signal is true;
	signal G18611: std_logic; attribute dont_touch of G18611: signal is true;
	signal G18612: std_logic; attribute dont_touch of G18612: signal is true;
	signal G18613: std_logic; attribute dont_touch of G18613: signal is true;
	signal G18614: std_logic; attribute dont_touch of G18614: signal is true;
	signal G18615: std_logic; attribute dont_touch of G18615: signal is true;
	signal G18616: std_logic; attribute dont_touch of G18616: signal is true;
	signal G18617: std_logic; attribute dont_touch of G18617: signal is true;
	signal G18618: std_logic; attribute dont_touch of G18618: signal is true;
	signal G18619: std_logic; attribute dont_touch of G18619: signal is true;
	signal G18620: std_logic; attribute dont_touch of G18620: signal is true;
	signal G18621: std_logic; attribute dont_touch of G18621: signal is true;
	signal G18622: std_logic; attribute dont_touch of G18622: signal is true;
	signal G18623: std_logic; attribute dont_touch of G18623: signal is true;
	signal G18624: std_logic; attribute dont_touch of G18624: signal is true;
	signal G18625: std_logic; attribute dont_touch of G18625: signal is true;
	signal G18626: std_logic; attribute dont_touch of G18626: signal is true;
	signal G18627: std_logic; attribute dont_touch of G18627: signal is true;
	signal G18628: std_logic; attribute dont_touch of G18628: signal is true;
	signal G18629: std_logic; attribute dont_touch of G18629: signal is true;
	signal G18630: std_logic; attribute dont_touch of G18630: signal is true;
	signal G18631: std_logic; attribute dont_touch of G18631: signal is true;
	signal G18632: std_logic; attribute dont_touch of G18632: signal is true;
	signal G18633: std_logic; attribute dont_touch of G18633: signal is true;
	signal G18634: std_logic; attribute dont_touch of G18634: signal is true;
	signal G18635: std_logic; attribute dont_touch of G18635: signal is true;
	signal G18636: std_logic; attribute dont_touch of G18636: signal is true;
	signal G18637: std_logic; attribute dont_touch of G18637: signal is true;
	signal G18638: std_logic; attribute dont_touch of G18638: signal is true;
	signal G18639: std_logic; attribute dont_touch of G18639: signal is true;
	signal G18640: std_logic; attribute dont_touch of G18640: signal is true;
	signal G18641: std_logic; attribute dont_touch of G18641: signal is true;
	signal G18642: std_logic; attribute dont_touch of G18642: signal is true;
	signal G18643: std_logic; attribute dont_touch of G18643: signal is true;
	signal G18644: std_logic; attribute dont_touch of G18644: signal is true;
	signal G18645: std_logic; attribute dont_touch of G18645: signal is true;
	signal G18646: std_logic; attribute dont_touch of G18646: signal is true;
	signal G18647: std_logic; attribute dont_touch of G18647: signal is true;
	signal G18648: std_logic; attribute dont_touch of G18648: signal is true;
	signal G18649: std_logic; attribute dont_touch of G18649: signal is true;
	signal G18650: std_logic; attribute dont_touch of G18650: signal is true;
	signal G18651: std_logic; attribute dont_touch of G18651: signal is true;
	signal G18652: std_logic; attribute dont_touch of G18652: signal is true;
	signal G18653: std_logic; attribute dont_touch of G18653: signal is true;
	signal G18654: std_logic; attribute dont_touch of G18654: signal is true;
	signal G18655: std_logic; attribute dont_touch of G18655: signal is true;
	signal G18656: std_logic; attribute dont_touch of G18656: signal is true;
	signal G18657: std_logic; attribute dont_touch of G18657: signal is true;
	signal G18658: std_logic; attribute dont_touch of G18658: signal is true;
	signal G18659: std_logic; attribute dont_touch of G18659: signal is true;
	signal G18660: std_logic; attribute dont_touch of G18660: signal is true;
	signal G18661: std_logic; attribute dont_touch of G18661: signal is true;
	signal G18662: std_logic; attribute dont_touch of G18662: signal is true;
	signal G18663: std_logic; attribute dont_touch of G18663: signal is true;
	signal G18664: std_logic; attribute dont_touch of G18664: signal is true;
	signal G18665: std_logic; attribute dont_touch of G18665: signal is true;
	signal G18666: std_logic; attribute dont_touch of G18666: signal is true;
	signal G18667: std_logic; attribute dont_touch of G18667: signal is true;
	signal G18668: std_logic; attribute dont_touch of G18668: signal is true;
	signal G18669: std_logic; attribute dont_touch of G18669: signal is true;
	signal G18670: std_logic; attribute dont_touch of G18670: signal is true;
	signal G18671: std_logic; attribute dont_touch of G18671: signal is true;
	signal G18672: std_logic; attribute dont_touch of G18672: signal is true;
	signal G18673: std_logic; attribute dont_touch of G18673: signal is true;
	signal G18674: std_logic; attribute dont_touch of G18674: signal is true;
	signal G18675: std_logic; attribute dont_touch of G18675: signal is true;
	signal G18676: std_logic; attribute dont_touch of G18676: signal is true;
	signal G18677: std_logic; attribute dont_touch of G18677: signal is true;
	signal G18678: std_logic; attribute dont_touch of G18678: signal is true;
	signal G18679: std_logic; attribute dont_touch of G18679: signal is true;
	signal G18680: std_logic; attribute dont_touch of G18680: signal is true;
	signal G18681: std_logic; attribute dont_touch of G18681: signal is true;
	signal G18682: std_logic; attribute dont_touch of G18682: signal is true;
	signal G18683: std_logic; attribute dont_touch of G18683: signal is true;
	signal G18684: std_logic; attribute dont_touch of G18684: signal is true;
	signal G18685: std_logic; attribute dont_touch of G18685: signal is true;
	signal G18686: std_logic; attribute dont_touch of G18686: signal is true;
	signal G18687: std_logic; attribute dont_touch of G18687: signal is true;
	signal G18688: std_logic; attribute dont_touch of G18688: signal is true;
	signal G18689: std_logic; attribute dont_touch of G18689: signal is true;
	signal G18690: std_logic; attribute dont_touch of G18690: signal is true;
	signal G18691: std_logic; attribute dont_touch of G18691: signal is true;
	signal G18692: std_logic; attribute dont_touch of G18692: signal is true;
	signal G18693: std_logic; attribute dont_touch of G18693: signal is true;
	signal G18694: std_logic; attribute dont_touch of G18694: signal is true;
	signal G18695: std_logic; attribute dont_touch of G18695: signal is true;
	signal G18696: std_logic; attribute dont_touch of G18696: signal is true;
	signal G18697: std_logic; attribute dont_touch of G18697: signal is true;
	signal G18698: std_logic; attribute dont_touch of G18698: signal is true;
	signal G18699: std_logic; attribute dont_touch of G18699: signal is true;
	signal G18700: std_logic; attribute dont_touch of G18700: signal is true;
	signal G18701: std_logic; attribute dont_touch of G18701: signal is true;
	signal G18702: std_logic; attribute dont_touch of G18702: signal is true;
	signal G18703: std_logic; attribute dont_touch of G18703: signal is true;
	signal G18704: std_logic; attribute dont_touch of G18704: signal is true;
	signal G18705: std_logic; attribute dont_touch of G18705: signal is true;
	signal G18706: std_logic; attribute dont_touch of G18706: signal is true;
	signal G18707: std_logic; attribute dont_touch of G18707: signal is true;
	signal G18708: std_logic; attribute dont_touch of G18708: signal is true;
	signal G18709: std_logic; attribute dont_touch of G18709: signal is true;
	signal G18710: std_logic; attribute dont_touch of G18710: signal is true;
	signal G18711: std_logic; attribute dont_touch of G18711: signal is true;
	signal G18712: std_logic; attribute dont_touch of G18712: signal is true;
	signal G18713: std_logic; attribute dont_touch of G18713: signal is true;
	signal G18714: std_logic; attribute dont_touch of G18714: signal is true;
	signal G18715: std_logic; attribute dont_touch of G18715: signal is true;
	signal G18716: std_logic; attribute dont_touch of G18716: signal is true;
	signal G18717: std_logic; attribute dont_touch of G18717: signal is true;
	signal G18718: std_logic; attribute dont_touch of G18718: signal is true;
	signal G18719: std_logic; attribute dont_touch of G18719: signal is true;
	signal G18720: std_logic; attribute dont_touch of G18720: signal is true;
	signal G18721: std_logic; attribute dont_touch of G18721: signal is true;
	signal G18722: std_logic; attribute dont_touch of G18722: signal is true;
	signal G18723: std_logic; attribute dont_touch of G18723: signal is true;
	signal G18724: std_logic; attribute dont_touch of G18724: signal is true;
	signal G18725: std_logic; attribute dont_touch of G18725: signal is true;
	signal G18726: std_logic; attribute dont_touch of G18726: signal is true;
	signal G18727: std_logic; attribute dont_touch of G18727: signal is true;
	signal G18728: std_logic; attribute dont_touch of G18728: signal is true;
	signal G18729: std_logic; attribute dont_touch of G18729: signal is true;
	signal G18730: std_logic; attribute dont_touch of G18730: signal is true;
	signal G18731: std_logic; attribute dont_touch of G18731: signal is true;
	signal G18732: std_logic; attribute dont_touch of G18732: signal is true;
	signal G18733: std_logic; attribute dont_touch of G18733: signal is true;
	signal G18734: std_logic; attribute dont_touch of G18734: signal is true;
	signal G18735: std_logic; attribute dont_touch of G18735: signal is true;
	signal G18736: std_logic; attribute dont_touch of G18736: signal is true;
	signal G18737: std_logic; attribute dont_touch of G18737: signal is true;
	signal G18738: std_logic; attribute dont_touch of G18738: signal is true;
	signal G18739: std_logic; attribute dont_touch of G18739: signal is true;
	signal G18740: std_logic; attribute dont_touch of G18740: signal is true;
	signal G18741: std_logic; attribute dont_touch of G18741: signal is true;
	signal G18742: std_logic; attribute dont_touch of G18742: signal is true;
	signal G18743: std_logic; attribute dont_touch of G18743: signal is true;
	signal G18744: std_logic; attribute dont_touch of G18744: signal is true;
	signal G18745: std_logic; attribute dont_touch of G18745: signal is true;
	signal G18746: std_logic; attribute dont_touch of G18746: signal is true;
	signal G18747: std_logic; attribute dont_touch of G18747: signal is true;
	signal G18748: std_logic; attribute dont_touch of G18748: signal is true;
	signal G18749: std_logic; attribute dont_touch of G18749: signal is true;
	signal G18750: std_logic; attribute dont_touch of G18750: signal is true;
	signal G18751: std_logic; attribute dont_touch of G18751: signal is true;
	signal G18752: std_logic; attribute dont_touch of G18752: signal is true;
	signal G18753: std_logic; attribute dont_touch of G18753: signal is true;
	signal G18754: std_logic; attribute dont_touch of G18754: signal is true;
	signal G18755: std_logic; attribute dont_touch of G18755: signal is true;
	signal G18756: std_logic; attribute dont_touch of G18756: signal is true;
	signal G18757: std_logic; attribute dont_touch of G18757: signal is true;
	signal G18758: std_logic; attribute dont_touch of G18758: signal is true;
	signal G18759: std_logic; attribute dont_touch of G18759: signal is true;
	signal G18760: std_logic; attribute dont_touch of G18760: signal is true;
	signal G18761: std_logic; attribute dont_touch of G18761: signal is true;
	signal G18762: std_logic; attribute dont_touch of G18762: signal is true;
	signal G18763: std_logic; attribute dont_touch of G18763: signal is true;
	signal G18764: std_logic; attribute dont_touch of G18764: signal is true;
	signal G18765: std_logic; attribute dont_touch of G18765: signal is true;
	signal G18766: std_logic; attribute dont_touch of G18766: signal is true;
	signal G18767: std_logic; attribute dont_touch of G18767: signal is true;
	signal G18768: std_logic; attribute dont_touch of G18768: signal is true;
	signal G18769: std_logic; attribute dont_touch of G18769: signal is true;
	signal G18770: std_logic; attribute dont_touch of G18770: signal is true;
	signal G18771: std_logic; attribute dont_touch of G18771: signal is true;
	signal G18772: std_logic; attribute dont_touch of G18772: signal is true;
	signal G18773: std_logic; attribute dont_touch of G18773: signal is true;
	signal G18774: std_logic; attribute dont_touch of G18774: signal is true;
	signal G18775: std_logic; attribute dont_touch of G18775: signal is true;
	signal G18776: std_logic; attribute dont_touch of G18776: signal is true;
	signal G18777: std_logic; attribute dont_touch of G18777: signal is true;
	signal G18778: std_logic; attribute dont_touch of G18778: signal is true;
	signal G18779: std_logic; attribute dont_touch of G18779: signal is true;
	signal G18780: std_logic; attribute dont_touch of G18780: signal is true;
	signal G18781: std_logic; attribute dont_touch of G18781: signal is true;
	signal G18782: std_logic; attribute dont_touch of G18782: signal is true;
	signal G18783: std_logic; attribute dont_touch of G18783: signal is true;
	signal G18784: std_logic; attribute dont_touch of G18784: signal is true;
	signal G18785: std_logic; attribute dont_touch of G18785: signal is true;
	signal G18786: std_logic; attribute dont_touch of G18786: signal is true;
	signal G18787: std_logic; attribute dont_touch of G18787: signal is true;
	signal G18788: std_logic; attribute dont_touch of G18788: signal is true;
	signal G18789: std_logic; attribute dont_touch of G18789: signal is true;
	signal G18790: std_logic; attribute dont_touch of G18790: signal is true;
	signal G18791: std_logic; attribute dont_touch of G18791: signal is true;
	signal G18792: std_logic; attribute dont_touch of G18792: signal is true;
	signal G18793: std_logic; attribute dont_touch of G18793: signal is true;
	signal G18794: std_logic; attribute dont_touch of G18794: signal is true;
	signal G18795: std_logic; attribute dont_touch of G18795: signal is true;
	signal G18796: std_logic; attribute dont_touch of G18796: signal is true;
	signal G18797: std_logic; attribute dont_touch of G18797: signal is true;
	signal G18798: std_logic; attribute dont_touch of G18798: signal is true;
	signal G18799: std_logic; attribute dont_touch of G18799: signal is true;
	signal G18800: std_logic; attribute dont_touch of G18800: signal is true;
	signal G18801: std_logic; attribute dont_touch of G18801: signal is true;
	signal G18802: std_logic; attribute dont_touch of G18802: signal is true;
	signal G18803: std_logic; attribute dont_touch of G18803: signal is true;
	signal G18804: std_logic; attribute dont_touch of G18804: signal is true;
	signal G18805: std_logic; attribute dont_touch of G18805: signal is true;
	signal G18806: std_logic; attribute dont_touch of G18806: signal is true;
	signal G18807: std_logic; attribute dont_touch of G18807: signal is true;
	signal G18808: std_logic; attribute dont_touch of G18808: signal is true;
	signal G18809: std_logic; attribute dont_touch of G18809: signal is true;
	signal G18810: std_logic; attribute dont_touch of G18810: signal is true;
	signal G18811: std_logic; attribute dont_touch of G18811: signal is true;
	signal G18812: std_logic; attribute dont_touch of G18812: signal is true;
	signal G18813: std_logic; attribute dont_touch of G18813: signal is true;
	signal G18814: std_logic; attribute dont_touch of G18814: signal is true;
	signal G18815: std_logic; attribute dont_touch of G18815: signal is true;
	signal G18816: std_logic; attribute dont_touch of G18816: signal is true;
	signal G18817: std_logic; attribute dont_touch of G18817: signal is true;
	signal G18818: std_logic; attribute dont_touch of G18818: signal is true;
	signal G18819: std_logic; attribute dont_touch of G18819: signal is true;
	signal G18820: std_logic; attribute dont_touch of G18820: signal is true;
	signal G18821: std_logic; attribute dont_touch of G18821: signal is true;
	signal G18822: std_logic; attribute dont_touch of G18822: signal is true;
	signal G18823: std_logic; attribute dont_touch of G18823: signal is true;
	signal G18824: std_logic; attribute dont_touch of G18824: signal is true;
	signal G18825: std_logic; attribute dont_touch of G18825: signal is true;
	signal G18826: std_logic; attribute dont_touch of G18826: signal is true;
	signal G18827: std_logic; attribute dont_touch of G18827: signal is true;
	signal G18828: std_logic; attribute dont_touch of G18828: signal is true;
	signal G18829: std_logic; attribute dont_touch of G18829: signal is true;
	signal G18830: std_logic; attribute dont_touch of G18830: signal is true;
	signal G18831: std_logic; attribute dont_touch of G18831: signal is true;
	signal G18832: std_logic; attribute dont_touch of G18832: signal is true;
	signal G18833: std_logic; attribute dont_touch of G18833: signal is true;
	signal G18874: std_logic; attribute dont_touch of G18874: signal is true;
	signal G18875: std_logic; attribute dont_touch of G18875: signal is true;
	signal G18876: std_logic; attribute dont_touch of G18876: signal is true;
	signal G18877: std_logic; attribute dont_touch of G18877: signal is true;
	signal G18878: std_logic; attribute dont_touch of G18878: signal is true;
	signal G18879: std_logic; attribute dont_touch of G18879: signal is true;
	signal G18880: std_logic; attribute dont_touch of G18880: signal is true;
	signal G18882: std_logic; attribute dont_touch of G18882: signal is true;
	signal G18883: std_logic; attribute dont_touch of G18883: signal is true;
	signal G18884: std_logic; attribute dont_touch of G18884: signal is true;
	signal G18885: std_logic; attribute dont_touch of G18885: signal is true;
	signal G18886: std_logic; attribute dont_touch of G18886: signal is true;
	signal G18887: std_logic; attribute dont_touch of G18887: signal is true;
	signal G18888: std_logic; attribute dont_touch of G18888: signal is true;
	signal G18889: std_logic; attribute dont_touch of G18889: signal is true;
	signal G18890: std_logic; attribute dont_touch of G18890: signal is true;
	signal G18891: std_logic; attribute dont_touch of G18891: signal is true;
	signal G18892: std_logic; attribute dont_touch of G18892: signal is true;
	signal G18893: std_logic; attribute dont_touch of G18893: signal is true;
	signal G18894: std_logic; attribute dont_touch of G18894: signal is true;
	signal G18895: std_logic; attribute dont_touch of G18895: signal is true;
	signal G18896: std_logic; attribute dont_touch of G18896: signal is true;
	signal G18897: std_logic; attribute dont_touch of G18897: signal is true;
	signal G18898: std_logic; attribute dont_touch of G18898: signal is true;
	signal G18903: std_logic; attribute dont_touch of G18903: signal is true;
	signal G18904: std_logic; attribute dont_touch of G18904: signal is true;
	signal G18905: std_logic; attribute dont_touch of G18905: signal is true;
	signal G18906: std_logic; attribute dont_touch of G18906: signal is true;
	signal G18907: std_logic; attribute dont_touch of G18907: signal is true;
	signal G18908: std_logic; attribute dont_touch of G18908: signal is true;
	signal G18909: std_logic; attribute dont_touch of G18909: signal is true;
	signal G18910: std_logic; attribute dont_touch of G18910: signal is true;
	signal G18911: std_logic; attribute dont_touch of G18911: signal is true;
	signal G18916: std_logic; attribute dont_touch of G18916: signal is true;
	signal G18917: std_logic; attribute dont_touch of G18917: signal is true;
	signal G18918: std_logic; attribute dont_touch of G18918: signal is true;
	signal G18926: std_logic; attribute dont_touch of G18926: signal is true;
	signal G18929: std_logic; attribute dont_touch of G18929: signal is true;
	signal G18930: std_logic; attribute dont_touch of G18930: signal is true;
	signal G18931: std_logic; attribute dont_touch of G18931: signal is true;
	signal G18932: std_logic; attribute dont_touch of G18932: signal is true;
	signal G18933: std_logic; attribute dont_touch of G18933: signal is true;
	signal G18934: std_logic; attribute dont_touch of G18934: signal is true;
	signal G18935: std_logic; attribute dont_touch of G18935: signal is true;
	signal G18938: std_logic; attribute dont_touch of G18938: signal is true;
	signal G18939: std_logic; attribute dont_touch of G18939: signal is true;
	signal G18940: std_logic; attribute dont_touch of G18940: signal is true;
	signal G18943: std_logic; attribute dont_touch of G18943: signal is true;
	signal G18944: std_logic; attribute dont_touch of G18944: signal is true;
	signal G18945: std_logic; attribute dont_touch of G18945: signal is true;
	signal G18946: std_logic; attribute dont_touch of G18946: signal is true;
	signal G18947: std_logic; attribute dont_touch of G18947: signal is true;
	signal G18948: std_logic; attribute dont_touch of G18948: signal is true;
	signal G18949: std_logic; attribute dont_touch of G18949: signal is true;
	signal G18950: std_logic; attribute dont_touch of G18950: signal is true;
	signal G18951: std_logic; attribute dont_touch of G18951: signal is true;
	signal G18952: std_logic; attribute dont_touch of G18952: signal is true;
	signal G18953: std_logic; attribute dont_touch of G18953: signal is true;
	signal G18954: std_logic; attribute dont_touch of G18954: signal is true;
	signal G18957: std_logic; attribute dont_touch of G18957: signal is true;
	signal G18974: std_logic; attribute dont_touch of G18974: signal is true;
	signal G18975: std_logic; attribute dont_touch of G18975: signal is true;
	signal G18976: std_logic; attribute dont_touch of G18976: signal is true;
	signal G18977: std_logic; attribute dont_touch of G18977: signal is true;
	signal G18978: std_logic; attribute dont_touch of G18978: signal is true;
	signal G18979: std_logic; attribute dont_touch of G18979: signal is true;
	signal G18980: std_logic; attribute dont_touch of G18980: signal is true;
	signal G18981: std_logic; attribute dont_touch of G18981: signal is true;
	signal G18982: std_logic; attribute dont_touch of G18982: signal is true;
	signal G18983: std_logic; attribute dont_touch of G18983: signal is true;
	signal G18984: std_logic; attribute dont_touch of G18984: signal is true;
	signal G18987: std_logic; attribute dont_touch of G18987: signal is true;
	signal G18988: std_logic; attribute dont_touch of G18988: signal is true;
	signal G18989: std_logic; attribute dont_touch of G18989: signal is true;
	signal G18990: std_logic; attribute dont_touch of G18990: signal is true;
	signal G18991: std_logic; attribute dont_touch of G18991: signal is true;
	signal G18992: std_logic; attribute dont_touch of G18992: signal is true;
	signal G18993: std_logic; attribute dont_touch of G18993: signal is true;
	signal G18994: std_logic; attribute dont_touch of G18994: signal is true;
	signal G18997: std_logic; attribute dont_touch of G18997: signal is true;
	signal G19050: std_logic; attribute dont_touch of G19050: signal is true;
	signal G19061: std_logic; attribute dont_touch of G19061: signal is true;
	signal G19062: std_logic; attribute dont_touch of G19062: signal is true;
	signal G19063: std_logic; attribute dont_touch of G19063: signal is true;
	signal G19067: std_logic; attribute dont_touch of G19067: signal is true;
	signal G19068: std_logic; attribute dont_touch of G19068: signal is true;
	signal G19069: std_logic; attribute dont_touch of G19069: signal is true;
	signal G19070: std_logic; attribute dont_touch of G19070: signal is true;
	signal G19071: std_logic; attribute dont_touch of G19071: signal is true;
	signal G19074: std_logic; attribute dont_touch of G19074: signal is true;
	signal G19127: std_logic; attribute dont_touch of G19127: signal is true;
	signal G19128: std_logic; attribute dont_touch of G19128: signal is true;
	signal G19139: std_logic; attribute dont_touch of G19139: signal is true;
	signal G19140: std_logic; attribute dont_touch of G19140: signal is true;
	signal G19144: std_logic; attribute dont_touch of G19144: signal is true;
	signal G19145: std_logic; attribute dont_touch of G19145: signal is true;
	signal G19146: std_logic; attribute dont_touch of G19146: signal is true;
	signal G19147: std_logic; attribute dont_touch of G19147: signal is true;
	signal G19200: std_logic; attribute dont_touch of G19200: signal is true;
	signal G19206: std_logic; attribute dont_touch of G19206: signal is true;
	signal G19207: std_logic; attribute dont_touch of G19207: signal is true;
	signal G19208: std_logic; attribute dont_touch of G19208: signal is true;
	signal G19209: std_logic; attribute dont_touch of G19209: signal is true;
	signal G19210: std_logic; attribute dont_touch of G19210: signal is true;
	signal G19263: std_logic; attribute dont_touch of G19263: signal is true;
	signal G19264: std_logic; attribute dont_touch of G19264: signal is true;
	signal G19265: std_logic; attribute dont_touch of G19265: signal is true;
	signal G19266: std_logic; attribute dont_touch of G19266: signal is true;
	signal G19267: std_logic; attribute dont_touch of G19267: signal is true;
	signal G19268: std_logic; attribute dont_touch of G19268: signal is true;
	signal G19273: std_logic; attribute dont_touch of G19273: signal is true;
	signal G19274: std_logic; attribute dont_touch of G19274: signal is true;
	signal G19275: std_logic; attribute dont_touch of G19275: signal is true;
	signal G19276: std_logic; attribute dont_touch of G19276: signal is true;
	signal G19277: std_logic; attribute dont_touch of G19277: signal is true;
	signal G19330: std_logic; attribute dont_touch of G19330: signal is true;
	signal G19333: std_logic; attribute dont_touch of G19333: signal is true;
	signal G19335: std_logic; attribute dont_touch of G19335: signal is true;
	signal G19336: std_logic; attribute dont_touch of G19336: signal is true;
	signal G19337: std_logic; attribute dont_touch of G19337: signal is true;
	signal G19338: std_logic; attribute dont_touch of G19338: signal is true;
	signal G19343: std_logic; attribute dont_touch of G19343: signal is true;
	signal G19344: std_logic; attribute dont_touch of G19344: signal is true;
	signal G19345: std_logic; attribute dont_touch of G19345: signal is true;
	signal G19350: std_logic; attribute dont_touch of G19350: signal is true;
	signal G19351: std_logic; attribute dont_touch of G19351: signal is true;
	signal G19352: std_logic; attribute dont_touch of G19352: signal is true;
	signal G19353: std_logic; attribute dont_touch of G19353: signal is true;
	signal G19354: std_logic; attribute dont_touch of G19354: signal is true;
	signal G19355: std_logic; attribute dont_touch of G19355: signal is true;
	signal G19356: std_logic; attribute dont_touch of G19356: signal is true;
	signal G19358: std_logic; attribute dont_touch of G19358: signal is true;
	signal G19359: std_logic; attribute dont_touch of G19359: signal is true;
	signal G19360: std_logic; attribute dont_touch of G19360: signal is true;
	signal G19361: std_logic; attribute dont_touch of G19361: signal is true;
	signal G19362: std_logic; attribute dont_touch of G19362: signal is true;
	signal G19363: std_logic; attribute dont_touch of G19363: signal is true;
	signal G19364: std_logic; attribute dont_touch of G19364: signal is true;
	signal G19365: std_logic; attribute dont_touch of G19365: signal is true;
	signal G19366: std_logic; attribute dont_touch of G19366: signal is true;
	signal G19367: std_logic; attribute dont_touch of G19367: signal is true;
	signal G19368: std_logic; attribute dont_touch of G19368: signal is true;
	signal G19369: std_logic; attribute dont_touch of G19369: signal is true;
	signal G19370: std_logic; attribute dont_touch of G19370: signal is true;
	signal G19371: std_logic; attribute dont_touch of G19371: signal is true;
	signal G19372: std_logic; attribute dont_touch of G19372: signal is true;
	signal G19373: std_logic; attribute dont_touch of G19373: signal is true;
	signal G19374: std_logic; attribute dont_touch of G19374: signal is true;
	signal G19375: std_logic; attribute dont_touch of G19375: signal is true;
	signal G19376: std_logic; attribute dont_touch of G19376: signal is true;
	signal G19379: std_logic; attribute dont_touch of G19379: signal is true;
	signal G19383: std_logic; attribute dont_touch of G19383: signal is true;
	signal G19384: std_logic; attribute dont_touch of G19384: signal is true;
	signal G19385: std_logic; attribute dont_touch of G19385: signal is true;
	signal G19386: std_logic; attribute dont_touch of G19386: signal is true;
	signal G19387: std_logic; attribute dont_touch of G19387: signal is true;
	signal G19388: std_logic; attribute dont_touch of G19388: signal is true;
	signal G19389: std_logic; attribute dont_touch of G19389: signal is true;
	signal G19393: std_logic; attribute dont_touch of G19393: signal is true;
	signal G19394: std_logic; attribute dont_touch of G19394: signal is true;
	signal G19395: std_logic; attribute dont_touch of G19395: signal is true;
	signal G19396: std_logic; attribute dont_touch of G19396: signal is true;
	signal G19397: std_logic; attribute dont_touch of G19397: signal is true;
	signal G19398: std_logic; attribute dont_touch of G19398: signal is true;
	signal G19399: std_logic; attribute dont_touch of G19399: signal is true;
	signal G19400: std_logic; attribute dont_touch of G19400: signal is true;
	signal G19401: std_logic; attribute dont_touch of G19401: signal is true;
	signal G19402: std_logic; attribute dont_touch of G19402: signal is true;
	signal G19407: std_logic; attribute dont_touch of G19407: signal is true;
	signal G19408: std_logic; attribute dont_touch of G19408: signal is true;
	signal G19409: std_logic; attribute dont_touch of G19409: signal is true;
	signal G19410: std_logic; attribute dont_touch of G19410: signal is true;
	signal G19411: std_logic; attribute dont_touch of G19411: signal is true;
	signal G19412: std_logic; attribute dont_touch of G19412: signal is true;
	signal G19413: std_logic; attribute dont_touch of G19413: signal is true;
	signal G19414: std_logic; attribute dont_touch of G19414: signal is true;
	signal G19415: std_logic; attribute dont_touch of G19415: signal is true;
	signal G19416: std_logic; attribute dont_touch of G19416: signal is true;
	signal G19417: std_logic; attribute dont_touch of G19417: signal is true;
	signal G19421: std_logic; attribute dont_touch of G19421: signal is true;
	signal G19422: std_logic; attribute dont_touch of G19422: signal is true;
	signal G19427: std_logic; attribute dont_touch of G19427: signal is true;
	signal G19428: std_logic; attribute dont_touch of G19428: signal is true;
	signal G19429: std_logic; attribute dont_touch of G19429: signal is true;
	signal G19430: std_logic; attribute dont_touch of G19430: signal is true;
	signal G19431: std_logic; attribute dont_touch of G19431: signal is true;
	signal G19432: std_logic; attribute dont_touch of G19432: signal is true;
	signal G19433: std_logic; attribute dont_touch of G19433: signal is true;
	signal G19434: std_logic; attribute dont_touch of G19434: signal is true;
	signal G19435: std_logic; attribute dont_touch of G19435: signal is true;
	signal G19436: std_logic; attribute dont_touch of G19436: signal is true;
	signal G19437: std_logic; attribute dont_touch of G19437: signal is true;
	signal G19438: std_logic; attribute dont_touch of G19438: signal is true;
	signal G19439: std_logic; attribute dont_touch of G19439: signal is true;
	signal G19440: std_logic; attribute dont_touch of G19440: signal is true;
	signal G19441: std_logic; attribute dont_touch of G19441: signal is true;
	signal G19442: std_logic; attribute dont_touch of G19442: signal is true;
	signal G19443: std_logic; attribute dont_touch of G19443: signal is true;
	signal G19444: std_logic; attribute dont_touch of G19444: signal is true;
	signal G19445: std_logic; attribute dont_touch of G19445: signal is true;
	signal G19446: std_logic; attribute dont_touch of G19446: signal is true;
	signal G19449: std_logic; attribute dont_touch of G19449: signal is true;
	signal G19450: std_logic; attribute dont_touch of G19450: signal is true;
	signal G19451: std_logic; attribute dont_touch of G19451: signal is true;
	signal G19452: std_logic; attribute dont_touch of G19452: signal is true;
	signal G19453: std_logic; attribute dont_touch of G19453: signal is true;
	signal G19454: std_logic; attribute dont_touch of G19454: signal is true;
	signal G19455: std_logic; attribute dont_touch of G19455: signal is true;
	signal G19458: std_logic; attribute dont_touch of G19458: signal is true;
	signal G19461: std_logic; attribute dont_touch of G19461: signal is true;
	signal G19462: std_logic; attribute dont_touch of G19462: signal is true;
	signal G19466: std_logic; attribute dont_touch of G19466: signal is true;
	signal G19467: std_logic; attribute dont_touch of G19467: signal is true;
	signal G19468: std_logic; attribute dont_touch of G19468: signal is true;
	signal G19469: std_logic; attribute dont_touch of G19469: signal is true;
	signal G19470: std_logic; attribute dont_touch of G19470: signal is true;
	signal G19471: std_logic; attribute dont_touch of G19471: signal is true;
	signal G19472: std_logic; attribute dont_touch of G19472: signal is true;
	signal G19473: std_logic; attribute dont_touch of G19473: signal is true;
	signal G19474: std_logic; attribute dont_touch of G19474: signal is true;
	signal G19475: std_logic; attribute dont_touch of G19475: signal is true;
	signal G19476: std_logic; attribute dont_touch of G19476: signal is true;
	signal G19477: std_logic; attribute dont_touch of G19477: signal is true;
	signal G19478: std_logic; attribute dont_touch of G19478: signal is true;
	signal G19479: std_logic; attribute dont_touch of G19479: signal is true;
	signal G19480: std_logic; attribute dont_touch of G19480: signal is true;
	signal G19481: std_logic; attribute dont_touch of G19481: signal is true;
	signal G19482: std_logic; attribute dont_touch of G19482: signal is true;
	signal G19483: std_logic; attribute dont_touch of G19483: signal is true;
	signal G19486: std_logic; attribute dont_touch of G19486: signal is true;
	signal G19487: std_logic; attribute dont_touch of G19487: signal is true;
	signal G19488: std_logic; attribute dont_touch of G19488: signal is true;
	signal G19489: std_logic; attribute dont_touch of G19489: signal is true;
	signal G19490: std_logic; attribute dont_touch of G19490: signal is true;
	signal G19491: std_logic; attribute dont_touch of G19491: signal is true;
	signal G19492: std_logic; attribute dont_touch of G19492: signal is true;
	signal G19493: std_logic; attribute dont_touch of G19493: signal is true;
	signal G19494: std_logic; attribute dont_touch of G19494: signal is true;
	signal G19495: std_logic; attribute dont_touch of G19495: signal is true;
	signal G19498: std_logic; attribute dont_touch of G19498: signal is true;
	signal G19499: std_logic; attribute dont_touch of G19499: signal is true;
	signal G19500: std_logic; attribute dont_touch of G19500: signal is true;
	signal G19501: std_logic; attribute dont_touch of G19501: signal is true;
	signal G19502: std_logic; attribute dont_touch of G19502: signal is true;
	signal G19503: std_logic; attribute dont_touch of G19503: signal is true;
	signal G19504: std_logic; attribute dont_touch of G19504: signal is true;
	signal G19505: std_logic; attribute dont_touch of G19505: signal is true;
	signal G19506: std_logic; attribute dont_touch of G19506: signal is true;
	signal G19510: std_logic; attribute dont_touch of G19510: signal is true;
	signal G19513: std_logic; attribute dont_touch of G19513: signal is true;
	signal G19516: std_logic; attribute dont_touch of G19516: signal is true;
	signal G19517: std_logic; attribute dont_touch of G19517: signal is true;
	signal G19518: std_logic; attribute dont_touch of G19518: signal is true;
	signal G19519: std_logic; attribute dont_touch of G19519: signal is true;
	signal G19520: std_logic; attribute dont_touch of G19520: signal is true;
	signal G19521: std_logic; attribute dont_touch of G19521: signal is true;
	signal G19522: std_logic; attribute dont_touch of G19522: signal is true;
	signal G19523: std_logic; attribute dont_touch of G19523: signal is true;
	signal G19524: std_logic; attribute dont_touch of G19524: signal is true;
	signal G19525: std_logic; attribute dont_touch of G19525: signal is true;
	signal G19526: std_logic; attribute dont_touch of G19526: signal is true;
	signal G19527: std_logic; attribute dont_touch of G19527: signal is true;
	signal G19528: std_logic; attribute dont_touch of G19528: signal is true;
	signal G19529: std_logic; attribute dont_touch of G19529: signal is true;
	signal G19530: std_logic; attribute dont_touch of G19530: signal is true;
	signal G19531: std_logic; attribute dont_touch of G19531: signal is true;
	signal G19532: std_logic; attribute dont_touch of G19532: signal is true;
	signal G19533: std_logic; attribute dont_touch of G19533: signal is true;
	signal G19534: std_logic; attribute dont_touch of G19534: signal is true;
	signal G19535: std_logic; attribute dont_touch of G19535: signal is true;
	signal G19536: std_logic; attribute dont_touch of G19536: signal is true;
	signal G19537: std_logic; attribute dont_touch of G19537: signal is true;
	signal G19538: std_logic; attribute dont_touch of G19538: signal is true;
	signal G19539: std_logic; attribute dont_touch of G19539: signal is true;
	signal G19540: std_logic; attribute dont_touch of G19540: signal is true;
	signal G19541: std_logic; attribute dont_touch of G19541: signal is true;
	signal G19542: std_logic; attribute dont_touch of G19542: signal is true;
	signal G19543: std_logic; attribute dont_touch of G19543: signal is true;
	signal G19544: std_logic; attribute dont_touch of G19544: signal is true;
	signal G19545: std_logic; attribute dont_touch of G19545: signal is true;
	signal G19546: std_logic; attribute dont_touch of G19546: signal is true;
	signal G19549: std_logic; attribute dont_touch of G19549: signal is true;
	signal G19552: std_logic; attribute dont_touch of G19552: signal is true;
	signal G19553: std_logic; attribute dont_touch of G19553: signal is true;
	signal G19554: std_logic; attribute dont_touch of G19554: signal is true;
	signal G19555: std_logic; attribute dont_touch of G19555: signal is true;
	signal G19556: std_logic; attribute dont_touch of G19556: signal is true;
	signal G19557: std_logic; attribute dont_touch of G19557: signal is true;
	signal G19558: std_logic; attribute dont_touch of G19558: signal is true;
	signal G19559: std_logic; attribute dont_touch of G19559: signal is true;
	signal G19560: std_logic; attribute dont_touch of G19560: signal is true;
	signal G19564: std_logic; attribute dont_touch of G19564: signal is true;
	signal G19565: std_logic; attribute dont_touch of G19565: signal is true;
	signal G19566: std_logic; attribute dont_touch of G19566: signal is true;
	signal G19567: std_logic; attribute dont_touch of G19567: signal is true;
	signal G19568: std_logic; attribute dont_touch of G19568: signal is true;
	signal G19569: std_logic; attribute dont_touch of G19569: signal is true;
	signal G19570: std_logic; attribute dont_touch of G19570: signal is true;
	signal G19571: std_logic; attribute dont_touch of G19571: signal is true;
	signal G19572: std_logic; attribute dont_touch of G19572: signal is true;
	signal G19573: std_logic; attribute dont_touch of G19573: signal is true;
	signal G19574: std_logic; attribute dont_touch of G19574: signal is true;
	signal G19575: std_logic; attribute dont_touch of G19575: signal is true;
	signal G19576: std_logic; attribute dont_touch of G19576: signal is true;
	signal G19577: std_logic; attribute dont_touch of G19577: signal is true;
	signal G19578: std_logic; attribute dont_touch of G19578: signal is true;
	signal G19579: std_logic; attribute dont_touch of G19579: signal is true;
	signal G19580: std_logic; attribute dont_touch of G19580: signal is true;
	signal G19581: std_logic; attribute dont_touch of G19581: signal is true;
	signal G19585: std_logic; attribute dont_touch of G19585: signal is true;
	signal G19586: std_logic; attribute dont_touch of G19586: signal is true;
	signal G19587: std_logic; attribute dont_touch of G19587: signal is true;
	signal G19588: std_logic; attribute dont_touch of G19588: signal is true;
	signal G19589: std_logic; attribute dont_touch of G19589: signal is true;
	signal G19592: std_logic; attribute dont_touch of G19592: signal is true;
	signal G19593: std_logic; attribute dont_touch of G19593: signal is true;
	signal G19594: std_logic; attribute dont_touch of G19594: signal is true;
	signal G19595: std_logic; attribute dont_touch of G19595: signal is true;
	signal G19596: std_logic; attribute dont_touch of G19596: signal is true;
	signal G19597: std_logic; attribute dont_touch of G19597: signal is true;
	signal G19600: std_logic; attribute dont_touch of G19600: signal is true;
	signal G19601: std_logic; attribute dont_touch of G19601: signal is true;
	signal G19602: std_logic; attribute dont_touch of G19602: signal is true;
	signal G19603: std_logic; attribute dont_touch of G19603: signal is true;
	signal G19604: std_logic; attribute dont_touch of G19604: signal is true;
	signal G19605: std_logic; attribute dont_touch of G19605: signal is true;
	signal G19606: std_logic; attribute dont_touch of G19606: signal is true;
	signal G19609: std_logic; attribute dont_touch of G19609: signal is true;
	signal G19610: std_logic; attribute dont_touch of G19610: signal is true;
	signal G19611: std_logic; attribute dont_touch of G19611: signal is true;
	signal G19612: std_logic; attribute dont_touch of G19612: signal is true;
	signal G19613: std_logic; attribute dont_touch of G19613: signal is true;
	signal G19614: std_logic; attribute dont_touch of G19614: signal is true;
	signal G19617: std_logic; attribute dont_touch of G19617: signal is true;
	signal G19618: std_logic; attribute dont_touch of G19618: signal is true;
	signal G19619: std_logic; attribute dont_touch of G19619: signal is true;
	signal G19620: std_logic; attribute dont_touch of G19620: signal is true;
	signal G19626: std_logic; attribute dont_touch of G19626: signal is true;
	signal G19629: std_logic; attribute dont_touch of G19629: signal is true;
	signal G19630: std_logic; attribute dont_touch of G19630: signal is true;
	signal G19631: std_logic; attribute dont_touch of G19631: signal is true;
	signal G19632: std_logic; attribute dont_touch of G19632: signal is true;
	signal G19633: std_logic; attribute dont_touch of G19633: signal is true;
	signal G19634: std_logic; attribute dont_touch of G19634: signal is true;
	signal G19635: std_logic; attribute dont_touch of G19635: signal is true;
	signal G19636: std_logic; attribute dont_touch of G19636: signal is true;
	signal G19637: std_logic; attribute dont_touch of G19637: signal is true;
	signal G19638: std_logic; attribute dont_touch of G19638: signal is true;
	signal G19644: std_logic; attribute dont_touch of G19644: signal is true;
	signal G19649: std_logic; attribute dont_touch of G19649: signal is true;
	signal G19650: std_logic; attribute dont_touch of G19650: signal is true;
	signal G19651: std_logic; attribute dont_touch of G19651: signal is true;
	signal G19652: std_logic; attribute dont_touch of G19652: signal is true;
	signal G19653: std_logic; attribute dont_touch of G19653: signal is true;
	signal G19654: std_logic; attribute dont_touch of G19654: signal is true;
	signal G19655: std_logic; attribute dont_touch of G19655: signal is true;
	signal G19656: std_logic; attribute dont_touch of G19656: signal is true;
	signal G19657: std_logic; attribute dont_touch of G19657: signal is true;
	signal G19658: std_logic; attribute dont_touch of G19658: signal is true;
	signal G19659: std_logic; attribute dont_touch of G19659: signal is true;
	signal G19660: std_logic; attribute dont_touch of G19660: signal is true;
	signal G19661: std_logic; attribute dont_touch of G19661: signal is true;
	signal G19662: std_logic; attribute dont_touch of G19662: signal is true;
	signal G19666: std_logic; attribute dont_touch of G19666: signal is true;
	signal G19670: std_logic; attribute dont_touch of G19670: signal is true;
	signal G19671: std_logic; attribute dont_touch of G19671: signal is true;
	signal G19672: std_logic; attribute dont_touch of G19672: signal is true;
	signal G19673: std_logic; attribute dont_touch of G19673: signal is true;
	signal G19674: std_logic; attribute dont_touch of G19674: signal is true;
	signal G19675: std_logic; attribute dont_touch of G19675: signal is true;
	signal G19676: std_logic; attribute dont_touch of G19676: signal is true;
	signal G19677: std_logic; attribute dont_touch of G19677: signal is true;
	signal G19678: std_logic; attribute dont_touch of G19678: signal is true;
	signal G19679: std_logic; attribute dont_touch of G19679: signal is true;
	signal G19680: std_logic; attribute dont_touch of G19680: signal is true;
	signal G19681: std_logic; attribute dont_touch of G19681: signal is true;
	signal G19682: std_logic; attribute dont_touch of G19682: signal is true;
	signal G19683: std_logic; attribute dont_touch of G19683: signal is true;
	signal G19684: std_logic; attribute dont_touch of G19684: signal is true;
	signal G19685: std_logic; attribute dont_touch of G19685: signal is true;
	signal G19686: std_logic; attribute dont_touch of G19686: signal is true;
	signal G19687: std_logic; attribute dont_touch of G19687: signal is true;
	signal G19688: std_logic; attribute dont_touch of G19688: signal is true;
	signal G19689: std_logic; attribute dont_touch of G19689: signal is true;
	signal G19690: std_logic; attribute dont_touch of G19690: signal is true;
	signal G19691: std_logic; attribute dont_touch of G19691: signal is true;
	signal G19692: std_logic; attribute dont_touch of G19692: signal is true;
	signal G19693: std_logic; attribute dont_touch of G19693: signal is true;
	signal G19694: std_logic; attribute dont_touch of G19694: signal is true;
	signal G19695: std_logic; attribute dont_touch of G19695: signal is true;
	signal G19696: std_logic; attribute dont_touch of G19696: signal is true;
	signal G19697: std_logic; attribute dont_touch of G19697: signal is true;
	signal G19698: std_logic; attribute dont_touch of G19698: signal is true;
	signal G19699: std_logic; attribute dont_touch of G19699: signal is true;
	signal G19709: std_logic; attribute dont_touch of G19709: signal is true;
	signal G19710: std_logic; attribute dont_touch of G19710: signal is true;
	signal G19711: std_logic; attribute dont_touch of G19711: signal is true;
	signal G19712: std_logic; attribute dont_touch of G19712: signal is true;
	signal G19713: std_logic; attribute dont_touch of G19713: signal is true;
	signal G19714: std_logic; attribute dont_touch of G19714: signal is true;
	signal G19715: std_logic; attribute dont_touch of G19715: signal is true;
	signal G19716: std_logic; attribute dont_touch of G19716: signal is true;
	signal G19717: std_logic; attribute dont_touch of G19717: signal is true;
	signal G19718: std_logic; attribute dont_touch of G19718: signal is true;
	signal G19719: std_logic; attribute dont_touch of G19719: signal is true;
	signal G19720: std_logic; attribute dont_touch of G19720: signal is true;
	signal G19730: std_logic; attribute dont_touch of G19730: signal is true;
	signal G19731: std_logic; attribute dont_touch of G19731: signal is true;
	signal G19732: std_logic; attribute dont_touch of G19732: signal is true;
	signal G19733: std_logic; attribute dont_touch of G19733: signal is true;
	signal G19734: std_logic; attribute dont_touch of G19734: signal is true;
	signal G19735: std_logic; attribute dont_touch of G19735: signal is true;
	signal G19736: std_logic; attribute dont_touch of G19736: signal is true;
	signal G19737: std_logic; attribute dont_touch of G19737: signal is true;
	signal G19738: std_logic; attribute dont_touch of G19738: signal is true;
	signal G19739: std_logic; attribute dont_touch of G19739: signal is true;
	signal G19740: std_logic; attribute dont_touch of G19740: signal is true;
	signal G19741: std_logic; attribute dont_touch of G19741: signal is true;
	signal G19742: std_logic; attribute dont_touch of G19742: signal is true;
	signal G19743: std_logic; attribute dont_touch of G19743: signal is true;
	signal G19744: std_logic; attribute dont_touch of G19744: signal is true;
	signal G19745: std_logic; attribute dont_touch of G19745: signal is true;
	signal G19746: std_logic; attribute dont_touch of G19746: signal is true;
	signal G19747: std_logic; attribute dont_touch of G19747: signal is true;
	signal G19748: std_logic; attribute dont_touch of G19748: signal is true;
	signal G19749: std_logic; attribute dont_touch of G19749: signal is true;
	signal G19750: std_logic; attribute dont_touch of G19750: signal is true;
	signal G19751: std_logic; attribute dont_touch of G19751: signal is true;
	signal G19752: std_logic; attribute dont_touch of G19752: signal is true;
	signal G19753: std_logic; attribute dont_touch of G19753: signal is true;
	signal G19754: std_logic; attribute dont_touch of G19754: signal is true;
	signal G19755: std_logic; attribute dont_touch of G19755: signal is true;
	signal G19756: std_logic; attribute dont_touch of G19756: signal is true;
	signal G19757: std_logic; attribute dont_touch of G19757: signal is true;
	signal G19760: std_logic; attribute dont_touch of G19760: signal is true;
	signal G19761: std_logic; attribute dont_touch of G19761: signal is true;
	signal G19762: std_logic; attribute dont_touch of G19762: signal is true;
	signal G19763: std_logic; attribute dont_touch of G19763: signal is true;
	signal G19764: std_logic; attribute dont_touch of G19764: signal is true;
	signal G19765: std_logic; attribute dont_touch of G19765: signal is true;
	signal G19766: std_logic; attribute dont_touch of G19766: signal is true;
	signal G19767: std_logic; attribute dont_touch of G19767: signal is true;
	signal G19768: std_logic; attribute dont_touch of G19768: signal is true;
	signal G19769: std_logic; attribute dont_touch of G19769: signal is true;
	signal G19770: std_logic; attribute dont_touch of G19770: signal is true;
	signal G19771: std_logic; attribute dont_touch of G19771: signal is true;
	signal G19772: std_logic; attribute dont_touch of G19772: signal is true;
	signal G19773: std_logic; attribute dont_touch of G19773: signal is true;
	signal G19776: std_logic; attribute dont_touch of G19776: signal is true;
	signal G19777: std_logic; attribute dont_touch of G19777: signal is true;
	signal G19778: std_logic; attribute dont_touch of G19778: signal is true;
	signal G19779: std_logic; attribute dont_touch of G19779: signal is true;
	signal G19780: std_logic; attribute dont_touch of G19780: signal is true;
	signal G19781: std_logic; attribute dont_touch of G19781: signal is true;
	signal G19782: std_logic; attribute dont_touch of G19782: signal is true;
	signal G19783: std_logic; attribute dont_touch of G19783: signal is true;
	signal G19784: std_logic; attribute dont_touch of G19784: signal is true;
	signal G19785: std_logic; attribute dont_touch of G19785: signal is true;
	signal G19786: std_logic; attribute dont_touch of G19786: signal is true;
	signal G19787: std_logic; attribute dont_touch of G19787: signal is true;
	signal G19788: std_logic; attribute dont_touch of G19788: signal is true;
	signal G19789: std_logic; attribute dont_touch of G19789: signal is true;
	signal G19790: std_logic; attribute dont_touch of G19790: signal is true;
	signal G19791: std_logic; attribute dont_touch of G19791: signal is true;
	signal G19792: std_logic; attribute dont_touch of G19792: signal is true;
	signal G19793: std_logic; attribute dont_touch of G19793: signal is true;
	signal G19794: std_logic; attribute dont_touch of G19794: signal is true;
	signal G19795: std_logic; attribute dont_touch of G19795: signal is true;
	signal G19798: std_logic; attribute dont_touch of G19798: signal is true;
	signal G19799: std_logic; attribute dont_touch of G19799: signal is true;
	signal G19800: std_logic; attribute dont_touch of G19800: signal is true;
	signal G19801: std_logic; attribute dont_touch of G19801: signal is true;
	signal G19852: std_logic; attribute dont_touch of G19852: signal is true;
	signal G19853: std_logic; attribute dont_touch of G19853: signal is true;
	signal G19854: std_logic; attribute dont_touch of G19854: signal is true;
	signal G19855: std_logic; attribute dont_touch of G19855: signal is true;
	signal G19856: std_logic; attribute dont_touch of G19856: signal is true;
	signal G19857: std_logic; attribute dont_touch of G19857: signal is true;
	signal G19860: std_logic; attribute dont_touch of G19860: signal is true;
	signal G19861: std_logic; attribute dont_touch of G19861: signal is true;
	signal G19862: std_logic; attribute dont_touch of G19862: signal is true;
	signal G19865: std_logic; attribute dont_touch of G19865: signal is true;
	signal G19866: std_logic; attribute dont_touch of G19866: signal is true;
	signal G19869: std_logic; attribute dont_touch of G19869: signal is true;
	signal G19872: std_logic; attribute dont_touch of G19872: signal is true;
	signal G19873: std_logic; attribute dont_touch of G19873: signal is true;
	signal G19874: std_logic; attribute dont_touch of G19874: signal is true;
	signal G19875: std_logic; attribute dont_touch of G19875: signal is true;
	signal G19878: std_logic; attribute dont_touch of G19878: signal is true;
	signal G19879: std_logic; attribute dont_touch of G19879: signal is true;
	signal G19880: std_logic; attribute dont_touch of G19880: signal is true;
	signal G19881: std_logic; attribute dont_touch of G19881: signal is true;
	signal G19882: std_logic; attribute dont_touch of G19882: signal is true;
	signal G19885: std_logic; attribute dont_touch of G19885: signal is true;
	signal G19886: std_logic; attribute dont_touch of G19886: signal is true;
	signal G19887: std_logic; attribute dont_touch of G19887: signal is true;
	signal G19890: std_logic; attribute dont_touch of G19890: signal is true;
	signal G19902: std_logic; attribute dont_touch of G19902: signal is true;
	signal G19903: std_logic; attribute dont_touch of G19903: signal is true;
	signal G19904: std_logic; attribute dont_touch of G19904: signal is true;
	signal G19905: std_logic; attribute dont_touch of G19905: signal is true;
	signal G19906: std_logic; attribute dont_touch of G19906: signal is true;
	signal G19907: std_logic; attribute dont_touch of G19907: signal is true;
	signal G19908: std_logic; attribute dont_touch of G19908: signal is true;
	signal G19911: std_logic; attribute dont_touch of G19911: signal is true;
	signal G19912: std_logic; attribute dont_touch of G19912: signal is true;
	signal G19913: std_logic; attribute dont_touch of G19913: signal is true;
	signal G19914: std_logic; attribute dont_touch of G19914: signal is true;
	signal G19915: std_logic; attribute dont_touch of G19915: signal is true;
	signal G19916: std_logic; attribute dont_touch of G19916: signal is true;
	signal G19919: std_logic; attribute dont_touch of G19919: signal is true;
	signal G19930: std_logic; attribute dont_touch of G19930: signal is true;
	signal G19931: std_logic; attribute dont_touch of G19931: signal is true;
	signal G19932: std_logic; attribute dont_touch of G19932: signal is true;
	signal G19935: std_logic; attribute dont_touch of G19935: signal is true;
	signal G19947: std_logic; attribute dont_touch of G19947: signal is true;
	signal G19948: std_logic; attribute dont_touch of G19948: signal is true;
	signal G19949: std_logic; attribute dont_touch of G19949: signal is true;
	signal G19950: std_logic; attribute dont_touch of G19950: signal is true;
	signal G19951: std_logic; attribute dont_touch of G19951: signal is true;
	signal G19952: std_logic; attribute dont_touch of G19952: signal is true;
	signal G19953: std_logic; attribute dont_touch of G19953: signal is true;
	signal G19954: std_logic; attribute dont_touch of G19954: signal is true;
	signal G19957: std_logic; attribute dont_touch of G19957: signal is true;
	signal G19960: std_logic; attribute dont_touch of G19960: signal is true;
	signal G19961: std_logic; attribute dont_touch of G19961: signal is true;
	signal G19962: std_logic; attribute dont_touch of G19962: signal is true;
	signal G19963: std_logic; attribute dont_touch of G19963: signal is true;
	signal G19964: std_logic; attribute dont_touch of G19964: signal is true;
	signal G19965: std_logic; attribute dont_touch of G19965: signal is true;
	signal G19968: std_logic; attribute dont_touch of G19968: signal is true;
	signal G19979: std_logic; attribute dont_touch of G19979: signal is true;
	signal G19980: std_logic; attribute dont_touch of G19980: signal is true;
	signal G19981: std_logic; attribute dont_touch of G19981: signal is true;
	signal G19984: std_logic; attribute dont_touch of G19984: signal is true;
	signal G19996: std_logic; attribute dont_touch of G19996: signal is true;
	signal G19997: std_logic; attribute dont_touch of G19997: signal is true;
	signal G19998: std_logic; attribute dont_touch of G19998: signal is true;
	signal G19999: std_logic; attribute dont_touch of G19999: signal is true;
	signal G20000: std_logic; attribute dont_touch of G20000: signal is true;
	signal G20004: std_logic; attribute dont_touch of G20004: signal is true;
	signal G20005: std_logic; attribute dont_touch of G20005: signal is true;
	signal G20006: std_logic; attribute dont_touch of G20006: signal is true;
	signal G20007: std_logic; attribute dont_touch of G20007: signal is true;
	signal G20008: std_logic; attribute dont_touch of G20008: signal is true;
	signal G20009: std_logic; attribute dont_touch of G20009: signal is true;
	signal G20010: std_logic; attribute dont_touch of G20010: signal is true;
	signal G20011: std_logic; attribute dont_touch of G20011: signal is true;
	signal G20014: std_logic; attribute dont_touch of G20014: signal is true;
	signal G20025: std_logic; attribute dont_touch of G20025: signal is true;
	signal G20026: std_logic; attribute dont_touch of G20026: signal is true;
	signal G20027: std_logic; attribute dont_touch of G20027: signal is true;
	signal G20028: std_logic; attribute dont_touch of G20028: signal is true;
	signal G20033: std_logic; attribute dont_touch of G20033: signal is true;
	signal G20034: std_logic; attribute dont_touch of G20034: signal is true;
	signal G20035: std_logic; attribute dont_touch of G20035: signal is true;
	signal G20036: std_logic; attribute dont_touch of G20036: signal is true;
	signal G20037: std_logic; attribute dont_touch of G20037: signal is true;
	signal G20038: std_logic; attribute dont_touch of G20038: signal is true;
	signal G20039: std_logic; attribute dont_touch of G20039: signal is true;
	signal G20040: std_logic; attribute dont_touch of G20040: signal is true;
	signal G20041: std_logic; attribute dont_touch of G20041: signal is true;
	signal G20046: std_logic; attribute dont_touch of G20046: signal is true;
	signal G20050: std_logic; attribute dont_touch of G20050: signal is true;
	signal G20051: std_logic; attribute dont_touch of G20051: signal is true;
	signal G20052: std_logic; attribute dont_touch of G20052: signal is true;
	signal G20053: std_logic; attribute dont_touch of G20053: signal is true;
	signal G20054: std_logic; attribute dont_touch of G20054: signal is true;
	signal G20055: std_logic; attribute dont_touch of G20055: signal is true;
	signal G20056: std_logic; attribute dont_touch of G20056: signal is true;
	signal G20057: std_logic; attribute dont_touch of G20057: signal is true;
	signal G20058: std_logic; attribute dont_touch of G20058: signal is true;
	signal G20059: std_logic; attribute dont_touch of G20059: signal is true;
	signal G20060: std_logic; attribute dont_touch of G20060: signal is true;
	signal G20063: std_logic; attribute dont_touch of G20063: signal is true;
	signal G20064: std_logic; attribute dont_touch of G20064: signal is true;
	signal G20065: std_logic; attribute dont_touch of G20065: signal is true;
	signal G20066: std_logic; attribute dont_touch of G20066: signal is true;
	signal G20067: std_logic; attribute dont_touch of G20067: signal is true;
	signal G20068: std_logic; attribute dont_touch of G20068: signal is true;
	signal G20069: std_logic; attribute dont_touch of G20069: signal is true;
	signal G20070: std_logic; attribute dont_touch of G20070: signal is true;
	signal G20071: std_logic; attribute dont_touch of G20071: signal is true;
	signal G20072: std_logic; attribute dont_touch of G20072: signal is true;
	signal G20073: std_logic; attribute dont_touch of G20073: signal is true;
	signal G20076: std_logic; attribute dont_touch of G20076: signal is true;
	signal G20077: std_logic; attribute dont_touch of G20077: signal is true;
	signal G20078: std_logic; attribute dont_touch of G20078: signal is true;
	signal G20079: std_logic; attribute dont_touch of G20079: signal is true;
	signal G20080: std_logic; attribute dont_touch of G20080: signal is true;
	signal G20081: std_logic; attribute dont_touch of G20081: signal is true;
	signal G20082: std_logic; attribute dont_touch of G20082: signal is true;
	signal G20083: std_logic; attribute dont_touch of G20083: signal is true;
	signal G20084: std_logic; attribute dont_touch of G20084: signal is true;
	signal G20085: std_logic; attribute dont_touch of G20085: signal is true;
	signal G20086: std_logic; attribute dont_touch of G20086: signal is true;
	signal G20087: std_logic; attribute dont_touch of G20087: signal is true;
	signal G20088: std_logic; attribute dont_touch of G20088: signal is true;
	signal G20089: std_logic; attribute dont_touch of G20089: signal is true;
	signal G20090: std_logic; attribute dont_touch of G20090: signal is true;
	signal G20091: std_logic; attribute dont_touch of G20091: signal is true;
	signal G20092: std_logic; attribute dont_touch of G20092: signal is true;
	signal G20093: std_logic; attribute dont_touch of G20093: signal is true;
	signal G20094: std_logic; attribute dont_touch of G20094: signal is true;
	signal G20095: std_logic; attribute dont_touch of G20095: signal is true;
	signal G20096: std_logic; attribute dont_touch of G20096: signal is true;
	signal G20097: std_logic; attribute dont_touch of G20097: signal is true;
	signal G20100: std_logic; attribute dont_touch of G20100: signal is true;
	signal G20101: std_logic; attribute dont_touch of G20101: signal is true;
	signal G20102: std_logic; attribute dont_touch of G20102: signal is true;
	signal G20103: std_logic; attribute dont_touch of G20103: signal is true;
	signal G20104: std_logic; attribute dont_touch of G20104: signal is true;
	signal G20105: std_logic; attribute dont_touch of G20105: signal is true;
	signal G20106: std_logic; attribute dont_touch of G20106: signal is true;
	signal G20107: std_logic; attribute dont_touch of G20107: signal is true;
	signal G20108: std_logic; attribute dont_touch of G20108: signal is true;
	signal G20109: std_logic; attribute dont_touch of G20109: signal is true;
	signal G20110: std_logic; attribute dont_touch of G20110: signal is true;
	signal G20111: std_logic; attribute dont_touch of G20111: signal is true;
	signal G20112: std_logic; attribute dont_touch of G20112: signal is true;
	signal G20113: std_logic; attribute dont_touch of G20113: signal is true;
	signal G20114: std_logic; attribute dont_touch of G20114: signal is true;
	signal G20127: std_logic; attribute dont_touch of G20127: signal is true;
	signal G20128: std_logic; attribute dont_touch of G20128: signal is true;
	signal G20129: std_logic; attribute dont_touch of G20129: signal is true;
	signal G20130: std_logic; attribute dont_touch of G20130: signal is true;
	signal G20131: std_logic; attribute dont_touch of G20131: signal is true;
	signal G20132: std_logic; attribute dont_touch of G20132: signal is true;
	signal G20133: std_logic; attribute dont_touch of G20133: signal is true;
	signal G20134: std_logic; attribute dont_touch of G20134: signal is true;
	signal G20135: std_logic; attribute dont_touch of G20135: signal is true;
	signal G20136: std_logic; attribute dont_touch of G20136: signal is true;
	signal G20144: std_logic; attribute dont_touch of G20144: signal is true;
	signal G20145: std_logic; attribute dont_touch of G20145: signal is true;
	signal G20146: std_logic; attribute dont_touch of G20146: signal is true;
	signal G20147: std_logic; attribute dont_touch of G20147: signal is true;
	signal G20148: std_logic; attribute dont_touch of G20148: signal is true;
	signal G20149: std_logic; attribute dont_touch of G20149: signal is true;
	signal G20150: std_logic; attribute dont_touch of G20150: signal is true;
	signal G20151: std_logic; attribute dont_touch of G20151: signal is true;
	signal G20152: std_logic; attribute dont_touch of G20152: signal is true;
	signal G20153: std_logic; attribute dont_touch of G20153: signal is true;
	signal G20154: std_logic; attribute dont_touch of G20154: signal is true;
	signal G20157: std_logic; attribute dont_touch of G20157: signal is true;
	signal G20158: std_logic; attribute dont_touch of G20158: signal is true;
	signal G20159: std_logic; attribute dont_touch of G20159: signal is true;
	signal G20160: std_logic; attribute dont_touch of G20160: signal is true;
	signal G20161: std_logic; attribute dont_touch of G20161: signal is true;
	signal G20162: std_logic; attribute dont_touch of G20162: signal is true;
	signal G20163: std_logic; attribute dont_touch of G20163: signal is true;
	signal G20164: std_logic; attribute dont_touch of G20164: signal is true;
	signal G20165: std_logic; attribute dont_touch of G20165: signal is true;
	signal G20166: std_logic; attribute dont_touch of G20166: signal is true;
	signal G20167: std_logic; attribute dont_touch of G20167: signal is true;
	signal G20168: std_logic; attribute dont_touch of G20168: signal is true;
	signal G20169: std_logic; attribute dont_touch of G20169: signal is true;
	signal G20170: std_logic; attribute dont_touch of G20170: signal is true;
	signal G20171: std_logic; attribute dont_touch of G20171: signal is true;
	signal G20172: std_logic; attribute dont_touch of G20172: signal is true;
	signal G20173: std_logic; attribute dont_touch of G20173: signal is true;
	signal G20174: std_logic; attribute dont_touch of G20174: signal is true;
	signal G20175: std_logic; attribute dont_touch of G20175: signal is true;
	signal G20178: std_logic; attribute dont_touch of G20178: signal is true;
	signal G20179: std_logic; attribute dont_touch of G20179: signal is true;
	signal G20180: std_logic; attribute dont_touch of G20180: signal is true;
	signal G20181: std_logic; attribute dont_touch of G20181: signal is true;
	signal G20182: std_logic; attribute dont_touch of G20182: signal is true;
	signal G20183: std_logic; attribute dont_touch of G20183: signal is true;
	signal G20184: std_logic; attribute dont_touch of G20184: signal is true;
	signal G20185: std_logic; attribute dont_touch of G20185: signal is true;
	signal G20186: std_logic; attribute dont_touch of G20186: signal is true;
	signal G20187: std_logic; attribute dont_touch of G20187: signal is true;
	signal G20188: std_logic; attribute dont_touch of G20188: signal is true;
	signal G20189: std_logic; attribute dont_touch of G20189: signal is true;
	signal G20190: std_logic; attribute dont_touch of G20190: signal is true;
	signal G20191: std_logic; attribute dont_touch of G20191: signal is true;
	signal G20192: std_logic; attribute dont_touch of G20192: signal is true;
	signal G20193: std_logic; attribute dont_touch of G20193: signal is true;
	signal G20194: std_logic; attribute dont_touch of G20194: signal is true;
	signal G20195: std_logic; attribute dont_touch of G20195: signal is true;
	signal G20196: std_logic; attribute dont_touch of G20196: signal is true;
	signal G20197: std_logic; attribute dont_touch of G20197: signal is true;
	signal G20198: std_logic; attribute dont_touch of G20198: signal is true;
	signal G20199: std_logic; attribute dont_touch of G20199: signal is true;
	signal G20200: std_logic; attribute dont_touch of G20200: signal is true;
	signal G20201: std_logic; attribute dont_touch of G20201: signal is true;
	signal G20202: std_logic; attribute dont_touch of G20202: signal is true;
	signal G20203: std_logic; attribute dont_touch of G20203: signal is true;
	signal G20204: std_logic; attribute dont_touch of G20204: signal is true;
	signal G20207: std_logic; attribute dont_touch of G20207: signal is true;
	signal G20208: std_logic; attribute dont_touch of G20208: signal is true;
	signal G20209: std_logic; attribute dont_touch of G20209: signal is true;
	signal G20210: std_logic; attribute dont_touch of G20210: signal is true;
	signal G20211: std_logic; attribute dont_touch of G20211: signal is true;
	signal G20212: std_logic; attribute dont_touch of G20212: signal is true;
	signal G20213: std_logic; attribute dont_touch of G20213: signal is true;
	signal G20214: std_logic; attribute dont_touch of G20214: signal is true;
	signal G20215: std_logic; attribute dont_touch of G20215: signal is true;
	signal G20216: std_logic; attribute dont_touch of G20216: signal is true;
	signal G20217: std_logic; attribute dont_touch of G20217: signal is true;
	signal G20218: std_logic; attribute dont_touch of G20218: signal is true;
	signal G20219: std_logic; attribute dont_touch of G20219: signal is true;
	signal G20229: std_logic; attribute dont_touch of G20229: signal is true;
	signal G20230: std_logic; attribute dont_touch of G20230: signal is true;
	signal G20231: std_logic; attribute dont_touch of G20231: signal is true;
	signal G20232: std_logic; attribute dont_touch of G20232: signal is true;
	signal G20233: std_logic; attribute dont_touch of G20233: signal is true;
	signal G20234: std_logic; attribute dont_touch of G20234: signal is true;
	signal G20235: std_logic; attribute dont_touch of G20235: signal is true;
	signal G20236: std_logic; attribute dont_touch of G20236: signal is true;
	signal G20237: std_logic; attribute dont_touch of G20237: signal is true;
	signal G20238: std_logic; attribute dont_touch of G20238: signal is true;
	signal G20239: std_logic; attribute dont_touch of G20239: signal is true;
	signal G20240: std_logic; attribute dont_touch of G20240: signal is true;
	signal G20241: std_logic; attribute dont_touch of G20241: signal is true;
	signal G20242: std_logic; attribute dont_touch of G20242: signal is true;
	signal G20247: std_logic; attribute dont_touch of G20247: signal is true;
	signal G20248: std_logic; attribute dont_touch of G20248: signal is true;
	signal G20265: std_logic; attribute dont_touch of G20265: signal is true;
	signal G20266: std_logic; attribute dont_touch of G20266: signal is true;
	signal G20267: std_logic; attribute dont_touch of G20267: signal is true;
	signal G20268: std_logic; attribute dont_touch of G20268: signal is true;
	signal G20269: std_logic; attribute dont_touch of G20269: signal is true;
	signal G20270: std_logic; attribute dont_touch of G20270: signal is true;
	signal G20271: std_logic; attribute dont_touch of G20271: signal is true;
	signal G20272: std_logic; attribute dont_touch of G20272: signal is true;
	signal G20273: std_logic; attribute dont_touch of G20273: signal is true;
	signal G20274: std_logic; attribute dont_touch of G20274: signal is true;
	signal G20275: std_logic; attribute dont_touch of G20275: signal is true;
	signal G20276: std_logic; attribute dont_touch of G20276: signal is true;
	signal G20277: std_logic; attribute dont_touch of G20277: signal is true;
	signal G20283: std_logic; attribute dont_touch of G20283: signal is true;
	signal G20320: std_logic; attribute dont_touch of G20320: signal is true;
	signal G20321: std_logic; attribute dont_touch of G20321: signal is true;
	signal G20322: std_logic; attribute dont_touch of G20322: signal is true;
	signal G20323: std_logic; attribute dont_touch of G20323: signal is true;
	signal G20324: std_logic; attribute dont_touch of G20324: signal is true;
	signal G20325: std_logic; attribute dont_touch of G20325: signal is true;
	signal G20326: std_logic; attribute dont_touch of G20326: signal is true;
	signal G20327: std_logic; attribute dont_touch of G20327: signal is true;
	signal G20328: std_logic; attribute dont_touch of G20328: signal is true;
	signal G20329: std_logic; attribute dont_touch of G20329: signal is true;
	signal G20330: std_logic; attribute dont_touch of G20330: signal is true;
	signal G20371: std_logic; attribute dont_touch of G20371: signal is true;
	signal G20372: std_logic; attribute dont_touch of G20372: signal is true;
	signal G20373: std_logic; attribute dont_touch of G20373: signal is true;
	signal G20374: std_logic; attribute dont_touch of G20374: signal is true;
	signal G20375: std_logic; attribute dont_touch of G20375: signal is true;
	signal G20379: std_logic; attribute dont_touch of G20379: signal is true;
	signal G20380: std_logic; attribute dont_touch of G20380: signal is true;
	signal G20381: std_logic; attribute dont_touch of G20381: signal is true;
	signal G20382: std_logic; attribute dont_touch of G20382: signal is true;
	signal G20383: std_logic; attribute dont_touch of G20383: signal is true;
	signal G20384: std_logic; attribute dont_touch of G20384: signal is true;
	signal G20385: std_logic; attribute dont_touch of G20385: signal is true;
	signal G20386: std_logic; attribute dont_touch of G20386: signal is true;
	signal G20387: std_logic; attribute dont_touch of G20387: signal is true;
	signal G20388: std_logic; attribute dont_touch of G20388: signal is true;
	signal G20389: std_logic; attribute dont_touch of G20389: signal is true;
	signal G20390: std_logic; attribute dont_touch of G20390: signal is true;
	signal G20391: std_logic; attribute dont_touch of G20391: signal is true;
	signal G20432: std_logic; attribute dont_touch of G20432: signal is true;
	signal G20433: std_logic; attribute dont_touch of G20433: signal is true;
	signal G20434: std_logic; attribute dont_touch of G20434: signal is true;
	signal G20435: std_logic; attribute dont_touch of G20435: signal is true;
	signal G20436: std_logic; attribute dont_touch of G20436: signal is true;
	signal G20441: std_logic; attribute dont_touch of G20441: signal is true;
	signal G20442: std_logic; attribute dont_touch of G20442: signal is true;
	signal G20443: std_logic; attribute dont_touch of G20443: signal is true;
	signal G20444: std_logic; attribute dont_touch of G20444: signal is true;
	signal G20445: std_logic; attribute dont_touch of G20445: signal is true;
	signal G20446: std_logic; attribute dont_touch of G20446: signal is true;
	signal G20447: std_logic; attribute dont_touch of G20447: signal is true;
	signal G20448: std_logic; attribute dont_touch of G20448: signal is true;
	signal G20449: std_logic; attribute dont_touch of G20449: signal is true;
	signal G20450: std_logic; attribute dont_touch of G20450: signal is true;
	signal G20451: std_logic; attribute dont_touch of G20451: signal is true;
	signal G20452: std_logic; attribute dont_touch of G20452: signal is true;
	signal G20453: std_logic; attribute dont_touch of G20453: signal is true;
	signal G20494: std_logic; attribute dont_touch of G20494: signal is true;
	signal G20495: std_logic; attribute dont_touch of G20495: signal is true;
	signal G20496: std_logic; attribute dont_touch of G20496: signal is true;
	signal G20497: std_logic; attribute dont_touch of G20497: signal is true;
	signal G20498: std_logic; attribute dont_touch of G20498: signal is true;
	signal G20499: std_logic; attribute dont_touch of G20499: signal is true;
	signal G20500: std_logic; attribute dont_touch of G20500: signal is true;
	signal G20501: std_logic; attribute dont_touch of G20501: signal is true;
	signal G20502: std_logic; attribute dont_touch of G20502: signal is true;
	signal G20503: std_logic; attribute dont_touch of G20503: signal is true;
	signal G20504: std_logic; attribute dont_touch of G20504: signal is true;
	signal G20505: std_logic; attribute dont_touch of G20505: signal is true;
	signal G20506: std_logic; attribute dont_touch of G20506: signal is true;
	signal G20507: std_logic; attribute dont_touch of G20507: signal is true;
	signal G20508: std_logic; attribute dont_touch of G20508: signal is true;
	signal G20509: std_logic; attribute dont_touch of G20509: signal is true;
	signal G20510: std_logic; attribute dont_touch of G20510: signal is true;
	signal G20511: std_logic; attribute dont_touch of G20511: signal is true;
	signal G20512: std_logic; attribute dont_touch of G20512: signal is true;
	signal G20513: std_logic; attribute dont_touch of G20513: signal is true;
	signal G20514: std_logic; attribute dont_touch of G20514: signal is true;
	signal G20515: std_logic; attribute dont_touch of G20515: signal is true;
	signal G20516: std_logic; attribute dont_touch of G20516: signal is true;
	signal G20522: std_logic; attribute dont_touch of G20522: signal is true;
	signal G20523: std_logic; attribute dont_touch of G20523: signal is true;
	signal G20524: std_logic; attribute dont_touch of G20524: signal is true;
	signal G20525: std_logic; attribute dont_touch of G20525: signal is true;
	signal G20526: std_logic; attribute dont_touch of G20526: signal is true;
	signal G20527: std_logic; attribute dont_touch of G20527: signal is true;
	signal G20528: std_logic; attribute dont_touch of G20528: signal is true;
	signal G20529: std_logic; attribute dont_touch of G20529: signal is true;
	signal G20530: std_logic; attribute dont_touch of G20530: signal is true;
	signal G20531: std_logic; attribute dont_touch of G20531: signal is true;
	signal G20532: std_logic; attribute dont_touch of G20532: signal is true;
	signal G20533: std_logic; attribute dont_touch of G20533: signal is true;
	signal G20534: std_logic; attribute dont_touch of G20534: signal is true;
	signal G20535: std_logic; attribute dont_touch of G20535: signal is true;
	signal G20536: std_logic; attribute dont_touch of G20536: signal is true;
	signal G20537: std_logic; attribute dont_touch of G20537: signal is true;
	signal G20538: std_logic; attribute dont_touch of G20538: signal is true;
	signal G20539: std_logic; attribute dont_touch of G20539: signal is true;
	signal G20540: std_logic; attribute dont_touch of G20540: signal is true;
	signal G20541: std_logic; attribute dont_touch of G20541: signal is true;
	signal G20542: std_logic; attribute dont_touch of G20542: signal is true;
	signal G20543: std_logic; attribute dont_touch of G20543: signal is true;
	signal G20544: std_logic; attribute dont_touch of G20544: signal is true;
	signal G20545: std_logic; attribute dont_touch of G20545: signal is true;
	signal G20546: std_logic; attribute dont_touch of G20546: signal is true;
	signal G20547: std_logic; attribute dont_touch of G20547: signal is true;
	signal G20548: std_logic; attribute dont_touch of G20548: signal is true;
	signal G20549: std_logic; attribute dont_touch of G20549: signal is true;
	signal G20550: std_logic; attribute dont_touch of G20550: signal is true;
	signal G20551: std_logic; attribute dont_touch of G20551: signal is true;
	signal G20552: std_logic; attribute dont_touch of G20552: signal is true;
	signal G20553: std_logic; attribute dont_touch of G20553: signal is true;
	signal G20554: std_logic; attribute dont_touch of G20554: signal is true;
	signal G20555: std_logic; attribute dont_touch of G20555: signal is true;
	signal G20556: std_logic; attribute dont_touch of G20556: signal is true;
	signal G20558: std_logic; attribute dont_touch of G20558: signal is true;
	signal G20559: std_logic; attribute dont_touch of G20559: signal is true;
	signal G20560: std_logic; attribute dont_touch of G20560: signal is true;
	signal G20561: std_logic; attribute dont_touch of G20561: signal is true;
	signal G20562: std_logic; attribute dont_touch of G20562: signal is true;
	signal G20563: std_logic; attribute dont_touch of G20563: signal is true;
	signal G20564: std_logic; attribute dont_touch of G20564: signal is true;
	signal G20565: std_logic; attribute dont_touch of G20565: signal is true;
	signal G20566: std_logic; attribute dont_touch of G20566: signal is true;
	signal G20567: std_logic; attribute dont_touch of G20567: signal is true;
	signal G20568: std_logic; attribute dont_touch of G20568: signal is true;
	signal G20569: std_logic; attribute dont_touch of G20569: signal is true;
	signal G20570: std_logic; attribute dont_touch of G20570: signal is true;
	signal G20571: std_logic; attribute dont_touch of G20571: signal is true;
	signal G20572: std_logic; attribute dont_touch of G20572: signal is true;
	signal G20573: std_logic; attribute dont_touch of G20573: signal is true;
	signal G20574: std_logic; attribute dont_touch of G20574: signal is true;
	signal G20575: std_logic; attribute dont_touch of G20575: signal is true;
	signal G20576: std_logic; attribute dont_touch of G20576: signal is true;
	signal G20577: std_logic; attribute dont_touch of G20577: signal is true;
	signal G20578: std_logic; attribute dont_touch of G20578: signal is true;
	signal G20579: std_logic; attribute dont_touch of G20579: signal is true;
	signal G20580: std_logic; attribute dont_touch of G20580: signal is true;
	signal G20581: std_logic; attribute dont_touch of G20581: signal is true;
	signal G20582: std_logic; attribute dont_touch of G20582: signal is true;
	signal G20583: std_logic; attribute dont_touch of G20583: signal is true;
	signal G20584: std_logic; attribute dont_touch of G20584: signal is true;
	signal G20585: std_logic; attribute dont_touch of G20585: signal is true;
	signal G20586: std_logic; attribute dont_touch of G20586: signal is true;
	signal G20587: std_logic; attribute dont_touch of G20587: signal is true;
	signal G20588: std_logic; attribute dont_touch of G20588: signal is true;
	signal G20589: std_logic; attribute dont_touch of G20589: signal is true;
	signal G20590: std_logic; attribute dont_touch of G20590: signal is true;
	signal G20591: std_logic; attribute dont_touch of G20591: signal is true;
	signal G20592: std_logic; attribute dont_touch of G20592: signal is true;
	signal G20593: std_logic; attribute dont_touch of G20593: signal is true;
	signal G20594: std_logic; attribute dont_touch of G20594: signal is true;
	signal G20595: std_logic; attribute dont_touch of G20595: signal is true;
	signal G20596: std_logic; attribute dont_touch of G20596: signal is true;
	signal G20597: std_logic; attribute dont_touch of G20597: signal is true;
	signal G20598: std_logic; attribute dont_touch of G20598: signal is true;
	signal G20599: std_logic; attribute dont_touch of G20599: signal is true;
	signal G20600: std_logic; attribute dont_touch of G20600: signal is true;
	signal G20601: std_logic; attribute dont_touch of G20601: signal is true;
	signal G20602: std_logic; attribute dont_touch of G20602: signal is true;
	signal G20603: std_logic; attribute dont_touch of G20603: signal is true;
	signal G20604: std_logic; attribute dont_touch of G20604: signal is true;
	signal G20605: std_logic; attribute dont_touch of G20605: signal is true;
	signal G20606: std_logic; attribute dont_touch of G20606: signal is true;
	signal G20607: std_logic; attribute dont_touch of G20607: signal is true;
	signal G20608: std_logic; attribute dont_touch of G20608: signal is true;
	signal G20609: std_logic; attribute dont_touch of G20609: signal is true;
	signal G20610: std_logic; attribute dont_touch of G20610: signal is true;
	signal G20611: std_logic; attribute dont_touch of G20611: signal is true;
	signal G20612: std_logic; attribute dont_touch of G20612: signal is true;
	signal G20613: std_logic; attribute dont_touch of G20613: signal is true;
	signal G20614: std_logic; attribute dont_touch of G20614: signal is true;
	signal G20615: std_logic; attribute dont_touch of G20615: signal is true;
	signal G20616: std_logic; attribute dont_touch of G20616: signal is true;
	signal G20617: std_logic; attribute dont_touch of G20617: signal is true;
	signal G20618: std_logic; attribute dont_touch of G20618: signal is true;
	signal G20619: std_logic; attribute dont_touch of G20619: signal is true;
	signal G20622: std_logic; attribute dont_touch of G20622: signal is true;
	signal G20623: std_logic; attribute dont_touch of G20623: signal is true;
	signal G20624: std_logic; attribute dont_touch of G20624: signal is true;
	signal G20625: std_logic; attribute dont_touch of G20625: signal is true;
	signal G20626: std_logic; attribute dont_touch of G20626: signal is true;
	signal G20627: std_logic; attribute dont_touch of G20627: signal is true;
	signal G20628: std_logic; attribute dont_touch of G20628: signal is true;
	signal G20629: std_logic; attribute dont_touch of G20629: signal is true;
	signal G20630: std_logic; attribute dont_touch of G20630: signal is true;
	signal G20631: std_logic; attribute dont_touch of G20631: signal is true;
	signal G20632: std_logic; attribute dont_touch of G20632: signal is true;
	signal G20633: std_logic; attribute dont_touch of G20633: signal is true;
	signal G20634: std_logic; attribute dont_touch of G20634: signal is true;
	signal G20635: std_logic; attribute dont_touch of G20635: signal is true;
	signal G20636: std_logic; attribute dont_touch of G20636: signal is true;
	signal G20637: std_logic; attribute dont_touch of G20637: signal is true;
	signal G20638: std_logic; attribute dont_touch of G20638: signal is true;
	signal G20639: std_logic; attribute dont_touch of G20639: signal is true;
	signal G20640: std_logic; attribute dont_touch of G20640: signal is true;
	signal G20641: std_logic; attribute dont_touch of G20641: signal is true;
	signal G20642: std_logic; attribute dont_touch of G20642: signal is true;
	signal G20643: std_logic; attribute dont_touch of G20643: signal is true;
	signal G20644: std_logic; attribute dont_touch of G20644: signal is true;
	signal G20645: std_logic; attribute dont_touch of G20645: signal is true;
	signal G20648: std_logic; attribute dont_touch of G20648: signal is true;
	signal G20649: std_logic; attribute dont_touch of G20649: signal is true;
	signal G20650: std_logic; attribute dont_touch of G20650: signal is true;
	signal G20651: std_logic; attribute dont_touch of G20651: signal is true;
	signal G20653: std_logic; attribute dont_touch of G20653: signal is true;
	signal G20655: std_logic; attribute dont_touch of G20655: signal is true;
	signal G20656: std_logic; attribute dont_touch of G20656: signal is true;
	signal G20657: std_logic; attribute dont_touch of G20657: signal is true;
	signal G20658: std_logic; attribute dont_touch of G20658: signal is true;
	signal G20659: std_logic; attribute dont_touch of G20659: signal is true;
	signal G20660: std_logic; attribute dont_touch of G20660: signal is true;
	signal G20661: std_logic; attribute dont_touch of G20661: signal is true;
	signal G20662: std_logic; attribute dont_touch of G20662: signal is true;
	signal G20663: std_logic; attribute dont_touch of G20663: signal is true;
	signal G20664: std_logic; attribute dont_touch of G20664: signal is true;
	signal G20665: std_logic; attribute dont_touch of G20665: signal is true;
	signal G20666: std_logic; attribute dont_touch of G20666: signal is true;
	signal G20667: std_logic; attribute dont_touch of G20667: signal is true;
	signal G20668: std_logic; attribute dont_touch of G20668: signal is true;
	signal G20669: std_logic; attribute dont_touch of G20669: signal is true;
	signal G20670: std_logic; attribute dont_touch of G20670: signal is true;
	signal G20671: std_logic; attribute dont_touch of G20671: signal is true;
	signal G20672: std_logic; attribute dont_touch of G20672: signal is true;
	signal G20673: std_logic; attribute dont_touch of G20673: signal is true;
	signal G20674: std_logic; attribute dont_touch of G20674: signal is true;
	signal G20675: std_logic; attribute dont_touch of G20675: signal is true;
	signal G20676: std_logic; attribute dont_touch of G20676: signal is true;
	signal G20679: std_logic; attribute dont_touch of G20679: signal is true;
	signal G20680: std_logic; attribute dont_touch of G20680: signal is true;
	signal G20681: std_logic; attribute dont_touch of G20681: signal is true;
	signal G20682: std_logic; attribute dont_touch of G20682: signal is true;
	signal G20695: std_logic; attribute dont_touch of G20695: signal is true;
	signal G20696: std_logic; attribute dont_touch of G20696: signal is true;
	signal G20697: std_logic; attribute dont_touch of G20697: signal is true;
	signal G20698: std_logic; attribute dont_touch of G20698: signal is true;
	signal G20699: std_logic; attribute dont_touch of G20699: signal is true;
	signal G20700: std_logic; attribute dont_touch of G20700: signal is true;
	signal G20701: std_logic; attribute dont_touch of G20701: signal is true;
	signal G20702: std_logic; attribute dont_touch of G20702: signal is true;
	signal G20703: std_logic; attribute dont_touch of G20703: signal is true;
	signal G20704: std_logic; attribute dont_touch of G20704: signal is true;
	signal G20705: std_logic; attribute dont_touch of G20705: signal is true;
	signal G20706: std_logic; attribute dont_touch of G20706: signal is true;
	signal G20707: std_logic; attribute dont_touch of G20707: signal is true;
	signal G20708: std_logic; attribute dont_touch of G20708: signal is true;
	signal G20709: std_logic; attribute dont_touch of G20709: signal is true;
	signal G20710: std_logic; attribute dont_touch of G20710: signal is true;
	signal G20711: std_logic; attribute dont_touch of G20711: signal is true;
	signal G20712: std_logic; attribute dont_touch of G20712: signal is true;
	signal G20713: std_logic; attribute dont_touch of G20713: signal is true;
	signal G20714: std_logic; attribute dont_touch of G20714: signal is true;
	signal G20715: std_logic; attribute dont_touch of G20715: signal is true;
	signal G20716: std_logic; attribute dont_touch of G20716: signal is true;
	signal G20717: std_logic; attribute dont_touch of G20717: signal is true;
	signal G20720: std_logic; attribute dont_touch of G20720: signal is true;
	signal G20732: std_logic; attribute dont_touch of G20732: signal is true;
	signal G20733: std_logic; attribute dont_touch of G20733: signal is true;
	signal G20734: std_logic; attribute dont_touch of G20734: signal is true;
	signal G20737: std_logic; attribute dont_touch of G20737: signal is true;
	signal G20738: std_logic; attribute dont_touch of G20738: signal is true;
	signal G20739: std_logic; attribute dont_touch of G20739: signal is true;
	signal G20751: std_logic; attribute dont_touch of G20751: signal is true;
	signal G20764: std_logic; attribute dont_touch of G20764: signal is true;
	signal G20765: std_logic; attribute dont_touch of G20765: signal is true;
	signal G20766: std_logic; attribute dont_touch of G20766: signal is true;
	signal G20767: std_logic; attribute dont_touch of G20767: signal is true;
	signal G20768: std_logic; attribute dont_touch of G20768: signal is true;
	signal G20769: std_logic; attribute dont_touch of G20769: signal is true;
	signal G20770: std_logic; attribute dont_touch of G20770: signal is true;
	signal G20771: std_logic; attribute dont_touch of G20771: signal is true;
	signal G20772: std_logic; attribute dont_touch of G20772: signal is true;
	signal G20773: std_logic; attribute dont_touch of G20773: signal is true;
	signal G20774: std_logic; attribute dont_touch of G20774: signal is true;
	signal G20775: std_logic; attribute dont_touch of G20775: signal is true;
	signal G20776: std_logic; attribute dont_touch of G20776: signal is true;
	signal G20777: std_logic; attribute dont_touch of G20777: signal is true;
	signal G20778: std_logic; attribute dont_touch of G20778: signal is true;
	signal G20779: std_logic; attribute dont_touch of G20779: signal is true;
	signal G20780: std_logic; attribute dont_touch of G20780: signal is true;
	signal G20781: std_logic; attribute dont_touch of G20781: signal is true;
	signal G20782: std_logic; attribute dont_touch of G20782: signal is true;
	signal G20783: std_logic; attribute dont_touch of G20783: signal is true;
	signal G20784: std_logic; attribute dont_touch of G20784: signal is true;
	signal G20785: std_logic; attribute dont_touch of G20785: signal is true;
	signal G20838: std_logic; attribute dont_touch of G20838: signal is true;
	signal G20841: std_logic; attribute dont_touch of G20841: signal is true;
	signal G20852: std_logic; attribute dont_touch of G20852: signal is true;
	signal G20853: std_logic; attribute dont_touch of G20853: signal is true;
	signal G20854: std_logic; attribute dont_touch of G20854: signal is true;
	signal G20857: std_logic; attribute dont_touch of G20857: signal is true;
	signal G20869: std_logic; attribute dont_touch of G20869: signal is true;
	signal G20870: std_logic; attribute dont_touch of G20870: signal is true;
	signal G20871: std_logic; attribute dont_touch of G20871: signal is true;
	signal G20874: std_logic; attribute dont_touch of G20874: signal is true;
	signal G20875: std_logic; attribute dont_touch of G20875: signal is true;
	signal G20887: std_logic; attribute dont_touch of G20887: signal is true;
	signal G20900: std_logic; attribute dont_touch of G20900: signal is true;
	signal G20902: std_logic; attribute dont_touch of G20902: signal is true;
	signal G20903: std_logic; attribute dont_touch of G20903: signal is true;
	signal G20904: std_logic; attribute dont_touch of G20904: signal is true;
	signal G20905: std_logic; attribute dont_touch of G20905: signal is true;
	signal G20909: std_logic; attribute dont_touch of G20909: signal is true;
	signal G20910: std_logic; attribute dont_touch of G20910: signal is true;
	signal G20911: std_logic; attribute dont_touch of G20911: signal is true;
	signal G20912: std_logic; attribute dont_touch of G20912: signal is true;
	signal G20913: std_logic; attribute dont_touch of G20913: signal is true;
	signal G20914: std_logic; attribute dont_touch of G20914: signal is true;
	signal G20915: std_logic; attribute dont_touch of G20915: signal is true;
	signal G20916: std_logic; attribute dont_touch of G20916: signal is true;
	signal G20917: std_logic; attribute dont_touch of G20917: signal is true;
	signal G20918: std_logic; attribute dont_touch of G20918: signal is true;
	signal G20919: std_logic; attribute dont_touch of G20919: signal is true;
	signal G20920: std_logic; attribute dont_touch of G20920: signal is true;
	signal G20921: std_logic; attribute dont_touch of G20921: signal is true;
	signal G20922: std_logic; attribute dont_touch of G20922: signal is true;
	signal G20923: std_logic; attribute dont_touch of G20923: signal is true;
	signal G20924: std_logic; attribute dont_touch of G20924: signal is true;
	signal G20977: std_logic; attribute dont_touch of G20977: signal is true;
	signal G20978: std_logic; attribute dont_touch of G20978: signal is true;
	signal G20979: std_logic; attribute dont_touch of G20979: signal is true;
	signal G20982: std_logic; attribute dont_touch of G20982: signal is true;
	signal G20993: std_logic; attribute dont_touch of G20993: signal is true;
	signal G20994: std_logic; attribute dont_touch of G20994: signal is true;
	signal G20995: std_logic; attribute dont_touch of G20995: signal is true;
	signal G20998: std_logic; attribute dont_touch of G20998: signal is true;
	signal G21010: std_logic; attribute dont_touch of G21010: signal is true;
	signal G21011: std_logic; attribute dont_touch of G21011: signal is true;
	signal G21012: std_logic; attribute dont_touch of G21012: signal is true;
	signal G21024: std_logic; attribute dont_touch of G21024: signal is true;
	signal G21036: std_logic; attribute dont_touch of G21036: signal is true;
	signal G21037: std_logic; attribute dont_touch of G21037: signal is true;
	signal G21048: std_logic; attribute dont_touch of G21048: signal is true;
	signal G21049: std_logic; attribute dont_touch of G21049: signal is true;
	signal G21050: std_logic; attribute dont_touch of G21050: signal is true;
	signal G21051: std_logic; attribute dont_touch of G21051: signal is true;
	signal G21052: std_logic; attribute dont_touch of G21052: signal is true;
	signal G21053: std_logic; attribute dont_touch of G21053: signal is true;
	signal G21054: std_logic; attribute dont_touch of G21054: signal is true;
	signal G21055: std_logic; attribute dont_touch of G21055: signal is true;
	signal G21056: std_logic; attribute dont_touch of G21056: signal is true;
	signal G21057: std_logic; attribute dont_touch of G21057: signal is true;
	signal G21058: std_logic; attribute dont_touch of G21058: signal is true;
	signal G21059: std_logic; attribute dont_touch of G21059: signal is true;
	signal G21060: std_logic; attribute dont_touch of G21060: signal is true;
	signal G21061: std_logic; attribute dont_touch of G21061: signal is true;
	signal G21062: std_logic; attribute dont_touch of G21062: signal is true;
	signal G21066: std_logic; attribute dont_touch of G21066: signal is true;
	signal G21067: std_logic; attribute dont_touch of G21067: signal is true;
	signal G21068: std_logic; attribute dont_touch of G21068: signal is true;
	signal G21069: std_logic; attribute dont_touch of G21069: signal is true;
	signal G21070: std_logic; attribute dont_touch of G21070: signal is true;
	signal G21123: std_logic; attribute dont_touch of G21123: signal is true;
	signal G21124: std_logic; attribute dont_touch of G21124: signal is true;
	signal G21127: std_logic; attribute dont_touch of G21127: signal is true;
	signal G21138: std_logic; attribute dont_touch of G21138: signal is true;
	signal G21139: std_logic; attribute dont_touch of G21139: signal is true;
	signal G21140: std_logic; attribute dont_touch of G21140: signal is true;
	signal G21143: std_logic; attribute dont_touch of G21143: signal is true;
	signal G21155: std_logic; attribute dont_touch of G21155: signal is true;
	signal G21156: std_logic; attribute dont_touch of G21156: signal is true;
	signal G21160: std_logic; attribute dont_touch of G21160: signal is true;
	signal G21163: std_logic; attribute dont_touch of G21163: signal is true;
	signal G21175: std_logic; attribute dont_touch of G21175: signal is true;
	signal G21177: std_logic; attribute dont_touch of G21177: signal is true;
	signal G21178: std_logic; attribute dont_touch of G21178: signal is true;
	signal G21179: std_logic; attribute dont_touch of G21179: signal is true;
	signal G21180: std_logic; attribute dont_touch of G21180: signal is true;
	signal G21181: std_logic; attribute dont_touch of G21181: signal is true;
	signal G21182: std_logic; attribute dont_touch of G21182: signal is true;
	signal G21183: std_logic; attribute dont_touch of G21183: signal is true;
	signal G21184: std_logic; attribute dont_touch of G21184: signal is true;
	signal G21185: std_logic; attribute dont_touch of G21185: signal is true;
	signal G21186: std_logic; attribute dont_touch of G21186: signal is true;
	signal G21187: std_logic; attribute dont_touch of G21187: signal is true;
	signal G21188: std_logic; attribute dont_touch of G21188: signal is true;
	signal G21189: std_logic; attribute dont_touch of G21189: signal is true;
	signal G21190: std_logic; attribute dont_touch of G21190: signal is true;
	signal G21193: std_logic; attribute dont_touch of G21193: signal is true;
	signal G21204: std_logic; attribute dont_touch of G21204: signal is true;
	signal G21205: std_logic; attribute dont_touch of G21205: signal is true;
	signal G21206: std_logic; attribute dont_touch of G21206: signal is true;
	signal G21209: std_logic; attribute dont_touch of G21209: signal is true;
	signal G21221: std_logic; attribute dont_touch of G21221: signal is true;
	signal G21222: std_logic; attribute dont_touch of G21222: signal is true;
	signal G21225: std_logic; attribute dont_touch of G21225: signal is true;
	signal G21228: std_logic; attribute dont_touch of G21228: signal is true;
	signal G21246: std_logic; attribute dont_touch of G21246: signal is true;
	signal G21247: std_logic; attribute dont_touch of G21247: signal is true;
	signal G21248: std_logic; attribute dont_touch of G21248: signal is true;
	signal G21249: std_logic; attribute dont_touch of G21249: signal is true;
	signal G21250: std_logic; attribute dont_touch of G21250: signal is true;
	signal G21251: std_logic; attribute dont_touch of G21251: signal is true;
	signal G21252: std_logic; attribute dont_touch of G21252: signal is true;
	signal G21253: std_logic; attribute dont_touch of G21253: signal is true;
	signal G21256: std_logic; attribute dont_touch of G21256: signal is true;
	signal G21267: std_logic; attribute dont_touch of G21267: signal is true;
	signal G21268: std_logic; attribute dont_touch of G21268: signal is true;
	signal G21269: std_logic; attribute dont_touch of G21269: signal is true;
	signal G21271: std_logic; attribute dont_touch of G21271: signal is true;
	signal G21272: std_logic; attribute dont_touch of G21272: signal is true;
	signal G21273: std_logic; attribute dont_touch of G21273: signal is true;
	signal G21274: std_logic; attribute dont_touch of G21274: signal is true;
	signal G21275: std_logic; attribute dont_touch of G21275: signal is true;
	signal G21276: std_logic; attribute dont_touch of G21276: signal is true;
	signal G21277: std_logic; attribute dont_touch of G21277: signal is true;
	signal G21278: std_logic; attribute dont_touch of G21278: signal is true;
	signal G21279: std_logic; attribute dont_touch of G21279: signal is true;
	signal G21280: std_logic; attribute dont_touch of G21280: signal is true;
	signal G21281: std_logic; attribute dont_touch of G21281: signal is true;
	signal G21282: std_logic; attribute dont_touch of G21282: signal is true;
	signal G21283: std_logic; attribute dont_touch of G21283: signal is true;
	signal G21284: std_logic; attribute dont_touch of G21284: signal is true;
	signal G21285: std_logic; attribute dont_touch of G21285: signal is true;
	signal G21286: std_logic; attribute dont_touch of G21286: signal is true;
	signal G21287: std_logic; attribute dont_touch of G21287: signal is true;
	signal G21288: std_logic; attribute dont_touch of G21288: signal is true;
	signal G21289: std_logic; attribute dont_touch of G21289: signal is true;
	signal G21290: std_logic; attribute dont_touch of G21290: signal is true;
	signal G21291: std_logic; attribute dont_touch of G21291: signal is true;
	signal G21293: std_logic; attribute dont_touch of G21293: signal is true;
	signal G21294: std_logic; attribute dont_touch of G21294: signal is true;
	signal G21295: std_logic; attribute dont_touch of G21295: signal is true;
	signal G21296: std_logic; attribute dont_touch of G21296: signal is true;
	signal G21297: std_logic; attribute dont_touch of G21297: signal is true;
	signal G21298: std_logic; attribute dont_touch of G21298: signal is true;
	signal G21299: std_logic; attribute dont_touch of G21299: signal is true;
	signal G21300: std_logic; attribute dont_touch of G21300: signal is true;
	signal G21301: std_logic; attribute dont_touch of G21301: signal is true;
	signal G21302: std_logic; attribute dont_touch of G21302: signal is true;
	signal G21303: std_logic; attribute dont_touch of G21303: signal is true;
	signal G21304: std_logic; attribute dont_touch of G21304: signal is true;
	signal G21305: std_logic; attribute dont_touch of G21305: signal is true;
	signal G21306: std_logic; attribute dont_touch of G21306: signal is true;
	signal G21307: std_logic; attribute dont_touch of G21307: signal is true;
	signal G21308: std_logic; attribute dont_touch of G21308: signal is true;
	signal G21326: std_logic; attribute dont_touch of G21326: signal is true;
	signal G21329: std_logic; attribute dont_touch of G21329: signal is true;
	signal G21330: std_logic; attribute dont_touch of G21330: signal is true;
	signal G21331: std_logic; attribute dont_touch of G21331: signal is true;
	signal G21332: std_logic; attribute dont_touch of G21332: signal is true;
	signal G21333: std_logic; attribute dont_touch of G21333: signal is true;
	signal G21334: std_logic; attribute dont_touch of G21334: signal is true;
	signal G21335: std_logic; attribute dont_touch of G21335: signal is true;
	signal G21336: std_logic; attribute dont_touch of G21336: signal is true;
	signal G21337: std_logic; attribute dont_touch of G21337: signal is true;
	signal G21338: std_logic; attribute dont_touch of G21338: signal is true;
	signal G21339: std_logic; attribute dont_touch of G21339: signal is true;
	signal G21340: std_logic; attribute dont_touch of G21340: signal is true;
	signal G21343: std_logic; attribute dont_touch of G21343: signal is true;
	signal G21344: std_logic; attribute dont_touch of G21344: signal is true;
	signal G21345: std_logic; attribute dont_touch of G21345: signal is true;
	signal G21346: std_logic; attribute dont_touch of G21346: signal is true;
	signal G21347: std_logic; attribute dont_touch of G21347: signal is true;
	signal G21348: std_logic; attribute dont_touch of G21348: signal is true;
	signal G21349: std_logic; attribute dont_touch of G21349: signal is true;
	signal G21350: std_logic; attribute dont_touch of G21350: signal is true;
	signal G21351: std_logic; attribute dont_touch of G21351: signal is true;
	signal G21352: std_logic; attribute dont_touch of G21352: signal is true;
	signal G21353: std_logic; attribute dont_touch of G21353: signal is true;
	signal G21354: std_logic; attribute dont_touch of G21354: signal is true;
	signal G21355: std_logic; attribute dont_touch of G21355: signal is true;
	signal G21356: std_logic; attribute dont_touch of G21356: signal is true;
	signal G21357: std_logic; attribute dont_touch of G21357: signal is true;
	signal G21358: std_logic; attribute dont_touch of G21358: signal is true;
	signal G21359: std_logic; attribute dont_touch of G21359: signal is true;
	signal G21360: std_logic; attribute dont_touch of G21360: signal is true;
	signal G21361: std_logic; attribute dont_touch of G21361: signal is true;
	signal G21362: std_logic; attribute dont_touch of G21362: signal is true;
	signal G21363: std_logic; attribute dont_touch of G21363: signal is true;
	signal G21364: std_logic; attribute dont_touch of G21364: signal is true;
	signal G21365: std_logic; attribute dont_touch of G21365: signal is true;
	signal G21366: std_logic; attribute dont_touch of G21366: signal is true;
	signal G21369: std_logic; attribute dont_touch of G21369: signal is true;
	signal G21370: std_logic; attribute dont_touch of G21370: signal is true;
	signal G21377: std_logic; attribute dont_touch of G21377: signal is true;
	signal G21378: std_logic; attribute dont_touch of G21378: signal is true;
	signal G21379: std_logic; attribute dont_touch of G21379: signal is true;
	signal G21380: std_logic; attribute dont_touch of G21380: signal is true;
	signal G21381: std_logic; attribute dont_touch of G21381: signal is true;
	signal G21382: std_logic; attribute dont_touch of G21382: signal is true;
	signal G21383: std_logic; attribute dont_touch of G21383: signal is true;
	signal G21384: std_logic; attribute dont_touch of G21384: signal is true;
	signal G21385: std_logic; attribute dont_touch of G21385: signal is true;
	signal G21386: std_logic; attribute dont_touch of G21386: signal is true;
	signal G21387: std_logic; attribute dont_touch of G21387: signal is true;
	signal G21388: std_logic; attribute dont_touch of G21388: signal is true;
	signal G21389: std_logic; attribute dont_touch of G21389: signal is true;
	signal G21393: std_logic; attribute dont_touch of G21393: signal is true;
	signal G21394: std_logic; attribute dont_touch of G21394: signal is true;
	signal G21395: std_logic; attribute dont_touch of G21395: signal is true;
	signal G21396: std_logic; attribute dont_touch of G21396: signal is true;
	signal G21397: std_logic; attribute dont_touch of G21397: signal is true;
	signal G21398: std_logic; attribute dont_touch of G21398: signal is true;
	signal G21399: std_logic; attribute dont_touch of G21399: signal is true;
	signal G21400: std_logic; attribute dont_touch of G21400: signal is true;
	signal G21401: std_logic; attribute dont_touch of G21401: signal is true;
	signal G21402: std_logic; attribute dont_touch of G21402: signal is true;
	signal G21403: std_logic; attribute dont_touch of G21403: signal is true;
	signal G21404: std_logic; attribute dont_touch of G21404: signal is true;
	signal G21405: std_logic; attribute dont_touch of G21405: signal is true;
	signal G21406: std_logic; attribute dont_touch of G21406: signal is true;
	signal G21407: std_logic; attribute dont_touch of G21407: signal is true;
	signal G21408: std_logic; attribute dont_touch of G21408: signal is true;
	signal G21409: std_logic; attribute dont_touch of G21409: signal is true;
	signal G21410: std_logic; attribute dont_touch of G21410: signal is true;
	signal G21411: std_logic; attribute dont_touch of G21411: signal is true;
	signal G21412: std_logic; attribute dont_touch of G21412: signal is true;
	signal G21413: std_logic; attribute dont_touch of G21413: signal is true;
	signal G21414: std_logic; attribute dont_touch of G21414: signal is true;
	signal G21415: std_logic; attribute dont_touch of G21415: signal is true;
	signal G21416: std_logic; attribute dont_touch of G21416: signal is true;
	signal G21417: std_logic; attribute dont_touch of G21417: signal is true;
	signal G21418: std_logic; attribute dont_touch of G21418: signal is true;
	signal G21419: std_logic; attribute dont_touch of G21419: signal is true;
	signal G21420: std_logic; attribute dont_touch of G21420: signal is true;
	signal G21421: std_logic; attribute dont_touch of G21421: signal is true;
	signal G21422: std_logic; attribute dont_touch of G21422: signal is true;
	signal G21423: std_logic; attribute dont_touch of G21423: signal is true;
	signal G21424: std_logic; attribute dont_touch of G21424: signal is true;
	signal G21425: std_logic; attribute dont_touch of G21425: signal is true;
	signal G21426: std_logic; attribute dont_touch of G21426: signal is true;
	signal G21427: std_logic; attribute dont_touch of G21427: signal is true;
	signal G21428: std_logic; attribute dont_touch of G21428: signal is true;
	signal G21429: std_logic; attribute dont_touch of G21429: signal is true;
	signal G21430: std_logic; attribute dont_touch of G21430: signal is true;
	signal G21431: std_logic; attribute dont_touch of G21431: signal is true;
	signal G21432: std_logic; attribute dont_touch of G21432: signal is true;
	signal G21433: std_logic; attribute dont_touch of G21433: signal is true;
	signal G21434: std_logic; attribute dont_touch of G21434: signal is true;
	signal G21451: std_logic; attribute dont_touch of G21451: signal is true;
	signal G21452: std_logic; attribute dont_touch of G21452: signal is true;
	signal G21453: std_logic; attribute dont_touch of G21453: signal is true;
	signal G21454: std_logic; attribute dont_touch of G21454: signal is true;
	signal G21455: std_logic; attribute dont_touch of G21455: signal is true;
	signal G21456: std_logic; attribute dont_touch of G21456: signal is true;
	signal G21457: std_logic; attribute dont_touch of G21457: signal is true;
	signal G21458: std_logic; attribute dont_touch of G21458: signal is true;
	signal G21459: std_logic; attribute dont_touch of G21459: signal is true;
	signal G21460: std_logic; attribute dont_touch of G21460: signal is true;
	signal G21461: std_logic; attribute dont_touch of G21461: signal is true;
	signal G21462: std_logic; attribute dont_touch of G21462: signal is true;
	signal G21463: std_logic; attribute dont_touch of G21463: signal is true;
	signal G21464: std_logic; attribute dont_touch of G21464: signal is true;
	signal G21465: std_logic; attribute dont_touch of G21465: signal is true;
	signal G21466: std_logic; attribute dont_touch of G21466: signal is true;
	signal G21467: std_logic; attribute dont_touch of G21467: signal is true;
	signal G21468: std_logic; attribute dont_touch of G21468: signal is true;
	signal G21509: std_logic; attribute dont_touch of G21509: signal is true;
	signal G21510: std_logic; attribute dont_touch of G21510: signal is true;
	signal G21511: std_logic; attribute dont_touch of G21511: signal is true;
	signal G21512: std_logic; attribute dont_touch of G21512: signal is true;
	signal G21513: std_logic; attribute dont_touch of G21513: signal is true;
	signal G21514: std_logic; attribute dont_touch of G21514: signal is true;
	signal G21555: std_logic; attribute dont_touch of G21555: signal is true;
	signal G21556: std_logic; attribute dont_touch of G21556: signal is true;
	signal G21557: std_logic; attribute dont_touch of G21557: signal is true;
	signal G21558: std_logic; attribute dont_touch of G21558: signal is true;
	signal G21559: std_logic; attribute dont_touch of G21559: signal is true;
	signal G21560: std_logic; attribute dont_touch of G21560: signal is true;
	signal G21561: std_logic; attribute dont_touch of G21561: signal is true;
	signal G21562: std_logic; attribute dont_touch of G21562: signal is true;
	signal G21603: std_logic; attribute dont_touch of G21603: signal is true;
	signal G21604: std_logic; attribute dont_touch of G21604: signal is true;
	signal G21605: std_logic; attribute dont_touch of G21605: signal is true;
	signal G21606: std_logic; attribute dont_touch of G21606: signal is true;
	signal G21607: std_logic; attribute dont_touch of G21607: signal is true;
	signal G21608: std_logic; attribute dont_touch of G21608: signal is true;
	signal G21609: std_logic; attribute dont_touch of G21609: signal is true;
	signal G21610: std_logic; attribute dont_touch of G21610: signal is true;
	signal G21611: std_logic; attribute dont_touch of G21611: signal is true;
	signal G21652: std_logic; attribute dont_touch of G21652: signal is true;
	signal G21653: std_logic; attribute dont_touch of G21653: signal is true;
	signal G21654: std_logic; attribute dont_touch of G21654: signal is true;
	signal G21655: std_logic; attribute dont_touch of G21655: signal is true;
	signal G21656: std_logic; attribute dont_touch of G21656: signal is true;
	signal G21657: std_logic; attribute dont_touch of G21657: signal is true;
	signal G21658: std_logic; attribute dont_touch of G21658: signal is true;
	signal G21659: std_logic; attribute dont_touch of G21659: signal is true;
	signal G21660: std_logic; attribute dont_touch of G21660: signal is true;
	signal G21661: std_logic; attribute dont_touch of G21661: signal is true;
	signal G21662: std_logic; attribute dont_touch of G21662: signal is true;
	signal G21665: std_logic; attribute dont_touch of G21665: signal is true;
	signal G21666: std_logic; attribute dont_touch of G21666: signal is true;
	signal G21669: std_logic; attribute dont_touch of G21669: signal is true;
	signal G21670: std_logic; attribute dont_touch of G21670: signal is true;
	signal G21673: std_logic; attribute dont_touch of G21673: signal is true;
	signal G21674: std_logic; attribute dont_touch of G21674: signal is true;
	signal G21677: std_logic; attribute dont_touch of G21677: signal is true;
	signal G21678: std_logic; attribute dont_touch of G21678: signal is true;
	signal G21681: std_logic; attribute dont_touch of G21681: signal is true;
	signal G21682: std_logic; attribute dont_touch of G21682: signal is true;
	signal G21685: std_logic; attribute dont_touch of G21685: signal is true;
	signal G21686: std_logic; attribute dont_touch of G21686: signal is true;
	signal G21689: std_logic; attribute dont_touch of G21689: signal is true;
	signal G21690: std_logic; attribute dont_touch of G21690: signal is true;
	signal G21693: std_logic; attribute dont_touch of G21693: signal is true;
	signal G21694: std_logic; attribute dont_touch of G21694: signal is true;
	signal G21697: std_logic; attribute dont_touch of G21697: signal is true;
	signal G21699: std_logic; attribute dont_touch of G21699: signal is true;
	signal G21700: std_logic; attribute dont_touch of G21700: signal is true;
	signal G21701: std_logic; attribute dont_touch of G21701: signal is true;
	signal G21702: std_logic; attribute dont_touch of G21702: signal is true;
	signal G21703: std_logic; attribute dont_touch of G21703: signal is true;
	signal G21704: std_logic; attribute dont_touch of G21704: signal is true;
	signal G21705: std_logic; attribute dont_touch of G21705: signal is true;
	signal G21706: std_logic; attribute dont_touch of G21706: signal is true;
	signal G21707: std_logic; attribute dont_touch of G21707: signal is true;
	signal G21708: std_logic; attribute dont_touch of G21708: signal is true;
	signal G21709: std_logic; attribute dont_touch of G21709: signal is true;
	signal G21710: std_logic; attribute dont_touch of G21710: signal is true;
	signal G21711: std_logic; attribute dont_touch of G21711: signal is true;
	signal G21712: std_logic; attribute dont_touch of G21712: signal is true;
	signal G21713: std_logic; attribute dont_touch of G21713: signal is true;
	signal G21714: std_logic; attribute dont_touch of G21714: signal is true;
	signal G21715: std_logic; attribute dont_touch of G21715: signal is true;
	signal G21716: std_logic; attribute dont_touch of G21716: signal is true;
	signal G21717: std_logic; attribute dont_touch of G21717: signal is true;
	signal G21718: std_logic; attribute dont_touch of G21718: signal is true;
	signal G21719: std_logic; attribute dont_touch of G21719: signal is true;
	signal G21720: std_logic; attribute dont_touch of G21720: signal is true;
	signal G21721: std_logic; attribute dont_touch of G21721: signal is true;
	signal G21722: std_logic; attribute dont_touch of G21722: signal is true;
	signal G21723: std_logic; attribute dont_touch of G21723: signal is true;
	signal G21724: std_logic; attribute dont_touch of G21724: signal is true;
	signal G21725: std_logic; attribute dont_touch of G21725: signal is true;
	signal G21726: std_logic; attribute dont_touch of G21726: signal is true;
	signal G21728: std_logic; attribute dont_touch of G21728: signal is true;
	signal G21729: std_logic; attribute dont_touch of G21729: signal is true;
	signal G21730: std_logic; attribute dont_touch of G21730: signal is true;
	signal G21731: std_logic; attribute dont_touch of G21731: signal is true;
	signal G21732: std_logic; attribute dont_touch of G21732: signal is true;
	signal G21733: std_logic; attribute dont_touch of G21733: signal is true;
	signal G21734: std_logic; attribute dont_touch of G21734: signal is true;
	signal G21735: std_logic; attribute dont_touch of G21735: signal is true;
	signal G21736: std_logic; attribute dont_touch of G21736: signal is true;
	signal G21737: std_logic; attribute dont_touch of G21737: signal is true;
	signal G21738: std_logic; attribute dont_touch of G21738: signal is true;
	signal G21739: std_logic; attribute dont_touch of G21739: signal is true;
	signal G21740: std_logic; attribute dont_touch of G21740: signal is true;
	signal G21741: std_logic; attribute dont_touch of G21741: signal is true;
	signal G21742: std_logic; attribute dont_touch of G21742: signal is true;
	signal G21743: std_logic; attribute dont_touch of G21743: signal is true;
	signal G21744: std_logic; attribute dont_touch of G21744: signal is true;
	signal G21745: std_logic; attribute dont_touch of G21745: signal is true;
	signal G21746: std_logic; attribute dont_touch of G21746: signal is true;
	signal G21747: std_logic; attribute dont_touch of G21747: signal is true;
	signal G21748: std_logic; attribute dont_touch of G21748: signal is true;
	signal G21749: std_logic; attribute dont_touch of G21749: signal is true;
	signal G21750: std_logic; attribute dont_touch of G21750: signal is true;
	signal G21751: std_logic; attribute dont_touch of G21751: signal is true;
	signal G21752: std_logic; attribute dont_touch of G21752: signal is true;
	signal G21753: std_logic; attribute dont_touch of G21753: signal is true;
	signal G21754: std_logic; attribute dont_touch of G21754: signal is true;
	signal G21755: std_logic; attribute dont_touch of G21755: signal is true;
	signal G21756: std_logic; attribute dont_touch of G21756: signal is true;
	signal G21757: std_logic; attribute dont_touch of G21757: signal is true;
	signal G21758: std_logic; attribute dont_touch of G21758: signal is true;
	signal G21759: std_logic; attribute dont_touch of G21759: signal is true;
	signal G21760: std_logic; attribute dont_touch of G21760: signal is true;
	signal G21761: std_logic; attribute dont_touch of G21761: signal is true;
	signal G21762: std_logic; attribute dont_touch of G21762: signal is true;
	signal G21763: std_logic; attribute dont_touch of G21763: signal is true;
	signal G21764: std_logic; attribute dont_touch of G21764: signal is true;
	signal G21765: std_logic; attribute dont_touch of G21765: signal is true;
	signal G21766: std_logic; attribute dont_touch of G21766: signal is true;
	signal G21767: std_logic; attribute dont_touch of G21767: signal is true;
	signal G21768: std_logic; attribute dont_touch of G21768: signal is true;
	signal G21769: std_logic; attribute dont_touch of G21769: signal is true;
	signal G21770: std_logic; attribute dont_touch of G21770: signal is true;
	signal G21771: std_logic; attribute dont_touch of G21771: signal is true;
	signal G21772: std_logic; attribute dont_touch of G21772: signal is true;
	signal G21773: std_logic; attribute dont_touch of G21773: signal is true;
	signal G21774: std_logic; attribute dont_touch of G21774: signal is true;
	signal G21775: std_logic; attribute dont_touch of G21775: signal is true;
	signal G21776: std_logic; attribute dont_touch of G21776: signal is true;
	signal G21777: std_logic; attribute dont_touch of G21777: signal is true;
	signal G21778: std_logic; attribute dont_touch of G21778: signal is true;
	signal G21779: std_logic; attribute dont_touch of G21779: signal is true;
	signal G21780: std_logic; attribute dont_touch of G21780: signal is true;
	signal G21781: std_logic; attribute dont_touch of G21781: signal is true;
	signal G21782: std_logic; attribute dont_touch of G21782: signal is true;
	signal G21783: std_logic; attribute dont_touch of G21783: signal is true;
	signal G21784: std_logic; attribute dont_touch of G21784: signal is true;
	signal G21785: std_logic; attribute dont_touch of G21785: signal is true;
	signal G21786: std_logic; attribute dont_touch of G21786: signal is true;
	signal G21787: std_logic; attribute dont_touch of G21787: signal is true;
	signal G21788: std_logic; attribute dont_touch of G21788: signal is true;
	signal G21789: std_logic; attribute dont_touch of G21789: signal is true;
	signal G21790: std_logic; attribute dont_touch of G21790: signal is true;
	signal G21791: std_logic; attribute dont_touch of G21791: signal is true;
	signal G21792: std_logic; attribute dont_touch of G21792: signal is true;
	signal G21793: std_logic; attribute dont_touch of G21793: signal is true;
	signal G21794: std_logic; attribute dont_touch of G21794: signal is true;
	signal G21795: std_logic; attribute dont_touch of G21795: signal is true;
	signal G21796: std_logic; attribute dont_touch of G21796: signal is true;
	signal G21797: std_logic; attribute dont_touch of G21797: signal is true;
	signal G21798: std_logic; attribute dont_touch of G21798: signal is true;
	signal G21799: std_logic; attribute dont_touch of G21799: signal is true;
	signal G21800: std_logic; attribute dont_touch of G21800: signal is true;
	signal G21801: std_logic; attribute dont_touch of G21801: signal is true;
	signal G21802: std_logic; attribute dont_touch of G21802: signal is true;
	signal G21803: std_logic; attribute dont_touch of G21803: signal is true;
	signal G21804: std_logic; attribute dont_touch of G21804: signal is true;
	signal G21805: std_logic; attribute dont_touch of G21805: signal is true;
	signal G21806: std_logic; attribute dont_touch of G21806: signal is true;
	signal G21807: std_logic; attribute dont_touch of G21807: signal is true;
	signal G21808: std_logic; attribute dont_touch of G21808: signal is true;
	signal G21809: std_logic; attribute dont_touch of G21809: signal is true;
	signal G21810: std_logic; attribute dont_touch of G21810: signal is true;
	signal G21811: std_logic; attribute dont_touch of G21811: signal is true;
	signal G21812: std_logic; attribute dont_touch of G21812: signal is true;
	signal G21813: std_logic; attribute dont_touch of G21813: signal is true;
	signal G21814: std_logic; attribute dont_touch of G21814: signal is true;
	signal G21815: std_logic; attribute dont_touch of G21815: signal is true;
	signal G21816: std_logic; attribute dont_touch of G21816: signal is true;
	signal G21817: std_logic; attribute dont_touch of G21817: signal is true;
	signal G21818: std_logic; attribute dont_touch of G21818: signal is true;
	signal G21819: std_logic; attribute dont_touch of G21819: signal is true;
	signal G21820: std_logic; attribute dont_touch of G21820: signal is true;
	signal G21821: std_logic; attribute dont_touch of G21821: signal is true;
	signal G21822: std_logic; attribute dont_touch of G21822: signal is true;
	signal G21823: std_logic; attribute dont_touch of G21823: signal is true;
	signal G21824: std_logic; attribute dont_touch of G21824: signal is true;
	signal G21825: std_logic; attribute dont_touch of G21825: signal is true;
	signal G21826: std_logic; attribute dont_touch of G21826: signal is true;
	signal G21827: std_logic; attribute dont_touch of G21827: signal is true;
	signal G21828: std_logic; attribute dont_touch of G21828: signal is true;
	signal G21829: std_logic; attribute dont_touch of G21829: signal is true;
	signal G21830: std_logic; attribute dont_touch of G21830: signal is true;
	signal G21831: std_logic; attribute dont_touch of G21831: signal is true;
	signal G21832: std_logic; attribute dont_touch of G21832: signal is true;
	signal G21833: std_logic; attribute dont_touch of G21833: signal is true;
	signal G21834: std_logic; attribute dont_touch of G21834: signal is true;
	signal G21835: std_logic; attribute dont_touch of G21835: signal is true;
	signal G21836: std_logic; attribute dont_touch of G21836: signal is true;
	signal G21837: std_logic; attribute dont_touch of G21837: signal is true;
	signal G21838: std_logic; attribute dont_touch of G21838: signal is true;
	signal G21839: std_logic; attribute dont_touch of G21839: signal is true;
	signal G21840: std_logic; attribute dont_touch of G21840: signal is true;
	signal G21841: std_logic; attribute dont_touch of G21841: signal is true;
	signal G21842: std_logic; attribute dont_touch of G21842: signal is true;
	signal G21843: std_logic; attribute dont_touch of G21843: signal is true;
	signal G21844: std_logic; attribute dont_touch of G21844: signal is true;
	signal G21845: std_logic; attribute dont_touch of G21845: signal is true;
	signal G21846: std_logic; attribute dont_touch of G21846: signal is true;
	signal G21847: std_logic; attribute dont_touch of G21847: signal is true;
	signal G21848: std_logic; attribute dont_touch of G21848: signal is true;
	signal G21849: std_logic; attribute dont_touch of G21849: signal is true;
	signal G21850: std_logic; attribute dont_touch of G21850: signal is true;
	signal G21851: std_logic; attribute dont_touch of G21851: signal is true;
	signal G21852: std_logic; attribute dont_touch of G21852: signal is true;
	signal G21853: std_logic; attribute dont_touch of G21853: signal is true;
	signal G21854: std_logic; attribute dont_touch of G21854: signal is true;
	signal G21855: std_logic; attribute dont_touch of G21855: signal is true;
	signal G21856: std_logic; attribute dont_touch of G21856: signal is true;
	signal G21857: std_logic; attribute dont_touch of G21857: signal is true;
	signal G21858: std_logic; attribute dont_touch of G21858: signal is true;
	signal G21859: std_logic; attribute dont_touch of G21859: signal is true;
	signal G21860: std_logic; attribute dont_touch of G21860: signal is true;
	signal G21861: std_logic; attribute dont_touch of G21861: signal is true;
	signal G21862: std_logic; attribute dont_touch of G21862: signal is true;
	signal G21863: std_logic; attribute dont_touch of G21863: signal is true;
	signal G21864: std_logic; attribute dont_touch of G21864: signal is true;
	signal G21865: std_logic; attribute dont_touch of G21865: signal is true;
	signal G21866: std_logic; attribute dont_touch of G21866: signal is true;
	signal G21867: std_logic; attribute dont_touch of G21867: signal is true;
	signal G21868: std_logic; attribute dont_touch of G21868: signal is true;
	signal G21869: std_logic; attribute dont_touch of G21869: signal is true;
	signal G21870: std_logic; attribute dont_touch of G21870: signal is true;
	signal G21871: std_logic; attribute dont_touch of G21871: signal is true;
	signal G21872: std_logic; attribute dont_touch of G21872: signal is true;
	signal G21873: std_logic; attribute dont_touch of G21873: signal is true;
	signal G21874: std_logic; attribute dont_touch of G21874: signal is true;
	signal G21875: std_logic; attribute dont_touch of G21875: signal is true;
	signal G21876: std_logic; attribute dont_touch of G21876: signal is true;
	signal G21877: std_logic; attribute dont_touch of G21877: signal is true;
	signal G21878: std_logic; attribute dont_touch of G21878: signal is true;
	signal G21879: std_logic; attribute dont_touch of G21879: signal is true;
	signal G21880: std_logic; attribute dont_touch of G21880: signal is true;
	signal G21881: std_logic; attribute dont_touch of G21881: signal is true;
	signal G21882: std_logic; attribute dont_touch of G21882: signal is true;
	signal G21883: std_logic; attribute dont_touch of G21883: signal is true;
	signal G21884: std_logic; attribute dont_touch of G21884: signal is true;
	signal G21885: std_logic; attribute dont_touch of G21885: signal is true;
	signal G21886: std_logic; attribute dont_touch of G21886: signal is true;
	signal G21887: std_logic; attribute dont_touch of G21887: signal is true;
	signal G21888: std_logic; attribute dont_touch of G21888: signal is true;
	signal G21889: std_logic; attribute dont_touch of G21889: signal is true;
	signal G21890: std_logic; attribute dont_touch of G21890: signal is true;
	signal G21891: std_logic; attribute dont_touch of G21891: signal is true;
	signal G21892: std_logic; attribute dont_touch of G21892: signal is true;
	signal G21893: std_logic; attribute dont_touch of G21893: signal is true;
	signal G21894: std_logic; attribute dont_touch of G21894: signal is true;
	signal G21895: std_logic; attribute dont_touch of G21895: signal is true;
	signal G21896: std_logic; attribute dont_touch of G21896: signal is true;
	signal G21897: std_logic; attribute dont_touch of G21897: signal is true;
	signal G21898: std_logic; attribute dont_touch of G21898: signal is true;
	signal G21899: std_logic; attribute dont_touch of G21899: signal is true;
	signal G21900: std_logic; attribute dont_touch of G21900: signal is true;
	signal G21901: std_logic; attribute dont_touch of G21901: signal is true;
	signal G21902: std_logic; attribute dont_touch of G21902: signal is true;
	signal G21903: std_logic; attribute dont_touch of G21903: signal is true;
	signal G21904: std_logic; attribute dont_touch of G21904: signal is true;
	signal G21905: std_logic; attribute dont_touch of G21905: signal is true;
	signal G21906: std_logic; attribute dont_touch of G21906: signal is true;
	signal G21907: std_logic; attribute dont_touch of G21907: signal is true;
	signal G21908: std_logic; attribute dont_touch of G21908: signal is true;
	signal G21909: std_logic; attribute dont_touch of G21909: signal is true;
	signal G21910: std_logic; attribute dont_touch of G21910: signal is true;
	signal G21911: std_logic; attribute dont_touch of G21911: signal is true;
	signal G21912: std_logic; attribute dont_touch of G21912: signal is true;
	signal G21913: std_logic; attribute dont_touch of G21913: signal is true;
	signal G21914: std_logic; attribute dont_touch of G21914: signal is true;
	signal G21915: std_logic; attribute dont_touch of G21915: signal is true;
	signal G21916: std_logic; attribute dont_touch of G21916: signal is true;
	signal G21917: std_logic; attribute dont_touch of G21917: signal is true;
	signal G21918: std_logic; attribute dont_touch of G21918: signal is true;
	signal G21919: std_logic; attribute dont_touch of G21919: signal is true;
	signal G21920: std_logic; attribute dont_touch of G21920: signal is true;
	signal G21921: std_logic; attribute dont_touch of G21921: signal is true;
	signal G21922: std_logic; attribute dont_touch of G21922: signal is true;
	signal G21923: std_logic; attribute dont_touch of G21923: signal is true;
	signal G21924: std_logic; attribute dont_touch of G21924: signal is true;
	signal G21925: std_logic; attribute dont_touch of G21925: signal is true;
	signal G21926: std_logic; attribute dont_touch of G21926: signal is true;
	signal G21927: std_logic; attribute dont_touch of G21927: signal is true;
	signal G21928: std_logic; attribute dont_touch of G21928: signal is true;
	signal G21929: std_logic; attribute dont_touch of G21929: signal is true;
	signal G21930: std_logic; attribute dont_touch of G21930: signal is true;
	signal G21931: std_logic; attribute dont_touch of G21931: signal is true;
	signal G21932: std_logic; attribute dont_touch of G21932: signal is true;
	signal G21933: std_logic; attribute dont_touch of G21933: signal is true;
	signal G21934: std_logic; attribute dont_touch of G21934: signal is true;
	signal G21935: std_logic; attribute dont_touch of G21935: signal is true;
	signal G21936: std_logic; attribute dont_touch of G21936: signal is true;
	signal G21937: std_logic; attribute dont_touch of G21937: signal is true;
	signal G21938: std_logic; attribute dont_touch of G21938: signal is true;
	signal G21939: std_logic; attribute dont_touch of G21939: signal is true;
	signal G21940: std_logic; attribute dont_touch of G21940: signal is true;
	signal G21941: std_logic; attribute dont_touch of G21941: signal is true;
	signal G21942: std_logic; attribute dont_touch of G21942: signal is true;
	signal G21943: std_logic; attribute dont_touch of G21943: signal is true;
	signal G21944: std_logic; attribute dont_touch of G21944: signal is true;
	signal G21945: std_logic; attribute dont_touch of G21945: signal is true;
	signal G21946: std_logic; attribute dont_touch of G21946: signal is true;
	signal G21947: std_logic; attribute dont_touch of G21947: signal is true;
	signal G21948: std_logic; attribute dont_touch of G21948: signal is true;
	signal G21949: std_logic; attribute dont_touch of G21949: signal is true;
	signal G21950: std_logic; attribute dont_touch of G21950: signal is true;
	signal G21951: std_logic; attribute dont_touch of G21951: signal is true;
	signal G21952: std_logic; attribute dont_touch of G21952: signal is true;
	signal G21953: std_logic; attribute dont_touch of G21953: signal is true;
	signal G21954: std_logic; attribute dont_touch of G21954: signal is true;
	signal G21955: std_logic; attribute dont_touch of G21955: signal is true;
	signal G21956: std_logic; attribute dont_touch of G21956: signal is true;
	signal G21957: std_logic; attribute dont_touch of G21957: signal is true;
	signal G21958: std_logic; attribute dont_touch of G21958: signal is true;
	signal G21959: std_logic; attribute dont_touch of G21959: signal is true;
	signal G21960: std_logic; attribute dont_touch of G21960: signal is true;
	signal G21961: std_logic; attribute dont_touch of G21961: signal is true;
	signal G21962: std_logic; attribute dont_touch of G21962: signal is true;
	signal G21963: std_logic; attribute dont_touch of G21963: signal is true;
	signal G21964: std_logic; attribute dont_touch of G21964: signal is true;
	signal G21965: std_logic; attribute dont_touch of G21965: signal is true;
	signal G21966: std_logic; attribute dont_touch of G21966: signal is true;
	signal G21967: std_logic; attribute dont_touch of G21967: signal is true;
	signal G21968: std_logic; attribute dont_touch of G21968: signal is true;
	signal G21969: std_logic; attribute dont_touch of G21969: signal is true;
	signal G21970: std_logic; attribute dont_touch of G21970: signal is true;
	signal G21971: std_logic; attribute dont_touch of G21971: signal is true;
	signal G21972: std_logic; attribute dont_touch of G21972: signal is true;
	signal G21973: std_logic; attribute dont_touch of G21973: signal is true;
	signal G21974: std_logic; attribute dont_touch of G21974: signal is true;
	signal G21975: std_logic; attribute dont_touch of G21975: signal is true;
	signal G21976: std_logic; attribute dont_touch of G21976: signal is true;
	signal G21977: std_logic; attribute dont_touch of G21977: signal is true;
	signal G21978: std_logic; attribute dont_touch of G21978: signal is true;
	signal G21979: std_logic; attribute dont_touch of G21979: signal is true;
	signal G21980: std_logic; attribute dont_touch of G21980: signal is true;
	signal G21981: std_logic; attribute dont_touch of G21981: signal is true;
	signal G21982: std_logic; attribute dont_touch of G21982: signal is true;
	signal G21983: std_logic; attribute dont_touch of G21983: signal is true;
	signal G21984: std_logic; attribute dont_touch of G21984: signal is true;
	signal G21985: std_logic; attribute dont_touch of G21985: signal is true;
	signal G21986: std_logic; attribute dont_touch of G21986: signal is true;
	signal G21987: std_logic; attribute dont_touch of G21987: signal is true;
	signal G21988: std_logic; attribute dont_touch of G21988: signal is true;
	signal G21989: std_logic; attribute dont_touch of G21989: signal is true;
	signal G21990: std_logic; attribute dont_touch of G21990: signal is true;
	signal G21991: std_logic; attribute dont_touch of G21991: signal is true;
	signal G21992: std_logic; attribute dont_touch of G21992: signal is true;
	signal G21993: std_logic; attribute dont_touch of G21993: signal is true;
	signal G21994: std_logic; attribute dont_touch of G21994: signal is true;
	signal G21995: std_logic; attribute dont_touch of G21995: signal is true;
	signal G21996: std_logic; attribute dont_touch of G21996: signal is true;
	signal G21997: std_logic; attribute dont_touch of G21997: signal is true;
	signal G21998: std_logic; attribute dont_touch of G21998: signal is true;
	signal G21999: std_logic; attribute dont_touch of G21999: signal is true;
	signal G22000: std_logic; attribute dont_touch of G22000: signal is true;
	signal G22001: std_logic; attribute dont_touch of G22001: signal is true;
	signal G22002: std_logic; attribute dont_touch of G22002: signal is true;
	signal G22003: std_logic; attribute dont_touch of G22003: signal is true;
	signal G22004: std_logic; attribute dont_touch of G22004: signal is true;
	signal G22005: std_logic; attribute dont_touch of G22005: signal is true;
	signal G22006: std_logic; attribute dont_touch of G22006: signal is true;
	signal G22007: std_logic; attribute dont_touch of G22007: signal is true;
	signal G22008: std_logic; attribute dont_touch of G22008: signal is true;
	signal G22009: std_logic; attribute dont_touch of G22009: signal is true;
	signal G22010: std_logic; attribute dont_touch of G22010: signal is true;
	signal G22011: std_logic; attribute dont_touch of G22011: signal is true;
	signal G22012: std_logic; attribute dont_touch of G22012: signal is true;
	signal G22013: std_logic; attribute dont_touch of G22013: signal is true;
	signal G22014: std_logic; attribute dont_touch of G22014: signal is true;
	signal G22015: std_logic; attribute dont_touch of G22015: signal is true;
	signal G22016: std_logic; attribute dont_touch of G22016: signal is true;
	signal G22017: std_logic; attribute dont_touch of G22017: signal is true;
	signal G22018: std_logic; attribute dont_touch of G22018: signal is true;
	signal G22019: std_logic; attribute dont_touch of G22019: signal is true;
	signal G22020: std_logic; attribute dont_touch of G22020: signal is true;
	signal G22021: std_logic; attribute dont_touch of G22021: signal is true;
	signal G22022: std_logic; attribute dont_touch of G22022: signal is true;
	signal G22023: std_logic; attribute dont_touch of G22023: signal is true;
	signal G22024: std_logic; attribute dont_touch of G22024: signal is true;
	signal G22025: std_logic; attribute dont_touch of G22025: signal is true;
	signal G22026: std_logic; attribute dont_touch of G22026: signal is true;
	signal G22027: std_logic; attribute dont_touch of G22027: signal is true;
	signal G22028: std_logic; attribute dont_touch of G22028: signal is true;
	signal G22029: std_logic; attribute dont_touch of G22029: signal is true;
	signal G22030: std_logic; attribute dont_touch of G22030: signal is true;
	signal G22031: std_logic; attribute dont_touch of G22031: signal is true;
	signal G22032: std_logic; attribute dont_touch of G22032: signal is true;
	signal G22033: std_logic; attribute dont_touch of G22033: signal is true;
	signal G22034: std_logic; attribute dont_touch of G22034: signal is true;
	signal G22035: std_logic; attribute dont_touch of G22035: signal is true;
	signal G22036: std_logic; attribute dont_touch of G22036: signal is true;
	signal G22037: std_logic; attribute dont_touch of G22037: signal is true;
	signal G22038: std_logic; attribute dont_touch of G22038: signal is true;
	signal G22039: std_logic; attribute dont_touch of G22039: signal is true;
	signal G22040: std_logic; attribute dont_touch of G22040: signal is true;
	signal G22041: std_logic; attribute dont_touch of G22041: signal is true;
	signal G22042: std_logic; attribute dont_touch of G22042: signal is true;
	signal G22043: std_logic; attribute dont_touch of G22043: signal is true;
	signal G22044: std_logic; attribute dont_touch of G22044: signal is true;
	signal G22045: std_logic; attribute dont_touch of G22045: signal is true;
	signal G22046: std_logic; attribute dont_touch of G22046: signal is true;
	signal G22047: std_logic; attribute dont_touch of G22047: signal is true;
	signal G22048: std_logic; attribute dont_touch of G22048: signal is true;
	signal G22049: std_logic; attribute dont_touch of G22049: signal is true;
	signal G22050: std_logic; attribute dont_touch of G22050: signal is true;
	signal G22051: std_logic; attribute dont_touch of G22051: signal is true;
	signal G22052: std_logic; attribute dont_touch of G22052: signal is true;
	signal G22053: std_logic; attribute dont_touch of G22053: signal is true;
	signal G22054: std_logic; attribute dont_touch of G22054: signal is true;
	signal G22055: std_logic; attribute dont_touch of G22055: signal is true;
	signal G22056: std_logic; attribute dont_touch of G22056: signal is true;
	signal G22057: std_logic; attribute dont_touch of G22057: signal is true;
	signal G22058: std_logic; attribute dont_touch of G22058: signal is true;
	signal G22059: std_logic; attribute dont_touch of G22059: signal is true;
	signal G22060: std_logic; attribute dont_touch of G22060: signal is true;
	signal G22061: std_logic; attribute dont_touch of G22061: signal is true;
	signal G22062: std_logic; attribute dont_touch of G22062: signal is true;
	signal G22063: std_logic; attribute dont_touch of G22063: signal is true;
	signal G22064: std_logic; attribute dont_touch of G22064: signal is true;
	signal G22065: std_logic; attribute dont_touch of G22065: signal is true;
	signal G22066: std_logic; attribute dont_touch of G22066: signal is true;
	signal G22067: std_logic; attribute dont_touch of G22067: signal is true;
	signal G22068: std_logic; attribute dont_touch of G22068: signal is true;
	signal G22069: std_logic; attribute dont_touch of G22069: signal is true;
	signal G22070: std_logic; attribute dont_touch of G22070: signal is true;
	signal G22071: std_logic; attribute dont_touch of G22071: signal is true;
	signal G22072: std_logic; attribute dont_touch of G22072: signal is true;
	signal G22073: std_logic; attribute dont_touch of G22073: signal is true;
	signal G22074: std_logic; attribute dont_touch of G22074: signal is true;
	signal G22075: std_logic; attribute dont_touch of G22075: signal is true;
	signal G22076: std_logic; attribute dont_touch of G22076: signal is true;
	signal G22077: std_logic; attribute dont_touch of G22077: signal is true;
	signal G22078: std_logic; attribute dont_touch of G22078: signal is true;
	signal G22079: std_logic; attribute dont_touch of G22079: signal is true;
	signal G22080: std_logic; attribute dont_touch of G22080: signal is true;
	signal G22081: std_logic; attribute dont_touch of G22081: signal is true;
	signal G22082: std_logic; attribute dont_touch of G22082: signal is true;
	signal G22083: std_logic; attribute dont_touch of G22083: signal is true;
	signal G22084: std_logic; attribute dont_touch of G22084: signal is true;
	signal G22085: std_logic; attribute dont_touch of G22085: signal is true;
	signal G22086: std_logic; attribute dont_touch of G22086: signal is true;
	signal G22087: std_logic; attribute dont_touch of G22087: signal is true;
	signal G22088: std_logic; attribute dont_touch of G22088: signal is true;
	signal G22089: std_logic; attribute dont_touch of G22089: signal is true;
	signal G22090: std_logic; attribute dont_touch of G22090: signal is true;
	signal G22091: std_logic; attribute dont_touch of G22091: signal is true;
	signal G22092: std_logic; attribute dont_touch of G22092: signal is true;
	signal G22093: std_logic; attribute dont_touch of G22093: signal is true;
	signal G22094: std_logic; attribute dont_touch of G22094: signal is true;
	signal G22095: std_logic; attribute dont_touch of G22095: signal is true;
	signal G22096: std_logic; attribute dont_touch of G22096: signal is true;
	signal G22097: std_logic; attribute dont_touch of G22097: signal is true;
	signal G22098: std_logic; attribute dont_touch of G22098: signal is true;
	signal G22099: std_logic; attribute dont_touch of G22099: signal is true;
	signal G22100: std_logic; attribute dont_touch of G22100: signal is true;
	signal G22101: std_logic; attribute dont_touch of G22101: signal is true;
	signal G22102: std_logic; attribute dont_touch of G22102: signal is true;
	signal G22103: std_logic; attribute dont_touch of G22103: signal is true;
	signal G22104: std_logic; attribute dont_touch of G22104: signal is true;
	signal G22105: std_logic; attribute dont_touch of G22105: signal is true;
	signal G22106: std_logic; attribute dont_touch of G22106: signal is true;
	signal G22107: std_logic; attribute dont_touch of G22107: signal is true;
	signal G22108: std_logic; attribute dont_touch of G22108: signal is true;
	signal G22109: std_logic; attribute dont_touch of G22109: signal is true;
	signal G22110: std_logic; attribute dont_touch of G22110: signal is true;
	signal G22111: std_logic; attribute dont_touch of G22111: signal is true;
	signal G22112: std_logic; attribute dont_touch of G22112: signal is true;
	signal G22113: std_logic; attribute dont_touch of G22113: signal is true;
	signal G22114: std_logic; attribute dont_touch of G22114: signal is true;
	signal G22115: std_logic; attribute dont_touch of G22115: signal is true;
	signal G22116: std_logic; attribute dont_touch of G22116: signal is true;
	signal G22117: std_logic; attribute dont_touch of G22117: signal is true;
	signal G22118: std_logic; attribute dont_touch of G22118: signal is true;
	signal G22119: std_logic; attribute dont_touch of G22119: signal is true;
	signal G22120: std_logic; attribute dont_touch of G22120: signal is true;
	signal G22121: std_logic; attribute dont_touch of G22121: signal is true;
	signal G22122: std_logic; attribute dont_touch of G22122: signal is true;
	signal G22123: std_logic; attribute dont_touch of G22123: signal is true;
	signal G22124: std_logic; attribute dont_touch of G22124: signal is true;
	signal G22125: std_logic; attribute dont_touch of G22125: signal is true;
	signal G22126: std_logic; attribute dont_touch of G22126: signal is true;
	signal G22127: std_logic; attribute dont_touch of G22127: signal is true;
	signal G22128: std_logic; attribute dont_touch of G22128: signal is true;
	signal G22129: std_logic; attribute dont_touch of G22129: signal is true;
	signal G22130: std_logic; attribute dont_touch of G22130: signal is true;
	signal G22131: std_logic; attribute dont_touch of G22131: signal is true;
	signal G22132: std_logic; attribute dont_touch of G22132: signal is true;
	signal G22133: std_logic; attribute dont_touch of G22133: signal is true;
	signal G22134: std_logic; attribute dont_touch of G22134: signal is true;
	signal G22135: std_logic; attribute dont_touch of G22135: signal is true;
	signal G22136: std_logic; attribute dont_touch of G22136: signal is true;
	signal G22137: std_logic; attribute dont_touch of G22137: signal is true;
	signal G22138: std_logic; attribute dont_touch of G22138: signal is true;
	signal G22139: std_logic; attribute dont_touch of G22139: signal is true;
	signal G22142: std_logic; attribute dont_touch of G22142: signal is true;
	signal G22143: std_logic; attribute dont_touch of G22143: signal is true;
	signal G22144: std_logic; attribute dont_touch of G22144: signal is true;
	signal G22145: std_logic; attribute dont_touch of G22145: signal is true;
	signal G22146: std_logic; attribute dont_touch of G22146: signal is true;
	signal G22147: std_logic; attribute dont_touch of G22147: signal is true;
	signal G22148: std_logic; attribute dont_touch of G22148: signal is true;
	signal G22149: std_logic; attribute dont_touch of G22149: signal is true;
	signal G22150: std_logic; attribute dont_touch of G22150: signal is true;
	signal G22151: std_logic; attribute dont_touch of G22151: signal is true;
	signal G22152: std_logic; attribute dont_touch of G22152: signal is true;
	signal G22153: std_logic; attribute dont_touch of G22153: signal is true;
	signal G22154: std_logic; attribute dont_touch of G22154: signal is true;
	signal G22155: std_logic; attribute dont_touch of G22155: signal is true;
	signal G22156: std_logic; attribute dont_touch of G22156: signal is true;
	signal G22157: std_logic; attribute dont_touch of G22157: signal is true;
	signal G22158: std_logic; attribute dont_touch of G22158: signal is true;
	signal G22159: std_logic; attribute dont_touch of G22159: signal is true;
	signal G22160: std_logic; attribute dont_touch of G22160: signal is true;
	signal G22161: std_logic; attribute dont_touch of G22161: signal is true;
	signal G22165: std_logic; attribute dont_touch of G22165: signal is true;
	signal G22166: std_logic; attribute dont_touch of G22166: signal is true;
	signal G22167: std_logic; attribute dont_touch of G22167: signal is true;
	signal G22168: std_logic; attribute dont_touch of G22168: signal is true;
	signal G22169: std_logic; attribute dont_touch of G22169: signal is true;
	signal G22170: std_logic; attribute dont_touch of G22170: signal is true;
	signal G22171: std_logic; attribute dont_touch of G22171: signal is true;
	signal G22172: std_logic; attribute dont_touch of G22172: signal is true;
	signal G22173: std_logic; attribute dont_touch of G22173: signal is true;
	signal G22176: std_logic; attribute dont_touch of G22176: signal is true;
	signal G22177: std_logic; attribute dont_touch of G22177: signal is true;
	signal G22178: std_logic; attribute dont_touch of G22178: signal is true;
	signal G22179: std_logic; attribute dont_touch of G22179: signal is true;
	signal G22180: std_logic; attribute dont_touch of G22180: signal is true;
	signal G22181: std_logic; attribute dont_touch of G22181: signal is true;
	signal G22182: std_logic; attribute dont_touch of G22182: signal is true;
	signal G22189: std_logic; attribute dont_touch of G22189: signal is true;
	signal G22190: std_logic; attribute dont_touch of G22190: signal is true;
	signal G22191: std_logic; attribute dont_touch of G22191: signal is true;
	signal G22192: std_logic; attribute dont_touch of G22192: signal is true;
	signal G22193: std_logic; attribute dont_touch of G22193: signal is true;
	signal G22194: std_logic; attribute dont_touch of G22194: signal is true;
	signal G22197: std_logic; attribute dont_touch of G22197: signal is true;
	signal G22198: std_logic; attribute dont_touch of G22198: signal is true;
	signal G22199: std_logic; attribute dont_touch of G22199: signal is true;
	signal G22200: std_logic; attribute dont_touch of G22200: signal is true;
	signal G22201: std_logic; attribute dont_touch of G22201: signal is true;
	signal G22202: std_logic; attribute dont_touch of G22202: signal is true;
	signal G22207: std_logic; attribute dont_touch of G22207: signal is true;
	signal G22208: std_logic; attribute dont_touch of G22208: signal is true;
	signal G22209: std_logic; attribute dont_touch of G22209: signal is true;
	signal G22210: std_logic; attribute dont_touch of G22210: signal is true;
	signal G22213: std_logic; attribute dont_touch of G22213: signal is true;
	signal G22214: std_logic; attribute dont_touch of G22214: signal is true;
	signal G22215: std_logic; attribute dont_touch of G22215: signal is true;
	signal G22216: std_logic; attribute dont_touch of G22216: signal is true;
	signal G22217: std_logic; attribute dont_touch of G22217: signal is true;
	signal G22218: std_logic; attribute dont_touch of G22218: signal is true;
	signal G22219: std_logic; attribute dont_touch of G22219: signal is true;
	signal G22220: std_logic; attribute dont_touch of G22220: signal is true;
	signal G22223: std_logic; attribute dont_touch of G22223: signal is true;
	signal G22224: std_logic; attribute dont_touch of G22224: signal is true;
	signal G22225: std_logic; attribute dont_touch of G22225: signal is true;
	signal G22226: std_logic; attribute dont_touch of G22226: signal is true;
	signal G22227: std_logic; attribute dont_touch of G22227: signal is true;
	signal G22228: std_logic; attribute dont_touch of G22228: signal is true;
	signal G22298: std_logic; attribute dont_touch of G22298: signal is true;
	signal G22299: std_logic; attribute dont_touch of G22299: signal is true;
	signal G22300: std_logic; attribute dont_touch of G22300: signal is true;
	signal G22303: std_logic; attribute dont_touch of G22303: signal is true;
	signal G22304: std_logic; attribute dont_touch of G22304: signal is true;
	signal G22305: std_logic; attribute dont_touch of G22305: signal is true;
	signal G22306: std_logic; attribute dont_touch of G22306: signal is true;
	signal G22307: std_logic; attribute dont_touch of G22307: signal is true;
	signal G22308: std_logic; attribute dont_touch of G22308: signal is true;
	signal G22309: std_logic; attribute dont_touch of G22309: signal is true;
	signal G22310: std_logic; attribute dont_touch of G22310: signal is true;
	signal G22311: std_logic; attribute dont_touch of G22311: signal is true;
	signal G22312: std_logic; attribute dont_touch of G22312: signal is true;
	signal G22316: std_logic; attribute dont_touch of G22316: signal is true;
	signal G22317: std_logic; attribute dont_touch of G22317: signal is true;
	signal G22318: std_logic; attribute dont_touch of G22318: signal is true;
	signal G22319: std_logic; attribute dont_touch of G22319: signal is true;
	signal G22325: std_logic; attribute dont_touch of G22325: signal is true;
	signal G22329: std_logic; attribute dont_touch of G22329: signal is true;
	signal G22330: std_logic; attribute dont_touch of G22330: signal is true;
	signal G22331: std_logic; attribute dont_touch of G22331: signal is true;
	signal G22332: std_logic; attribute dont_touch of G22332: signal is true;
	signal G22338: std_logic; attribute dont_touch of G22338: signal is true;
	signal G22339: std_logic; attribute dont_touch of G22339: signal is true;
	signal G22340: std_logic; attribute dont_touch of G22340: signal is true;
	signal G22341: std_logic; attribute dont_touch of G22341: signal is true;
	signal G22342: std_logic; attribute dont_touch of G22342: signal is true;
	signal G22357: std_logic; attribute dont_touch of G22357: signal is true;
	signal G22358: std_logic; attribute dont_touch of G22358: signal is true;
	signal G22359: std_logic; attribute dont_touch of G22359: signal is true;
	signal G22360: std_logic; attribute dont_touch of G22360: signal is true;
	signal G22369: std_logic; attribute dont_touch of G22369: signal is true;
	signal G22384: std_logic; attribute dont_touch of G22384: signal is true;
	signal G22399: std_logic; attribute dont_touch of G22399: signal is true;
	signal G22400: std_logic; attribute dont_touch of G22400: signal is true;
	signal G22405: std_logic; attribute dont_touch of G22405: signal is true;
	signal G22406: std_logic; attribute dont_touch of G22406: signal is true;
	signal G22407: std_logic; attribute dont_touch of G22407: signal is true;
	signal G22408: std_logic; attribute dont_touch of G22408: signal is true;
	signal G22409: std_logic; attribute dont_touch of G22409: signal is true;
	signal G22417: std_logic; attribute dont_touch of G22417: signal is true;
	signal G22432: std_logic; attribute dont_touch of G22432: signal is true;
	signal G22447: std_logic; attribute dont_touch of G22447: signal is true;
	signal G22448: std_logic; attribute dont_touch of G22448: signal is true;
	signal G22449: std_logic; attribute dont_touch of G22449: signal is true;
	signal G22450: std_logic; attribute dont_touch of G22450: signal is true;
	signal G22455: std_logic; attribute dont_touch of G22455: signal is true;
	signal G22456: std_logic; attribute dont_touch of G22456: signal is true;
	signal G22457: std_logic; attribute dont_touch of G22457: signal is true;
	signal G22472: std_logic; attribute dont_touch of G22472: signal is true;
	signal G22487: std_logic; attribute dont_touch of G22487: signal is true;
	signal G22488: std_logic; attribute dont_touch of G22488: signal is true;
	signal G22489: std_logic; attribute dont_touch of G22489: signal is true;
	signal G22490: std_logic; attribute dont_touch of G22490: signal is true;
	signal G22491: std_logic; attribute dont_touch of G22491: signal is true;
	signal G22492: std_logic; attribute dont_touch of G22492: signal is true;
	signal G22493: std_logic; attribute dont_touch of G22493: signal is true;
	signal G22494: std_logic; attribute dont_touch of G22494: signal is true;
	signal G22495: std_logic; attribute dont_touch of G22495: signal is true;
	signal G22496: std_logic; attribute dont_touch of G22496: signal is true;
	signal G22497: std_logic; attribute dont_touch of G22497: signal is true;
	signal G22498: std_logic; attribute dont_touch of G22498: signal is true;
	signal G22513: std_logic; attribute dont_touch of G22513: signal is true;
	signal G22514: std_logic; attribute dont_touch of G22514: signal is true;
	signal G22515: std_logic; attribute dont_touch of G22515: signal is true;
	signal G22516: std_logic; attribute dont_touch of G22516: signal is true;
	signal G22517: std_logic; attribute dont_touch of G22517: signal is true;
	signal G22518: std_logic; attribute dont_touch of G22518: signal is true;
	signal G22519: std_logic; attribute dont_touch of G22519: signal is true;
	signal G22520: std_logic; attribute dont_touch of G22520: signal is true;
	signal G22521: std_logic; attribute dont_touch of G22521: signal is true;
	signal G22522: std_logic; attribute dont_touch of G22522: signal is true;
	signal G22523: std_logic; attribute dont_touch of G22523: signal is true;
	signal G22524: std_logic; attribute dont_touch of G22524: signal is true;
	signal G22525: std_logic; attribute dont_touch of G22525: signal is true;
	signal G22526: std_logic; attribute dont_touch of G22526: signal is true;
	signal G22527: std_logic; attribute dont_touch of G22527: signal is true;
	signal G22528: std_logic; attribute dont_touch of G22528: signal is true;
	signal G22529: std_logic; attribute dont_touch of G22529: signal is true;
	signal G22530: std_logic; attribute dont_touch of G22530: signal is true;
	signal G22531: std_logic; attribute dont_touch of G22531: signal is true;
	signal G22534: std_logic; attribute dont_touch of G22534: signal is true;
	signal G22535: std_logic; attribute dont_touch of G22535: signal is true;
	signal G22536: std_logic; attribute dont_touch of G22536: signal is true;
	signal G22537: std_logic; attribute dont_touch of G22537: signal is true;
	signal G22538: std_logic; attribute dont_touch of G22538: signal is true;
	signal G22539: std_logic; attribute dont_touch of G22539: signal is true;
	signal G22540: std_logic; attribute dont_touch of G22540: signal is true;
	signal G22541: std_logic; attribute dont_touch of G22541: signal is true;
	signal G22542: std_logic; attribute dont_touch of G22542: signal is true;
	signal G22543: std_logic; attribute dont_touch of G22543: signal is true;
	signal G22544: std_logic; attribute dont_touch of G22544: signal is true;
	signal G22545: std_logic; attribute dont_touch of G22545: signal is true;
	signal G22546: std_logic; attribute dont_touch of G22546: signal is true;
	signal G22547: std_logic; attribute dont_touch of G22547: signal is true;
	signal G22550: std_logic; attribute dont_touch of G22550: signal is true;
	signal G22585: std_logic; attribute dont_touch of G22585: signal is true;
	signal G22588: std_logic; attribute dont_touch of G22588: signal is true;
	signal G22589: std_logic; attribute dont_touch of G22589: signal is true;
	signal G22590: std_logic; attribute dont_touch of G22590: signal is true;
	signal G22591: std_logic; attribute dont_touch of G22591: signal is true;
	signal G22592: std_logic; attribute dont_touch of G22592: signal is true;
	signal G22593: std_logic; attribute dont_touch of G22593: signal is true;
	signal G22594: std_logic; attribute dont_touch of G22594: signal is true;
	signal G22622: std_logic; attribute dont_touch of G22622: signal is true;
	signal G22623: std_logic; attribute dont_touch of G22623: signal is true;
	signal G22624: std_logic; attribute dont_touch of G22624: signal is true;
	signal G22625: std_logic; attribute dont_touch of G22625: signal is true;
	signal G22626: std_logic; attribute dont_touch of G22626: signal is true;
	signal G22632: std_logic; attribute dont_touch of G22632: signal is true;
	signal G22633: std_logic; attribute dont_touch of G22633: signal is true;
	signal G22634: std_logic; attribute dont_touch of G22634: signal is true;
	signal G22635: std_logic; attribute dont_touch of G22635: signal is true;
	signal G22636: std_logic; attribute dont_touch of G22636: signal is true;
	signal G22637: std_logic; attribute dont_touch of G22637: signal is true;
	signal G22638: std_logic; attribute dont_touch of G22638: signal is true;
	signal G22639: std_logic; attribute dont_touch of G22639: signal is true;
	signal G22640: std_logic; attribute dont_touch of G22640: signal is true;
	signal G22641: std_logic; attribute dont_touch of G22641: signal is true;
	signal G22642: std_logic; attribute dont_touch of G22642: signal is true;
	signal G22643: std_logic; attribute dont_touch of G22643: signal is true;
	signal G22644: std_logic; attribute dont_touch of G22644: signal is true;
	signal G22645: std_logic; attribute dont_touch of G22645: signal is true;
	signal G22646: std_logic; attribute dont_touch of G22646: signal is true;
	signal G22647: std_logic; attribute dont_touch of G22647: signal is true;
	signal G22648: std_logic; attribute dont_touch of G22648: signal is true;
	signal G22649: std_logic; attribute dont_touch of G22649: signal is true;
	signal G22650: std_logic; attribute dont_touch of G22650: signal is true;
	signal G22651: std_logic; attribute dont_touch of G22651: signal is true;
	signal G22652: std_logic; attribute dont_touch of G22652: signal is true;
	signal G22653: std_logic; attribute dont_touch of G22653: signal is true;
	signal G22654: std_logic; attribute dont_touch of G22654: signal is true;
	signal G22658: std_logic; attribute dont_touch of G22658: signal is true;
	signal G22659: std_logic; attribute dont_touch of G22659: signal is true;
	signal G22660: std_logic; attribute dont_touch of G22660: signal is true;
	signal G22661: std_logic; attribute dont_touch of G22661: signal is true;
	signal G22662: std_logic; attribute dont_touch of G22662: signal is true;
	signal G22663: std_logic; attribute dont_touch of G22663: signal is true;
	signal G22664: std_logic; attribute dont_touch of G22664: signal is true;
	signal G22665: std_logic; attribute dont_touch of G22665: signal is true;
	signal G22666: std_logic; attribute dont_touch of G22666: signal is true;
	signal G22667: std_logic; attribute dont_touch of G22667: signal is true;
	signal G22668: std_logic; attribute dont_touch of G22668: signal is true;
	signal G22669: std_logic; attribute dont_touch of G22669: signal is true;
	signal G22670: std_logic; attribute dont_touch of G22670: signal is true;
	signal G22679: std_logic; attribute dont_touch of G22679: signal is true;
	signal G22680: std_logic; attribute dont_touch of G22680: signal is true;
	signal G22681: std_logic; attribute dont_touch of G22681: signal is true;
	signal G22682: std_logic; attribute dont_touch of G22682: signal is true;
	signal G22683: std_logic; attribute dont_touch of G22683: signal is true;
	signal G22684: std_logic; attribute dont_touch of G22684: signal is true;
	signal G22685: std_logic; attribute dont_touch of G22685: signal is true;
	signal G22686: std_logic; attribute dont_touch of G22686: signal is true;
	signal G22687: std_logic; attribute dont_touch of G22687: signal is true;
	signal G22688: std_logic; attribute dont_touch of G22688: signal is true;
	signal G22689: std_logic; attribute dont_touch of G22689: signal is true;
	signal G22698: std_logic; attribute dont_touch of G22698: signal is true;
	signal G22707: std_logic; attribute dont_touch of G22707: signal is true;
	signal G22708: std_logic; attribute dont_touch of G22708: signal is true;
	signal G22709: std_logic; attribute dont_touch of G22709: signal is true;
	signal G22710: std_logic; attribute dont_touch of G22710: signal is true;
	signal G22711: std_logic; attribute dont_touch of G22711: signal is true;
	signal G22712: std_logic; attribute dont_touch of G22712: signal is true;
	signal G22713: std_logic; attribute dont_touch of G22713: signal is true;
	signal G22714: std_logic; attribute dont_touch of G22714: signal is true;
	signal G22715: std_logic; attribute dont_touch of G22715: signal is true;
	signal G22716: std_logic; attribute dont_touch of G22716: signal is true;
	signal G22717: std_logic; attribute dont_touch of G22717: signal is true;
	signal G22718: std_logic; attribute dont_touch of G22718: signal is true;
	signal G22719: std_logic; attribute dont_touch of G22719: signal is true;
	signal G22720: std_logic; attribute dont_touch of G22720: signal is true;
	signal G22721: std_logic; attribute dont_touch of G22721: signal is true;
	signal G22722: std_logic; attribute dont_touch of G22722: signal is true;
	signal G22751: std_logic; attribute dont_touch of G22751: signal is true;
	signal G22752: std_logic; attribute dont_touch of G22752: signal is true;
	signal G22753: std_logic; attribute dont_touch of G22753: signal is true;
	signal G22754: std_logic; attribute dont_touch of G22754: signal is true;
	signal G22755: std_logic; attribute dont_touch of G22755: signal is true;
	signal G22756: std_logic; attribute dont_touch of G22756: signal is true;
	signal G22757: std_logic; attribute dont_touch of G22757: signal is true;
	signal G22758: std_logic; attribute dont_touch of G22758: signal is true;
	signal G22759: std_logic; attribute dont_touch of G22759: signal is true;
	signal G22760: std_logic; attribute dont_touch of G22760: signal is true;
	signal G22761: std_logic; attribute dont_touch of G22761: signal is true;
	signal G22762: std_logic; attribute dont_touch of G22762: signal is true;
	signal G22763: std_logic; attribute dont_touch of G22763: signal is true;
	signal G22830: std_logic; attribute dont_touch of G22830: signal is true;
	signal G22831: std_logic; attribute dont_touch of G22831: signal is true;
	signal G22832: std_logic; attribute dont_touch of G22832: signal is true;
	signal G22833: std_logic; attribute dont_touch of G22833: signal is true;
	signal G22834: std_logic; attribute dont_touch of G22834: signal is true;
	signal G22835: std_logic; attribute dont_touch of G22835: signal is true;
	signal G22836: std_logic; attribute dont_touch of G22836: signal is true;
	signal G22837: std_logic; attribute dont_touch of G22837: signal is true;
	signal G22838: std_logic; attribute dont_touch of G22838: signal is true;
	signal G22839: std_logic; attribute dont_touch of G22839: signal is true;
	signal G22840: std_logic; attribute dont_touch of G22840: signal is true;
	signal G22841: std_logic; attribute dont_touch of G22841: signal is true;
	signal G22842: std_logic; attribute dont_touch of G22842: signal is true;
	signal G22843: std_logic; attribute dont_touch of G22843: signal is true;
	signal G22844: std_logic; attribute dont_touch of G22844: signal is true;
	signal G22845: std_logic; attribute dont_touch of G22845: signal is true;
	signal G22846: std_logic; attribute dont_touch of G22846: signal is true;
	signal G22847: std_logic; attribute dont_touch of G22847: signal is true;
	signal G22848: std_logic; attribute dont_touch of G22848: signal is true;
	signal G22849: std_logic; attribute dont_touch of G22849: signal is true;
	signal G22850: std_logic; attribute dont_touch of G22850: signal is true;
	signal G22851: std_logic; attribute dont_touch of G22851: signal is true;
	signal G22852: std_logic; attribute dont_touch of G22852: signal is true;
	signal G22853: std_logic; attribute dont_touch of G22853: signal is true;
	signal G22854: std_logic; attribute dont_touch of G22854: signal is true;
	signal G22855: std_logic; attribute dont_touch of G22855: signal is true;
	signal G22856: std_logic; attribute dont_touch of G22856: signal is true;
	signal G22857: std_logic; attribute dont_touch of G22857: signal is true;
	signal G22858: std_logic; attribute dont_touch of G22858: signal is true;
	signal G22859: std_logic; attribute dont_touch of G22859: signal is true;
	signal G22860: std_logic; attribute dont_touch of G22860: signal is true;
	signal G22861: std_logic; attribute dont_touch of G22861: signal is true;
	signal G22862: std_logic; attribute dont_touch of G22862: signal is true;
	signal G22863: std_logic; attribute dont_touch of G22863: signal is true;
	signal G22864: std_logic; attribute dont_touch of G22864: signal is true;
	signal G22865: std_logic; attribute dont_touch of G22865: signal is true;
	signal G22866: std_logic; attribute dont_touch of G22866: signal is true;
	signal G22867: std_logic; attribute dont_touch of G22867: signal is true;
	signal G22868: std_logic; attribute dont_touch of G22868: signal is true;
	signal G22869: std_logic; attribute dont_touch of G22869: signal is true;
	signal G22870: std_logic; attribute dont_touch of G22870: signal is true;
	signal G22871: std_logic; attribute dont_touch of G22871: signal is true;
	signal G22872: std_logic; attribute dont_touch of G22872: signal is true;
	signal G22873: std_logic; attribute dont_touch of G22873: signal is true;
	signal G22874: std_logic; attribute dont_touch of G22874: signal is true;
	signal G22875: std_logic; attribute dont_touch of G22875: signal is true;
	signal G22876: std_logic; attribute dont_touch of G22876: signal is true;
	signal G22881: std_logic; attribute dont_touch of G22881: signal is true;
	signal G22882: std_logic; attribute dont_touch of G22882: signal is true;
	signal G22883: std_logic; attribute dont_touch of G22883: signal is true;
	signal G22884: std_logic; attribute dont_touch of G22884: signal is true;
	signal G22885: std_logic; attribute dont_touch of G22885: signal is true;
	signal G22896: std_logic; attribute dont_touch of G22896: signal is true;
	signal G22897: std_logic; attribute dont_touch of G22897: signal is true;
	signal G22898: std_logic; attribute dont_touch of G22898: signal is true;
	signal G22899: std_logic; attribute dont_touch of G22899: signal is true;
	signal G22900: std_logic; attribute dont_touch of G22900: signal is true;
	signal G22901: std_logic; attribute dont_touch of G22901: signal is true;
	signal G22902: std_logic; attribute dont_touch of G22902: signal is true;
	signal G22903: std_logic; attribute dont_touch of G22903: signal is true;
	signal G22904: std_logic; attribute dont_touch of G22904: signal is true;
	signal G22905: std_logic; attribute dont_touch of G22905: signal is true;
	signal G22906: std_logic; attribute dont_touch of G22906: signal is true;
	signal G22907: std_logic; attribute dont_touch of G22907: signal is true;
	signal G22908: std_logic; attribute dont_touch of G22908: signal is true;
	signal G22919: std_logic; attribute dont_touch of G22919: signal is true;
	signal G22920: std_logic; attribute dont_touch of G22920: signal is true;
	signal G22921: std_logic; attribute dont_touch of G22921: signal is true;
	signal G22922: std_logic; attribute dont_touch of G22922: signal is true;
	signal G22923: std_logic; attribute dont_touch of G22923: signal is true;
	signal G22926: std_logic; attribute dont_touch of G22926: signal is true;
	signal G22927: std_logic; attribute dont_touch of G22927: signal is true;
	signal G22928: std_logic; attribute dont_touch of G22928: signal is true;
	signal G22929: std_logic; attribute dont_touch of G22929: signal is true;
	signal G22935: std_logic; attribute dont_touch of G22935: signal is true;
	signal G22936: std_logic; attribute dont_touch of G22936: signal is true;
	signal G22937: std_logic; attribute dont_touch of G22937: signal is true;
	signal G22938: std_logic; attribute dont_touch of G22938: signal is true;
	signal G22939: std_logic; attribute dont_touch of G22939: signal is true;
	signal G22940: std_logic; attribute dont_touch of G22940: signal is true;
	signal G22941: std_logic; attribute dont_touch of G22941: signal is true;
	signal G22942: std_logic; attribute dont_touch of G22942: signal is true;
	signal G22957: std_logic; attribute dont_touch of G22957: signal is true;
	signal G22973: std_logic; attribute dont_touch of G22973: signal is true;
	signal G22974: std_logic; attribute dont_touch of G22974: signal is true;
	signal G22975: std_logic; attribute dont_touch of G22975: signal is true;
	signal G22976: std_logic; attribute dont_touch of G22976: signal is true;
	signal G22979: std_logic; attribute dont_touch of G22979: signal is true;
	signal G22980: std_logic; attribute dont_touch of G22980: signal is true;
	signal G22981: std_logic; attribute dont_touch of G22981: signal is true;
	signal G22982: std_logic; attribute dont_touch of G22982: signal is true;
	signal G22983: std_logic; attribute dont_touch of G22983: signal is true;
	signal G22984: std_logic; attribute dont_touch of G22984: signal is true;
	signal G22985: std_logic; attribute dont_touch of G22985: signal is true;
	signal G22986: std_logic; attribute dont_touch of G22986: signal is true;
	signal G22987: std_logic; attribute dont_touch of G22987: signal is true;
	signal G22988: std_logic; attribute dont_touch of G22988: signal is true;
	signal G22989: std_logic; attribute dont_touch of G22989: signal is true;
	signal G22990: std_logic; attribute dont_touch of G22990: signal is true;
	signal G22991: std_logic; attribute dont_touch of G22991: signal is true;
	signal G22992: std_logic; attribute dont_touch of G22992: signal is true;
	signal G22993: std_logic; attribute dont_touch of G22993: signal is true;
	signal G22994: std_logic; attribute dont_touch of G22994: signal is true;
	signal G22995: std_logic; attribute dont_touch of G22995: signal is true;
	signal G22996: std_logic; attribute dont_touch of G22996: signal is true;
	signal G22997: std_logic; attribute dont_touch of G22997: signal is true;
	signal G22998: std_logic; attribute dont_touch of G22998: signal is true;
	signal G22999: std_logic; attribute dont_touch of G22999: signal is true;
	signal G23000: std_logic; attribute dont_touch of G23000: signal is true;
	signal G23001: std_logic; attribute dont_touch of G23001: signal is true;
	signal G23003: std_logic; attribute dont_touch of G23003: signal is true;
	signal G23004: std_logic; attribute dont_touch of G23004: signal is true;
	signal G23005: std_logic; attribute dont_touch of G23005: signal is true;
	signal G23006: std_logic; attribute dont_touch of G23006: signal is true;
	signal G23007: std_logic; attribute dont_touch of G23007: signal is true;
	signal G23008: std_logic; attribute dont_touch of G23008: signal is true;
	signal G23009: std_logic; attribute dont_touch of G23009: signal is true;
	signal G23010: std_logic; attribute dont_touch of G23010: signal is true;
	signal G23011: std_logic; attribute dont_touch of G23011: signal is true;
	signal G23012: std_logic; attribute dont_touch of G23012: signal is true;
	signal G23013: std_logic; attribute dont_touch of G23013: signal is true;
	signal G23014: std_logic; attribute dont_touch of G23014: signal is true;
	signal G23015: std_logic; attribute dont_touch of G23015: signal is true;
	signal G23016: std_logic; attribute dont_touch of G23016: signal is true;
	signal G23017: std_logic; attribute dont_touch of G23017: signal is true;
	signal G23018: std_logic; attribute dont_touch of G23018: signal is true;
	signal G23019: std_logic; attribute dont_touch of G23019: signal is true;
	signal G23020: std_logic; attribute dont_touch of G23020: signal is true;
	signal G23021: std_logic; attribute dont_touch of G23021: signal is true;
	signal G23022: std_logic; attribute dont_touch of G23022: signal is true;
	signal G23023: std_logic; attribute dont_touch of G23023: signal is true;
	signal G23024: std_logic; attribute dont_touch of G23024: signal is true;
	signal G23025: std_logic; attribute dont_touch of G23025: signal is true;
	signal G23026: std_logic; attribute dont_touch of G23026: signal is true;
	signal G23027: std_logic; attribute dont_touch of G23027: signal is true;
	signal G23028: std_logic; attribute dont_touch of G23028: signal is true;
	signal G23029: std_logic; attribute dont_touch of G23029: signal is true;
	signal G23030: std_logic; attribute dont_touch of G23030: signal is true;
	signal G23031: std_logic; attribute dont_touch of G23031: signal is true;
	signal G23032: std_logic; attribute dont_touch of G23032: signal is true;
	signal G23041: std_logic; attribute dont_touch of G23041: signal is true;
	signal G23042: std_logic; attribute dont_touch of G23042: signal is true;
	signal G23046: std_logic; attribute dont_touch of G23046: signal is true;
	signal G23047: std_logic; attribute dont_touch of G23047: signal is true;
	signal G23050: std_logic; attribute dont_touch of G23050: signal is true;
	signal G23051: std_logic; attribute dont_touch of G23051: signal is true;
	signal G23052: std_logic; attribute dont_touch of G23052: signal is true;
	signal G23055: std_logic; attribute dont_touch of G23055: signal is true;
	signal G23056: std_logic; attribute dont_touch of G23056: signal is true;
	signal G23057: std_logic; attribute dont_touch of G23057: signal is true;
	signal G23058: std_logic; attribute dont_touch of G23058: signal is true;
	signal G23059: std_logic; attribute dont_touch of G23059: signal is true;
	signal G23060: std_logic; attribute dont_touch of G23060: signal is true;
	signal G23061: std_logic; attribute dont_touch of G23061: signal is true;
	signal G23062: std_logic; attribute dont_touch of G23062: signal is true;
	signal G23063: std_logic; attribute dont_touch of G23063: signal is true;
	signal G23066: std_logic; attribute dont_touch of G23066: signal is true;
	signal G23067: std_logic; attribute dont_touch of G23067: signal is true;
	signal G23076: std_logic; attribute dont_touch of G23076: signal is true;
	signal G23079: std_logic; attribute dont_touch of G23079: signal is true;
	signal G23082: std_logic; attribute dont_touch of G23082: signal is true;
	signal G23083: std_logic; attribute dont_touch of G23083: signal is true;
	signal G23084: std_logic; attribute dont_touch of G23084: signal is true;
	signal G23085: std_logic; attribute dont_touch of G23085: signal is true;
	signal G23086: std_logic; attribute dont_touch of G23086: signal is true;
	signal G23087: std_logic; attribute dont_touch of G23087: signal is true;
	signal G23088: std_logic; attribute dont_touch of G23088: signal is true;
	signal G23103: std_logic; attribute dont_touch of G23103: signal is true;
	signal G23104: std_logic; attribute dont_touch of G23104: signal is true;
	signal G23105: std_logic; attribute dont_touch of G23105: signal is true;
	signal G23108: std_logic; attribute dont_touch of G23108: signal is true;
	signal G23111: std_logic; attribute dont_touch of G23111: signal is true;
	signal G23112: std_logic; attribute dont_touch of G23112: signal is true;
	signal G23121: std_logic; attribute dont_touch of G23121: signal is true;
	signal G23124: std_logic; attribute dont_touch of G23124: signal is true;
	signal G23127: std_logic; attribute dont_touch of G23127: signal is true;
	signal G23128: std_logic; attribute dont_touch of G23128: signal is true;
	signal G23129: std_logic; attribute dont_touch of G23129: signal is true;
	signal G23130: std_logic; attribute dont_touch of G23130: signal is true;
	signal G23131: std_logic; attribute dont_touch of G23131: signal is true;
	signal G23132: std_logic; attribute dont_touch of G23132: signal is true;
	signal G23135: std_logic; attribute dont_touch of G23135: signal is true;
	signal G23138: std_logic; attribute dont_touch of G23138: signal is true;
	signal G23139: std_logic; attribute dont_touch of G23139: signal is true;
	signal G23148: std_logic; attribute dont_touch of G23148: signal is true;
	signal G23151: std_logic; attribute dont_touch of G23151: signal is true;
	signal G23152: std_logic; attribute dont_touch of G23152: signal is true;
	signal G23153: std_logic; attribute dont_touch of G23153: signal is true;
	signal G23154: std_logic; attribute dont_touch of G23154: signal is true;
	signal G23162: std_logic; attribute dont_touch of G23162: signal is true;
	signal G23165: std_logic; attribute dont_touch of G23165: signal is true;
	signal G23166: std_logic; attribute dont_touch of G23166: signal is true;
	signal G23167: std_logic; attribute dont_touch of G23167: signal is true;
	signal G23170: std_logic; attribute dont_touch of G23170: signal is true;
	signal G23171: std_logic; attribute dont_touch of G23171: signal is true;
	signal G23172: std_logic; attribute dont_touch of G23172: signal is true;
	signal G23182: std_logic; attribute dont_touch of G23182: signal is true;
	signal G23183: std_logic; attribute dont_touch of G23183: signal is true;
	signal G23184: std_logic; attribute dont_touch of G23184: signal is true;
	signal G23187: std_logic; attribute dont_touch of G23187: signal is true;
	signal G23188: std_logic; attribute dont_touch of G23188: signal is true;
	signal G23189: std_logic; attribute dont_touch of G23189: signal is true;
	signal G23191: std_logic; attribute dont_touch of G23191: signal is true;
	signal G23192: std_logic; attribute dont_touch of G23192: signal is true;
	signal G23193: std_logic; attribute dont_touch of G23193: signal is true;
	signal G23194: std_logic; attribute dont_touch of G23194: signal is true;
	signal G23195: std_logic; attribute dont_touch of G23195: signal is true;
	signal G23196: std_logic; attribute dont_touch of G23196: signal is true;
	signal G23197: std_logic; attribute dont_touch of G23197: signal is true;
	signal G23198: std_logic; attribute dont_touch of G23198: signal is true;
	signal G23201: std_logic; attribute dont_touch of G23201: signal is true;
	signal G23202: std_logic; attribute dont_touch of G23202: signal is true;
	signal G23203: std_logic; attribute dont_touch of G23203: signal is true;
	signal G23204: std_logic; attribute dont_touch of G23204: signal is true;
	signal G23208: std_logic; attribute dont_touch of G23208: signal is true;
	signal G23209: std_logic; attribute dont_touch of G23209: signal is true;
	signal G23210: std_logic; attribute dont_touch of G23210: signal is true;
	signal G23211: std_logic; attribute dont_touch of G23211: signal is true;
	signal G23214: std_logic; attribute dont_touch of G23214: signal is true;
	signal G23215: std_logic; attribute dont_touch of G23215: signal is true;
	signal G23216: std_logic; attribute dont_touch of G23216: signal is true;
	signal G23217: std_logic; attribute dont_touch of G23217: signal is true;
	signal G23218: std_logic; attribute dont_touch of G23218: signal is true;
	signal G23219: std_logic; attribute dont_touch of G23219: signal is true;
	signal G23220: std_logic; attribute dont_touch of G23220: signal is true;
	signal G23221: std_logic; attribute dont_touch of G23221: signal is true;
	signal G23222: std_logic; attribute dont_touch of G23222: signal is true;
	signal G23223: std_logic; attribute dont_touch of G23223: signal is true;
	signal G23226: std_logic; attribute dont_touch of G23226: signal is true;
	signal G23227: std_logic; attribute dont_touch of G23227: signal is true;
	signal G23228: std_logic; attribute dont_touch of G23228: signal is true;
	signal G23229: std_logic; attribute dont_touch of G23229: signal is true;
	signal G23230: std_logic; attribute dont_touch of G23230: signal is true;
	signal G23231: std_logic; attribute dont_touch of G23231: signal is true;
	signal G23232: std_logic; attribute dont_touch of G23232: signal is true;
	signal G23233: std_logic; attribute dont_touch of G23233: signal is true;
	signal G23234: std_logic; attribute dont_touch of G23234: signal is true;
	signal G23235: std_logic; attribute dont_touch of G23235: signal is true;
	signal G23236: std_logic; attribute dont_touch of G23236: signal is true;
	signal G23237: std_logic; attribute dont_touch of G23237: signal is true;
	signal G23238: std_logic; attribute dont_touch of G23238: signal is true;
	signal G23239: std_logic; attribute dont_touch of G23239: signal is true;
	signal G23242: std_logic; attribute dont_touch of G23242: signal is true;
	signal G23243: std_logic; attribute dont_touch of G23243: signal is true;
	signal G23244: std_logic; attribute dont_touch of G23244: signal is true;
	signal G23245: std_logic; attribute dont_touch of G23245: signal is true;
	signal G23246: std_logic; attribute dont_touch of G23246: signal is true;
	signal G23247: std_logic; attribute dont_touch of G23247: signal is true;
	signal G23248: std_logic; attribute dont_touch of G23248: signal is true;
	signal G23249: std_logic; attribute dont_touch of G23249: signal is true;
	signal G23250: std_logic; attribute dont_touch of G23250: signal is true;
	signal G23251: std_logic; attribute dont_touch of G23251: signal is true;
	signal G23252: std_logic; attribute dont_touch of G23252: signal is true;
	signal G23253: std_logic; attribute dont_touch of G23253: signal is true;
	signal G23254: std_logic; attribute dont_touch of G23254: signal is true;
	signal G23255: std_logic; attribute dont_touch of G23255: signal is true;
	signal G23256: std_logic; attribute dont_touch of G23256: signal is true;
	signal G23257: std_logic; attribute dont_touch of G23257: signal is true;
	signal G23258: std_logic; attribute dont_touch of G23258: signal is true;
	signal G23259: std_logic; attribute dont_touch of G23259: signal is true;
	signal G23260: std_logic; attribute dont_touch of G23260: signal is true;
	signal G23261: std_logic; attribute dont_touch of G23261: signal is true;
	signal G23262: std_logic; attribute dont_touch of G23262: signal is true;
	signal G23263: std_logic; attribute dont_touch of G23263: signal is true;
	signal G23264: std_logic; attribute dont_touch of G23264: signal is true;
	signal G23265: std_logic; attribute dont_touch of G23265: signal is true;
	signal G23266: std_logic; attribute dont_touch of G23266: signal is true;
	signal G23267: std_logic; attribute dont_touch of G23267: signal is true;
	signal G23270: std_logic; attribute dont_touch of G23270: signal is true;
	signal G23271: std_logic; attribute dont_touch of G23271: signal is true;
	signal G23272: std_logic; attribute dont_touch of G23272: signal is true;
	signal G23273: std_logic; attribute dont_touch of G23273: signal is true;
	signal G23274: std_logic; attribute dont_touch of G23274: signal is true;
	signal G23275: std_logic; attribute dont_touch of G23275: signal is true;
	signal G23276: std_logic; attribute dont_touch of G23276: signal is true;
	signal G23277: std_logic; attribute dont_touch of G23277: signal is true;
	signal G23278: std_logic; attribute dont_touch of G23278: signal is true;
	signal G23279: std_logic; attribute dont_touch of G23279: signal is true;
	signal G23280: std_logic; attribute dont_touch of G23280: signal is true;
	signal G23281: std_logic; attribute dont_touch of G23281: signal is true;
	signal G23282: std_logic; attribute dont_touch of G23282: signal is true;
	signal G23283: std_logic; attribute dont_touch of G23283: signal is true;
	signal G23284: std_logic; attribute dont_touch of G23284: signal is true;
	signal G23285: std_logic; attribute dont_touch of G23285: signal is true;
	signal G23286: std_logic; attribute dont_touch of G23286: signal is true;
	signal G23289: std_logic; attribute dont_touch of G23289: signal is true;
	signal G23290: std_logic; attribute dont_touch of G23290: signal is true;
	signal G23291: std_logic; attribute dont_touch of G23291: signal is true;
	signal G23292: std_logic; attribute dont_touch of G23292: signal is true;
	signal G23293: std_logic; attribute dont_touch of G23293: signal is true;
	signal G23296: std_logic; attribute dont_touch of G23296: signal is true;
	signal G23297: std_logic; attribute dont_touch of G23297: signal is true;
	signal G23298: std_logic; attribute dont_touch of G23298: signal is true;
	signal G23299: std_logic; attribute dont_touch of G23299: signal is true;
	signal G23300: std_logic; attribute dont_touch of G23300: signal is true;
	signal G23301: std_logic; attribute dont_touch of G23301: signal is true;
	signal G23302: std_logic; attribute dont_touch of G23302: signal is true;
	signal G23303: std_logic; attribute dont_touch of G23303: signal is true;
	signal G23304: std_logic; attribute dont_touch of G23304: signal is true;
	signal G23305: std_logic; attribute dont_touch of G23305: signal is true;
	signal G23306: std_logic; attribute dont_touch of G23306: signal is true;
	signal G23307: std_logic; attribute dont_touch of G23307: signal is true;
	signal G23308: std_logic; attribute dont_touch of G23308: signal is true;
	signal G23309: std_logic; attribute dont_touch of G23309: signal is true;
	signal G23312: std_logic; attribute dont_touch of G23312: signal is true;
	signal G23313: std_logic; attribute dont_touch of G23313: signal is true;
	signal G23314: std_logic; attribute dont_touch of G23314: signal is true;
	signal G23317: std_logic; attribute dont_touch of G23317: signal is true;
	signal G23318: std_logic; attribute dont_touch of G23318: signal is true;
	signal G23319: std_logic; attribute dont_touch of G23319: signal is true;
	signal G23320: std_logic; attribute dont_touch of G23320: signal is true;
	signal G23321: std_logic; attribute dont_touch of G23321: signal is true;
	signal G23322: std_logic; attribute dont_touch of G23322: signal is true;
	signal G23323: std_logic; attribute dont_touch of G23323: signal is true;
	signal G23324: std_logic; attribute dont_touch of G23324: signal is true;
	signal G23331: std_logic; attribute dont_touch of G23331: signal is true;
	signal G23332: std_logic; attribute dont_touch of G23332: signal is true;
	signal G23333: std_logic; attribute dont_touch of G23333: signal is true;
	signal G23334: std_logic; attribute dont_touch of G23334: signal is true;
	signal G23335: std_logic; attribute dont_touch of G23335: signal is true;
	signal G23336: std_logic; attribute dont_touch of G23336: signal is true;
	signal G23337: std_logic; attribute dont_touch of G23337: signal is true;
	signal G23338: std_logic; attribute dont_touch of G23338: signal is true;
	signal G23339: std_logic; attribute dont_touch of G23339: signal is true;
	signal G23340: std_logic; attribute dont_touch of G23340: signal is true;
	signal G23341: std_logic; attribute dont_touch of G23341: signal is true;
	signal G23342: std_logic; attribute dont_touch of G23342: signal is true;
	signal G23345: std_logic; attribute dont_touch of G23345: signal is true;
	signal G23346: std_logic; attribute dont_touch of G23346: signal is true;
	signal G23347: std_logic; attribute dont_touch of G23347: signal is true;
	signal G23348: std_logic; attribute dont_touch of G23348: signal is true;
	signal G23349: std_logic; attribute dont_touch of G23349: signal is true;
	signal G23350: std_logic; attribute dont_touch of G23350: signal is true;
	signal G23351: std_logic; attribute dont_touch of G23351: signal is true;
	signal G23352: std_logic; attribute dont_touch of G23352: signal is true;
	signal G23353: std_logic; attribute dont_touch of G23353: signal is true;
	signal G23354: std_logic; attribute dont_touch of G23354: signal is true;
	signal G23355: std_logic; attribute dont_touch of G23355: signal is true;
	signal G23356: std_logic; attribute dont_touch of G23356: signal is true;
	signal G23357: std_logic; attribute dont_touch of G23357: signal is true;
	signal G23358: std_logic; attribute dont_touch of G23358: signal is true;
	signal G23359: std_logic; attribute dont_touch of G23359: signal is true;
	signal G23360: std_logic; attribute dont_touch of G23360: signal is true;
	signal G23361: std_logic; attribute dont_touch of G23361: signal is true;
	signal G23362: std_logic; attribute dont_touch of G23362: signal is true;
	signal G23363: std_logic; attribute dont_touch of G23363: signal is true;
	signal G23372: std_logic; attribute dont_touch of G23372: signal is true;
	signal G23373: std_logic; attribute dont_touch of G23373: signal is true;
	signal G23374: std_logic; attribute dont_touch of G23374: signal is true;
	signal G23375: std_logic; attribute dont_touch of G23375: signal is true;
	signal G23376: std_logic; attribute dont_touch of G23376: signal is true;
	signal G23377: std_logic; attribute dont_touch of G23377: signal is true;
	signal G23378: std_logic; attribute dont_touch of G23378: signal is true;
	signal G23379: std_logic; attribute dont_touch of G23379: signal is true;
	signal G23380: std_logic; attribute dont_touch of G23380: signal is true;
	signal G23381: std_logic; attribute dont_touch of G23381: signal is true;
	signal G23382: std_logic; attribute dont_touch of G23382: signal is true;
	signal G23383: std_logic; attribute dont_touch of G23383: signal is true;
	signal G23384: std_logic; attribute dont_touch of G23384: signal is true;
	signal G23385: std_logic; attribute dont_touch of G23385: signal is true;
	signal G23386: std_logic; attribute dont_touch of G23386: signal is true;
	signal G23387: std_logic; attribute dont_touch of G23387: signal is true;
	signal G23388: std_logic; attribute dont_touch of G23388: signal is true;
	signal G23389: std_logic; attribute dont_touch of G23389: signal is true;
	signal G23390: std_logic; attribute dont_touch of G23390: signal is true;
	signal G23391: std_logic; attribute dont_touch of G23391: signal is true;
	signal G23392: std_logic; attribute dont_touch of G23392: signal is true;
	signal G23393: std_logic; attribute dont_touch of G23393: signal is true;
	signal G23394: std_logic; attribute dont_touch of G23394: signal is true;
	signal G23395: std_logic; attribute dont_touch of G23395: signal is true;
	signal G23396: std_logic; attribute dont_touch of G23396: signal is true;
	signal G23397: std_logic; attribute dont_touch of G23397: signal is true;
	signal G23398: std_logic; attribute dont_touch of G23398: signal is true;
	signal G23399: std_logic; attribute dont_touch of G23399: signal is true;
	signal G23400: std_logic; attribute dont_touch of G23400: signal is true;
	signal G23401: std_logic; attribute dont_touch of G23401: signal is true;
	signal G23402: std_logic; attribute dont_touch of G23402: signal is true;
	signal G23403: std_logic; attribute dont_touch of G23403: signal is true;
	signal G23404: std_logic; attribute dont_touch of G23404: signal is true;
	signal G23405: std_logic; attribute dont_touch of G23405: signal is true;
	signal G23406: std_logic; attribute dont_touch of G23406: signal is true;
	signal G23407: std_logic; attribute dont_touch of G23407: signal is true;
	signal G23408: std_logic; attribute dont_touch of G23408: signal is true;
	signal G23409: std_logic; attribute dont_touch of G23409: signal is true;
	signal G23410: std_logic; attribute dont_touch of G23410: signal is true;
	signal G23411: std_logic; attribute dont_touch of G23411: signal is true;
	signal G23412: std_logic; attribute dont_touch of G23412: signal is true;
	signal G23413: std_logic; attribute dont_touch of G23413: signal is true;
	signal G23414: std_logic; attribute dont_touch of G23414: signal is true;
	signal G23415: std_logic; attribute dont_touch of G23415: signal is true;
	signal G23416: std_logic; attribute dont_touch of G23416: signal is true;
	signal G23417: std_logic; attribute dont_touch of G23417: signal is true;
	signal G23418: std_logic; attribute dont_touch of G23418: signal is true;
	signal G23419: std_logic; attribute dont_touch of G23419: signal is true;
	signal G23420: std_logic; attribute dont_touch of G23420: signal is true;
	signal G23421: std_logic; attribute dont_touch of G23421: signal is true;
	signal G23422: std_logic; attribute dont_touch of G23422: signal is true;
	signal G23423: std_logic; attribute dont_touch of G23423: signal is true;
	signal G23424: std_logic; attribute dont_touch of G23424: signal is true;
	signal G23425: std_logic; attribute dont_touch of G23425: signal is true;
	signal G23426: std_logic; attribute dont_touch of G23426: signal is true;
	signal G23427: std_logic; attribute dont_touch of G23427: signal is true;
	signal G23428: std_logic; attribute dont_touch of G23428: signal is true;
	signal G23429: std_logic; attribute dont_touch of G23429: signal is true;
	signal G23430: std_logic; attribute dont_touch of G23430: signal is true;
	signal G23431: std_logic; attribute dont_touch of G23431: signal is true;
	signal G23432: std_logic; attribute dont_touch of G23432: signal is true;
	signal G23433: std_logic; attribute dont_touch of G23433: signal is true;
	signal G23434: std_logic; attribute dont_touch of G23434: signal is true;
	signal G23435: std_logic; attribute dont_touch of G23435: signal is true;
	signal G23436: std_logic; attribute dont_touch of G23436: signal is true;
	signal G23439: std_logic; attribute dont_touch of G23439: signal is true;
	signal G23440: std_logic; attribute dont_touch of G23440: signal is true;
	signal G23443: std_logic; attribute dont_touch of G23443: signal is true;
	signal G23444: std_logic; attribute dont_touch of G23444: signal is true;
	signal G23445: std_logic; attribute dont_touch of G23445: signal is true;
	signal G23446: std_logic; attribute dont_touch of G23446: signal is true;
	signal G23447: std_logic; attribute dont_touch of G23447: signal is true;
	signal G23448: std_logic; attribute dont_touch of G23448: signal is true;
	signal G23449: std_logic; attribute dont_touch of G23449: signal is true;
	signal G23450: std_logic; attribute dont_touch of G23450: signal is true;
	signal G23451: std_logic; attribute dont_touch of G23451: signal is true;
	signal G23452: std_logic; attribute dont_touch of G23452: signal is true;
	signal G23453: std_logic; attribute dont_touch of G23453: signal is true;
	signal G23456: std_logic; attribute dont_touch of G23456: signal is true;
	signal G23457: std_logic; attribute dont_touch of G23457: signal is true;
	signal G23458: std_logic; attribute dont_touch of G23458: signal is true;
	signal G23459: std_logic; attribute dont_touch of G23459: signal is true;
	signal G23460: std_logic; attribute dont_touch of G23460: signal is true;
	signal G23461: std_logic; attribute dont_touch of G23461: signal is true;
	signal G23462: std_logic; attribute dont_touch of G23462: signal is true;
	signal G23471: std_logic; attribute dont_touch of G23471: signal is true;
	signal G23472: std_logic; attribute dont_touch of G23472: signal is true;
	signal G23473: std_logic; attribute dont_touch of G23473: signal is true;
	signal G23474: std_logic; attribute dont_touch of G23474: signal is true;
	signal G23475: std_logic; attribute dont_touch of G23475: signal is true;
	signal G23476: std_logic; attribute dont_touch of G23476: signal is true;
	signal G23477: std_logic; attribute dont_touch of G23477: signal is true;
	signal G23478: std_logic; attribute dont_touch of G23478: signal is true;
	signal G23479: std_logic; attribute dont_touch of G23479: signal is true;
	signal G23480: std_logic; attribute dont_touch of G23480: signal is true;
	signal G23481: std_logic; attribute dont_touch of G23481: signal is true;
	signal G23482: std_logic; attribute dont_touch of G23482: signal is true;
	signal G23483: std_logic; attribute dont_touch of G23483: signal is true;
	signal G23484: std_logic; attribute dont_touch of G23484: signal is true;
	signal G23485: std_logic; attribute dont_touch of G23485: signal is true;
	signal G23486: std_logic; attribute dont_touch of G23486: signal is true;
	signal G23487: std_logic; attribute dont_touch of G23487: signal is true;
	signal G23488: std_logic; attribute dont_touch of G23488: signal is true;
	signal G23489: std_logic; attribute dont_touch of G23489: signal is true;
	signal G23490: std_logic; attribute dont_touch of G23490: signal is true;
	signal G23491: std_logic; attribute dont_touch of G23491: signal is true;
	signal G23492: std_logic; attribute dont_touch of G23492: signal is true;
	signal G23493: std_logic; attribute dont_touch of G23493: signal is true;
	signal G23494: std_logic; attribute dont_touch of G23494: signal is true;
	signal G23495: std_logic; attribute dont_touch of G23495: signal is true;
	signal G23496: std_logic; attribute dont_touch of G23496: signal is true;
	signal G23497: std_logic; attribute dont_touch of G23497: signal is true;
	signal G23498: std_logic; attribute dont_touch of G23498: signal is true;
	signal G23499: std_logic; attribute dont_touch of G23499: signal is true;
	signal G23500: std_logic; attribute dont_touch of G23500: signal is true;
	signal G23501: std_logic; attribute dont_touch of G23501: signal is true;
	signal G23502: std_logic; attribute dont_touch of G23502: signal is true;
	signal G23503: std_logic; attribute dont_touch of G23503: signal is true;
	signal G23504: std_logic; attribute dont_touch of G23504: signal is true;
	signal G23505: std_logic; attribute dont_touch of G23505: signal is true;
	signal G23506: std_logic; attribute dont_touch of G23506: signal is true;
	signal G23507: std_logic; attribute dont_touch of G23507: signal is true;
	signal G23508: std_logic; attribute dont_touch of G23508: signal is true;
	signal G23509: std_logic; attribute dont_touch of G23509: signal is true;
	signal G23510: std_logic; attribute dont_touch of G23510: signal is true;
	signal G23511: std_logic; attribute dont_touch of G23511: signal is true;
	signal G23512: std_logic; attribute dont_touch of G23512: signal is true;
	signal G23513: std_logic; attribute dont_touch of G23513: signal is true;
	signal G23514: std_logic; attribute dont_touch of G23514: signal is true;
	signal G23515: std_logic; attribute dont_touch of G23515: signal is true;
	signal G23516: std_logic; attribute dont_touch of G23516: signal is true;
	signal G23517: std_logic; attribute dont_touch of G23517: signal is true;
	signal G23518: std_logic; attribute dont_touch of G23518: signal is true;
	signal G23519: std_logic; attribute dont_touch of G23519: signal is true;
	signal G23520: std_logic; attribute dont_touch of G23520: signal is true;
	signal G23521: std_logic; attribute dont_touch of G23521: signal is true;
	signal G23522: std_logic; attribute dont_touch of G23522: signal is true;
	signal G23523: std_logic; attribute dont_touch of G23523: signal is true;
	signal G23524: std_logic; attribute dont_touch of G23524: signal is true;
	signal G23525: std_logic; attribute dont_touch of G23525: signal is true;
	signal G23526: std_logic; attribute dont_touch of G23526: signal is true;
	signal G23527: std_logic; attribute dont_touch of G23527: signal is true;
	signal G23528: std_logic; attribute dont_touch of G23528: signal is true;
	signal G23529: std_logic; attribute dont_touch of G23529: signal is true;
	signal G23530: std_logic; attribute dont_touch of G23530: signal is true;
	signal G23531: std_logic; attribute dont_touch of G23531: signal is true;
	signal G23532: std_logic; attribute dont_touch of G23532: signal is true;
	signal G23533: std_logic; attribute dont_touch of G23533: signal is true;
	signal G23534: std_logic; attribute dont_touch of G23534: signal is true;
	signal G23537: std_logic; attribute dont_touch of G23537: signal is true;
	signal G23538: std_logic; attribute dont_touch of G23538: signal is true;
	signal G23539: std_logic; attribute dont_touch of G23539: signal is true;
	signal G23540: std_logic; attribute dont_touch of G23540: signal is true;
	signal G23541: std_logic; attribute dont_touch of G23541: signal is true;
	signal G23542: std_logic; attribute dont_touch of G23542: signal is true;
	signal G23543: std_logic; attribute dont_touch of G23543: signal is true;
	signal G23544: std_logic; attribute dont_touch of G23544: signal is true;
	signal G23545: std_logic; attribute dont_touch of G23545: signal is true;
	signal G23546: std_logic; attribute dont_touch of G23546: signal is true;
	signal G23547: std_logic; attribute dont_touch of G23547: signal is true;
	signal G23548: std_logic; attribute dont_touch of G23548: signal is true;
	signal G23549: std_logic; attribute dont_touch of G23549: signal is true;
	signal G23550: std_logic; attribute dont_touch of G23550: signal is true;
	signal G23551: std_logic; attribute dont_touch of G23551: signal is true;
	signal G23552: std_logic; attribute dont_touch of G23552: signal is true;
	signal G23553: std_logic; attribute dont_touch of G23553: signal is true;
	signal G23554: std_logic; attribute dont_touch of G23554: signal is true;
	signal G23555: std_logic; attribute dont_touch of G23555: signal is true;
	signal G23558: std_logic; attribute dont_touch of G23558: signal is true;
	signal G23559: std_logic; attribute dont_touch of G23559: signal is true;
	signal G23560: std_logic; attribute dont_touch of G23560: signal is true;
	signal G23563: std_logic; attribute dont_touch of G23563: signal is true;
	signal G23564: std_logic; attribute dont_touch of G23564: signal is true;
	signal G23565: std_logic; attribute dont_touch of G23565: signal is true;
	signal G23566: std_logic; attribute dont_touch of G23566: signal is true;
	signal G23567: std_logic; attribute dont_touch of G23567: signal is true;
	signal G23568: std_logic; attribute dont_touch of G23568: signal is true;
	signal G23569: std_logic; attribute dont_touch of G23569: signal is true;
	signal G23570: std_logic; attribute dont_touch of G23570: signal is true;
	signal G23571: std_logic; attribute dont_touch of G23571: signal is true;
	signal G23572: std_logic; attribute dont_touch of G23572: signal is true;
	signal G23573: std_logic; attribute dont_touch of G23573: signal is true;
	signal G23574: std_logic; attribute dont_touch of G23574: signal is true;
	signal G23575: std_logic; attribute dont_touch of G23575: signal is true;
	signal G23576: std_logic; attribute dont_touch of G23576: signal is true;
	signal G23577: std_logic; attribute dont_touch of G23577: signal is true;
	signal G23578: std_logic; attribute dont_touch of G23578: signal is true;
	signal G23581: std_logic; attribute dont_touch of G23581: signal is true;
	signal G23582: std_logic; attribute dont_touch of G23582: signal is true;
	signal G23585: std_logic; attribute dont_touch of G23585: signal is true;
	signal G23586: std_logic; attribute dont_touch of G23586: signal is true;
	signal G23589: std_logic; attribute dont_touch of G23589: signal is true;
	signal G23590: std_logic; attribute dont_touch of G23590: signal is true;
	signal G23599: std_logic; attribute dont_touch of G23599: signal is true;
	signal G23602: std_logic; attribute dont_touch of G23602: signal is true;
	signal G23605: std_logic; attribute dont_touch of G23605: signal is true;
	signal G23606: std_logic; attribute dont_touch of G23606: signal is true;
	signal G23607: std_logic; attribute dont_touch of G23607: signal is true;
	signal G23608: std_logic; attribute dont_touch of G23608: signal is true;
	signal G23609: std_logic; attribute dont_touch of G23609: signal is true;
	signal G23610: std_logic; attribute dont_touch of G23610: signal is true;
	signal G23611: std_logic; attribute dont_touch of G23611: signal is true;
	signal G23613: std_logic; attribute dont_touch of G23613: signal is true;
	signal G23614: std_logic; attribute dont_touch of G23614: signal is true;
	signal G23615: std_logic; attribute dont_touch of G23615: signal is true;
	signal G23616: std_logic; attribute dont_touch of G23616: signal is true;
	signal G23617: std_logic; attribute dont_touch of G23617: signal is true;
	signal G23618: std_logic; attribute dont_touch of G23618: signal is true;
	signal G23619: std_logic; attribute dont_touch of G23619: signal is true;
	signal G23620: std_logic; attribute dont_touch of G23620: signal is true;
	signal G23623: std_logic; attribute dont_touch of G23623: signal is true;
	signal G23626: std_logic; attribute dont_touch of G23626: signal is true;
	signal G23629: std_logic; attribute dont_touch of G23629: signal is true;
	signal G23630: std_logic; attribute dont_touch of G23630: signal is true;
	signal G23639: std_logic; attribute dont_touch of G23639: signal is true;
	signal G23642: std_logic; attribute dont_touch of G23642: signal is true;
	signal G23645: std_logic; attribute dont_touch of G23645: signal is true;
	signal G23646: std_logic; attribute dont_touch of G23646: signal is true;
	signal G23647: std_logic; attribute dont_touch of G23647: signal is true;
	signal G23648: std_logic; attribute dont_touch of G23648: signal is true;
	signal G23649: std_logic; attribute dont_touch of G23649: signal is true;
	signal G23650: std_logic; attribute dont_touch of G23650: signal is true;
	signal G23651: std_logic; attribute dont_touch of G23651: signal is true;
	signal G23653: std_logic; attribute dont_touch of G23653: signal is true;
	signal G23654: std_logic; attribute dont_touch of G23654: signal is true;
	signal G23655: std_logic; attribute dont_touch of G23655: signal is true;
	signal G23656: std_logic; attribute dont_touch of G23656: signal is true;
	signal G23657: std_logic; attribute dont_touch of G23657: signal is true;
	signal G23658: std_logic; attribute dont_touch of G23658: signal is true;
	signal G23659: std_logic; attribute dont_touch of G23659: signal is true;
	signal G23662: std_logic; attribute dont_touch of G23662: signal is true;
	signal G23665: std_logic; attribute dont_touch of G23665: signal is true;
	signal G23666: std_logic; attribute dont_touch of G23666: signal is true;
	signal G23675: std_logic; attribute dont_touch of G23675: signal is true;
	signal G23678: std_logic; attribute dont_touch of G23678: signal is true;
	signal G23681: std_logic; attribute dont_touch of G23681: signal is true;
	signal G23682: std_logic; attribute dont_touch of G23682: signal is true;
	signal G23684: std_logic; attribute dont_touch of G23684: signal is true;
	signal G23685: std_logic; attribute dont_touch of G23685: signal is true;
	signal G23686: std_logic; attribute dont_touch of G23686: signal is true;
	signal G23687: std_logic; attribute dont_touch of G23687: signal is true;
	signal G23690: std_logic; attribute dont_touch of G23690: signal is true;
	signal G23691: std_logic; attribute dont_touch of G23691: signal is true;
	signal G23692: std_logic; attribute dont_touch of G23692: signal is true;
	signal G23695: std_logic; attribute dont_touch of G23695: signal is true;
	signal G23698: std_logic; attribute dont_touch of G23698: signal is true;
	signal G23699: std_logic; attribute dont_touch of G23699: signal is true;
	signal G23708: std_logic; attribute dont_touch of G23708: signal is true;
	signal G23711: std_logic; attribute dont_touch of G23711: signal is true;
	signal G23714: std_logic; attribute dont_touch of G23714: signal is true;
	signal G23715: std_logic; attribute dont_touch of G23715: signal is true;
	signal G23716: std_logic; attribute dont_touch of G23716: signal is true;
	signal G23719: std_logic; attribute dont_touch of G23719: signal is true;
	signal G23720: std_logic; attribute dont_touch of G23720: signal is true;
	signal G23721: std_logic; attribute dont_touch of G23721: signal is true;
	signal G23724: std_logic; attribute dont_touch of G23724: signal is true;
	signal G23725: std_logic; attribute dont_touch of G23725: signal is true;
	signal G23726: std_logic; attribute dont_touch of G23726: signal is true;
	signal G23729: std_logic; attribute dont_touch of G23729: signal is true;
	signal G23732: std_logic; attribute dont_touch of G23732: signal is true;
	signal G23733: std_logic; attribute dont_touch of G23733: signal is true;
	signal G23742: std_logic; attribute dont_touch of G23742: signal is true;
	signal G23745: std_logic; attribute dont_touch of G23745: signal is true;
	signal G23746: std_logic; attribute dont_touch of G23746: signal is true;
	signal G23747: std_logic; attribute dont_touch of G23747: signal is true;
	signal G23748: std_logic; attribute dont_touch of G23748: signal is true;
	signal G23749: std_logic; attribute dont_touch of G23749: signal is true;
	signal G23750: std_logic; attribute dont_touch of G23750: signal is true;
	signal G23751: std_logic; attribute dont_touch of G23751: signal is true;
	signal G23754: std_logic; attribute dont_touch of G23754: signal is true;
	signal G23755: std_logic; attribute dont_touch of G23755: signal is true;
	signal G23756: std_logic; attribute dont_touch of G23756: signal is true;
	signal G23760: std_logic; attribute dont_touch of G23760: signal is true;
	signal G23761: std_logic; attribute dont_touch of G23761: signal is true;
	signal G23762: std_logic; attribute dont_touch of G23762: signal is true;
	signal G23763: std_logic; attribute dont_touch of G23763: signal is true;
	signal G23764: std_logic; attribute dont_touch of G23764: signal is true;
	signal G23767: std_logic; attribute dont_touch of G23767: signal is true;
	signal G23768: std_logic; attribute dont_touch of G23768: signal is true;
	signal G23769: std_logic; attribute dont_touch of G23769: signal is true;
	signal G23770: std_logic; attribute dont_touch of G23770: signal is true;
	signal G23771: std_logic; attribute dont_touch of G23771: signal is true;
	signal G23774: std_logic; attribute dont_touch of G23774: signal is true;
	signal G23775: std_logic; attribute dont_touch of G23775: signal is true;
	signal G23776: std_logic; attribute dont_touch of G23776: signal is true;
	signal G23777: std_logic; attribute dont_touch of G23777: signal is true;
	signal G23778: std_logic; attribute dont_touch of G23778: signal is true;
	signal G23779: std_logic; attribute dont_touch of G23779: signal is true;
	signal G23780: std_logic; attribute dont_touch of G23780: signal is true;
	signal G23781: std_logic; attribute dont_touch of G23781: signal is true;
	signal G23782: std_logic; attribute dont_touch of G23782: signal is true;
	signal G23786: std_logic; attribute dont_touch of G23786: signal is true;
	signal G23787: std_logic; attribute dont_touch of G23787: signal is true;
	signal G23788: std_logic; attribute dont_touch of G23788: signal is true;
	signal G23789: std_logic; attribute dont_touch of G23789: signal is true;
	signal G23792: std_logic; attribute dont_touch of G23792: signal is true;
	signal G23793: std_logic; attribute dont_touch of G23793: signal is true;
	signal G23794: std_logic; attribute dont_touch of G23794: signal is true;
	signal G23795: std_logic; attribute dont_touch of G23795: signal is true;
	signal G23796: std_logic; attribute dont_touch of G23796: signal is true;
	signal G23799: std_logic; attribute dont_touch of G23799: signal is true;
	signal G23800: std_logic; attribute dont_touch of G23800: signal is true;
	signal G23801: std_logic; attribute dont_touch of G23801: signal is true;
	signal G23802: std_logic; attribute dont_touch of G23802: signal is true;
	signal G23809: std_logic; attribute dont_touch of G23809: signal is true;
	signal G23810: std_logic; attribute dont_touch of G23810: signal is true;
	signal G23811: std_logic; attribute dont_touch of G23811: signal is true;
	signal G23812: std_logic; attribute dont_touch of G23812: signal is true;
	signal G23813: std_logic; attribute dont_touch of G23813: signal is true;
	signal G23814: std_logic; attribute dont_touch of G23814: signal is true;
	signal G23815: std_logic; attribute dont_touch of G23815: signal is true;
	signal G23816: std_logic; attribute dont_touch of G23816: signal is true;
	signal G23819: std_logic; attribute dont_touch of G23819: signal is true;
	signal G23820: std_logic; attribute dont_touch of G23820: signal is true;
	signal G23821: std_logic; attribute dont_touch of G23821: signal is true;
	signal G23822: std_logic; attribute dont_touch of G23822: signal is true;
	signal G23823: std_logic; attribute dont_touch of G23823: signal is true;
	signal G23824: std_logic; attribute dont_touch of G23824: signal is true;
	signal G23825: std_logic; attribute dont_touch of G23825: signal is true;
	signal G23828: std_logic; attribute dont_touch of G23828: signal is true;
	signal G23835: std_logic; attribute dont_touch of G23835: signal is true;
	signal G23836: std_logic; attribute dont_touch of G23836: signal is true;
	signal G23837: std_logic; attribute dont_touch of G23837: signal is true;
	signal G23838: std_logic; attribute dont_touch of G23838: signal is true;
	signal G23839: std_logic; attribute dont_touch of G23839: signal is true;
	signal G23840: std_logic; attribute dont_touch of G23840: signal is true;
	signal G23841: std_logic; attribute dont_touch of G23841: signal is true;
	signal G23842: std_logic; attribute dont_touch of G23842: signal is true;
	signal G23843: std_logic; attribute dont_touch of G23843: signal is true;
	signal G23844: std_logic; attribute dont_touch of G23844: signal is true;
	signal G23847: std_logic; attribute dont_touch of G23847: signal is true;
	signal G23848: std_logic; attribute dont_touch of G23848: signal is true;
	signal G23849: std_logic; attribute dont_touch of G23849: signal is true;
	signal G23850: std_logic; attribute dont_touch of G23850: signal is true;
	signal G23854: std_logic; attribute dont_touch of G23854: signal is true;
	signal G23855: std_logic; attribute dont_touch of G23855: signal is true;
	signal G23856: std_logic; attribute dont_touch of G23856: signal is true;
	signal G23857: std_logic; attribute dont_touch of G23857: signal is true;
	signal G23858: std_logic; attribute dont_touch of G23858: signal is true;
	signal G23859: std_logic; attribute dont_touch of G23859: signal is true;
	signal G23860: std_logic; attribute dont_touch of G23860: signal is true;
	signal G23861: std_logic; attribute dont_touch of G23861: signal is true;
	signal G23862: std_logic; attribute dont_touch of G23862: signal is true;
	signal G23863: std_logic; attribute dont_touch of G23863: signal is true;
	signal G23864: std_logic; attribute dont_touch of G23864: signal is true;
	signal G23865: std_logic; attribute dont_touch of G23865: signal is true;
	signal G23868: std_logic; attribute dont_touch of G23868: signal is true;
	signal G23869: std_logic; attribute dont_touch of G23869: signal is true;
	signal G23870: std_logic; attribute dont_touch of G23870: signal is true;
	signal G23871: std_logic; attribute dont_touch of G23871: signal is true;
	signal G23872: std_logic; attribute dont_touch of G23872: signal is true;
	signal G23873: std_logic; attribute dont_touch of G23873: signal is true;
	signal G23874: std_logic; attribute dont_touch of G23874: signal is true;
	signal G23875: std_logic; attribute dont_touch of G23875: signal is true;
	signal G23876: std_logic; attribute dont_touch of G23876: signal is true;
	signal G23877: std_logic; attribute dont_touch of G23877: signal is true;
	signal G23878: std_logic; attribute dont_touch of G23878: signal is true;
	signal G23879: std_logic; attribute dont_touch of G23879: signal is true;
	signal G23880: std_logic; attribute dont_touch of G23880: signal is true;
	signal G23881: std_logic; attribute dont_touch of G23881: signal is true;
	signal G23882: std_logic; attribute dont_touch of G23882: signal is true;
	signal G23883: std_logic; attribute dont_touch of G23883: signal is true;
	signal G23884: std_logic; attribute dont_touch of G23884: signal is true;
	signal G23885: std_logic; attribute dont_touch of G23885: signal is true;
	signal G23886: std_logic; attribute dont_touch of G23886: signal is true;
	signal G23887: std_logic; attribute dont_touch of G23887: signal is true;
	signal G23888: std_logic; attribute dont_touch of G23888: signal is true;
	signal G23889: std_logic; attribute dont_touch of G23889: signal is true;
	signal G23890: std_logic; attribute dont_touch of G23890: signal is true;
	signal G23893: std_logic; attribute dont_touch of G23893: signal is true;
	signal G23894: std_logic; attribute dont_touch of G23894: signal is true;
	signal G23895: std_logic; attribute dont_touch of G23895: signal is true;
	signal G23896: std_logic; attribute dont_touch of G23896: signal is true;
	signal G23897: std_logic; attribute dont_touch of G23897: signal is true;
	signal G23898: std_logic; attribute dont_touch of G23898: signal is true;
	signal G23899: std_logic; attribute dont_touch of G23899: signal is true;
	signal G23900: std_logic; attribute dont_touch of G23900: signal is true;
	signal G23901: std_logic; attribute dont_touch of G23901: signal is true;
	signal G23902: std_logic; attribute dont_touch of G23902: signal is true;
	signal G23903: std_logic; attribute dont_touch of G23903: signal is true;
	signal G23904: std_logic; attribute dont_touch of G23904: signal is true;
	signal G23905: std_logic; attribute dont_touch of G23905: signal is true;
	signal G23906: std_logic; attribute dont_touch of G23906: signal is true;
	signal G23907: std_logic; attribute dont_touch of G23907: signal is true;
	signal G23908: std_logic; attribute dont_touch of G23908: signal is true;
	signal G23909: std_logic; attribute dont_touch of G23909: signal is true;
	signal G23912: std_logic; attribute dont_touch of G23912: signal is true;
	signal G23913: std_logic; attribute dont_touch of G23913: signal is true;
	signal G23914: std_logic; attribute dont_touch of G23914: signal is true;
	signal G23915: std_logic; attribute dont_touch of G23915: signal is true;
	signal G23916: std_logic; attribute dont_touch of G23916: signal is true;
	signal G23917: std_logic; attribute dont_touch of G23917: signal is true;
	signal G23918: std_logic; attribute dont_touch of G23918: signal is true;
	signal G23919: std_logic; attribute dont_touch of G23919: signal is true;
	signal G23920: std_logic; attribute dont_touch of G23920: signal is true;
	signal G23921: std_logic; attribute dont_touch of G23921: signal is true;
	signal G23922: std_logic; attribute dont_touch of G23922: signal is true;
	signal G23923: std_logic; attribute dont_touch of G23923: signal is true;
	signal G23924: std_logic; attribute dont_touch of G23924: signal is true;
	signal G23925: std_logic; attribute dont_touch of G23925: signal is true;
	signal G23926: std_logic; attribute dont_touch of G23926: signal is true;
	signal G23927: std_logic; attribute dont_touch of G23927: signal is true;
	signal G23928: std_logic; attribute dont_touch of G23928: signal is true;
	signal G23929: std_logic; attribute dont_touch of G23929: signal is true;
	signal G23930: std_logic; attribute dont_touch of G23930: signal is true;
	signal G23931: std_logic; attribute dont_touch of G23931: signal is true;
	signal G23932: std_logic; attribute dont_touch of G23932: signal is true;
	signal G23935: std_logic; attribute dont_touch of G23935: signal is true;
	signal G23936: std_logic; attribute dont_touch of G23936: signal is true;
	signal G23937: std_logic; attribute dont_touch of G23937: signal is true;
	signal G23938: std_logic; attribute dont_touch of G23938: signal is true;
	signal G23939: std_logic; attribute dont_touch of G23939: signal is true;
	signal G23940: std_logic; attribute dont_touch of G23940: signal is true;
	signal G23941: std_logic; attribute dont_touch of G23941: signal is true;
	signal G23942: std_logic; attribute dont_touch of G23942: signal is true;
	signal G23943: std_logic; attribute dont_touch of G23943: signal is true;
	signal G23944: std_logic; attribute dont_touch of G23944: signal is true;
	signal G23945: std_logic; attribute dont_touch of G23945: signal is true;
	signal G23946: std_logic; attribute dont_touch of G23946: signal is true;
	signal G23947: std_logic; attribute dont_touch of G23947: signal is true;
	signal G23948: std_logic; attribute dont_touch of G23948: signal is true;
	signal G23949: std_logic; attribute dont_touch of G23949: signal is true;
	signal G23952: std_logic; attribute dont_touch of G23952: signal is true;
	signal G23953: std_logic; attribute dont_touch of G23953: signal is true;
	signal G23954: std_logic; attribute dont_touch of G23954: signal is true;
	signal G23955: std_logic; attribute dont_touch of G23955: signal is true;
	signal G23956: std_logic; attribute dont_touch of G23956: signal is true;
	signal G23957: std_logic; attribute dont_touch of G23957: signal is true;
	signal G23958: std_logic; attribute dont_touch of G23958: signal is true;
	signal G23961: std_logic; attribute dont_touch of G23961: signal is true;
	signal G23962: std_logic; attribute dont_touch of G23962: signal is true;
	signal G23963: std_logic; attribute dont_touch of G23963: signal is true;
	signal G23964: std_logic; attribute dont_touch of G23964: signal is true;
	signal G23965: std_logic; attribute dont_touch of G23965: signal is true;
	signal G23966: std_logic; attribute dont_touch of G23966: signal is true;
	signal G23967: std_logic; attribute dont_touch of G23967: signal is true;
	signal G23968: std_logic; attribute dont_touch of G23968: signal is true;
	signal G23969: std_logic; attribute dont_touch of G23969: signal is true;
	signal G23970: std_logic; attribute dont_touch of G23970: signal is true;
	signal G23971: std_logic; attribute dont_touch of G23971: signal is true;
	signal G23972: std_logic; attribute dont_touch of G23972: signal is true;
	signal G23975: std_logic; attribute dont_touch of G23975: signal is true;
	signal G23978: std_logic; attribute dont_touch of G23978: signal is true;
	signal G23982: std_logic; attribute dont_touch of G23982: signal is true;
	signal G23983: std_logic; attribute dont_touch of G23983: signal is true;
	signal G23984: std_logic; attribute dont_touch of G23984: signal is true;
	signal G23985: std_logic; attribute dont_touch of G23985: signal is true;
	signal G23986: std_logic; attribute dont_touch of G23986: signal is true;
	signal G23987: std_logic; attribute dont_touch of G23987: signal is true;
	signal G23988: std_logic; attribute dont_touch of G23988: signal is true;
	signal G23989: std_logic; attribute dont_touch of G23989: signal is true;
	signal G23990: std_logic; attribute dont_touch of G23990: signal is true;
	signal G23991: std_logic; attribute dont_touch of G23991: signal is true;
	signal G23992: std_logic; attribute dont_touch of G23992: signal is true;
	signal G23993: std_logic; attribute dont_touch of G23993: signal is true;
	signal G23994: std_logic; attribute dont_touch of G23994: signal is true;
	signal G23995: std_logic; attribute dont_touch of G23995: signal is true;
	signal G23996: std_logic; attribute dont_touch of G23996: signal is true;
	signal G23997: std_logic; attribute dont_touch of G23997: signal is true;
	signal G23998: std_logic; attribute dont_touch of G23998: signal is true;
	signal G23999: std_logic; attribute dont_touch of G23999: signal is true;
	signal G24000: std_logic; attribute dont_touch of G24000: signal is true;
	signal G24001: std_logic; attribute dont_touch of G24001: signal is true;
	signal G24002: std_logic; attribute dont_touch of G24002: signal is true;
	signal G24003: std_logic; attribute dont_touch of G24003: signal is true;
	signal G24004: std_logic; attribute dont_touch of G24004: signal is true;
	signal G24005: std_logic; attribute dont_touch of G24005: signal is true;
	signal G24008: std_logic; attribute dont_touch of G24008: signal is true;
	signal G24009: std_logic; attribute dont_touch of G24009: signal is true;
	signal G24010: std_logic; attribute dont_touch of G24010: signal is true;
	signal G24011: std_logic; attribute dont_touch of G24011: signal is true;
	signal G24012: std_logic; attribute dont_touch of G24012: signal is true;
	signal G24013: std_logic; attribute dont_touch of G24013: signal is true;
	signal G24014: std_logic; attribute dont_touch of G24014: signal is true;
	signal G24015: std_logic; attribute dont_touch of G24015: signal is true;
	signal G24016: std_logic; attribute dont_touch of G24016: signal is true;
	signal G24017: std_logic; attribute dont_touch of G24017: signal is true;
	signal G24018: std_logic; attribute dont_touch of G24018: signal is true;
	signal G24019: std_logic; attribute dont_touch of G24019: signal is true;
	signal G24020: std_logic; attribute dont_touch of G24020: signal is true;
	signal G24021: std_logic; attribute dont_touch of G24021: signal is true;
	signal G24022: std_logic; attribute dont_touch of G24022: signal is true;
	signal G24023: std_logic; attribute dont_touch of G24023: signal is true;
	signal G24024: std_logic; attribute dont_touch of G24024: signal is true;
	signal G24025: std_logic; attribute dont_touch of G24025: signal is true;
	signal G24026: std_logic; attribute dont_touch of G24026: signal is true;
	signal G24027: std_logic; attribute dont_touch of G24027: signal is true;
	signal G24028: std_logic; attribute dont_touch of G24028: signal is true;
	signal G24029: std_logic; attribute dont_touch of G24029: signal is true;
	signal G24030: std_logic; attribute dont_touch of G24030: signal is true;
	signal G24031: std_logic; attribute dont_touch of G24031: signal is true;
	signal G24032: std_logic; attribute dont_touch of G24032: signal is true;
	signal G24033: std_logic; attribute dont_touch of G24033: signal is true;
	signal G24034: std_logic; attribute dont_touch of G24034: signal is true;
	signal G24035: std_logic; attribute dont_touch of G24035: signal is true;
	signal G24036: std_logic; attribute dont_touch of G24036: signal is true;
	signal G24037: std_logic; attribute dont_touch of G24037: signal is true;
	signal G24038: std_logic; attribute dont_touch of G24038: signal is true;
	signal G24039: std_logic; attribute dont_touch of G24039: signal is true;
	signal G24040: std_logic; attribute dont_touch of G24040: signal is true;
	signal G24041: std_logic; attribute dont_touch of G24041: signal is true;
	signal G24042: std_logic; attribute dont_touch of G24042: signal is true;
	signal G24043: std_logic; attribute dont_touch of G24043: signal is true;
	signal G24044: std_logic; attribute dont_touch of G24044: signal is true;
	signal G24045: std_logic; attribute dont_touch of G24045: signal is true;
	signal G24046: std_logic; attribute dont_touch of G24046: signal is true;
	signal G24047: std_logic; attribute dont_touch of G24047: signal is true;
	signal G24048: std_logic; attribute dont_touch of G24048: signal is true;
	signal G24049: std_logic; attribute dont_touch of G24049: signal is true;
	signal G24050: std_logic; attribute dont_touch of G24050: signal is true;
	signal G24051: std_logic; attribute dont_touch of G24051: signal is true;
	signal G24052: std_logic; attribute dont_touch of G24052: signal is true;
	signal G24053: std_logic; attribute dont_touch of G24053: signal is true;
	signal G24054: std_logic; attribute dont_touch of G24054: signal is true;
	signal G24055: std_logic; attribute dont_touch of G24055: signal is true;
	signal G24056: std_logic; attribute dont_touch of G24056: signal is true;
	signal G24057: std_logic; attribute dont_touch of G24057: signal is true;
	signal G24058: std_logic; attribute dont_touch of G24058: signal is true;
	signal G24059: std_logic; attribute dont_touch of G24059: signal is true;
	signal G24060: std_logic; attribute dont_touch of G24060: signal is true;
	signal G24061: std_logic; attribute dont_touch of G24061: signal is true;
	signal G24062: std_logic; attribute dont_touch of G24062: signal is true;
	signal G24063: std_logic; attribute dont_touch of G24063: signal is true;
	signal G24064: std_logic; attribute dont_touch of G24064: signal is true;
	signal G24065: std_logic; attribute dont_touch of G24065: signal is true;
	signal G24066: std_logic; attribute dont_touch of G24066: signal is true;
	signal G24067: std_logic; attribute dont_touch of G24067: signal is true;
	signal G24068: std_logic; attribute dont_touch of G24068: signal is true;
	signal G24069: std_logic; attribute dont_touch of G24069: signal is true;
	signal G24070: std_logic; attribute dont_touch of G24070: signal is true;
	signal G24071: std_logic; attribute dont_touch of G24071: signal is true;
	signal G24072: std_logic; attribute dont_touch of G24072: signal is true;
	signal G24073: std_logic; attribute dont_touch of G24073: signal is true;
	signal G24074: std_logic; attribute dont_touch of G24074: signal is true;
	signal G24075: std_logic; attribute dont_touch of G24075: signal is true;
	signal G24076: std_logic; attribute dont_touch of G24076: signal is true;
	signal G24077: std_logic; attribute dont_touch of G24077: signal is true;
	signal G24078: std_logic; attribute dont_touch of G24078: signal is true;
	signal G24079: std_logic; attribute dont_touch of G24079: signal is true;
	signal G24080: std_logic; attribute dont_touch of G24080: signal is true;
	signal G24081: std_logic; attribute dont_touch of G24081: signal is true;
	signal G24082: std_logic; attribute dont_touch of G24082: signal is true;
	signal G24083: std_logic; attribute dont_touch of G24083: signal is true;
	signal G24084: std_logic; attribute dont_touch of G24084: signal is true;
	signal G24085: std_logic; attribute dont_touch of G24085: signal is true;
	signal G24086: std_logic; attribute dont_touch of G24086: signal is true;
	signal G24087: std_logic; attribute dont_touch of G24087: signal is true;
	signal G24088: std_logic; attribute dont_touch of G24088: signal is true;
	signal G24089: std_logic; attribute dont_touch of G24089: signal is true;
	signal G24090: std_logic; attribute dont_touch of G24090: signal is true;
	signal G24091: std_logic; attribute dont_touch of G24091: signal is true;
	signal G24092: std_logic; attribute dont_touch of G24092: signal is true;
	signal G24093: std_logic; attribute dont_touch of G24093: signal is true;
	signal G24094: std_logic; attribute dont_touch of G24094: signal is true;
	signal G24095: std_logic; attribute dont_touch of G24095: signal is true;
	signal G24096: std_logic; attribute dont_touch of G24096: signal is true;
	signal G24097: std_logic; attribute dont_touch of G24097: signal is true;
	signal G24098: std_logic; attribute dont_touch of G24098: signal is true;
	signal G24099: std_logic; attribute dont_touch of G24099: signal is true;
	signal G24100: std_logic; attribute dont_touch of G24100: signal is true;
	signal G24101: std_logic; attribute dont_touch of G24101: signal is true;
	signal G24102: std_logic; attribute dont_touch of G24102: signal is true;
	signal G24103: std_logic; attribute dont_touch of G24103: signal is true;
	signal G24104: std_logic; attribute dont_touch of G24104: signal is true;
	signal G24105: std_logic; attribute dont_touch of G24105: signal is true;
	signal G24106: std_logic; attribute dont_touch of G24106: signal is true;
	signal G24107: std_logic; attribute dont_touch of G24107: signal is true;
	signal G24108: std_logic; attribute dont_touch of G24108: signal is true;
	signal G24109: std_logic; attribute dont_touch of G24109: signal is true;
	signal G24110: std_logic; attribute dont_touch of G24110: signal is true;
	signal G24111: std_logic; attribute dont_touch of G24111: signal is true;
	signal G24112: std_logic; attribute dont_touch of G24112: signal is true;
	signal G24113: std_logic; attribute dont_touch of G24113: signal is true;
	signal G24114: std_logic; attribute dont_touch of G24114: signal is true;
	signal G24115: std_logic; attribute dont_touch of G24115: signal is true;
	signal G24116: std_logic; attribute dont_touch of G24116: signal is true;
	signal G24117: std_logic; attribute dont_touch of G24117: signal is true;
	signal G24118: std_logic; attribute dont_touch of G24118: signal is true;
	signal G24119: std_logic; attribute dont_touch of G24119: signal is true;
	signal G24120: std_logic; attribute dont_touch of G24120: signal is true;
	signal G24121: std_logic; attribute dont_touch of G24121: signal is true;
	signal G24122: std_logic; attribute dont_touch of G24122: signal is true;
	signal G24123: std_logic; attribute dont_touch of G24123: signal is true;
	signal G24124: std_logic; attribute dont_touch of G24124: signal is true;
	signal G24125: std_logic; attribute dont_touch of G24125: signal is true;
	signal G24126: std_logic; attribute dont_touch of G24126: signal is true;
	signal G24127: std_logic; attribute dont_touch of G24127: signal is true;
	signal G24128: std_logic; attribute dont_touch of G24128: signal is true;
	signal G24129: std_logic; attribute dont_touch of G24129: signal is true;
	signal G24130: std_logic; attribute dont_touch of G24130: signal is true;
	signal G24131: std_logic; attribute dont_touch of G24131: signal is true;
	signal G24132: std_logic; attribute dont_touch of G24132: signal is true;
	signal G24133: std_logic; attribute dont_touch of G24133: signal is true;
	signal G24134: std_logic; attribute dont_touch of G24134: signal is true;
	signal G24135: std_logic; attribute dont_touch of G24135: signal is true;
	signal G24136: std_logic; attribute dont_touch of G24136: signal is true;
	signal G24137: std_logic; attribute dont_touch of G24137: signal is true;
	signal G24138: std_logic; attribute dont_touch of G24138: signal is true;
	signal G24139: std_logic; attribute dont_touch of G24139: signal is true;
	signal G24140: std_logic; attribute dont_touch of G24140: signal is true;
	signal G24141: std_logic; attribute dont_touch of G24141: signal is true;
	signal G24142: std_logic; attribute dont_touch of G24142: signal is true;
	signal G24143: std_logic; attribute dont_touch of G24143: signal is true;
	signal G24144: std_logic; attribute dont_touch of G24144: signal is true;
	signal G24145: std_logic; attribute dont_touch of G24145: signal is true;
	signal G24146: std_logic; attribute dont_touch of G24146: signal is true;
	signal G24147: std_logic; attribute dont_touch of G24147: signal is true;
	signal G24148: std_logic; attribute dont_touch of G24148: signal is true;
	signal G24149: std_logic; attribute dont_touch of G24149: signal is true;
	signal G24150: std_logic; attribute dont_touch of G24150: signal is true;
	signal G24152: std_logic; attribute dont_touch of G24152: signal is true;
	signal G24153: std_logic; attribute dont_touch of G24153: signal is true;
	signal G24154: std_logic; attribute dont_touch of G24154: signal is true;
	signal G24155: std_logic; attribute dont_touch of G24155: signal is true;
	signal G24156: std_logic; attribute dont_touch of G24156: signal is true;
	signal G24157: std_logic; attribute dont_touch of G24157: signal is true;
	signal G24158: std_logic; attribute dont_touch of G24158: signal is true;
	signal G24159: std_logic; attribute dont_touch of G24159: signal is true;
	signal G24160: std_logic; attribute dont_touch of G24160: signal is true;
	signal G24186: std_logic; attribute dont_touch of G24186: signal is true;
	signal G24187: std_logic; attribute dont_touch of G24187: signal is true;
	signal G24188: std_logic; attribute dont_touch of G24188: signal is true;
	signal G24189: std_logic; attribute dont_touch of G24189: signal is true;
	signal G24190: std_logic; attribute dont_touch of G24190: signal is true;
	signal G24191: std_logic; attribute dont_touch of G24191: signal is true;
	signal G24192: std_logic; attribute dont_touch of G24192: signal is true;
	signal G24193: std_logic; attribute dont_touch of G24193: signal is true;
	signal G24194: std_logic; attribute dont_touch of G24194: signal is true;
	signal G24195: std_logic; attribute dont_touch of G24195: signal is true;
	signal G24196: std_logic; attribute dont_touch of G24196: signal is true;
	signal G24197: std_logic; attribute dont_touch of G24197: signal is true;
	signal G24198: std_logic; attribute dont_touch of G24198: signal is true;
	signal G24199: std_logic; attribute dont_touch of G24199: signal is true;
	signal G24200: std_logic; attribute dont_touch of G24200: signal is true;
	signal G24201: std_logic; attribute dont_touch of G24201: signal is true;
	signal G24202: std_logic; attribute dont_touch of G24202: signal is true;
	signal G24203: std_logic; attribute dont_touch of G24203: signal is true;
	signal G24204: std_logic; attribute dont_touch of G24204: signal is true;
	signal G24205: std_logic; attribute dont_touch of G24205: signal is true;
	signal G24206: std_logic; attribute dont_touch of G24206: signal is true;
	signal G24207: std_logic; attribute dont_touch of G24207: signal is true;
	signal G24208: std_logic; attribute dont_touch of G24208: signal is true;
	signal G24209: std_logic; attribute dont_touch of G24209: signal is true;
	signal G24210: std_logic; attribute dont_touch of G24210: signal is true;
	signal G24211: std_logic; attribute dont_touch of G24211: signal is true;
	signal G24212: std_logic; attribute dont_touch of G24212: signal is true;
	signal G24213: std_logic; attribute dont_touch of G24213: signal is true;
	signal G24214: std_logic; attribute dont_touch of G24214: signal is true;
	signal G24215: std_logic; attribute dont_touch of G24215: signal is true;
	signal G24216: std_logic; attribute dont_touch of G24216: signal is true;
	signal G24217: std_logic; attribute dont_touch of G24217: signal is true;
	signal G24218: std_logic; attribute dont_touch of G24218: signal is true;
	signal G24219: std_logic; attribute dont_touch of G24219: signal is true;
	signal G24220: std_logic; attribute dont_touch of G24220: signal is true;
	signal G24221: std_logic; attribute dont_touch of G24221: signal is true;
	signal G24222: std_logic; attribute dont_touch of G24222: signal is true;
	signal G24223: std_logic; attribute dont_touch of G24223: signal is true;
	signal G24224: std_logic; attribute dont_touch of G24224: signal is true;
	signal G24225: std_logic; attribute dont_touch of G24225: signal is true;
	signal G24226: std_logic; attribute dont_touch of G24226: signal is true;
	signal G24227: std_logic; attribute dont_touch of G24227: signal is true;
	signal G24228: std_logic; attribute dont_touch of G24228: signal is true;
	signal G24229: std_logic; attribute dont_touch of G24229: signal is true;
	signal G24230: std_logic; attribute dont_touch of G24230: signal is true;
	signal G24231: std_logic; attribute dont_touch of G24231: signal is true;
	signal G24232: std_logic; attribute dont_touch of G24232: signal is true;
	signal G24233: std_logic; attribute dont_touch of G24233: signal is true;
	signal G24234: std_logic; attribute dont_touch of G24234: signal is true;
	signal G24235: std_logic; attribute dont_touch of G24235: signal is true;
	signal G24236: std_logic; attribute dont_touch of G24236: signal is true;
	signal G24237: std_logic; attribute dont_touch of G24237: signal is true;
	signal G24238: std_logic; attribute dont_touch of G24238: signal is true;
	signal G24239: std_logic; attribute dont_touch of G24239: signal is true;
	signal G24240: std_logic; attribute dont_touch of G24240: signal is true;
	signal G24241: std_logic; attribute dont_touch of G24241: signal is true;
	signal G24242: std_logic; attribute dont_touch of G24242: signal is true;
	signal G24243: std_logic; attribute dont_touch of G24243: signal is true;
	signal G24244: std_logic; attribute dont_touch of G24244: signal is true;
	signal G24245: std_logic; attribute dont_touch of G24245: signal is true;
	signal G24246: std_logic; attribute dont_touch of G24246: signal is true;
	signal G24247: std_logic; attribute dont_touch of G24247: signal is true;
	signal G24248: std_logic; attribute dont_touch of G24248: signal is true;
	signal G24249: std_logic; attribute dont_touch of G24249: signal is true;
	signal G24250: std_logic; attribute dont_touch of G24250: signal is true;
	signal G24251: std_logic; attribute dont_touch of G24251: signal is true;
	signal G24252: std_logic; attribute dont_touch of G24252: signal is true;
	signal G24253: std_logic; attribute dont_touch of G24253: signal is true;
	signal G24254: std_logic; attribute dont_touch of G24254: signal is true;
	signal G24255: std_logic; attribute dont_touch of G24255: signal is true;
	signal G24256: std_logic; attribute dont_touch of G24256: signal is true;
	signal G24257: std_logic; attribute dont_touch of G24257: signal is true;
	signal G24258: std_logic; attribute dont_touch of G24258: signal is true;
	signal G24259: std_logic; attribute dont_touch of G24259: signal is true;
	signal G24260: std_logic; attribute dont_touch of G24260: signal is true;
	signal G24261: std_logic; attribute dont_touch of G24261: signal is true;
	signal G24262: std_logic; attribute dont_touch of G24262: signal is true;
	signal G24263: std_logic; attribute dont_touch of G24263: signal is true;
	signal G24264: std_logic; attribute dont_touch of G24264: signal is true;
	signal G24265: std_logic; attribute dont_touch of G24265: signal is true;
	signal G24266: std_logic; attribute dont_touch of G24266: signal is true;
	signal G24267: std_logic; attribute dont_touch of G24267: signal is true;
	signal G24268: std_logic; attribute dont_touch of G24268: signal is true;
	signal G24269: std_logic; attribute dont_touch of G24269: signal is true;
	signal G24270: std_logic; attribute dont_touch of G24270: signal is true;
	signal G24271: std_logic; attribute dont_touch of G24271: signal is true;
	signal G24272: std_logic; attribute dont_touch of G24272: signal is true;
	signal G24273: std_logic; attribute dont_touch of G24273: signal is true;
	signal G24274: std_logic; attribute dont_touch of G24274: signal is true;
	signal G24275: std_logic; attribute dont_touch of G24275: signal is true;
	signal G24276: std_logic; attribute dont_touch of G24276: signal is true;
	signal G24277: std_logic; attribute dont_touch of G24277: signal is true;
	signal G24278: std_logic; attribute dont_touch of G24278: signal is true;
	signal G24279: std_logic; attribute dont_touch of G24279: signal is true;
	signal G24280: std_logic; attribute dont_touch of G24280: signal is true;
	signal G24281: std_logic; attribute dont_touch of G24281: signal is true;
	signal G24282: std_logic; attribute dont_touch of G24282: signal is true;
	signal G24283: std_logic; attribute dont_touch of G24283: signal is true;
	signal G24284: std_logic; attribute dont_touch of G24284: signal is true;
	signal G24285: std_logic; attribute dont_touch of G24285: signal is true;
	signal G24286: std_logic; attribute dont_touch of G24286: signal is true;
	signal G24287: std_logic; attribute dont_touch of G24287: signal is true;
	signal G24288: std_logic; attribute dont_touch of G24288: signal is true;
	signal G24289: std_logic; attribute dont_touch of G24289: signal is true;
	signal G24290: std_logic; attribute dont_touch of G24290: signal is true;
	signal G24291: std_logic; attribute dont_touch of G24291: signal is true;
	signal G24292: std_logic; attribute dont_touch of G24292: signal is true;
	signal G24293: std_logic; attribute dont_touch of G24293: signal is true;
	signal G24294: std_logic; attribute dont_touch of G24294: signal is true;
	signal G24295: std_logic; attribute dont_touch of G24295: signal is true;
	signal G24296: std_logic; attribute dont_touch of G24296: signal is true;
	signal G24297: std_logic; attribute dont_touch of G24297: signal is true;
	signal G24298: std_logic; attribute dont_touch of G24298: signal is true;
	signal G24299: std_logic; attribute dont_touch of G24299: signal is true;
	signal G24300: std_logic; attribute dont_touch of G24300: signal is true;
	signal G24301: std_logic; attribute dont_touch of G24301: signal is true;
	signal G24302: std_logic; attribute dont_touch of G24302: signal is true;
	signal G24303: std_logic; attribute dont_touch of G24303: signal is true;
	signal G24304: std_logic; attribute dont_touch of G24304: signal is true;
	signal G24305: std_logic; attribute dont_touch of G24305: signal is true;
	signal G24306: std_logic; attribute dont_touch of G24306: signal is true;
	signal G24307: std_logic; attribute dont_touch of G24307: signal is true;
	signal G24308: std_logic; attribute dont_touch of G24308: signal is true;
	signal G24309: std_logic; attribute dont_touch of G24309: signal is true;
	signal G24310: std_logic; attribute dont_touch of G24310: signal is true;
	signal G24311: std_logic; attribute dont_touch of G24311: signal is true;
	signal G24312: std_logic; attribute dont_touch of G24312: signal is true;
	signal G24313: std_logic; attribute dont_touch of G24313: signal is true;
	signal G24314: std_logic; attribute dont_touch of G24314: signal is true;
	signal G24315: std_logic; attribute dont_touch of G24315: signal is true;
	signal G24316: std_logic; attribute dont_touch of G24316: signal is true;
	signal G24317: std_logic; attribute dont_touch of G24317: signal is true;
	signal G24318: std_logic; attribute dont_touch of G24318: signal is true;
	signal G24319: std_logic; attribute dont_touch of G24319: signal is true;
	signal G24320: std_logic; attribute dont_touch of G24320: signal is true;
	signal G24321: std_logic; attribute dont_touch of G24321: signal is true;
	signal G24322: std_logic; attribute dont_touch of G24322: signal is true;
	signal G24323: std_logic; attribute dont_touch of G24323: signal is true;
	signal G24324: std_logic; attribute dont_touch of G24324: signal is true;
	signal G24325: std_logic; attribute dont_touch of G24325: signal is true;
	signal G24326: std_logic; attribute dont_touch of G24326: signal is true;
	signal G24327: std_logic; attribute dont_touch of G24327: signal is true;
	signal G24328: std_logic; attribute dont_touch of G24328: signal is true;
	signal G24329: std_logic; attribute dont_touch of G24329: signal is true;
	signal G24330: std_logic; attribute dont_touch of G24330: signal is true;
	signal G24331: std_logic; attribute dont_touch of G24331: signal is true;
	signal G24332: std_logic; attribute dont_touch of G24332: signal is true;
	signal G24333: std_logic; attribute dont_touch of G24333: signal is true;
	signal G24334: std_logic; attribute dont_touch of G24334: signal is true;
	signal G24335: std_logic; attribute dont_touch of G24335: signal is true;
	signal G24336: std_logic; attribute dont_touch of G24336: signal is true;
	signal G24337: std_logic; attribute dont_touch of G24337: signal is true;
	signal G24338: std_logic; attribute dont_touch of G24338: signal is true;
	signal G24339: std_logic; attribute dont_touch of G24339: signal is true;
	signal G24340: std_logic; attribute dont_touch of G24340: signal is true;
	signal G24341: std_logic; attribute dont_touch of G24341: signal is true;
	signal G24342: std_logic; attribute dont_touch of G24342: signal is true;
	signal G24343: std_logic; attribute dont_touch of G24343: signal is true;
	signal G24344: std_logic; attribute dont_touch of G24344: signal is true;
	signal G24345: std_logic; attribute dont_touch of G24345: signal is true;
	signal G24346: std_logic; attribute dont_touch of G24346: signal is true;
	signal G24347: std_logic; attribute dont_touch of G24347: signal is true;
	signal G24348: std_logic; attribute dont_touch of G24348: signal is true;
	signal G24349: std_logic; attribute dont_touch of G24349: signal is true;
	signal G24350: std_logic; attribute dont_touch of G24350: signal is true;
	signal G24351: std_logic; attribute dont_touch of G24351: signal is true;
	signal G24352: std_logic; attribute dont_touch of G24352: signal is true;
	signal G24353: std_logic; attribute dont_touch of G24353: signal is true;
	signal G24354: std_logic; attribute dont_touch of G24354: signal is true;
	signal G24355: std_logic; attribute dont_touch of G24355: signal is true;
	signal G24356: std_logic; attribute dont_touch of G24356: signal is true;
	signal G24357: std_logic; attribute dont_touch of G24357: signal is true;
	signal G24358: std_logic; attribute dont_touch of G24358: signal is true;
	signal G24359: std_logic; attribute dont_touch of G24359: signal is true;
	signal G24360: std_logic; attribute dont_touch of G24360: signal is true;
	signal G24361: std_logic; attribute dont_touch of G24361: signal is true;
	signal G24362: std_logic; attribute dont_touch of G24362: signal is true;
	signal G24363: std_logic; attribute dont_touch of G24363: signal is true;
	signal G24364: std_logic; attribute dont_touch of G24364: signal is true;
	signal G24365: std_logic; attribute dont_touch of G24365: signal is true;
	signal G24366: std_logic; attribute dont_touch of G24366: signal is true;
	signal G24367: std_logic; attribute dont_touch of G24367: signal is true;
	signal G24368: std_logic; attribute dont_touch of G24368: signal is true;
	signal G24369: std_logic; attribute dont_touch of G24369: signal is true;
	signal G24372: std_logic; attribute dont_touch of G24372: signal is true;
	signal G24373: std_logic; attribute dont_touch of G24373: signal is true;
	signal G24374: std_logic; attribute dont_touch of G24374: signal is true;
	signal G24375: std_logic; attribute dont_touch of G24375: signal is true;
	signal G24376: std_logic; attribute dont_touch of G24376: signal is true;
	signal G24377: std_logic; attribute dont_touch of G24377: signal is true;
	signal G24378: std_logic; attribute dont_touch of G24378: signal is true;
	signal G24379: std_logic; attribute dont_touch of G24379: signal is true;
	signal G24380: std_logic; attribute dont_touch of G24380: signal is true;
	signal G24383: std_logic; attribute dont_touch of G24383: signal is true;
	signal G24384: std_logic; attribute dont_touch of G24384: signal is true;
	signal G24385: std_logic; attribute dont_touch of G24385: signal is true;
	signal G24386: std_logic; attribute dont_touch of G24386: signal is true;
	signal G24387: std_logic; attribute dont_touch of G24387: signal is true;
	signal G24388: std_logic; attribute dont_touch of G24388: signal is true;
	signal G24389: std_logic; attribute dont_touch of G24389: signal is true;
	signal G24390: std_logic; attribute dont_touch of G24390: signal is true;
	signal G24391: std_logic; attribute dont_touch of G24391: signal is true;
	signal G24392: std_logic; attribute dont_touch of G24392: signal is true;
	signal G24393: std_logic; attribute dont_touch of G24393: signal is true;
	signal G24394: std_logic; attribute dont_touch of G24394: signal is true;
	signal G24395: std_logic; attribute dont_touch of G24395: signal is true;
	signal G24396: std_logic; attribute dont_touch of G24396: signal is true;
	signal G24397: std_logic; attribute dont_touch of G24397: signal is true;
	signal G24398: std_logic; attribute dont_touch of G24398: signal is true;
	signal G24399: std_logic; attribute dont_touch of G24399: signal is true;
	signal G24400: std_logic; attribute dont_touch of G24400: signal is true;
	signal G24401: std_logic; attribute dont_touch of G24401: signal is true;
	signal G24402: std_logic; attribute dont_touch of G24402: signal is true;
	signal G24403: std_logic; attribute dont_touch of G24403: signal is true;
	signal G24404: std_logic; attribute dont_touch of G24404: signal is true;
	signal G24405: std_logic; attribute dont_touch of G24405: signal is true;
	signal G24406: std_logic; attribute dont_touch of G24406: signal is true;
	signal G24407: std_logic; attribute dont_touch of G24407: signal is true;
	signal G24408: std_logic; attribute dont_touch of G24408: signal is true;
	signal G24409: std_logic; attribute dont_touch of G24409: signal is true;
	signal G24410: std_logic; attribute dont_touch of G24410: signal is true;
	signal G24411: std_logic; attribute dont_touch of G24411: signal is true;
	signal G24415: std_logic; attribute dont_touch of G24415: signal is true;
	signal G24416: std_logic; attribute dont_touch of G24416: signal is true;
	signal G24417: std_logic; attribute dont_touch of G24417: signal is true;
	signal G24418: std_logic; attribute dont_touch of G24418: signal is true;
	signal G24419: std_logic; attribute dont_touch of G24419: signal is true;
	signal G24420: std_logic; attribute dont_touch of G24420: signal is true;
	signal G24421: std_logic; attribute dont_touch of G24421: signal is true;
	signal G24422: std_logic; attribute dont_touch of G24422: signal is true;
	signal G24423: std_logic; attribute dont_touch of G24423: signal is true;
	signal G24424: std_logic; attribute dont_touch of G24424: signal is true;
	signal G24425: std_logic; attribute dont_touch of G24425: signal is true;
	signal G24426: std_logic; attribute dont_touch of G24426: signal is true;
	signal G24427: std_logic; attribute dont_touch of G24427: signal is true;
	signal G24428: std_logic; attribute dont_touch of G24428: signal is true;
	signal G24429: std_logic; attribute dont_touch of G24429: signal is true;
	signal G24430: std_logic; attribute dont_touch of G24430: signal is true;
	signal G24431: std_logic; attribute dont_touch of G24431: signal is true;
	signal G24432: std_logic; attribute dont_touch of G24432: signal is true;
	signal G24433: std_logic; attribute dont_touch of G24433: signal is true;
	signal G24436: std_logic; attribute dont_touch of G24436: signal is true;
	signal G24437: std_logic; attribute dont_touch of G24437: signal is true;
	signal G24438: std_logic; attribute dont_touch of G24438: signal is true;
	signal G24439: std_logic; attribute dont_touch of G24439: signal is true;
	signal G24443: std_logic; attribute dont_touch of G24443: signal is true;
	signal G24444: std_logic; attribute dont_touch of G24444: signal is true;
	signal G24447: std_logic; attribute dont_touch of G24447: signal is true;
	signal G24450: std_logic; attribute dont_touch of G24450: signal is true;
	signal G24451: std_logic; attribute dont_touch of G24451: signal is true;
	signal G24452: std_logic; attribute dont_touch of G24452: signal is true;
	signal G24453: std_logic; attribute dont_touch of G24453: signal is true;
	signal G24457: std_logic; attribute dont_touch of G24457: signal is true;
	signal G24460: std_logic; attribute dont_touch of G24460: signal is true;
	signal G24463: std_logic; attribute dont_touch of G24463: signal is true;
	signal G24464: std_logic; attribute dont_touch of G24464: signal is true;
	signal G24465: std_logic; attribute dont_touch of G24465: signal is true;
	signal G24466: std_logic; attribute dont_touch of G24466: signal is true;
	signal G24467: std_logic; attribute dont_touch of G24467: signal is true;
	signal G24468: std_logic; attribute dont_touch of G24468: signal is true;
	signal G24471: std_logic; attribute dont_touch of G24471: signal is true;
	signal G24474: std_logic; attribute dont_touch of G24474: signal is true;
	signal G24475: std_logic; attribute dont_touch of G24475: signal is true;
	signal G24476: std_logic; attribute dont_touch of G24476: signal is true;
	signal G24477: std_logic; attribute dont_touch of G24477: signal is true;
	signal G24478: std_logic; attribute dont_touch of G24478: signal is true;
	signal G24481: std_logic; attribute dont_touch of G24481: signal is true;
	signal G24482: std_logic; attribute dont_touch of G24482: signal is true;
	signal G24483: std_logic; attribute dont_touch of G24483: signal is true;
	signal G24484: std_logic; attribute dont_touch of G24484: signal is true;
	signal G24485: std_logic; attribute dont_touch of G24485: signal is true;
	signal G24488: std_logic; attribute dont_touch of G24488: signal is true;
	signal G24489: std_logic; attribute dont_touch of G24489: signal is true;
	signal G24490: std_logic; attribute dont_touch of G24490: signal is true;
	signal G24491: std_logic; attribute dont_touch of G24491: signal is true;
	signal G24494: std_logic; attribute dont_touch of G24494: signal is true;
	signal G24495: std_logic; attribute dont_touch of G24495: signal is true;
	signal G24496: std_logic; attribute dont_touch of G24496: signal is true;
	signal G24497: std_logic; attribute dont_touch of G24497: signal is true;
	signal G24498: std_logic; attribute dont_touch of G24498: signal is true;
	signal G24499: std_logic; attribute dont_touch of G24499: signal is true;
	signal G24500: std_logic; attribute dont_touch of G24500: signal is true;
	signal G24501: std_logic; attribute dont_touch of G24501: signal is true;
	signal G24502: std_logic; attribute dont_touch of G24502: signal is true;
	signal G24503: std_logic; attribute dont_touch of G24503: signal is true;
	signal G24504: std_logic; attribute dont_touch of G24504: signal is true;
	signal G24505: std_logic; attribute dont_touch of G24505: signal is true;
	signal G24506: std_logic; attribute dont_touch of G24506: signal is true;
	signal G24507: std_logic; attribute dont_touch of G24507: signal is true;
	signal G24508: std_logic; attribute dont_touch of G24508: signal is true;
	signal G24509: std_logic; attribute dont_touch of G24509: signal is true;
	signal G24510: std_logic; attribute dont_touch of G24510: signal is true;
	signal G24514: std_logic; attribute dont_touch of G24514: signal is true;
	signal G24515: std_logic; attribute dont_touch of G24515: signal is true;
	signal G24516: std_logic; attribute dont_touch of G24516: signal is true;
	signal G24517: std_logic; attribute dont_touch of G24517: signal is true;
	signal G24518: std_logic; attribute dont_touch of G24518: signal is true;
	signal G24522: std_logic; attribute dont_touch of G24522: signal is true;
	signal G24523: std_logic; attribute dont_touch of G24523: signal is true;
	signal G24524: std_logic; attribute dont_touch of G24524: signal is true;
	signal G24525: std_logic; attribute dont_touch of G24525: signal is true;
	signal G24526: std_logic; attribute dont_touch of G24526: signal is true;
	signal G24527: std_logic; attribute dont_touch of G24527: signal is true;
	signal G24528: std_logic; attribute dont_touch of G24528: signal is true;
	signal G24532: std_logic; attribute dont_touch of G24532: signal is true;
	signal G24533: std_logic; attribute dont_touch of G24533: signal is true;
	signal G24534: std_logic; attribute dont_touch of G24534: signal is true;
	signal G24535: std_logic; attribute dont_touch of G24535: signal is true;
	signal G24536: std_logic; attribute dont_touch of G24536: signal is true;
	signal G24537: std_logic; attribute dont_touch of G24537: signal is true;
	signal G24540: std_logic; attribute dont_touch of G24540: signal is true;
	signal G24541: std_logic; attribute dont_touch of G24541: signal is true;
	signal G24544: std_logic; attribute dont_touch of G24544: signal is true;
	signal G24545: std_logic; attribute dont_touch of G24545: signal is true;
	signal G24546: std_logic; attribute dont_touch of G24546: signal is true;
	signal G24547: std_logic; attribute dont_touch of G24547: signal is true;
	signal G24548: std_logic; attribute dont_touch of G24548: signal is true;
	signal G24549: std_logic; attribute dont_touch of G24549: signal is true;
	signal G24550: std_logic; attribute dont_touch of G24550: signal is true;
	signal G24551: std_logic; attribute dont_touch of G24551: signal is true;
	signal G24552: std_logic; attribute dont_touch of G24552: signal is true;
	signal G24553: std_logic; attribute dont_touch of G24553: signal is true;
	signal G24554: std_logic; attribute dont_touch of G24554: signal is true;
	signal G24555: std_logic; attribute dont_touch of G24555: signal is true;
	signal G24556: std_logic; attribute dont_touch of G24556: signal is true;
	signal G24557: std_logic; attribute dont_touch of G24557: signal is true;
	signal G24558: std_logic; attribute dont_touch of G24558: signal is true;
	signal G24559: std_logic; attribute dont_touch of G24559: signal is true;
	signal G24560: std_logic; attribute dont_touch of G24560: signal is true;
	signal G24561: std_logic; attribute dont_touch of G24561: signal is true;
	signal G24564: std_logic; attribute dont_touch of G24564: signal is true;
	signal G24565: std_logic; attribute dont_touch of G24565: signal is true;
	signal G24566: std_logic; attribute dont_touch of G24566: signal is true;
	signal G24567: std_logic; attribute dont_touch of G24567: signal is true;
	signal G24568: std_logic; attribute dont_touch of G24568: signal is true;
	signal G24569: std_logic; attribute dont_touch of G24569: signal is true;
	signal G24570: std_logic; attribute dont_touch of G24570: signal is true;
	signal G24571: std_logic; attribute dont_touch of G24571: signal is true;
	signal G24572: std_logic; attribute dont_touch of G24572: signal is true;
	signal G24573: std_logic; attribute dont_touch of G24573: signal is true;
	signal G24574: std_logic; attribute dont_touch of G24574: signal is true;
	signal G24575: std_logic; attribute dont_touch of G24575: signal is true;
	signal G24576: std_logic; attribute dont_touch of G24576: signal is true;
	signal G24577: std_logic; attribute dont_touch of G24577: signal is true;
	signal G24578: std_logic; attribute dont_touch of G24578: signal is true;
	signal G24579: std_logic; attribute dont_touch of G24579: signal is true;
	signal G24580: std_logic; attribute dont_touch of G24580: signal is true;
	signal G24581: std_logic; attribute dont_touch of G24581: signal is true;
	signal G24582: std_logic; attribute dont_touch of G24582: signal is true;
	signal G24583: std_logic; attribute dont_touch of G24583: signal is true;
	signal G24584: std_logic; attribute dont_touch of G24584: signal is true;
	signal G24585: std_logic; attribute dont_touch of G24585: signal is true;
	signal G24586: std_logic; attribute dont_touch of G24586: signal is true;
	signal G24587: std_logic; attribute dont_touch of G24587: signal is true;
	signal G24588: std_logic; attribute dont_touch of G24588: signal is true;
	signal G24589: std_logic; attribute dont_touch of G24589: signal is true;
	signal G24590: std_logic; attribute dont_touch of G24590: signal is true;
	signal G24591: std_logic; attribute dont_touch of G24591: signal is true;
	signal G24600: std_logic; attribute dont_touch of G24600: signal is true;
	signal G24601: std_logic; attribute dont_touch of G24601: signal is true;
	signal G24602: std_logic; attribute dont_touch of G24602: signal is true;
	signal G24603: std_logic; attribute dont_touch of G24603: signal is true;
	signal G24604: std_logic; attribute dont_touch of G24604: signal is true;
	signal G24605: std_logic; attribute dont_touch of G24605: signal is true;
	signal G24606: std_logic; attribute dont_touch of G24606: signal is true;
	signal G24607: std_logic; attribute dont_touch of G24607: signal is true;
	signal G24608: std_logic; attribute dont_touch of G24608: signal is true;
	signal G24609: std_logic; attribute dont_touch of G24609: signal is true;
	signal G24618: std_logic; attribute dont_touch of G24618: signal is true;
	signal G24619: std_logic; attribute dont_touch of G24619: signal is true;
	signal G24620: std_logic; attribute dont_touch of G24620: signal is true;
	signal G24621: std_logic; attribute dont_touch of G24621: signal is true;
	signal G24622: std_logic; attribute dont_touch of G24622: signal is true;
	signal G24623: std_logic; attribute dont_touch of G24623: signal is true;
	signal G24624: std_logic; attribute dont_touch of G24624: signal is true;
	signal G24625: std_logic; attribute dont_touch of G24625: signal is true;
	signal G24626: std_logic; attribute dont_touch of G24626: signal is true;
	signal G24627: std_logic; attribute dont_touch of G24627: signal is true;
	signal G24628: std_logic; attribute dont_touch of G24628: signal is true;
	signal G24629: std_logic; attribute dont_touch of G24629: signal is true;
	signal G24630: std_logic; attribute dont_touch of G24630: signal is true;
	signal G24631: std_logic; attribute dont_touch of G24631: signal is true;
	signal G24634: std_logic; attribute dont_touch of G24634: signal is true;
	signal G24635: std_logic; attribute dont_touch of G24635: signal is true;
	signal G24636: std_logic; attribute dont_touch of G24636: signal is true;
	signal G24637: std_logic; attribute dont_touch of G24637: signal is true;
	signal G24638: std_logic; attribute dont_touch of G24638: signal is true;
	signal G24639: std_logic; attribute dont_touch of G24639: signal is true;
	signal G24640: std_logic; attribute dont_touch of G24640: signal is true;
	signal G24641: std_logic; attribute dont_touch of G24641: signal is true;
	signal G24642: std_logic; attribute dont_touch of G24642: signal is true;
	signal G24643: std_logic; attribute dont_touch of G24643: signal is true;
	signal G24644: std_logic; attribute dont_touch of G24644: signal is true;
	signal G24645: std_logic; attribute dont_touch of G24645: signal is true;
	signal G24646: std_logic; attribute dont_touch of G24646: signal is true;
	signal G24647: std_logic; attribute dont_touch of G24647: signal is true;
	signal G24648: std_logic; attribute dont_touch of G24648: signal is true;
	signal G24649: std_logic; attribute dont_touch of G24649: signal is true;
	signal G24650: std_logic; attribute dont_touch of G24650: signal is true;
	signal G24651: std_logic; attribute dont_touch of G24651: signal is true;
	signal G24652: std_logic; attribute dont_touch of G24652: signal is true;
	signal G24653: std_logic; attribute dont_touch of G24653: signal is true;
	signal G24654: std_logic; attribute dont_touch of G24654: signal is true;
	signal G24655: std_logic; attribute dont_touch of G24655: signal is true;
	signal G24656: std_logic; attribute dont_touch of G24656: signal is true;
	signal G24657: std_logic; attribute dont_touch of G24657: signal is true;
	signal G24658: std_logic; attribute dont_touch of G24658: signal is true;
	signal G24659: std_logic; attribute dont_touch of G24659: signal is true;
	signal G24660: std_logic; attribute dont_touch of G24660: signal is true;
	signal G24661: std_logic; attribute dont_touch of G24661: signal is true;
	signal G24662: std_logic; attribute dont_touch of G24662: signal is true;
	signal G24663: std_logic; attribute dont_touch of G24663: signal is true;
	signal G24664: std_logic; attribute dont_touch of G24664: signal is true;
	signal G24665: std_logic; attribute dont_touch of G24665: signal is true;
	signal G24666: std_logic; attribute dont_touch of G24666: signal is true;
	signal G24667: std_logic; attribute dont_touch of G24667: signal is true;
	signal G24668: std_logic; attribute dont_touch of G24668: signal is true;
	signal G24669: std_logic; attribute dont_touch of G24669: signal is true;
	signal G24670: std_logic; attribute dont_touch of G24670: signal is true;
	signal G24671: std_logic; attribute dont_touch of G24671: signal is true;
	signal G24672: std_logic; attribute dont_touch of G24672: signal is true;
	signal G24673: std_logic; attribute dont_touch of G24673: signal is true;
	signal G24674: std_logic; attribute dont_touch of G24674: signal is true;
	signal G24675: std_logic; attribute dont_touch of G24675: signal is true;
	signal G24676: std_logic; attribute dont_touch of G24676: signal is true;
	signal G24677: std_logic; attribute dont_touch of G24677: signal is true;
	signal G24678: std_logic; attribute dont_touch of G24678: signal is true;
	signal G24679: std_logic; attribute dont_touch of G24679: signal is true;
	signal G24680: std_logic; attribute dont_touch of G24680: signal is true;
	signal G24681: std_logic; attribute dont_touch of G24681: signal is true;
	signal G24682: std_logic; attribute dont_touch of G24682: signal is true;
	signal G24683: std_logic; attribute dont_touch of G24683: signal is true;
	signal G24684: std_logic; attribute dont_touch of G24684: signal is true;
	signal G24685: std_logic; attribute dont_touch of G24685: signal is true;
	signal G24686: std_logic; attribute dont_touch of G24686: signal is true;
	signal G24687: std_logic; attribute dont_touch of G24687: signal is true;
	signal G24688: std_logic; attribute dont_touch of G24688: signal is true;
	signal G24698: std_logic; attribute dont_touch of G24698: signal is true;
	signal G24699: std_logic; attribute dont_touch of G24699: signal is true;
	signal G24700: std_logic; attribute dont_touch of G24700: signal is true;
	signal G24701: std_logic; attribute dont_touch of G24701: signal is true;
	signal G24702: std_logic; attribute dont_touch of G24702: signal is true;
	signal G24703: std_logic; attribute dont_touch of G24703: signal is true;
	signal G24704: std_logic; attribute dont_touch of G24704: signal is true;
	signal G24705: std_logic; attribute dont_touch of G24705: signal is true;
	signal G24706: std_logic; attribute dont_touch of G24706: signal is true;
	signal G24707: std_logic; attribute dont_touch of G24707: signal is true;
	signal G24708: std_logic; attribute dont_touch of G24708: signal is true;
	signal G24709: std_logic; attribute dont_touch of G24709: signal is true;
	signal G24710: std_logic; attribute dont_touch of G24710: signal is true;
	signal G24711: std_logic; attribute dont_touch of G24711: signal is true;
	signal G24712: std_logic; attribute dont_touch of G24712: signal is true;
	signal G24713: std_logic; attribute dont_touch of G24713: signal is true;
	signal G24714: std_logic; attribute dont_touch of G24714: signal is true;
	signal G24715: std_logic; attribute dont_touch of G24715: signal is true;
	signal G24716: std_logic; attribute dont_touch of G24716: signal is true;
	signal G24717: std_logic; attribute dont_touch of G24717: signal is true;
	signal G24718: std_logic; attribute dont_touch of G24718: signal is true;
	signal G24719: std_logic; attribute dont_touch of G24719: signal is true;
	signal G24720: std_logic; attribute dont_touch of G24720: signal is true;
	signal G24721: std_logic; attribute dont_touch of G24721: signal is true;
	signal G24722: std_logic; attribute dont_touch of G24722: signal is true;
	signal G24723: std_logic; attribute dont_touch of G24723: signal is true;
	signal G24724: std_logic; attribute dont_touch of G24724: signal is true;
	signal G24725: std_logic; attribute dont_touch of G24725: signal is true;
	signal G24726: std_logic; attribute dont_touch of G24726: signal is true;
	signal G24727: std_logic; attribute dont_touch of G24727: signal is true;
	signal G24728: std_logic; attribute dont_touch of G24728: signal is true;
	signal G24729: std_logic; attribute dont_touch of G24729: signal is true;
	signal G24730: std_logic; attribute dont_touch of G24730: signal is true;
	signal G24731: std_logic; attribute dont_touch of G24731: signal is true;
	signal G24732: std_logic; attribute dont_touch of G24732: signal is true;
	signal G24743: std_logic; attribute dont_touch of G24743: signal is true;
	signal G24744: std_logic; attribute dont_touch of G24744: signal is true;
	signal G24745: std_logic; attribute dont_touch of G24745: signal is true;
	signal G24746: std_logic; attribute dont_touch of G24746: signal is true;
	signal G24747: std_logic; attribute dont_touch of G24747: signal is true;
	signal G24748: std_logic; attribute dont_touch of G24748: signal is true;
	signal G24749: std_logic; attribute dont_touch of G24749: signal is true;
	signal G24750: std_logic; attribute dont_touch of G24750: signal is true;
	signal G24751: std_logic; attribute dont_touch of G24751: signal is true;
	signal G24754: std_logic; attribute dont_touch of G24754: signal is true;
	signal G24755: std_logic; attribute dont_touch of G24755: signal is true;
	signal G24756: std_logic; attribute dont_touch of G24756: signal is true;
	signal G24757: std_logic; attribute dont_touch of G24757: signal is true;
	signal G24758: std_logic; attribute dont_touch of G24758: signal is true;
	signal G24759: std_logic; attribute dont_touch of G24759: signal is true;
	signal G24760: std_logic; attribute dont_touch of G24760: signal is true;
	signal G24761: std_logic; attribute dont_touch of G24761: signal is true;
	signal G24762: std_logic; attribute dont_touch of G24762: signal is true;
	signal G24763: std_logic; attribute dont_touch of G24763: signal is true;
	signal G24764: std_logic; attribute dont_touch of G24764: signal is true;
	signal G24765: std_logic; attribute dont_touch of G24765: signal is true;
	signal G24766: std_logic; attribute dont_touch of G24766: signal is true;
	signal G24769: std_logic; attribute dont_touch of G24769: signal is true;
	signal G24770: std_logic; attribute dont_touch of G24770: signal is true;
	signal G24771: std_logic; attribute dont_touch of G24771: signal is true;
	signal G24772: std_logic; attribute dont_touch of G24772: signal is true;
	signal G24773: std_logic; attribute dont_touch of G24773: signal is true;
	signal G24774: std_logic; attribute dont_touch of G24774: signal is true;
	signal G24775: std_logic; attribute dont_touch of G24775: signal is true;
	signal G24776: std_logic; attribute dont_touch of G24776: signal is true;
	signal G24777: std_logic; attribute dont_touch of G24777: signal is true;
	signal G24778: std_logic; attribute dont_touch of G24778: signal is true;
	signal G24779: std_logic; attribute dont_touch of G24779: signal is true;
	signal G24782: std_logic; attribute dont_touch of G24782: signal is true;
	signal G24785: std_logic; attribute dont_touch of G24785: signal is true;
	signal G24786: std_logic; attribute dont_touch of G24786: signal is true;
	signal G24787: std_logic; attribute dont_touch of G24787: signal is true;
	signal G24788: std_logic; attribute dont_touch of G24788: signal is true;
	signal G24789: std_logic; attribute dont_touch of G24789: signal is true;
	signal G24790: std_logic; attribute dont_touch of G24790: signal is true;
	signal G24791: std_logic; attribute dont_touch of G24791: signal is true;
	signal G24792: std_logic; attribute dont_touch of G24792: signal is true;
	signal G24793: std_logic; attribute dont_touch of G24793: signal is true;
	signal G24794: std_logic; attribute dont_touch of G24794: signal is true;
	signal G24795: std_logic; attribute dont_touch of G24795: signal is true;
	signal G24796: std_logic; attribute dont_touch of G24796: signal is true;
	signal G24797: std_logic; attribute dont_touch of G24797: signal is true;
	signal G24798: std_logic; attribute dont_touch of G24798: signal is true;
	signal G24799: std_logic; attribute dont_touch of G24799: signal is true;
	signal G24802: std_logic; attribute dont_touch of G24802: signal is true;
	signal G24803: std_logic; attribute dont_touch of G24803: signal is true;
	signal G24804: std_logic; attribute dont_touch of G24804: signal is true;
	signal G24807: std_logic; attribute dont_touch of G24807: signal is true;
	signal G24808: std_logic; attribute dont_touch of G24808: signal is true;
	signal G24809: std_logic; attribute dont_touch of G24809: signal is true;
	signal G24812: std_logic; attribute dont_touch of G24812: signal is true;
	signal G24813: std_logic; attribute dont_touch of G24813: signal is true;
	signal G24814: std_logic; attribute dont_touch of G24814: signal is true;
	signal G24817: std_logic; attribute dont_touch of G24817: signal is true;
	signal G24818: std_logic; attribute dont_touch of G24818: signal is true;
	signal G24819: std_logic; attribute dont_touch of G24819: signal is true;
	signal G24820: std_logic; attribute dont_touch of G24820: signal is true;
	signal G24821: std_logic; attribute dont_touch of G24821: signal is true;
	signal G24822: std_logic; attribute dont_touch of G24822: signal is true;
	signal G24825: std_logic; attribute dont_touch of G24825: signal is true;
	signal G24835: std_logic; attribute dont_touch of G24835: signal is true;
	signal G24836: std_logic; attribute dont_touch of G24836: signal is true;
	signal G24839: std_logic; attribute dont_touch of G24839: signal is true;
	signal G24840: std_logic; attribute dont_touch of G24840: signal is true;
	signal G24841: std_logic; attribute dont_touch of G24841: signal is true;
	signal G24842: std_logic; attribute dont_touch of G24842: signal is true;
	signal G24843: std_logic; attribute dont_touch of G24843: signal is true;
	signal G24846: std_logic; attribute dont_touch of G24846: signal is true;
	signal G24849: std_logic; attribute dont_touch of G24849: signal is true;
	signal G24850: std_logic; attribute dont_touch of G24850: signal is true;
	signal G24853: std_logic; attribute dont_touch of G24853: signal is true;
	signal G24854: std_logic; attribute dont_touch of G24854: signal is true;
	signal G24855: std_logic; attribute dont_touch of G24855: signal is true;
	signal G24858: std_logic; attribute dont_touch of G24858: signal is true;
	signal G24861: std_logic; attribute dont_touch of G24861: signal is true;
	signal G24864: std_logic; attribute dont_touch of G24864: signal is true;
	signal G24865: std_logic; attribute dont_touch of G24865: signal is true;
	signal G24866: std_logic; attribute dont_touch of G24866: signal is true;
	signal G24869: std_logic; attribute dont_touch of G24869: signal is true;
	signal G24872: std_logic; attribute dont_touch of G24872: signal is true;
	signal G24875: std_logic; attribute dont_touch of G24875: signal is true;
	signal G24879: std_logic; attribute dont_touch of G24879: signal is true;
	signal G24880: std_logic; attribute dont_touch of G24880: signal is true;
	signal G24881: std_logic; attribute dont_touch of G24881: signal is true;
	signal G24884: std_logic; attribute dont_touch of G24884: signal is true;
	signal G24887: std_logic; attribute dont_touch of G24887: signal is true;
	signal G24890: std_logic; attribute dont_touch of G24890: signal is true;
	signal G24891: std_logic; attribute dont_touch of G24891: signal is true;
	signal G24892: std_logic; attribute dont_touch of G24892: signal is true;
	signal G24893: std_logic; attribute dont_touch of G24893: signal is true;
	signal G24896: std_logic; attribute dont_touch of G24896: signal is true;
	signal G24897: std_logic; attribute dont_touch of G24897: signal is true;
	signal G24900: std_logic; attribute dont_touch of G24900: signal is true;
	signal G24903: std_logic; attribute dont_touch of G24903: signal is true;
	signal G24904: std_logic; attribute dont_touch of G24904: signal is true;
	signal G24905: std_logic; attribute dont_touch of G24905: signal is true;
	signal G24906: std_logic; attribute dont_touch of G24906: signal is true;
	signal G24907: std_logic; attribute dont_touch of G24907: signal is true;
	signal G24908: std_logic; attribute dont_touch of G24908: signal is true;
	signal G24911: std_logic; attribute dont_touch of G24911: signal is true;
	signal G24912: std_logic; attribute dont_touch of G24912: signal is true;
	signal G24913: std_logic; attribute dont_touch of G24913: signal is true;
	signal G24914: std_logic; attribute dont_touch of G24914: signal is true;
	signal G24915: std_logic; attribute dont_touch of G24915: signal is true;
	signal G24916: std_logic; attribute dont_touch of G24916: signal is true;
	signal G24917: std_logic; attribute dont_touch of G24917: signal is true;
	signal G24918: std_logic; attribute dont_touch of G24918: signal is true;
	signal G24919: std_logic; attribute dont_touch of G24919: signal is true;
	signal G24920: std_logic; attribute dont_touch of G24920: signal is true;
	signal G24921: std_logic; attribute dont_touch of G24921: signal is true;
	signal G24922: std_logic; attribute dont_touch of G24922: signal is true;
	signal G24923: std_logic; attribute dont_touch of G24923: signal is true;
	signal G24924: std_logic; attribute dont_touch of G24924: signal is true;
	signal G24925: std_logic; attribute dont_touch of G24925: signal is true;
	signal G24926: std_logic; attribute dont_touch of G24926: signal is true;
	signal G24929: std_logic; attribute dont_touch of G24929: signal is true;
	signal G24930: std_logic; attribute dont_touch of G24930: signal is true;
	signal G24931: std_logic; attribute dont_touch of G24931: signal is true;
	signal G24932: std_logic; attribute dont_touch of G24932: signal is true;
	signal G24933: std_logic; attribute dont_touch of G24933: signal is true;
	signal G24934: std_logic; attribute dont_touch of G24934: signal is true;
	signal G24935: std_logic; attribute dont_touch of G24935: signal is true;
	signal G24936: std_logic; attribute dont_touch of G24936: signal is true;
	signal G24939: std_logic; attribute dont_touch of G24939: signal is true;
	signal G24940: std_logic; attribute dont_touch of G24940: signal is true;
	signal G24941: std_logic; attribute dont_touch of G24941: signal is true;
	signal G24942: std_logic; attribute dont_touch of G24942: signal is true;
	signal G24943: std_logic; attribute dont_touch of G24943: signal is true;
	signal G24944: std_logic; attribute dont_touch of G24944: signal is true;
	signal G24945: std_logic; attribute dont_touch of G24945: signal is true;
	signal G24946: std_logic; attribute dont_touch of G24946: signal is true;
	signal G24949: std_logic; attribute dont_touch of G24949: signal is true;
	signal G24950: std_logic; attribute dont_touch of G24950: signal is true;
	signal G24951: std_logic; attribute dont_touch of G24951: signal is true;
	signal G24952: std_logic; attribute dont_touch of G24952: signal is true;
	signal G24953: std_logic; attribute dont_touch of G24953: signal is true;
	signal G24957: std_logic; attribute dont_touch of G24957: signal is true;
	signal G24958: std_logic; attribute dont_touch of G24958: signal is true;
	signal G24959: std_logic; attribute dont_touch of G24959: signal is true;
	signal G24960: std_logic; attribute dont_touch of G24960: signal is true;
	signal G24961: std_logic; attribute dont_touch of G24961: signal is true;
	signal G24962: std_logic; attribute dont_touch of G24962: signal is true;
	signal G24963: std_logic; attribute dont_touch of G24963: signal is true;
	signal G24964: std_logic; attribute dont_touch of G24964: signal is true;
	signal G24965: std_logic; attribute dont_touch of G24965: signal is true;
	signal G24966: std_logic; attribute dont_touch of G24966: signal is true;
	signal G24967: std_logic; attribute dont_touch of G24967: signal is true;
	signal G24968: std_logic; attribute dont_touch of G24968: signal is true;
	signal G24971: std_logic; attribute dont_touch of G24971: signal is true;
	signal G24972: std_logic; attribute dont_touch of G24972: signal is true;
	signal G24973: std_logic; attribute dont_touch of G24973: signal is true;
	signal G24974: std_logic; attribute dont_touch of G24974: signal is true;
	signal G24975: std_logic; attribute dont_touch of G24975: signal is true;
	signal G24976: std_logic; attribute dont_touch of G24976: signal is true;
	signal G24977: std_logic; attribute dont_touch of G24977: signal is true;
	signal G24978: std_logic; attribute dont_touch of G24978: signal is true;
	signal G24979: std_logic; attribute dont_touch of G24979: signal is true;
	signal G24980: std_logic; attribute dont_touch of G24980: signal is true;
	signal G24981: std_logic; attribute dont_touch of G24981: signal is true;
	signal G24982: std_logic; attribute dont_touch of G24982: signal is true;
	signal G24983: std_logic; attribute dont_touch of G24983: signal is true;
	signal G24984: std_logic; attribute dont_touch of G24984: signal is true;
	signal G24985: std_logic; attribute dont_touch of G24985: signal is true;
	signal G24986: std_logic; attribute dont_touch of G24986: signal is true;
	signal G24987: std_logic; attribute dont_touch of G24987: signal is true;
	signal G24988: std_logic; attribute dont_touch of G24988: signal is true;
	signal G24989: std_logic; attribute dont_touch of G24989: signal is true;
	signal G24990: std_logic; attribute dont_touch of G24990: signal is true;
	signal G24991: std_logic; attribute dont_touch of G24991: signal is true;
	signal G24992: std_logic; attribute dont_touch of G24992: signal is true;
	signal G24993: std_logic; attribute dont_touch of G24993: signal is true;
	signal G24994: std_logic; attribute dont_touch of G24994: signal is true;
	signal G24995: std_logic; attribute dont_touch of G24995: signal is true;
	signal G24996: std_logic; attribute dont_touch of G24996: signal is true;
	signal G24997: std_logic; attribute dont_touch of G24997: signal is true;
	signal G24998: std_logic; attribute dont_touch of G24998: signal is true;
	signal G24999: std_logic; attribute dont_touch of G24999: signal is true;
	signal G25000: std_logic; attribute dont_touch of G25000: signal is true;
	signal G25001: std_logic; attribute dont_touch of G25001: signal is true;
	signal G25002: std_logic; attribute dont_touch of G25002: signal is true;
	signal G25003: std_logic; attribute dont_touch of G25003: signal is true;
	signal G25004: std_logic; attribute dont_touch of G25004: signal is true;
	signal G25005: std_logic; attribute dont_touch of G25005: signal is true;
	signal G25006: std_logic; attribute dont_touch of G25006: signal is true;
	signal G25007: std_logic; attribute dont_touch of G25007: signal is true;
	signal G25008: std_logic; attribute dont_touch of G25008: signal is true;
	signal G25009: std_logic; attribute dont_touch of G25009: signal is true;
	signal G25010: std_logic; attribute dont_touch of G25010: signal is true;
	signal G25011: std_logic; attribute dont_touch of G25011: signal is true;
	signal G25012: std_logic; attribute dont_touch of G25012: signal is true;
	signal G25013: std_logic; attribute dont_touch of G25013: signal is true;
	signal G25014: std_logic; attribute dont_touch of G25014: signal is true;
	signal G25015: std_logic; attribute dont_touch of G25015: signal is true;
	signal G25016: std_logic; attribute dont_touch of G25016: signal is true;
	signal G25017: std_logic; attribute dont_touch of G25017: signal is true;
	signal G25018: std_logic; attribute dont_touch of G25018: signal is true;
	signal G25019: std_logic; attribute dont_touch of G25019: signal is true;
	signal G25020: std_logic; attribute dont_touch of G25020: signal is true;
	signal G25021: std_logic; attribute dont_touch of G25021: signal is true;
	signal G25022: std_logic; attribute dont_touch of G25022: signal is true;
	signal G25023: std_logic; attribute dont_touch of G25023: signal is true;
	signal G25024: std_logic; attribute dont_touch of G25024: signal is true;
	signal G25025: std_logic; attribute dont_touch of G25025: signal is true;
	signal G25026: std_logic; attribute dont_touch of G25026: signal is true;
	signal G25027: std_logic; attribute dont_touch of G25027: signal is true;
	signal G25030: std_logic; attribute dont_touch of G25030: signal is true;
	signal G25031: std_logic; attribute dont_touch of G25031: signal is true;
	signal G25032: std_logic; attribute dont_touch of G25032: signal is true;
	signal G25033: std_logic; attribute dont_touch of G25033: signal is true;
	signal G25034: std_logic; attribute dont_touch of G25034: signal is true;
	signal G25035: std_logic; attribute dont_touch of G25035: signal is true;
	signal G25036: std_logic; attribute dont_touch of G25036: signal is true;
	signal G25037: std_logic; attribute dont_touch of G25037: signal is true;
	signal G25038: std_logic; attribute dont_touch of G25038: signal is true;
	signal G25039: std_logic; attribute dont_touch of G25039: signal is true;
	signal G25040: std_logic; attribute dont_touch of G25040: signal is true;
	signal G25041: std_logic; attribute dont_touch of G25041: signal is true;
	signal G25042: std_logic; attribute dont_touch of G25042: signal is true;
	signal G25043: std_logic; attribute dont_touch of G25043: signal is true;
	signal G25044: std_logic; attribute dont_touch of G25044: signal is true;
	signal G25045: std_logic; attribute dont_touch of G25045: signal is true;
	signal G25046: std_logic; attribute dont_touch of G25046: signal is true;
	signal G25047: std_logic; attribute dont_touch of G25047: signal is true;
	signal G25048: std_logic; attribute dont_touch of G25048: signal is true;
	signal G25049: std_logic; attribute dont_touch of G25049: signal is true;
	signal G25050: std_logic; attribute dont_touch of G25050: signal is true;
	signal G25051: std_logic; attribute dont_touch of G25051: signal is true;
	signal G25054: std_logic; attribute dont_touch of G25054: signal is true;
	signal G25055: std_logic; attribute dont_touch of G25055: signal is true;
	signal G25056: std_logic; attribute dont_touch of G25056: signal is true;
	signal G25057: std_logic; attribute dont_touch of G25057: signal is true;
	signal G25058: std_logic; attribute dont_touch of G25058: signal is true;
	signal G25059: std_logic; attribute dont_touch of G25059: signal is true;
	signal G25060: std_logic; attribute dont_touch of G25060: signal is true;
	signal G25061: std_logic; attribute dont_touch of G25061: signal is true;
	signal G25062: std_logic; attribute dont_touch of G25062: signal is true;
	signal G25063: std_logic; attribute dont_touch of G25063: signal is true;
	signal G25064: std_logic; attribute dont_touch of G25064: signal is true;
	signal G25067: std_logic; attribute dont_touch of G25067: signal is true;
	signal G25068: std_logic; attribute dont_touch of G25068: signal is true;
	signal G25069: std_logic; attribute dont_touch of G25069: signal is true;
	signal G25070: std_logic; attribute dont_touch of G25070: signal is true;
	signal G25071: std_logic; attribute dont_touch of G25071: signal is true;
	signal G25072: std_logic; attribute dont_touch of G25072: signal is true;
	signal G25073: std_logic; attribute dont_touch of G25073: signal is true;
	signal G25076: std_logic; attribute dont_touch of G25076: signal is true;
	signal G25077: std_logic; attribute dont_touch of G25077: signal is true;
	signal G25078: std_logic; attribute dont_touch of G25078: signal is true;
	signal G25079: std_logic; attribute dont_touch of G25079: signal is true;
	signal G25080: std_logic; attribute dont_touch of G25080: signal is true;
	signal G25081: std_logic; attribute dont_touch of G25081: signal is true;
	signal G25082: std_logic; attribute dont_touch of G25082: signal is true;
	signal G25083: std_logic; attribute dont_touch of G25083: signal is true;
	signal G25084: std_logic; attribute dont_touch of G25084: signal is true;
	signal G25085: std_logic; attribute dont_touch of G25085: signal is true;
	signal G25086: std_logic; attribute dont_touch of G25086: signal is true;
	signal G25087: std_logic; attribute dont_touch of G25087: signal is true;
	signal G25088: std_logic; attribute dont_touch of G25088: signal is true;
	signal G25089: std_logic; attribute dont_touch of G25089: signal is true;
	signal G25090: std_logic; attribute dont_touch of G25090: signal is true;
	signal G25091: std_logic; attribute dont_touch of G25091: signal is true;
	signal G25092: std_logic; attribute dont_touch of G25092: signal is true;
	signal G25093: std_logic; attribute dont_touch of G25093: signal is true;
	signal G25094: std_logic; attribute dont_touch of G25094: signal is true;
	signal G25095: std_logic; attribute dont_touch of G25095: signal is true;
	signal G25096: std_logic; attribute dont_touch of G25096: signal is true;
	signal G25097: std_logic; attribute dont_touch of G25097: signal is true;
	signal G25098: std_logic; attribute dont_touch of G25098: signal is true;
	signal G25099: std_logic; attribute dont_touch of G25099: signal is true;
	signal G25100: std_logic; attribute dont_touch of G25100: signal is true;
	signal G25101: std_logic; attribute dont_touch of G25101: signal is true;
	signal G25102: std_logic; attribute dont_touch of G25102: signal is true;
	signal G25103: std_logic; attribute dont_touch of G25103: signal is true;
	signal G25104: std_logic; attribute dont_touch of G25104: signal is true;
	signal G25105: std_logic; attribute dont_touch of G25105: signal is true;
	signal G25106: std_logic; attribute dont_touch of G25106: signal is true;
	signal G25107: std_logic; attribute dont_touch of G25107: signal is true;
	signal G25108: std_logic; attribute dont_touch of G25108: signal is true;
	signal G25109: std_logic; attribute dont_touch of G25109: signal is true;
	signal G25110: std_logic; attribute dont_touch of G25110: signal is true;
	signal G25111: std_logic; attribute dont_touch of G25111: signal is true;
	signal G25112: std_logic; attribute dont_touch of G25112: signal is true;
	signal G25113: std_logic; attribute dont_touch of G25113: signal is true;
	signal G25115: std_logic; attribute dont_touch of G25115: signal is true;
	signal G25116: std_logic; attribute dont_touch of G25116: signal is true;
	signal G25117: std_logic; attribute dont_touch of G25117: signal is true;
	signal G25118: std_logic; attribute dont_touch of G25118: signal is true;
	signal G25119: std_logic; attribute dont_touch of G25119: signal is true;
	signal G25120: std_logic; attribute dont_touch of G25120: signal is true;
	signal G25121: std_logic; attribute dont_touch of G25121: signal is true;
	signal G25122: std_logic; attribute dont_touch of G25122: signal is true;
	signal G25123: std_logic; attribute dont_touch of G25123: signal is true;
	signal G25124: std_logic; attribute dont_touch of G25124: signal is true;
	signal G25125: std_logic; attribute dont_touch of G25125: signal is true;
	signal G25126: std_logic; attribute dont_touch of G25126: signal is true;
	signal G25127: std_logic; attribute dont_touch of G25127: signal is true;
	signal G25128: std_logic; attribute dont_touch of G25128: signal is true;
	signal G25129: std_logic; attribute dont_touch of G25129: signal is true;
	signal G25130: std_logic; attribute dont_touch of G25130: signal is true;
	signal G25131: std_logic; attribute dont_touch of G25131: signal is true;
	signal G25132: std_logic; attribute dont_touch of G25132: signal is true;
	signal G25133: std_logic; attribute dont_touch of G25133: signal is true;
	signal G25134: std_logic; attribute dont_touch of G25134: signal is true;
	signal G25135: std_logic; attribute dont_touch of G25135: signal is true;
	signal G25136: std_logic; attribute dont_touch of G25136: signal is true;
	signal G25137: std_logic; attribute dont_touch of G25137: signal is true;
	signal G25138: std_logic; attribute dont_touch of G25138: signal is true;
	signal G25139: std_logic; attribute dont_touch of G25139: signal is true;
	signal G25140: std_logic; attribute dont_touch of G25140: signal is true;
	signal G25141: std_logic; attribute dont_touch of G25141: signal is true;
	signal G25142: std_logic; attribute dont_touch of G25142: signal is true;
	signal G25143: std_logic; attribute dont_touch of G25143: signal is true;
	signal G25144: std_logic; attribute dont_touch of G25144: signal is true;
	signal G25147: std_logic; attribute dont_touch of G25147: signal is true;
	signal G25148: std_logic; attribute dont_touch of G25148: signal is true;
	signal G25149: std_logic; attribute dont_touch of G25149: signal is true;
	signal G25150: std_logic; attribute dont_touch of G25150: signal is true;
	signal G25151: std_logic; attribute dont_touch of G25151: signal is true;
	signal G25152: std_logic; attribute dont_touch of G25152: signal is true;
	signal G25153: std_logic; attribute dont_touch of G25153: signal is true;
	signal G25154: std_logic; attribute dont_touch of G25154: signal is true;
	signal G25155: std_logic; attribute dont_touch of G25155: signal is true;
	signal G25156: std_logic; attribute dont_touch of G25156: signal is true;
	signal G25157: std_logic; attribute dont_touch of G25157: signal is true;
	signal G25158: std_logic; attribute dont_touch of G25158: signal is true;
	signal G25159: std_logic; attribute dont_touch of G25159: signal is true;
	signal G25160: std_logic; attribute dont_touch of G25160: signal is true;
	signal G25163: std_logic; attribute dont_touch of G25163: signal is true;
	signal G25164: std_logic; attribute dont_touch of G25164: signal is true;
	signal G25165: std_logic; attribute dont_touch of G25165: signal is true;
	signal G25166: std_logic; attribute dont_touch of G25166: signal is true;
	signal G25168: std_logic; attribute dont_touch of G25168: signal is true;
	signal G25169: std_logic; attribute dont_touch of G25169: signal is true;
	signal G25170: std_logic; attribute dont_touch of G25170: signal is true;
	signal G25171: std_logic; attribute dont_touch of G25171: signal is true;
	signal G25172: std_logic; attribute dont_touch of G25172: signal is true;
	signal G25173: std_logic; attribute dont_touch of G25173: signal is true;
	signal G25174: std_logic; attribute dont_touch of G25174: signal is true;
	signal G25175: std_logic; attribute dont_touch of G25175: signal is true;
	signal G25178: std_logic; attribute dont_touch of G25178: signal is true;
	signal G25179: std_logic; attribute dont_touch of G25179: signal is true;
	signal G25180: std_logic; attribute dont_touch of G25180: signal is true;
	signal G25181: std_logic; attribute dont_touch of G25181: signal is true;
	signal G25182: std_logic; attribute dont_touch of G25182: signal is true;
	signal G25183: std_logic; attribute dont_touch of G25183: signal is true;
	signal G25184: std_logic; attribute dont_touch of G25184: signal is true;
	signal G25185: std_logic; attribute dont_touch of G25185: signal is true;
	signal G25186: std_logic; attribute dont_touch of G25186: signal is true;
	signal G25187: std_logic; attribute dont_touch of G25187: signal is true;
	signal G25188: std_logic; attribute dont_touch of G25188: signal is true;
	signal G25189: std_logic; attribute dont_touch of G25189: signal is true;
	signal G25192: std_logic; attribute dont_touch of G25192: signal is true;
	signal G25193: std_logic; attribute dont_touch of G25193: signal is true;
	signal G25194: std_logic; attribute dont_touch of G25194: signal is true;
	signal G25195: std_logic; attribute dont_touch of G25195: signal is true;
	signal G25196: std_logic; attribute dont_touch of G25196: signal is true;
	signal G25197: std_logic; attribute dont_touch of G25197: signal is true;
	signal G25198: std_logic; attribute dont_touch of G25198: signal is true;
	signal G25199: std_logic; attribute dont_touch of G25199: signal is true;
	signal G25200: std_logic; attribute dont_touch of G25200: signal is true;
	signal G25201: std_logic; attribute dont_touch of G25201: signal is true;
	signal G25202: std_logic; attribute dont_touch of G25202: signal is true;
	signal G25203: std_logic; attribute dont_touch of G25203: signal is true;
	signal G25206: std_logic; attribute dont_touch of G25206: signal is true;
	signal G25207: std_logic; attribute dont_touch of G25207: signal is true;
	signal G25208: std_logic; attribute dont_touch of G25208: signal is true;
	signal G25209: std_logic; attribute dont_touch of G25209: signal is true;
	signal G25210: std_logic; attribute dont_touch of G25210: signal is true;
	signal G25211: std_logic; attribute dont_touch of G25211: signal is true;
	signal G25212: std_logic; attribute dont_touch of G25212: signal is true;
	signal G25213: std_logic; attribute dont_touch of G25213: signal is true;
	signal G25214: std_logic; attribute dont_touch of G25214: signal is true;
	signal G25215: std_logic; attribute dont_touch of G25215: signal is true;
	signal G25216: std_logic; attribute dont_touch of G25216: signal is true;
	signal G25217: std_logic; attribute dont_touch of G25217: signal is true;
	signal G25218: std_logic; attribute dont_touch of G25218: signal is true;
	signal G25220: std_logic; attribute dont_touch of G25220: signal is true;
	signal G25221: std_logic; attribute dont_touch of G25221: signal is true;
	signal G25222: std_logic; attribute dont_touch of G25222: signal is true;
	signal G25223: std_logic; attribute dont_touch of G25223: signal is true;
	signal G25224: std_logic; attribute dont_touch of G25224: signal is true;
	signal G25225: std_logic; attribute dont_touch of G25225: signal is true;
	signal G25226: std_logic; attribute dont_touch of G25226: signal is true;
	signal G25227: std_logic; attribute dont_touch of G25227: signal is true;
	signal G25228: std_logic; attribute dont_touch of G25228: signal is true;
	signal G25229: std_logic; attribute dont_touch of G25229: signal is true;
	signal G25230: std_logic; attribute dont_touch of G25230: signal is true;
	signal G25231: std_logic; attribute dont_touch of G25231: signal is true;
	signal G25232: std_logic; attribute dont_touch of G25232: signal is true;
	signal G25233: std_logic; attribute dont_touch of G25233: signal is true;
	signal G25236: std_logic; attribute dont_touch of G25236: signal is true;
	signal G25237: std_logic; attribute dont_touch of G25237: signal is true;
	signal G25238: std_logic; attribute dont_touch of G25238: signal is true;
	signal G25239: std_logic; attribute dont_touch of G25239: signal is true;
	signal G25240: std_logic; attribute dont_touch of G25240: signal is true;
	signal G25241: std_logic; attribute dont_touch of G25241: signal is true;
	signal G25242: std_logic; attribute dont_touch of G25242: signal is true;
	signal G25243: std_logic; attribute dont_touch of G25243: signal is true;
	signal G25244: std_logic; attribute dont_touch of G25244: signal is true;
	signal G25245: std_logic; attribute dont_touch of G25245: signal is true;
	signal G25246: std_logic; attribute dont_touch of G25246: signal is true;
	signal G25247: std_logic; attribute dont_touch of G25247: signal is true;
	signal G25248: std_logic; attribute dont_touch of G25248: signal is true;
	signal G25249: std_logic; attribute dont_touch of G25249: signal is true;
	signal G25250: std_logic; attribute dont_touch of G25250: signal is true;
	signal G25255: std_logic; attribute dont_touch of G25255: signal is true;
	signal G25258: std_logic; attribute dont_touch of G25258: signal is true;
	signal G25260: std_logic; attribute dont_touch of G25260: signal is true;
	signal G25261: std_logic; attribute dont_touch of G25261: signal is true;
	signal G25262: std_logic; attribute dont_touch of G25262: signal is true;
	signal G25263: std_logic; attribute dont_touch of G25263: signal is true;
	signal G25264: std_logic; attribute dont_touch of G25264: signal is true;
	signal G25265: std_logic; attribute dont_touch of G25265: signal is true;
	signal G25266: std_logic; attribute dont_touch of G25266: signal is true;
	signal G25267: std_logic; attribute dont_touch of G25267: signal is true;
	signal G25268: std_logic; attribute dont_touch of G25268: signal is true;
	signal G25271: std_logic; attribute dont_touch of G25271: signal is true;
	signal G25272: std_logic; attribute dont_touch of G25272: signal is true;
	signal G25273: std_logic; attribute dont_touch of G25273: signal is true;
	signal G25274: std_logic; attribute dont_touch of G25274: signal is true;
	signal G25275: std_logic; attribute dont_touch of G25275: signal is true;
	signal G25282: std_logic; attribute dont_touch of G25282: signal is true;
	signal G25283: std_logic; attribute dont_touch of G25283: signal is true;
	signal G25284: std_logic; attribute dont_touch of G25284: signal is true;
	signal G25285: std_logic; attribute dont_touch of G25285: signal is true;
	signal G25286: std_logic; attribute dont_touch of G25286: signal is true;
	signal G25287: std_logic; attribute dont_touch of G25287: signal is true;
	signal G25288: std_logic; attribute dont_touch of G25288: signal is true;
	signal G25289: std_logic; attribute dont_touch of G25289: signal is true;
	signal G25290: std_logic; attribute dont_touch of G25290: signal is true;
	signal G25293: std_logic; attribute dont_touch of G25293: signal is true;
	signal G25296: std_logic; attribute dont_touch of G25296: signal is true;
	signal G25297: std_logic; attribute dont_touch of G25297: signal is true;
	signal G25298: std_logic; attribute dont_touch of G25298: signal is true;
	signal G25299: std_logic; attribute dont_touch of G25299: signal is true;
	signal G25300: std_logic; attribute dont_touch of G25300: signal is true;
	signal G25307: std_logic; attribute dont_touch of G25307: signal is true;
	signal G25308: std_logic; attribute dont_touch of G25308: signal is true;
	signal G25309: std_logic; attribute dont_touch of G25309: signal is true;
	signal G25316: std_logic; attribute dont_touch of G25316: signal is true;
	signal G25317: std_logic; attribute dont_touch of G25317: signal is true;
	signal G25321: std_logic; attribute dont_touch of G25321: signal is true;
	signal G25322: std_logic; attribute dont_touch of G25322: signal is true;
	signal G25323: std_logic; attribute dont_touch of G25323: signal is true;
	signal G25324: std_logic; attribute dont_touch of G25324: signal is true;
	signal G25325: std_logic; attribute dont_touch of G25325: signal is true;
	signal G25326: std_logic; attribute dont_touch of G25326: signal is true;
	signal G25327: std_logic; attribute dont_touch of G25327: signal is true;
	signal G25328: std_logic; attribute dont_touch of G25328: signal is true;
	signal G25331: std_logic; attribute dont_touch of G25331: signal is true;
	signal G25334: std_logic; attribute dont_touch of G25334: signal is true;
	signal G25337: std_logic; attribute dont_touch of G25337: signal is true;
	signal G25340: std_logic; attribute dont_touch of G25340: signal is true;
	signal G25341: std_logic; attribute dont_touch of G25341: signal is true;
	signal G25348: std_logic; attribute dont_touch of G25348: signal is true;
	signal G25349: std_logic; attribute dont_touch of G25349: signal is true;
	signal G25356: std_logic; attribute dont_touch of G25356: signal is true;
	signal G25357: std_logic; attribute dont_touch of G25357: signal is true;
	signal G25366: std_logic; attribute dont_touch of G25366: signal is true;
	signal G25367: std_logic; attribute dont_touch of G25367: signal is true;
	signal G25368: std_logic; attribute dont_touch of G25368: signal is true;
	signal G25369: std_logic; attribute dont_touch of G25369: signal is true;
	signal G25370: std_logic; attribute dont_touch of G25370: signal is true;
	signal G25371: std_logic; attribute dont_touch of G25371: signal is true;
	signal G25374: std_logic; attribute dont_touch of G25374: signal is true;
	signal G25377: std_logic; attribute dont_touch of G25377: signal is true;
	signal G25380: std_logic; attribute dont_touch of G25380: signal is true;
	signal G25381: std_logic; attribute dont_touch of G25381: signal is true;
	signal G25382: std_logic; attribute dont_touch of G25382: signal is true;
	signal G25385: std_logic; attribute dont_touch of G25385: signal is true;
	signal G25388: std_logic; attribute dont_touch of G25388: signal is true;
	signal G25389: std_logic; attribute dont_touch of G25389: signal is true;
	signal G25396: std_logic; attribute dont_touch of G25396: signal is true;
	signal G25399: std_logic; attribute dont_touch of G25399: signal is true;
	signal G25400: std_logic; attribute dont_touch of G25400: signal is true;
	signal G25407: std_logic; attribute dont_touch of G25407: signal is true;
	signal G25408: std_logic; attribute dont_touch of G25408: signal is true;
	signal G25409: std_logic; attribute dont_touch of G25409: signal is true;
	signal G25410: std_logic; attribute dont_touch of G25410: signal is true;
	signal G25411: std_logic; attribute dont_touch of G25411: signal is true;
	signal G25414: std_logic; attribute dont_touch of G25414: signal is true;
	signal G25417: std_logic; attribute dont_touch of G25417: signal is true;
	signal G25420: std_logic; attribute dont_touch of G25420: signal is true;
	signal G25423: std_logic; attribute dont_touch of G25423: signal is true;
	signal G25424: std_logic; attribute dont_touch of G25424: signal is true;
	signal G25425: std_logic; attribute dont_touch of G25425: signal is true;
	signal G25426: std_logic; attribute dont_touch of G25426: signal is true;
	signal G25429: std_logic; attribute dont_touch of G25429: signal is true;
	signal G25432: std_logic; attribute dont_touch of G25432: signal is true;
	signal G25435: std_logic; attribute dont_touch of G25435: signal is true;
	signal G25438: std_logic; attribute dont_touch of G25438: signal is true;
	signal G25439: std_logic; attribute dont_touch of G25439: signal is true;
	signal G25446: std_logic; attribute dont_touch of G25446: signal is true;
	signal G25447: std_logic; attribute dont_touch of G25447: signal is true;
	signal G25448: std_logic; attribute dont_touch of G25448: signal is true;
	signal G25449: std_logic; attribute dont_touch of G25449: signal is true;
	signal G25450: std_logic; attribute dont_touch of G25450: signal is true;
	signal G25451: std_logic; attribute dont_touch of G25451: signal is true;
	signal G25452: std_logic; attribute dont_touch of G25452: signal is true;
	signal G25453: std_logic; attribute dont_touch of G25453: signal is true;
	signal G25456: std_logic; attribute dont_touch of G25456: signal is true;
	signal G25459: std_logic; attribute dont_touch of G25459: signal is true;
	signal G25462: std_logic; attribute dont_touch of G25462: signal is true;
	signal G25465: std_logic; attribute dont_touch of G25465: signal is true;
	signal G25466: std_logic; attribute dont_touch of G25466: signal is true;
	signal G25467: std_logic; attribute dont_touch of G25467: signal is true;
	signal G25470: std_logic; attribute dont_touch of G25470: signal is true;
	signal G25473: std_logic; attribute dont_touch of G25473: signal is true;
	signal G25476: std_logic; attribute dont_touch of G25476: signal is true;
	signal G25479: std_logic; attribute dont_touch of G25479: signal is true;
	signal G25480: std_logic; attribute dont_touch of G25480: signal is true;
	signal G25481: std_logic; attribute dont_touch of G25481: signal is true;
	signal G25482: std_logic; attribute dont_touch of G25482: signal is true;
	signal G25485: std_logic; attribute dont_touch of G25485: signal is true;
	signal G25488: std_logic; attribute dont_touch of G25488: signal is true;
	signal G25491: std_logic; attribute dont_touch of G25491: signal is true;
	signal G25492: std_logic; attribute dont_touch of G25492: signal is true;
	signal G25495: std_logic; attribute dont_touch of G25495: signal is true;
	signal G25498: std_logic; attribute dont_touch of G25498: signal is true;
	signal G25501: std_logic; attribute dont_touch of G25501: signal is true;
	signal G25502: std_logic; attribute dont_touch of G25502: signal is true;
	signal G25503: std_logic; attribute dont_touch of G25503: signal is true;
	signal G25504: std_logic; attribute dont_touch of G25504: signal is true;
	signal G25505: std_logic; attribute dont_touch of G25505: signal is true;
	signal G25506: std_logic; attribute dont_touch of G25506: signal is true;
	signal G25507: std_logic; attribute dont_touch of G25507: signal is true;
	signal G25510: std_logic; attribute dont_touch of G25510: signal is true;
	signal G25513: std_logic; attribute dont_touch of G25513: signal is true;
	signal G25514: std_logic; attribute dont_touch of G25514: signal is true;
	signal G25517: std_logic; attribute dont_touch of G25517: signal is true;
	signal G25518: std_logic; attribute dont_touch of G25518: signal is true;
	signal G25521: std_logic; attribute dont_touch of G25521: signal is true;
	signal G25522: std_logic; attribute dont_touch of G25522: signal is true;
	signal G25523: std_logic; attribute dont_touch of G25523: signal is true;
	signal G25524: std_logic; attribute dont_touch of G25524: signal is true;
	signal G25525: std_logic; attribute dont_touch of G25525: signal is true;
	signal G25526: std_logic; attribute dont_touch of G25526: signal is true;
	signal G25527: std_logic; attribute dont_touch of G25527: signal is true;
	signal G25528: std_logic; attribute dont_touch of G25528: signal is true;
	signal G25529: std_logic; attribute dont_touch of G25529: signal is true;
	signal G25530: std_logic; attribute dont_touch of G25530: signal is true;
	signal G25531: std_logic; attribute dont_touch of G25531: signal is true;
	signal G25532: std_logic; attribute dont_touch of G25532: signal is true;
	signal G25533: std_logic; attribute dont_touch of G25533: signal is true;
	signal G25534: std_logic; attribute dont_touch of G25534: signal is true;
	signal G25535: std_logic; attribute dont_touch of G25535: signal is true;
	signal G25536: std_logic; attribute dont_touch of G25536: signal is true;
	signal G25537: std_logic; attribute dont_touch of G25537: signal is true;
	signal G25538: std_logic; attribute dont_touch of G25538: signal is true;
	signal G25539: std_logic; attribute dont_touch of G25539: signal is true;
	signal G25540: std_logic; attribute dont_touch of G25540: signal is true;
	signal G25541: std_logic; attribute dont_touch of G25541: signal is true;
	signal G25542: std_logic; attribute dont_touch of G25542: signal is true;
	signal G25543: std_logic; attribute dont_touch of G25543: signal is true;
	signal G25544: std_logic; attribute dont_touch of G25544: signal is true;
	signal G25545: std_logic; attribute dont_touch of G25545: signal is true;
	signal G25546: std_logic; attribute dont_touch of G25546: signal is true;
	signal G25547: std_logic; attribute dont_touch of G25547: signal is true;
	signal G25548: std_logic; attribute dont_touch of G25548: signal is true;
	signal G25549: std_logic; attribute dont_touch of G25549: signal is true;
	signal G25550: std_logic; attribute dont_touch of G25550: signal is true;
	signal G25551: std_logic; attribute dont_touch of G25551: signal is true;
	signal G25552: std_logic; attribute dont_touch of G25552: signal is true;
	signal G25553: std_logic; attribute dont_touch of G25553: signal is true;
	signal G25554: std_logic; attribute dont_touch of G25554: signal is true;
	signal G25555: std_logic; attribute dont_touch of G25555: signal is true;
	signal G25556: std_logic; attribute dont_touch of G25556: signal is true;
	signal G25557: std_logic; attribute dont_touch of G25557: signal is true;
	signal G25558: std_logic; attribute dont_touch of G25558: signal is true;
	signal G25559: std_logic; attribute dont_touch of G25559: signal is true;
	signal G25560: std_logic; attribute dont_touch of G25560: signal is true;
	signal G25561: std_logic; attribute dont_touch of G25561: signal is true;
	signal G25562: std_logic; attribute dont_touch of G25562: signal is true;
	signal G25563: std_logic; attribute dont_touch of G25563: signal is true;
	signal G25564: std_logic; attribute dont_touch of G25564: signal is true;
	signal G25565: std_logic; attribute dont_touch of G25565: signal is true;
	signal G25566: std_logic; attribute dont_touch of G25566: signal is true;
	signal G25567: std_logic; attribute dont_touch of G25567: signal is true;
	signal G25568: std_logic; attribute dont_touch of G25568: signal is true;
	signal G25569: std_logic; attribute dont_touch of G25569: signal is true;
	signal G25570: std_logic; attribute dont_touch of G25570: signal is true;
	signal G25571: std_logic; attribute dont_touch of G25571: signal is true;
	signal G25572: std_logic; attribute dont_touch of G25572: signal is true;
	signal G25573: std_logic; attribute dont_touch of G25573: signal is true;
	signal G25574: std_logic; attribute dont_touch of G25574: signal is true;
	signal G25575: std_logic; attribute dont_touch of G25575: signal is true;
	signal G25576: std_logic; attribute dont_touch of G25576: signal is true;
	signal G25577: std_logic; attribute dont_touch of G25577: signal is true;
	signal G25578: std_logic; attribute dont_touch of G25578: signal is true;
	signal G25579: std_logic; attribute dont_touch of G25579: signal is true;
	signal G25580: std_logic; attribute dont_touch of G25580: signal is true;
	signal G25581: std_logic; attribute dont_touch of G25581: signal is true;
	signal G25591: std_logic; attribute dont_touch of G25591: signal is true;
	signal G25592: std_logic; attribute dont_touch of G25592: signal is true;
	signal G25593: std_logic; attribute dont_touch of G25593: signal is true;
	signal G25594: std_logic; attribute dont_touch of G25594: signal is true;
	signal G25595: std_logic; attribute dont_touch of G25595: signal is true;
	signal G25596: std_logic; attribute dont_touch of G25596: signal is true;
	signal G25597: std_logic; attribute dont_touch of G25597: signal is true;
	signal G25598: std_logic; attribute dont_touch of G25598: signal is true;
	signal G25599: std_logic; attribute dont_touch of G25599: signal is true;
	signal G25600: std_logic; attribute dont_touch of G25600: signal is true;
	signal G25601: std_logic; attribute dont_touch of G25601: signal is true;
	signal G25602: std_logic; attribute dont_touch of G25602: signal is true;
	signal G25603: std_logic; attribute dont_touch of G25603: signal is true;
	signal G25604: std_logic; attribute dont_touch of G25604: signal is true;
	signal G25605: std_logic; attribute dont_touch of G25605: signal is true;
	signal G25606: std_logic; attribute dont_touch of G25606: signal is true;
	signal G25607: std_logic; attribute dont_touch of G25607: signal is true;
	signal G25608: std_logic; attribute dont_touch of G25608: signal is true;
	signal G25609: std_logic; attribute dont_touch of G25609: signal is true;
	signal G25610: std_logic; attribute dont_touch of G25610: signal is true;
	signal G25611: std_logic; attribute dont_touch of G25611: signal is true;
	signal G25612: std_logic; attribute dont_touch of G25612: signal is true;
	signal G25613: std_logic; attribute dont_touch of G25613: signal is true;
	signal G25614: std_logic; attribute dont_touch of G25614: signal is true;
	signal G25615: std_logic; attribute dont_touch of G25615: signal is true;
	signal G25616: std_logic; attribute dont_touch of G25616: signal is true;
	signal G25617: std_logic; attribute dont_touch of G25617: signal is true;
	signal G25618: std_logic; attribute dont_touch of G25618: signal is true;
	signal G25619: std_logic; attribute dont_touch of G25619: signal is true;
	signal G25620: std_logic; attribute dont_touch of G25620: signal is true;
	signal G25621: std_logic; attribute dont_touch of G25621: signal is true;
	signal G25622: std_logic; attribute dont_touch of G25622: signal is true;
	signal G25623: std_logic; attribute dont_touch of G25623: signal is true;
	signal G25624: std_logic; attribute dont_touch of G25624: signal is true;
	signal G25625: std_logic; attribute dont_touch of G25625: signal is true;
	signal G25626: std_logic; attribute dont_touch of G25626: signal is true;
	signal G25627: std_logic; attribute dont_touch of G25627: signal is true;
	signal G25628: std_logic; attribute dont_touch of G25628: signal is true;
	signal G25629: std_logic; attribute dont_touch of G25629: signal is true;
	signal G25630: std_logic; attribute dont_touch of G25630: signal is true;
	signal G25631: std_logic; attribute dont_touch of G25631: signal is true;
	signal G25632: std_logic; attribute dont_touch of G25632: signal is true;
	signal G25633: std_logic; attribute dont_touch of G25633: signal is true;
	signal G25634: std_logic; attribute dont_touch of G25634: signal is true;
	signal G25635: std_logic; attribute dont_touch of G25635: signal is true;
	signal G25636: std_logic; attribute dont_touch of G25636: signal is true;
	signal G25637: std_logic; attribute dont_touch of G25637: signal is true;
	signal G25638: std_logic; attribute dont_touch of G25638: signal is true;
	signal G25639: std_logic; attribute dont_touch of G25639: signal is true;
	signal G25640: std_logic; attribute dont_touch of G25640: signal is true;
	signal G25641: std_logic; attribute dont_touch of G25641: signal is true;
	signal G25642: std_logic; attribute dont_touch of G25642: signal is true;
	signal G25643: std_logic; attribute dont_touch of G25643: signal is true;
	signal G25644: std_logic; attribute dont_touch of G25644: signal is true;
	signal G25645: std_logic; attribute dont_touch of G25645: signal is true;
	signal G25646: std_logic; attribute dont_touch of G25646: signal is true;
	signal G25647: std_logic; attribute dont_touch of G25647: signal is true;
	signal G25648: std_logic; attribute dont_touch of G25648: signal is true;
	signal G25649: std_logic; attribute dont_touch of G25649: signal is true;
	signal G25650: std_logic; attribute dont_touch of G25650: signal is true;
	signal G25651: std_logic; attribute dont_touch of G25651: signal is true;
	signal G25652: std_logic; attribute dont_touch of G25652: signal is true;
	signal G25653: std_logic; attribute dont_touch of G25653: signal is true;
	signal G25654: std_logic; attribute dont_touch of G25654: signal is true;
	signal G25655: std_logic; attribute dont_touch of G25655: signal is true;
	signal G25656: std_logic; attribute dont_touch of G25656: signal is true;
	signal G25657: std_logic; attribute dont_touch of G25657: signal is true;
	signal G25658: std_logic; attribute dont_touch of G25658: signal is true;
	signal G25659: std_logic; attribute dont_touch of G25659: signal is true;
	signal G25660: std_logic; attribute dont_touch of G25660: signal is true;
	signal G25661: std_logic; attribute dont_touch of G25661: signal is true;
	signal G25662: std_logic; attribute dont_touch of G25662: signal is true;
	signal G25663: std_logic; attribute dont_touch of G25663: signal is true;
	signal G25664: std_logic; attribute dont_touch of G25664: signal is true;
	signal G25665: std_logic; attribute dont_touch of G25665: signal is true;
	signal G25666: std_logic; attribute dont_touch of G25666: signal is true;
	signal G25667: std_logic; attribute dont_touch of G25667: signal is true;
	signal G25668: std_logic; attribute dont_touch of G25668: signal is true;
	signal G25669: std_logic; attribute dont_touch of G25669: signal is true;
	signal G25670: std_logic; attribute dont_touch of G25670: signal is true;
	signal G25671: std_logic; attribute dont_touch of G25671: signal is true;
	signal G25672: std_logic; attribute dont_touch of G25672: signal is true;
	signal G25673: std_logic; attribute dont_touch of G25673: signal is true;
	signal G25674: std_logic; attribute dont_touch of G25674: signal is true;
	signal G25675: std_logic; attribute dont_touch of G25675: signal is true;
	signal G25676: std_logic; attribute dont_touch of G25676: signal is true;
	signal G25677: std_logic; attribute dont_touch of G25677: signal is true;
	signal G25678: std_logic; attribute dont_touch of G25678: signal is true;
	signal G25679: std_logic; attribute dont_touch of G25679: signal is true;
	signal G25680: std_logic; attribute dont_touch of G25680: signal is true;
	signal G25681: std_logic; attribute dont_touch of G25681: signal is true;
	signal G25682: std_logic; attribute dont_touch of G25682: signal is true;
	signal G25683: std_logic; attribute dont_touch of G25683: signal is true;
	signal G25684: std_logic; attribute dont_touch of G25684: signal is true;
	signal G25685: std_logic; attribute dont_touch of G25685: signal is true;
	signal G25686: std_logic; attribute dont_touch of G25686: signal is true;
	signal G25687: std_logic; attribute dont_touch of G25687: signal is true;
	signal G25688: std_logic; attribute dont_touch of G25688: signal is true;
	signal G25689: std_logic; attribute dont_touch of G25689: signal is true;
	signal G25690: std_logic; attribute dont_touch of G25690: signal is true;
	signal G25691: std_logic; attribute dont_touch of G25691: signal is true;
	signal G25692: std_logic; attribute dont_touch of G25692: signal is true;
	signal G25693: std_logic; attribute dont_touch of G25693: signal is true;
	signal G25694: std_logic; attribute dont_touch of G25694: signal is true;
	signal G25695: std_logic; attribute dont_touch of G25695: signal is true;
	signal G25696: std_logic; attribute dont_touch of G25696: signal is true;
	signal G25697: std_logic; attribute dont_touch of G25697: signal is true;
	signal G25698: std_logic; attribute dont_touch of G25698: signal is true;
	signal G25699: std_logic; attribute dont_touch of G25699: signal is true;
	signal G25700: std_logic; attribute dont_touch of G25700: signal is true;
	signal G25701: std_logic; attribute dont_touch of G25701: signal is true;
	signal G25702: std_logic; attribute dont_touch of G25702: signal is true;
	signal G25703: std_logic; attribute dont_touch of G25703: signal is true;
	signal G25704: std_logic; attribute dont_touch of G25704: signal is true;
	signal G25705: std_logic; attribute dont_touch of G25705: signal is true;
	signal G25706: std_logic; attribute dont_touch of G25706: signal is true;
	signal G25707: std_logic; attribute dont_touch of G25707: signal is true;
	signal G25708: std_logic; attribute dont_touch of G25708: signal is true;
	signal G25709: std_logic; attribute dont_touch of G25709: signal is true;
	signal G25710: std_logic; attribute dont_touch of G25710: signal is true;
	signal G25711: std_logic; attribute dont_touch of G25711: signal is true;
	signal G25712: std_logic; attribute dont_touch of G25712: signal is true;
	signal G25713: std_logic; attribute dont_touch of G25713: signal is true;
	signal G25714: std_logic; attribute dont_touch of G25714: signal is true;
	signal G25715: std_logic; attribute dont_touch of G25715: signal is true;
	signal G25716: std_logic; attribute dont_touch of G25716: signal is true;
	signal G25717: std_logic; attribute dont_touch of G25717: signal is true;
	signal G25718: std_logic; attribute dont_touch of G25718: signal is true;
	signal G25719: std_logic; attribute dont_touch of G25719: signal is true;
	signal G25720: std_logic; attribute dont_touch of G25720: signal is true;
	signal G25721: std_logic; attribute dont_touch of G25721: signal is true;
	signal G25722: std_logic; attribute dont_touch of G25722: signal is true;
	signal G25723: std_logic; attribute dont_touch of G25723: signal is true;
	signal G25724: std_logic; attribute dont_touch of G25724: signal is true;
	signal G25725: std_logic; attribute dont_touch of G25725: signal is true;
	signal G25726: std_logic; attribute dont_touch of G25726: signal is true;
	signal G25727: std_logic; attribute dont_touch of G25727: signal is true;
	signal G25728: std_logic; attribute dont_touch of G25728: signal is true;
	signal G25729: std_logic; attribute dont_touch of G25729: signal is true;
	signal G25730: std_logic; attribute dont_touch of G25730: signal is true;
	signal G25731: std_logic; attribute dont_touch of G25731: signal is true;
	signal G25732: std_logic; attribute dont_touch of G25732: signal is true;
	signal G25733: std_logic; attribute dont_touch of G25733: signal is true;
	signal G25734: std_logic; attribute dont_touch of G25734: signal is true;
	signal G25735: std_logic; attribute dont_touch of G25735: signal is true;
	signal G25736: std_logic; attribute dont_touch of G25736: signal is true;
	signal G25737: std_logic; attribute dont_touch of G25737: signal is true;
	signal G25738: std_logic; attribute dont_touch of G25738: signal is true;
	signal G25739: std_logic; attribute dont_touch of G25739: signal is true;
	signal G25740: std_logic; attribute dont_touch of G25740: signal is true;
	signal G25741: std_logic; attribute dont_touch of G25741: signal is true;
	signal G25742: std_logic; attribute dont_touch of G25742: signal is true;
	signal G25743: std_logic; attribute dont_touch of G25743: signal is true;
	signal G25744: std_logic; attribute dont_touch of G25744: signal is true;
	signal G25745: std_logic; attribute dont_touch of G25745: signal is true;
	signal G25746: std_logic; attribute dont_touch of G25746: signal is true;
	signal G25747: std_logic; attribute dont_touch of G25747: signal is true;
	signal G25748: std_logic; attribute dont_touch of G25748: signal is true;
	signal G25749: std_logic; attribute dont_touch of G25749: signal is true;
	signal G25750: std_logic; attribute dont_touch of G25750: signal is true;
	signal G25751: std_logic; attribute dont_touch of G25751: signal is true;
	signal G25752: std_logic; attribute dont_touch of G25752: signal is true;
	signal G25753: std_logic; attribute dont_touch of G25753: signal is true;
	signal G25754: std_logic; attribute dont_touch of G25754: signal is true;
	signal G25755: std_logic; attribute dont_touch of G25755: signal is true;
	signal G25756: std_logic; attribute dont_touch of G25756: signal is true;
	signal G25757: std_logic; attribute dont_touch of G25757: signal is true;
	signal G25758: std_logic; attribute dont_touch of G25758: signal is true;
	signal G25759: std_logic; attribute dont_touch of G25759: signal is true;
	signal G25760: std_logic; attribute dont_touch of G25760: signal is true;
	signal G25761: std_logic; attribute dont_touch of G25761: signal is true;
	signal G25762: std_logic; attribute dont_touch of G25762: signal is true;
	signal G25763: std_logic; attribute dont_touch of G25763: signal is true;
	signal G25764: std_logic; attribute dont_touch of G25764: signal is true;
	signal G25765: std_logic; attribute dont_touch of G25765: signal is true;
	signal G25766: std_logic; attribute dont_touch of G25766: signal is true;
	signal G25767: std_logic; attribute dont_touch of G25767: signal is true;
	signal G25768: std_logic; attribute dont_touch of G25768: signal is true;
	signal G25769: std_logic; attribute dont_touch of G25769: signal is true;
	signal G25770: std_logic; attribute dont_touch of G25770: signal is true;
	signal G25771: std_logic; attribute dont_touch of G25771: signal is true;
	signal G25772: std_logic; attribute dont_touch of G25772: signal is true;
	signal G25773: std_logic; attribute dont_touch of G25773: signal is true;
	signal G25774: std_logic; attribute dont_touch of G25774: signal is true;
	signal G25775: std_logic; attribute dont_touch of G25775: signal is true;
	signal G25776: std_logic; attribute dont_touch of G25776: signal is true;
	signal G25777: std_logic; attribute dont_touch of G25777: signal is true;
	signal G25778: std_logic; attribute dont_touch of G25778: signal is true;
	signal G25779: std_logic; attribute dont_touch of G25779: signal is true;
	signal G25780: std_logic; attribute dont_touch of G25780: signal is true;
	signal G25781: std_logic; attribute dont_touch of G25781: signal is true;
	signal G25782: std_logic; attribute dont_touch of G25782: signal is true;
	signal G25783: std_logic; attribute dont_touch of G25783: signal is true;
	signal G25784: std_logic; attribute dont_touch of G25784: signal is true;
	signal G25785: std_logic; attribute dont_touch of G25785: signal is true;
	signal G25786: std_logic; attribute dont_touch of G25786: signal is true;
	signal G25787: std_logic; attribute dont_touch of G25787: signal is true;
	signal G25788: std_logic; attribute dont_touch of G25788: signal is true;
	signal G25789: std_logic; attribute dont_touch of G25789: signal is true;
	signal G25790: std_logic; attribute dont_touch of G25790: signal is true;
	signal G25791: std_logic; attribute dont_touch of G25791: signal is true;
	signal G25800: std_logic; attribute dont_touch of G25800: signal is true;
	signal G25801: std_logic; attribute dont_touch of G25801: signal is true;
	signal G25802: std_logic; attribute dont_touch of G25802: signal is true;
	signal G25803: std_logic; attribute dont_touch of G25803: signal is true;
	signal G25804: std_logic; attribute dont_touch of G25804: signal is true;
	signal G25805: std_logic; attribute dont_touch of G25805: signal is true;
	signal G25814: std_logic; attribute dont_touch of G25814: signal is true;
	signal G25815: std_logic; attribute dont_touch of G25815: signal is true;
	signal G25816: std_logic; attribute dont_touch of G25816: signal is true;
	signal G25817: std_logic; attribute dont_touch of G25817: signal is true;
	signal G25818: std_logic; attribute dont_touch of G25818: signal is true;
	signal G25819: std_logic; attribute dont_touch of G25819: signal is true;
	signal G25820: std_logic; attribute dont_touch of G25820: signal is true;
	signal G25821: std_logic; attribute dont_touch of G25821: signal is true;
	signal G25830: std_logic; attribute dont_touch of G25830: signal is true;
	signal G25831: std_logic; attribute dont_touch of G25831: signal is true;
	signal G25832: std_logic; attribute dont_touch of G25832: signal is true;
	signal G25833: std_logic; attribute dont_touch of G25833: signal is true;
	signal G25834: std_logic; attribute dont_touch of G25834: signal is true;
	signal G25835: std_logic; attribute dont_touch of G25835: signal is true;
	signal G25836: std_logic; attribute dont_touch of G25836: signal is true;
	signal G25837: std_logic; attribute dont_touch of G25837: signal is true;
	signal G25838: std_logic; attribute dont_touch of G25838: signal is true;
	signal G25839: std_logic; attribute dont_touch of G25839: signal is true;
	signal G25848: std_logic; attribute dont_touch of G25848: signal is true;
	signal G25849: std_logic; attribute dont_touch of G25849: signal is true;
	signal G25850: std_logic; attribute dont_touch of G25850: signal is true;
	signal G25851: std_logic; attribute dont_touch of G25851: signal is true;
	signal G25852: std_logic; attribute dont_touch of G25852: signal is true;
	signal G25856: std_logic; attribute dont_touch of G25856: signal is true;
	signal G25865: std_logic; attribute dont_touch of G25865: signal is true;
	signal G25866: std_logic; attribute dont_touch of G25866: signal is true;
	signal G25867: std_logic; attribute dont_touch of G25867: signal is true;
	signal G25868: std_logic; attribute dont_touch of G25868: signal is true;
	signal G25869: std_logic; attribute dont_touch of G25869: signal is true;
	signal G25870: std_logic; attribute dont_touch of G25870: signal is true;
	signal G25871: std_logic; attribute dont_touch of G25871: signal is true;
	signal G25872: std_logic; attribute dont_touch of G25872: signal is true;
	signal G25873: std_logic; attribute dont_touch of G25873: signal is true;
	signal G25874: std_logic; attribute dont_touch of G25874: signal is true;
	signal G25875: std_logic; attribute dont_touch of G25875: signal is true;
	signal G25876: std_logic; attribute dont_touch of G25876: signal is true;
	signal G25877: std_logic; attribute dont_touch of G25877: signal is true;
	signal G25878: std_logic; attribute dont_touch of G25878: signal is true;
	signal G25879: std_logic; attribute dont_touch of G25879: signal is true;
	signal G25880: std_logic; attribute dont_touch of G25880: signal is true;
	signal G25881: std_logic; attribute dont_touch of G25881: signal is true;
	signal G25882: std_logic; attribute dont_touch of G25882: signal is true;
	signal G25883: std_logic; attribute dont_touch of G25883: signal is true;
	signal G25884: std_logic; attribute dont_touch of G25884: signal is true;
	signal G25885: std_logic; attribute dont_touch of G25885: signal is true;
	signal G25886: std_logic; attribute dont_touch of G25886: signal is true;
	signal G25887: std_logic; attribute dont_touch of G25887: signal is true;
	signal G25888: std_logic; attribute dont_touch of G25888: signal is true;
	signal G25892: std_logic; attribute dont_touch of G25892: signal is true;
	signal G25893: std_logic; attribute dont_touch of G25893: signal is true;
	signal G25894: std_logic; attribute dont_touch of G25894: signal is true;
	signal G25895: std_logic; attribute dont_touch of G25895: signal is true;
	signal G25899: std_logic; attribute dont_touch of G25899: signal is true;
	signal G25900: std_logic; attribute dont_touch of G25900: signal is true;
	signal G25901: std_logic; attribute dont_touch of G25901: signal is true;
	signal G25902: std_logic; attribute dont_touch of G25902: signal is true;
	signal G25903: std_logic; attribute dont_touch of G25903: signal is true;
	signal G25904: std_logic; attribute dont_touch of G25904: signal is true;
	signal G25905: std_logic; attribute dont_touch of G25905: signal is true;
	signal G25906: std_logic; attribute dont_touch of G25906: signal is true;
	signal G25907: std_logic; attribute dont_touch of G25907: signal is true;
	signal G25908: std_logic; attribute dont_touch of G25908: signal is true;
	signal G25909: std_logic; attribute dont_touch of G25909: signal is true;
	signal G25910: std_logic; attribute dont_touch of G25910: signal is true;
	signal G25911: std_logic; attribute dont_touch of G25911: signal is true;
	signal G25915: std_logic; attribute dont_touch of G25915: signal is true;
	signal G25916: std_logic; attribute dont_touch of G25916: signal is true;
	signal G25917: std_logic; attribute dont_touch of G25917: signal is true;
	signal G25921: std_logic; attribute dont_touch of G25921: signal is true;
	signal G25922: std_logic; attribute dont_touch of G25922: signal is true;
	signal G25923: std_logic; attribute dont_touch of G25923: signal is true;
	signal G25924: std_logic; attribute dont_touch of G25924: signal is true;
	signal G25925: std_logic; attribute dont_touch of G25925: signal is true;
	signal G25926: std_logic; attribute dont_touch of G25926: signal is true;
	signal G25927: std_logic; attribute dont_touch of G25927: signal is true;
	signal G25928: std_logic; attribute dont_touch of G25928: signal is true;
	signal G25929: std_logic; attribute dont_touch of G25929: signal is true;
	signal G25930: std_logic; attribute dont_touch of G25930: signal is true;
	signal G25931: std_logic; attribute dont_touch of G25931: signal is true;
	signal G25932: std_logic; attribute dont_touch of G25932: signal is true;
	signal G25935: std_logic; attribute dont_touch of G25935: signal is true;
	signal G25936: std_logic; attribute dont_touch of G25936: signal is true;
	signal G25937: std_logic; attribute dont_touch of G25937: signal is true;
	signal G25938: std_logic; attribute dont_touch of G25938: signal is true;
	signal G25939: std_logic; attribute dont_touch of G25939: signal is true;
	signal G25940: std_logic; attribute dont_touch of G25940: signal is true;
	signal G25941: std_logic; attribute dont_touch of G25941: signal is true;
	signal G25942: std_logic; attribute dont_touch of G25942: signal is true;
	signal G25943: std_logic; attribute dont_touch of G25943: signal is true;
	signal G25944: std_logic; attribute dont_touch of G25944: signal is true;
	signal G25945: std_logic; attribute dont_touch of G25945: signal is true;
	signal G25946: std_logic; attribute dont_touch of G25946: signal is true;
	signal G25947: std_logic; attribute dont_touch of G25947: signal is true;
	signal G25948: std_logic; attribute dont_touch of G25948: signal is true;
	signal G25949: std_logic; attribute dont_touch of G25949: signal is true;
	signal G25950: std_logic; attribute dont_touch of G25950: signal is true;
	signal G25951: std_logic; attribute dont_touch of G25951: signal is true;
	signal G25952: std_logic; attribute dont_touch of G25952: signal is true;
	signal G25953: std_logic; attribute dont_touch of G25953: signal is true;
	signal G25954: std_logic; attribute dont_touch of G25954: signal is true;
	signal G25955: std_logic; attribute dont_touch of G25955: signal is true;
	signal G25956: std_logic; attribute dont_touch of G25956: signal is true;
	signal G25957: std_logic; attribute dont_touch of G25957: signal is true;
	signal G25958: std_logic; attribute dont_touch of G25958: signal is true;
	signal G25959: std_logic; attribute dont_touch of G25959: signal is true;
	signal G25960: std_logic; attribute dont_touch of G25960: signal is true;
	signal G25961: std_logic; attribute dont_touch of G25961: signal is true;
	signal G25962: std_logic; attribute dont_touch of G25962: signal is true;
	signal G25963: std_logic; attribute dont_touch of G25963: signal is true;
	signal G25964: std_logic; attribute dont_touch of G25964: signal is true;
	signal G25965: std_logic; attribute dont_touch of G25965: signal is true;
	signal G25966: std_logic; attribute dont_touch of G25966: signal is true;
	signal G25967: std_logic; attribute dont_touch of G25967: signal is true;
	signal G25968: std_logic; attribute dont_touch of G25968: signal is true;
	signal G25969: std_logic; attribute dont_touch of G25969: signal is true;
	signal G25970: std_logic; attribute dont_touch of G25970: signal is true;
	signal G25971: std_logic; attribute dont_touch of G25971: signal is true;
	signal G25972: std_logic; attribute dont_touch of G25972: signal is true;
	signal G25973: std_logic; attribute dont_touch of G25973: signal is true;
	signal G25974: std_logic; attribute dont_touch of G25974: signal is true;
	signal G25975: std_logic; attribute dont_touch of G25975: signal is true;
	signal G25976: std_logic; attribute dont_touch of G25976: signal is true;
	signal G25977: std_logic; attribute dont_touch of G25977: signal is true;
	signal G25978: std_logic; attribute dont_touch of G25978: signal is true;
	signal G25979: std_logic; attribute dont_touch of G25979: signal is true;
	signal G25980: std_logic; attribute dont_touch of G25980: signal is true;
	signal G25981: std_logic; attribute dont_touch of G25981: signal is true;
	signal G25982: std_logic; attribute dont_touch of G25982: signal is true;
	signal G25983: std_logic; attribute dont_touch of G25983: signal is true;
	signal G25984: std_logic; attribute dont_touch of G25984: signal is true;
	signal G25985: std_logic; attribute dont_touch of G25985: signal is true;
	signal G25986: std_logic; attribute dont_touch of G25986: signal is true;
	signal G25987: std_logic; attribute dont_touch of G25987: signal is true;
	signal G25988: std_logic; attribute dont_touch of G25988: signal is true;
	signal G25989: std_logic; attribute dont_touch of G25989: signal is true;
	signal G25990: std_logic; attribute dont_touch of G25990: signal is true;
	signal G25991: std_logic; attribute dont_touch of G25991: signal is true;
	signal G25992: std_logic; attribute dont_touch of G25992: signal is true;
	signal G25993: std_logic; attribute dont_touch of G25993: signal is true;
	signal G25994: std_logic; attribute dont_touch of G25994: signal is true;
	signal G25995: std_logic; attribute dont_touch of G25995: signal is true;
	signal G25996: std_logic; attribute dont_touch of G25996: signal is true;
	signal G25997: std_logic; attribute dont_touch of G25997: signal is true;
	signal G26019: std_logic; attribute dont_touch of G26019: signal is true;
	signal G26020: std_logic; attribute dont_touch of G26020: signal is true;
	signal G26021: std_logic; attribute dont_touch of G26021: signal is true;
	signal G26022: std_logic; attribute dont_touch of G26022: signal is true;
	signal G26023: std_logic; attribute dont_touch of G26023: signal is true;
	signal G26024: std_logic; attribute dont_touch of G26024: signal is true;
	signal G26025: std_logic; attribute dont_touch of G26025: signal is true;
	signal G26026: std_logic; attribute dont_touch of G26026: signal is true;
	signal G26048: std_logic; attribute dont_touch of G26048: signal is true;
	signal G26049: std_logic; attribute dont_touch of G26049: signal is true;
	signal G26050: std_logic; attribute dont_touch of G26050: signal is true;
	signal G26051: std_logic; attribute dont_touch of G26051: signal is true;
	signal G26052: std_logic; attribute dont_touch of G26052: signal is true;
	signal G26053: std_logic; attribute dont_touch of G26053: signal is true;
	signal G26054: std_logic; attribute dont_touch of G26054: signal is true;
	signal G26055: std_logic; attribute dont_touch of G26055: signal is true;
	signal G26077: std_logic; attribute dont_touch of G26077: signal is true;
	signal G26078: std_logic; attribute dont_touch of G26078: signal is true;
	signal G26079: std_logic; attribute dont_touch of G26079: signal is true;
	signal G26080: std_logic; attribute dont_touch of G26080: signal is true;
	signal G26081: std_logic; attribute dont_touch of G26081: signal is true;
	signal G26082: std_logic; attribute dont_touch of G26082: signal is true;
	signal G26083: std_logic; attribute dont_touch of G26083: signal is true;
	signal G26084: std_logic; attribute dont_touch of G26084: signal is true;
	signal G26085: std_logic; attribute dont_touch of G26085: signal is true;
	signal G26086: std_logic; attribute dont_touch of G26086: signal is true;
	signal G26087: std_logic; attribute dont_touch of G26087: signal is true;
	signal G26088: std_logic; attribute dont_touch of G26088: signal is true;
	signal G26089: std_logic; attribute dont_touch of G26089: signal is true;
	signal G26090: std_logic; attribute dont_touch of G26090: signal is true;
	signal G26091: std_logic; attribute dont_touch of G26091: signal is true;
	signal G26092: std_logic; attribute dont_touch of G26092: signal is true;
	signal G26093: std_logic; attribute dont_touch of G26093: signal is true;
	signal G26094: std_logic; attribute dont_touch of G26094: signal is true;
	signal G26095: std_logic; attribute dont_touch of G26095: signal is true;
	signal G26096: std_logic; attribute dont_touch of G26096: signal is true;
	signal G26097: std_logic; attribute dont_touch of G26097: signal is true;
	signal G26098: std_logic; attribute dont_touch of G26098: signal is true;
	signal G26099: std_logic; attribute dont_touch of G26099: signal is true;
	signal G26100: std_logic; attribute dont_touch of G26100: signal is true;
	signal G26101: std_logic; attribute dont_touch of G26101: signal is true;
	signal G26102: std_logic; attribute dont_touch of G26102: signal is true;
	signal G26103: std_logic; attribute dont_touch of G26103: signal is true;
	signal G26104: std_logic; attribute dont_touch of G26104: signal is true;
	signal G26105: std_logic; attribute dont_touch of G26105: signal is true;
	signal G26119: std_logic; attribute dont_touch of G26119: signal is true;
	signal G26120: std_logic; attribute dont_touch of G26120: signal is true;
	signal G26121: std_logic; attribute dont_touch of G26121: signal is true;
	signal G26122: std_logic; attribute dont_touch of G26122: signal is true;
	signal G26123: std_logic; attribute dont_touch of G26123: signal is true;
	signal G26124: std_logic; attribute dont_touch of G26124: signal is true;
	signal G26125: std_logic; attribute dont_touch of G26125: signal is true;
	signal G26126: std_logic; attribute dont_touch of G26126: signal is true;
	signal G26127: std_logic; attribute dont_touch of G26127: signal is true;
	signal G26128: std_logic; attribute dont_touch of G26128: signal is true;
	signal G26129: std_logic; attribute dont_touch of G26129: signal is true;
	signal G26130: std_logic; attribute dont_touch of G26130: signal is true;
	signal G26131: std_logic; attribute dont_touch of G26131: signal is true;
	signal G26145: std_logic; attribute dont_touch of G26145: signal is true;
	signal G26146: std_logic; attribute dont_touch of G26146: signal is true;
	signal G26147: std_logic; attribute dont_touch of G26147: signal is true;
	signal G26148: std_logic; attribute dont_touch of G26148: signal is true;
	signal G26153: std_logic; attribute dont_touch of G26153: signal is true;
	signal G26154: std_logic; attribute dont_touch of G26154: signal is true;
	signal G26155: std_logic; attribute dont_touch of G26155: signal is true;
	signal G26156: std_logic; attribute dont_touch of G26156: signal is true;
	signal G26157: std_logic; attribute dont_touch of G26157: signal is true;
	signal G26158: std_logic; attribute dont_touch of G26158: signal is true;
	signal G26159: std_logic; attribute dont_touch of G26159: signal is true;
	signal G26160: std_logic; attribute dont_touch of G26160: signal is true;
	signal G26161: std_logic; attribute dont_touch of G26161: signal is true;
	signal G26162: std_logic; attribute dont_touch of G26162: signal is true;
	signal G26165: std_logic; attribute dont_touch of G26165: signal is true;
	signal G26166: std_logic; attribute dont_touch of G26166: signal is true;
	signal G26171: std_logic; attribute dont_touch of G26171: signal is true;
	signal G26176: std_logic; attribute dont_touch of G26176: signal is true;
	signal G26177: std_logic; attribute dont_touch of G26177: signal is true;
	signal G26178: std_logic; attribute dont_touch of G26178: signal is true;
	signal G26179: std_logic; attribute dont_touch of G26179: signal is true;
	signal G26180: std_logic; attribute dont_touch of G26180: signal is true;
	signal G26181: std_logic; attribute dont_touch of G26181: signal is true;
	signal G26182: std_logic; attribute dont_touch of G26182: signal is true;
	signal G26183: std_logic; attribute dont_touch of G26183: signal is true;
	signal G26186: std_logic; attribute dont_touch of G26186: signal is true;
	signal G26187: std_logic; attribute dont_touch of G26187: signal is true;
	signal G26190: std_logic; attribute dont_touch of G26190: signal is true;
	signal G26195: std_logic; attribute dont_touch of G26195: signal is true;
	signal G26200: std_logic; attribute dont_touch of G26200: signal is true;
	signal G26203: std_logic; attribute dont_touch of G26203: signal is true;
	signal G26204: std_logic; attribute dont_touch of G26204: signal is true;
	signal G26205: std_logic; attribute dont_touch of G26205: signal is true;
	signal G26206: std_logic; attribute dont_touch of G26206: signal is true;
	signal G26207: std_logic; attribute dont_touch of G26207: signal is true;
	signal G26208: std_logic; attribute dont_touch of G26208: signal is true;
	signal G26209: std_logic; attribute dont_touch of G26209: signal is true;
	signal G26212: std_logic; attribute dont_touch of G26212: signal is true;
	signal G26213: std_logic; attribute dont_touch of G26213: signal is true;
	signal G26218: std_logic; attribute dont_touch of G26218: signal is true;
	signal G26223: std_logic; attribute dont_touch of G26223: signal is true;
	signal G26226: std_logic; attribute dont_touch of G26226: signal is true;
	signal G26229: std_logic; attribute dont_touch of G26229: signal is true;
	signal G26230: std_logic; attribute dont_touch of G26230: signal is true;
	signal G26231: std_logic; attribute dont_touch of G26231: signal is true;
	signal G26232: std_logic; attribute dont_touch of G26232: signal is true;
	signal G26233: std_logic; attribute dont_touch of G26233: signal is true;
	signal G26234: std_logic; attribute dont_touch of G26234: signal is true;
	signal G26235: std_logic; attribute dont_touch of G26235: signal is true;
	signal G26236: std_logic; attribute dont_touch of G26236: signal is true;
	signal G26241: std_logic; attribute dont_touch of G26241: signal is true;
	signal G26244: std_logic; attribute dont_touch of G26244: signal is true;
	signal G26247: std_logic; attribute dont_touch of G26247: signal is true;
	signal G26248: std_logic; attribute dont_touch of G26248: signal is true;
	signal G26249: std_logic; attribute dont_touch of G26249: signal is true;
	signal G26250: std_logic; attribute dont_touch of G26250: signal is true;
	signal G26251: std_logic; attribute dont_touch of G26251: signal is true;
	signal G26252: std_logic; attribute dont_touch of G26252: signal is true;
	signal G26253: std_logic; attribute dont_touch of G26253: signal is true;
	signal G26254: std_logic; attribute dont_touch of G26254: signal is true;
	signal G26255: std_logic; attribute dont_touch of G26255: signal is true;
	signal G26256: std_logic; attribute dont_touch of G26256: signal is true;
	signal G26257: std_logic; attribute dont_touch of G26257: signal is true;
	signal G26258: std_logic; attribute dont_touch of G26258: signal is true;
	signal G26259: std_logic; attribute dont_touch of G26259: signal is true;
	signal G26260: std_logic; attribute dont_touch of G26260: signal is true;
	signal G26261: std_logic; attribute dont_touch of G26261: signal is true;
	signal G26264: std_logic; attribute dont_touch of G26264: signal is true;
	signal G26267: std_logic; attribute dont_touch of G26267: signal is true;
	signal G26268: std_logic; attribute dont_touch of G26268: signal is true;
	signal G26269: std_logic; attribute dont_touch of G26269: signal is true;
	signal G26270: std_logic; attribute dont_touch of G26270: signal is true;
	signal G26271: std_logic; attribute dont_touch of G26271: signal is true;
	signal G26272: std_logic; attribute dont_touch of G26272: signal is true;
	signal G26273: std_logic; attribute dont_touch of G26273: signal is true;
	signal G26274: std_logic; attribute dont_touch of G26274: signal is true;
	signal G26275: std_logic; attribute dont_touch of G26275: signal is true;
	signal G26276: std_logic; attribute dont_touch of G26276: signal is true;
	signal G26277: std_logic; attribute dont_touch of G26277: signal is true;
	signal G26278: std_logic; attribute dont_touch of G26278: signal is true;
	signal G26279: std_logic; attribute dont_touch of G26279: signal is true;
	signal G26280: std_logic; attribute dont_touch of G26280: signal is true;
	signal G26281: std_logic; attribute dont_touch of G26281: signal is true;
	signal G26284: std_logic; attribute dont_touch of G26284: signal is true;
	signal G26285: std_logic; attribute dont_touch of G26285: signal is true;
	signal G26286: std_logic; attribute dont_touch of G26286: signal is true;
	signal G26287: std_logic; attribute dont_touch of G26287: signal is true;
	signal G26288: std_logic; attribute dont_touch of G26288: signal is true;
	signal G26289: std_logic; attribute dont_touch of G26289: signal is true;
	signal G26290: std_logic; attribute dont_touch of G26290: signal is true;
	signal G26291: std_logic; attribute dont_touch of G26291: signal is true;
	signal G26292: std_logic; attribute dont_touch of G26292: signal is true;
	signal G26293: std_logic; attribute dont_touch of G26293: signal is true;
	signal G26294: std_logic; attribute dont_touch of G26294: signal is true;
	signal G26295: std_logic; attribute dont_touch of G26295: signal is true;
	signal G26296: std_logic; attribute dont_touch of G26296: signal is true;
	signal G26297: std_logic; attribute dont_touch of G26297: signal is true;
	signal G26298: std_logic; attribute dont_touch of G26298: signal is true;
	signal G26299: std_logic; attribute dont_touch of G26299: signal is true;
	signal G26300: std_logic; attribute dont_touch of G26300: signal is true;
	signal G26301: std_logic; attribute dont_touch of G26301: signal is true;
	signal G26302: std_logic; attribute dont_touch of G26302: signal is true;
	signal G26303: std_logic; attribute dont_touch of G26303: signal is true;
	signal G26304: std_logic; attribute dont_touch of G26304: signal is true;
	signal G26305: std_logic; attribute dont_touch of G26305: signal is true;
	signal G26306: std_logic; attribute dont_touch of G26306: signal is true;
	signal G26307: std_logic; attribute dont_touch of G26307: signal is true;
	signal G26308: std_logic; attribute dont_touch of G26308: signal is true;
	signal G26309: std_logic; attribute dont_touch of G26309: signal is true;
	signal G26310: std_logic; attribute dont_touch of G26310: signal is true;
	signal G26311: std_logic; attribute dont_touch of G26311: signal is true;
	signal G26312: std_logic; attribute dont_touch of G26312: signal is true;
	signal G26313: std_logic; attribute dont_touch of G26313: signal is true;
	signal G26314: std_logic; attribute dont_touch of G26314: signal is true;
	signal G26323: std_logic; attribute dont_touch of G26323: signal is true;
	signal G26324: std_logic; attribute dont_touch of G26324: signal is true;
	signal G26325: std_logic; attribute dont_touch of G26325: signal is true;
	signal G26326: std_logic; attribute dont_touch of G26326: signal is true;
	signal G26327: std_logic; attribute dont_touch of G26327: signal is true;
	signal G26328: std_logic; attribute dont_touch of G26328: signal is true;
	signal G26329: std_logic; attribute dont_touch of G26329: signal is true;
	signal G26330: std_logic; attribute dont_touch of G26330: signal is true;
	signal G26334: std_logic; attribute dont_touch of G26334: signal is true;
	signal G26335: std_logic; attribute dont_touch of G26335: signal is true;
	signal G26336: std_logic; attribute dont_touch of G26336: signal is true;
	signal G26337: std_logic; attribute dont_touch of G26337: signal is true;
	signal G26338: std_logic; attribute dont_touch of G26338: signal is true;
	signal G26339: std_logic; attribute dont_touch of G26339: signal is true;
	signal G26340: std_logic; attribute dont_touch of G26340: signal is true;
	signal G26341: std_logic; attribute dont_touch of G26341: signal is true;
	signal G26342: std_logic; attribute dont_touch of G26342: signal is true;
	signal G26343: std_logic; attribute dont_touch of G26343: signal is true;
	signal G26344: std_logic; attribute dont_touch of G26344: signal is true;
	signal G26345: std_logic; attribute dont_touch of G26345: signal is true;
	signal G26346: std_logic; attribute dont_touch of G26346: signal is true;
	signal G26347: std_logic; attribute dont_touch of G26347: signal is true;
	signal G26348: std_logic; attribute dont_touch of G26348: signal is true;
	signal G26349: std_logic; attribute dont_touch of G26349: signal is true;
	signal G26350: std_logic; attribute dont_touch of G26350: signal is true;
	signal G26351: std_logic; attribute dont_touch of G26351: signal is true;
	signal G26352: std_logic; attribute dont_touch of G26352: signal is true;
	signal G26356: std_logic; attribute dont_touch of G26356: signal is true;
	signal G26357: std_logic; attribute dont_touch of G26357: signal is true;
	signal G26358: std_logic; attribute dont_touch of G26358: signal is true;
	signal G26359: std_logic; attribute dont_touch of G26359: signal is true;
	signal G26360: std_logic; attribute dont_touch of G26360: signal is true;
	signal G26361: std_logic; attribute dont_touch of G26361: signal is true;
	signal G26362: std_logic; attribute dont_touch of G26362: signal is true;
	signal G26363: std_logic; attribute dont_touch of G26363: signal is true;
	signal G26364: std_logic; attribute dont_touch of G26364: signal is true;
	signal G26365: std_logic; attribute dont_touch of G26365: signal is true;
	signal G26377: std_logic; attribute dont_touch of G26377: signal is true;
	signal G26378: std_logic; attribute dont_touch of G26378: signal is true;
	signal G26379: std_logic; attribute dont_touch of G26379: signal is true;
	signal G26380: std_logic; attribute dont_touch of G26380: signal is true;
	signal G26381: std_logic; attribute dont_touch of G26381: signal is true;
	signal G26382: std_logic; attribute dont_touch of G26382: signal is true;
	signal G26386: std_logic; attribute dont_touch of G26386: signal is true;
	signal G26387: std_logic; attribute dont_touch of G26387: signal is true;
	signal G26388: std_logic; attribute dont_touch of G26388: signal is true;
	signal G26389: std_logic; attribute dont_touch of G26389: signal is true;
	signal G26390: std_logic; attribute dont_touch of G26390: signal is true;
	signal G26391: std_logic; attribute dont_touch of G26391: signal is true;
	signal G26392: std_logic; attribute dont_touch of G26392: signal is true;
	signal G26393: std_logic; attribute dont_touch of G26393: signal is true;
	signal G26394: std_logic; attribute dont_touch of G26394: signal is true;
	signal G26395: std_logic; attribute dont_touch of G26395: signal is true;
	signal G26396: std_logic; attribute dont_touch of G26396: signal is true;
	signal G26397: std_logic; attribute dont_touch of G26397: signal is true;
	signal G26398: std_logic; attribute dont_touch of G26398: signal is true;
	signal G26399: std_logic; attribute dont_touch of G26399: signal is true;
	signal G26400: std_logic; attribute dont_touch of G26400: signal is true;
	signal G26422: std_logic; attribute dont_touch of G26422: signal is true;
	signal G26423: std_logic; attribute dont_touch of G26423: signal is true;
	signal G26424: std_logic; attribute dont_touch of G26424: signal is true;
	signal G26483: std_logic; attribute dont_touch of G26483: signal is true;
	signal G26484: std_logic; attribute dont_touch of G26484: signal is true;
	signal G26485: std_logic; attribute dont_touch of G26485: signal is true;
	signal G26486: std_logic; attribute dont_touch of G26486: signal is true;
	signal G26487: std_logic; attribute dont_touch of G26487: signal is true;
	signal G26488: std_logic; attribute dont_touch of G26488: signal is true;
	signal G26510: std_logic; attribute dont_touch of G26510: signal is true;
	signal G26511: std_logic; attribute dont_touch of G26511: signal is true;
	signal G26512: std_logic; attribute dont_touch of G26512: signal is true;
	signal G26513: std_logic; attribute dont_touch of G26513: signal is true;
	signal G26514: std_logic; attribute dont_touch of G26514: signal is true;
	signal G26515: std_logic; attribute dont_touch of G26515: signal is true;
	signal G26516: std_logic; attribute dont_touch of G26516: signal is true;
	signal G26517: std_logic; attribute dont_touch of G26517: signal is true;
	signal G26518: std_logic; attribute dont_touch of G26518: signal is true;
	signal G26519: std_logic; attribute dont_touch of G26519: signal is true;
	signal G26541: std_logic; attribute dont_touch of G26541: signal is true;
	signal G26542: std_logic; attribute dont_touch of G26542: signal is true;
	signal G26543: std_logic; attribute dont_touch of G26543: signal is true;
	signal G26544: std_logic; attribute dont_touch of G26544: signal is true;
	signal G26545: std_logic; attribute dont_touch of G26545: signal is true;
	signal G26546: std_logic; attribute dont_touch of G26546: signal is true;
	signal G26547: std_logic; attribute dont_touch of G26547: signal is true;
	signal G26548: std_logic; attribute dont_touch of G26548: signal is true;
	signal G26549: std_logic; attribute dont_touch of G26549: signal is true;
	signal G26571: std_logic; attribute dont_touch of G26571: signal is true;
	signal G26572: std_logic; attribute dont_touch of G26572: signal is true;
	signal G26573: std_logic; attribute dont_touch of G26573: signal is true;
	signal G26574: std_logic; attribute dont_touch of G26574: signal is true;
	signal G26575: std_logic; attribute dont_touch of G26575: signal is true;
	signal G26576: std_logic; attribute dont_touch of G26576: signal is true;
	signal G26598: std_logic; attribute dont_touch of G26598: signal is true;
	signal G26602: std_logic; attribute dont_touch of G26602: signal is true;
	signal G26603: std_logic; attribute dont_touch of G26603: signal is true;
	signal G26604: std_logic; attribute dont_touch of G26604: signal is true;
	signal G26605: std_logic; attribute dont_touch of G26605: signal is true;
	signal G26606: std_logic; attribute dont_touch of G26606: signal is true;
	signal G26607: std_logic; attribute dont_touch of G26607: signal is true;
	signal G26608: std_logic; attribute dont_touch of G26608: signal is true;
	signal G26609: std_logic; attribute dont_touch of G26609: signal is true;
	signal G26610: std_logic; attribute dont_touch of G26610: signal is true;
	signal G26611: std_logic; attribute dont_touch of G26611: signal is true;
	signal G26612: std_logic; attribute dont_touch of G26612: signal is true;
	signal G26613: std_logic; attribute dont_touch of G26613: signal is true;
	signal G26614: std_logic; attribute dont_touch of G26614: signal is true;
	signal G26615: std_logic; attribute dont_touch of G26615: signal is true;
	signal G26616: std_logic; attribute dont_touch of G26616: signal is true;
	signal G26625: std_logic; attribute dont_touch of G26625: signal is true;
	signal G26628: std_logic; attribute dont_touch of G26628: signal is true;
	signal G26629: std_logic; attribute dont_touch of G26629: signal is true;
	signal G26630: std_logic; attribute dont_touch of G26630: signal is true;
	signal G26631: std_logic; attribute dont_touch of G26631: signal is true;
	signal G26632: std_logic; attribute dont_touch of G26632: signal is true;
	signal G26633: std_logic; attribute dont_touch of G26633: signal is true;
	signal G26634: std_logic; attribute dont_touch of G26634: signal is true;
	signal G26635: std_logic; attribute dont_touch of G26635: signal is true;
	signal G26636: std_logic; attribute dont_touch of G26636: signal is true;
	signal G26645: std_logic; attribute dont_touch of G26645: signal is true;
	signal G26648: std_logic; attribute dont_touch of G26648: signal is true;
	signal G26649: std_logic; attribute dont_touch of G26649: signal is true;
	signal G26650: std_logic; attribute dont_touch of G26650: signal is true;
	signal G26651: std_logic; attribute dont_touch of G26651: signal is true;
	signal G26652: std_logic; attribute dont_touch of G26652: signal is true;
	signal G26653: std_logic; attribute dont_touch of G26653: signal is true;
	signal G26654: std_logic; attribute dont_touch of G26654: signal is true;
	signal G26655: std_logic; attribute dont_touch of G26655: signal is true;
	signal G26656: std_logic; attribute dont_touch of G26656: signal is true;
	signal G26657: std_logic; attribute dont_touch of G26657: signal is true;
	signal G26666: std_logic; attribute dont_touch of G26666: signal is true;
	signal G26667: std_logic; attribute dont_touch of G26667: signal is true;
	signal G26670: std_logic; attribute dont_touch of G26670: signal is true;
	signal G26671: std_logic; attribute dont_touch of G26671: signal is true;
	signal G26672: std_logic; attribute dont_touch of G26672: signal is true;
	signal G26673: std_logic; attribute dont_touch of G26673: signal is true;
	signal G26679: std_logic; attribute dont_touch of G26679: signal is true;
	signal G26680: std_logic; attribute dont_touch of G26680: signal is true;
	signal G26681: std_logic; attribute dont_touch of G26681: signal is true;
	signal G26682: std_logic; attribute dont_touch of G26682: signal is true;
	signal G26683: std_logic; attribute dont_touch of G26683: signal is true;
	signal G26684: std_logic; attribute dont_touch of G26684: signal is true;
	signal G26685: std_logic; attribute dont_touch of G26685: signal is true;
	signal G26686: std_logic; attribute dont_touch of G26686: signal is true;
	signal G26689: std_logic; attribute dont_touch of G26689: signal is true;
	signal G26690: std_logic; attribute dont_touch of G26690: signal is true;
	signal G26693: std_logic; attribute dont_touch of G26693: signal is true;
	signal G26694: std_logic; attribute dont_touch of G26694: signal is true;
	signal G26700: std_logic; attribute dont_touch of G26700: signal is true;
	signal G26701: std_logic; attribute dont_touch of G26701: signal is true;
	signal G26702: std_logic; attribute dont_touch of G26702: signal is true;
	signal G26703: std_logic; attribute dont_touch of G26703: signal is true;
	signal G26709: std_logic; attribute dont_touch of G26709: signal is true;
	signal G26710: std_logic; attribute dont_touch of G26710: signal is true;
	signal G26711: std_logic; attribute dont_touch of G26711: signal is true;
	signal G26712: std_logic; attribute dont_touch of G26712: signal is true;
	signal G26713: std_logic; attribute dont_touch of G26713: signal is true;
	signal G26714: std_logic; attribute dont_touch of G26714: signal is true;
	signal G26715: std_logic; attribute dont_touch of G26715: signal is true;
	signal G26718: std_logic; attribute dont_touch of G26718: signal is true;
	signal G26719: std_logic; attribute dont_touch of G26719: signal is true;
	signal G26720: std_logic; attribute dont_touch of G26720: signal is true;
	signal G26721: std_logic; attribute dont_touch of G26721: signal is true;
	signal G26724: std_logic; attribute dont_touch of G26724: signal is true;
	signal G26725: std_logic; attribute dont_touch of G26725: signal is true;
	signal G26731: std_logic; attribute dont_touch of G26731: signal is true;
	signal G26732: std_logic; attribute dont_touch of G26732: signal is true;
	signal G26733: std_logic; attribute dont_touch of G26733: signal is true;
	signal G26736: std_logic; attribute dont_touch of G26736: signal is true;
	signal G26737: std_logic; attribute dont_touch of G26737: signal is true;
	signal G26743: std_logic; attribute dont_touch of G26743: signal is true;
	signal G26744: std_logic; attribute dont_touch of G26744: signal is true;
	signal G26745: std_logic; attribute dont_touch of G26745: signal is true;
	signal G26749: std_logic; attribute dont_touch of G26749: signal is true;
	signal G26750: std_logic; attribute dont_touch of G26750: signal is true;
	signal G26751: std_logic; attribute dont_touch of G26751: signal is true;
	signal G26752: std_logic; attribute dont_touch of G26752: signal is true;
	signal G26753: std_logic; attribute dont_touch of G26753: signal is true;
	signal G26754: std_logic; attribute dont_touch of G26754: signal is true;
	signal G26755: std_logic; attribute dont_touch of G26755: signal is true;
	signal G26758: std_logic; attribute dont_touch of G26758: signal is true;
	signal G26759: std_logic; attribute dont_touch of G26759: signal is true;
	signal G26765: std_logic; attribute dont_touch of G26765: signal is true;
	signal G26766: std_logic; attribute dont_touch of G26766: signal is true;
	signal G26769: std_logic; attribute dont_touch of G26769: signal is true;
	signal G26770: std_logic; attribute dont_touch of G26770: signal is true;
	signal G26776: std_logic; attribute dont_touch of G26776: signal is true;
	signal G26777: std_logic; attribute dont_touch of G26777: signal is true;
	signal G26778: std_logic; attribute dont_touch of G26778: signal is true;
	signal G26779: std_logic; attribute dont_touch of G26779: signal is true;
	signal G26780: std_logic; attribute dont_touch of G26780: signal is true;
	signal G26781: std_logic; attribute dont_touch of G26781: signal is true;
	signal G26782: std_logic; attribute dont_touch of G26782: signal is true;
	signal G26783: std_logic; attribute dont_touch of G26783: signal is true;
	signal G26784: std_logic; attribute dont_touch of G26784: signal is true;
	signal G26785: std_logic; attribute dont_touch of G26785: signal is true;
	signal G26788: std_logic; attribute dont_touch of G26788: signal is true;
	signal G26789: std_logic; attribute dont_touch of G26789: signal is true;
	signal G26792: std_logic; attribute dont_touch of G26792: signal is true;
	signal G26793: std_logic; attribute dont_touch of G26793: signal is true;
	signal G26799: std_logic; attribute dont_touch of G26799: signal is true;
	signal G26800: std_logic; attribute dont_touch of G26800: signal is true;
	signal G26802: std_logic; attribute dont_touch of G26802: signal is true;
	signal G26803: std_logic; attribute dont_touch of G26803: signal is true;
	signal G26804: std_logic; attribute dont_touch of G26804: signal is true;
	signal G26805: std_logic; attribute dont_touch of G26805: signal is true;
	signal G26808: std_logic; attribute dont_touch of G26808: signal is true;
	signal G26809: std_logic; attribute dont_touch of G26809: signal is true;
	signal G26810: std_logic; attribute dont_touch of G26810: signal is true;
	signal G26811: std_logic; attribute dont_touch of G26811: signal is true;
	signal G26812: std_logic; attribute dont_touch of G26812: signal is true;
	signal G26813: std_logic; attribute dont_touch of G26813: signal is true;
	signal G26814: std_logic; attribute dont_touch of G26814: signal is true;
	signal G26815: std_logic; attribute dont_touch of G26815: signal is true;
	signal G26816: std_logic; attribute dont_touch of G26816: signal is true;
	signal G26817: std_logic; attribute dont_touch of G26817: signal is true;
	signal G26818: std_logic; attribute dont_touch of G26818: signal is true;
	signal G26819: std_logic; attribute dont_touch of G26819: signal is true;
	signal G26820: std_logic; attribute dont_touch of G26820: signal is true;
	signal G26821: std_logic; attribute dont_touch of G26821: signal is true;
	signal G26822: std_logic; attribute dont_touch of G26822: signal is true;
	signal G26823: std_logic; attribute dont_touch of G26823: signal is true;
	signal G26824: std_logic; attribute dont_touch of G26824: signal is true;
	signal G26825: std_logic; attribute dont_touch of G26825: signal is true;
	signal G26826: std_logic; attribute dont_touch of G26826: signal is true;
	signal G26827: std_logic; attribute dont_touch of G26827: signal is true;
	signal G26828: std_logic; attribute dont_touch of G26828: signal is true;
	signal G26829: std_logic; attribute dont_touch of G26829: signal is true;
	signal G26830: std_logic; attribute dont_touch of G26830: signal is true;
	signal G26831: std_logic; attribute dont_touch of G26831: signal is true;
	signal G26832: std_logic; attribute dont_touch of G26832: signal is true;
	signal G26833: std_logic; attribute dont_touch of G26833: signal is true;
	signal G26834: std_logic; attribute dont_touch of G26834: signal is true;
	signal G26835: std_logic; attribute dont_touch of G26835: signal is true;
	signal G26836: std_logic; attribute dont_touch of G26836: signal is true;
	signal G26837: std_logic; attribute dont_touch of G26837: signal is true;
	signal G26838: std_logic; attribute dont_touch of G26838: signal is true;
	signal G26839: std_logic; attribute dont_touch of G26839: signal is true;
	signal G26840: std_logic; attribute dont_touch of G26840: signal is true;
	signal G26841: std_logic; attribute dont_touch of G26841: signal is true;
	signal G26842: std_logic; attribute dont_touch of G26842: signal is true;
	signal G26843: std_logic; attribute dont_touch of G26843: signal is true;
	signal G26844: std_logic; attribute dont_touch of G26844: signal is true;
	signal G26845: std_logic; attribute dont_touch of G26845: signal is true;
	signal G26846: std_logic; attribute dont_touch of G26846: signal is true;
	signal G26847: std_logic; attribute dont_touch of G26847: signal is true;
	signal G26848: std_logic; attribute dont_touch of G26848: signal is true;
	signal G26849: std_logic; attribute dont_touch of G26849: signal is true;
	signal G26850: std_logic; attribute dont_touch of G26850: signal is true;
	signal G26851: std_logic; attribute dont_touch of G26851: signal is true;
	signal G26852: std_logic; attribute dont_touch of G26852: signal is true;
	signal G26853: std_logic; attribute dont_touch of G26853: signal is true;
	signal G26854: std_logic; attribute dont_touch of G26854: signal is true;
	signal G26855: std_logic; attribute dont_touch of G26855: signal is true;
	signal G26856: std_logic; attribute dont_touch of G26856: signal is true;
	signal G26857: std_logic; attribute dont_touch of G26857: signal is true;
	signal G26858: std_logic; attribute dont_touch of G26858: signal is true;
	signal G26859: std_logic; attribute dont_touch of G26859: signal is true;
	signal G26860: std_logic; attribute dont_touch of G26860: signal is true;
	signal G26861: std_logic; attribute dont_touch of G26861: signal is true;
	signal G26862: std_logic; attribute dont_touch of G26862: signal is true;
	signal G26863: std_logic; attribute dont_touch of G26863: signal is true;
	signal G26864: std_logic; attribute dont_touch of G26864: signal is true;
	signal G26865: std_logic; attribute dont_touch of G26865: signal is true;
	signal G26866: std_logic; attribute dont_touch of G26866: signal is true;
	signal G26869: std_logic; attribute dont_touch of G26869: signal is true;
	signal G26870: std_logic; attribute dont_touch of G26870: signal is true;
	signal G26871: std_logic; attribute dont_touch of G26871: signal is true;
	signal G26872: std_logic; attribute dont_touch of G26872: signal is true;
	signal G26873: std_logic; attribute dont_touch of G26873: signal is true;
	signal G26874: std_logic; attribute dont_touch of G26874: signal is true;
	signal G26878: std_logic; attribute dont_touch of G26878: signal is true;
	signal G26879: std_logic; attribute dont_touch of G26879: signal is true;
	signal G26880: std_logic; attribute dont_touch of G26880: signal is true;
	signal G26881: std_logic; attribute dont_touch of G26881: signal is true;
	signal G26882: std_logic; attribute dont_touch of G26882: signal is true;
	signal G26883: std_logic; attribute dont_touch of G26883: signal is true;
	signal G26884: std_logic; attribute dont_touch of G26884: signal is true;
	signal G26885: std_logic; attribute dont_touch of G26885: signal is true;
	signal G26886: std_logic; attribute dont_touch of G26886: signal is true;
	signal G26887: std_logic; attribute dont_touch of G26887: signal is true;
	signal G26888: std_logic; attribute dont_touch of G26888: signal is true;
	signal G26889: std_logic; attribute dont_touch of G26889: signal is true;
	signal G26890: std_logic; attribute dont_touch of G26890: signal is true;
	signal G26891: std_logic; attribute dont_touch of G26891: signal is true;
	signal G26892: std_logic; attribute dont_touch of G26892: signal is true;
	signal G26893: std_logic; attribute dont_touch of G26893: signal is true;
	signal G26894: std_logic; attribute dont_touch of G26894: signal is true;
	signal G26895: std_logic; attribute dont_touch of G26895: signal is true;
	signal G26896: std_logic; attribute dont_touch of G26896: signal is true;
	signal G26897: std_logic; attribute dont_touch of G26897: signal is true;
	signal G26898: std_logic; attribute dont_touch of G26898: signal is true;
	signal G26899: std_logic; attribute dont_touch of G26899: signal is true;
	signal G26900: std_logic; attribute dont_touch of G26900: signal is true;
	signal G26901: std_logic; attribute dont_touch of G26901: signal is true;
	signal G26902: std_logic; attribute dont_touch of G26902: signal is true;
	signal G26903: std_logic; attribute dont_touch of G26903: signal is true;
	signal G26904: std_logic; attribute dont_touch of G26904: signal is true;
	signal G26905: std_logic; attribute dont_touch of G26905: signal is true;
	signal G26906: std_logic; attribute dont_touch of G26906: signal is true;
	signal G26907: std_logic; attribute dont_touch of G26907: signal is true;
	signal G26908: std_logic; attribute dont_touch of G26908: signal is true;
	signal G26909: std_logic; attribute dont_touch of G26909: signal is true;
	signal G26910: std_logic; attribute dont_touch of G26910: signal is true;
	signal G26911: std_logic; attribute dont_touch of G26911: signal is true;
	signal G26912: std_logic; attribute dont_touch of G26912: signal is true;
	signal G26913: std_logic; attribute dont_touch of G26913: signal is true;
	signal G26914: std_logic; attribute dont_touch of G26914: signal is true;
	signal G26915: std_logic; attribute dont_touch of G26915: signal is true;
	signal G26916: std_logic; attribute dont_touch of G26916: signal is true;
	signal G26917: std_logic; attribute dont_touch of G26917: signal is true;
	signal G26918: std_logic; attribute dont_touch of G26918: signal is true;
	signal G26919: std_logic; attribute dont_touch of G26919: signal is true;
	signal G26920: std_logic; attribute dont_touch of G26920: signal is true;
	signal G26921: std_logic; attribute dont_touch of G26921: signal is true;
	signal G26922: std_logic; attribute dont_touch of G26922: signal is true;
	signal G26923: std_logic; attribute dont_touch of G26923: signal is true;
	signal G26924: std_logic; attribute dont_touch of G26924: signal is true;
	signal G26925: std_logic; attribute dont_touch of G26925: signal is true;
	signal G26926: std_logic; attribute dont_touch of G26926: signal is true;
	signal G26927: std_logic; attribute dont_touch of G26927: signal is true;
	signal G26928: std_logic; attribute dont_touch of G26928: signal is true;
	signal G26929: std_logic; attribute dont_touch of G26929: signal is true;
	signal G26930: std_logic; attribute dont_touch of G26930: signal is true;
	signal G26931: std_logic; attribute dont_touch of G26931: signal is true;
	signal G26932: std_logic; attribute dont_touch of G26932: signal is true;
	signal G26933: std_logic; attribute dont_touch of G26933: signal is true;
	signal G26934: std_logic; attribute dont_touch of G26934: signal is true;
	signal G26935: std_logic; attribute dont_touch of G26935: signal is true;
	signal G26936: std_logic; attribute dont_touch of G26936: signal is true;
	signal G26937: std_logic; attribute dont_touch of G26937: signal is true;
	signal G26938: std_logic; attribute dont_touch of G26938: signal is true;
	signal G26939: std_logic; attribute dont_touch of G26939: signal is true;
	signal G26940: std_logic; attribute dont_touch of G26940: signal is true;
	signal G26941: std_logic; attribute dont_touch of G26941: signal is true;
	signal G26942: std_logic; attribute dont_touch of G26942: signal is true;
	signal G26943: std_logic; attribute dont_touch of G26943: signal is true;
	signal G26944: std_logic; attribute dont_touch of G26944: signal is true;
	signal G26945: std_logic; attribute dont_touch of G26945: signal is true;
	signal G26946: std_logic; attribute dont_touch of G26946: signal is true;
	signal G26947: std_logic; attribute dont_touch of G26947: signal is true;
	signal G26948: std_logic; attribute dont_touch of G26948: signal is true;
	signal G26949: std_logic; attribute dont_touch of G26949: signal is true;
	signal G26950: std_logic; attribute dont_touch of G26950: signal is true;
	signal G26951: std_logic; attribute dont_touch of G26951: signal is true;
	signal G26952: std_logic; attribute dont_touch of G26952: signal is true;
	signal G26953: std_logic; attribute dont_touch of G26953: signal is true;
	signal G26954: std_logic; attribute dont_touch of G26954: signal is true;
	signal G26955: std_logic; attribute dont_touch of G26955: signal is true;
	signal G26956: std_logic; attribute dont_touch of G26956: signal is true;
	signal G26957: std_logic; attribute dont_touch of G26957: signal is true;
	signal G26958: std_logic; attribute dont_touch of G26958: signal is true;
	signal G26959: std_logic; attribute dont_touch of G26959: signal is true;
	signal G26960: std_logic; attribute dont_touch of G26960: signal is true;
	signal G26961: std_logic; attribute dont_touch of G26961: signal is true;
	signal G26962: std_logic; attribute dont_touch of G26962: signal is true;
	signal G26963: std_logic; attribute dont_touch of G26963: signal is true;
	signal G26964: std_logic; attribute dont_touch of G26964: signal is true;
	signal G26965: std_logic; attribute dont_touch of G26965: signal is true;
	signal G26966: std_logic; attribute dont_touch of G26966: signal is true;
	signal G26967: std_logic; attribute dont_touch of G26967: signal is true;
	signal G26968: std_logic; attribute dont_touch of G26968: signal is true;
	signal G26969: std_logic; attribute dont_touch of G26969: signal is true;
	signal G26970: std_logic; attribute dont_touch of G26970: signal is true;
	signal G26971: std_logic; attribute dont_touch of G26971: signal is true;
	signal G26972: std_logic; attribute dont_touch of G26972: signal is true;
	signal G26973: std_logic; attribute dont_touch of G26973: signal is true;
	signal G26976: std_logic; attribute dont_touch of G26976: signal is true;
	signal G26977: std_logic; attribute dont_touch of G26977: signal is true;
	signal G26987: std_logic; attribute dont_touch of G26987: signal is true;
	signal G26990: std_logic; attribute dont_touch of G26990: signal is true;
	signal G26993: std_logic; attribute dont_touch of G26993: signal is true;
	signal G26994: std_logic; attribute dont_touch of G26994: signal is true;
	signal G27004: std_logic; attribute dont_touch of G27004: signal is true;
	signal G27007: std_logic; attribute dont_touch of G27007: signal is true;
	signal G27008: std_logic; attribute dont_touch of G27008: signal is true;
	signal G27009: std_logic; attribute dont_touch of G27009: signal is true;
	signal G27010: std_logic; attribute dont_touch of G27010: signal is true;
	signal G27011: std_logic; attribute dont_touch of G27011: signal is true;
	signal G27012: std_logic; attribute dont_touch of G27012: signal is true;
	signal G27013: std_logic; attribute dont_touch of G27013: signal is true;
	signal G27014: std_logic; attribute dont_touch of G27014: signal is true;
	signal G27015: std_logic; attribute dont_touch of G27015: signal is true;
	signal G27016: std_logic; attribute dont_touch of G27016: signal is true;
	signal G27017: std_logic; attribute dont_touch of G27017: signal is true;
	signal G27018: std_logic; attribute dont_touch of G27018: signal is true;
	signal G27019: std_logic; attribute dont_touch of G27019: signal is true;
	signal G27020: std_logic; attribute dont_touch of G27020: signal is true;
	signal G27024: std_logic; attribute dont_touch of G27024: signal is true;
	signal G27025: std_logic; attribute dont_touch of G27025: signal is true;
	signal G27026: std_logic; attribute dont_touch of G27026: signal is true;
	signal G27027: std_logic; attribute dont_touch of G27027: signal is true;
	signal G27028: std_logic; attribute dont_touch of G27028: signal is true;
	signal G27029: std_logic; attribute dont_touch of G27029: signal is true;
	signal G27030: std_logic; attribute dont_touch of G27030: signal is true;
	signal G27031: std_logic; attribute dont_touch of G27031: signal is true;
	signal G27032: std_logic; attribute dont_touch of G27032: signal is true;
	signal G27033: std_logic; attribute dont_touch of G27033: signal is true;
	signal G27034: std_logic; attribute dont_touch of G27034: signal is true;
	signal G27035: std_logic; attribute dont_touch of G27035: signal is true;
	signal G27036: std_logic; attribute dont_touch of G27036: signal is true;
	signal G27037: std_logic; attribute dont_touch of G27037: signal is true;
	signal G27038: std_logic; attribute dont_touch of G27038: signal is true;
	signal G27039: std_logic; attribute dont_touch of G27039: signal is true;
	signal G27040: std_logic; attribute dont_touch of G27040: signal is true;
	signal G27041: std_logic; attribute dont_touch of G27041: signal is true;
	signal G27042: std_logic; attribute dont_touch of G27042: signal is true;
	signal G27043: std_logic; attribute dont_touch of G27043: signal is true;
	signal G27044: std_logic; attribute dont_touch of G27044: signal is true;
	signal G27045: std_logic; attribute dont_touch of G27045: signal is true;
	signal G27046: std_logic; attribute dont_touch of G27046: signal is true;
	signal G27050: std_logic; attribute dont_touch of G27050: signal is true;
	signal G27051: std_logic; attribute dont_touch of G27051: signal is true;
	signal G27057: std_logic; attribute dont_touch of G27057: signal is true;
	signal G27058: std_logic; attribute dont_touch of G27058: signal is true;
	signal G27059: std_logic; attribute dont_touch of G27059: signal is true;
	signal G27063: std_logic; attribute dont_touch of G27063: signal is true;
	signal G27064: std_logic; attribute dont_touch of G27064: signal is true;
	signal G27073: std_logic; attribute dont_touch of G27073: signal is true;
	signal G27074: std_logic; attribute dont_touch of G27074: signal is true;
	signal G27083: std_logic; attribute dont_touch of G27083: signal is true;
	signal G27084: std_logic; attribute dont_touch of G27084: signal is true;
	signal G27085: std_logic; attribute dont_touch of G27085: signal is true;
	signal G27086: std_logic; attribute dont_touch of G27086: signal is true;
	signal G27087: std_logic; attribute dont_touch of G27087: signal is true;
	signal G27088: std_logic; attribute dont_touch of G27088: signal is true;
	signal G27089: std_logic; attribute dont_touch of G27089: signal is true;
	signal G27090: std_logic; attribute dont_touch of G27090: signal is true;
	signal G27091: std_logic; attribute dont_touch of G27091: signal is true;
	signal G27092: std_logic; attribute dont_touch of G27092: signal is true;
	signal G27093: std_logic; attribute dont_touch of G27093: signal is true;
	signal G27094: std_logic; attribute dont_touch of G27094: signal is true;
	signal G27095: std_logic; attribute dont_touch of G27095: signal is true;
	signal G27096: std_logic; attribute dont_touch of G27096: signal is true;
	signal G27097: std_logic; attribute dont_touch of G27097: signal is true;
	signal G27098: std_logic; attribute dont_touch of G27098: signal is true;
	signal G27099: std_logic; attribute dont_touch of G27099: signal is true;
	signal G27100: std_logic; attribute dont_touch of G27100: signal is true;
	signal G27101: std_logic; attribute dont_touch of G27101: signal is true;
	signal G27102: std_logic; attribute dont_touch of G27102: signal is true;
	signal G27103: std_logic; attribute dont_touch of G27103: signal is true;
	signal G27104: std_logic; attribute dont_touch of G27104: signal is true;
	signal G27105: std_logic; attribute dont_touch of G27105: signal is true;
	signal G27106: std_logic; attribute dont_touch of G27106: signal is true;
	signal G27107: std_logic; attribute dont_touch of G27107: signal is true;
	signal G27108: std_logic; attribute dont_touch of G27108: signal is true;
	signal G27112: std_logic; attribute dont_touch of G27112: signal is true;
	signal G27113: std_logic; attribute dont_touch of G27113: signal is true;
	signal G27114: std_logic; attribute dont_touch of G27114: signal is true;
	signal G27115: std_logic; attribute dont_touch of G27115: signal is true;
	signal G27116: std_logic; attribute dont_touch of G27116: signal is true;
	signal G27117: std_logic; attribute dont_touch of G27117: signal is true;
	signal G27118: std_logic; attribute dont_touch of G27118: signal is true;
	signal G27119: std_logic; attribute dont_touch of G27119: signal is true;
	signal G27120: std_logic; attribute dont_touch of G27120: signal is true;
	signal G27121: std_logic; attribute dont_touch of G27121: signal is true;
	signal G27122: std_logic; attribute dont_touch of G27122: signal is true;
	signal G27126: std_logic; attribute dont_touch of G27126: signal is true;
	signal G27127: std_logic; attribute dont_touch of G27127: signal is true;
	signal G27128: std_logic; attribute dont_touch of G27128: signal is true;
	signal G27129: std_logic; attribute dont_touch of G27129: signal is true;
	signal G27130: std_logic; attribute dont_touch of G27130: signal is true;
	signal G27131: std_logic; attribute dont_touch of G27131: signal is true;
	signal G27132: std_logic; attribute dont_touch of G27132: signal is true;
	signal G27133: std_logic; attribute dont_touch of G27133: signal is true;
	signal G27134: std_logic; attribute dont_touch of G27134: signal is true;
	signal G27135: std_logic; attribute dont_touch of G27135: signal is true;
	signal G27136: std_logic; attribute dont_touch of G27136: signal is true;
	signal G27137: std_logic; attribute dont_touch of G27137: signal is true;
	signal G27138: std_logic; attribute dont_touch of G27138: signal is true;
	signal G27139: std_logic; attribute dont_touch of G27139: signal is true;
	signal G27140: std_logic; attribute dont_touch of G27140: signal is true;
	signal G27141: std_logic; attribute dont_touch of G27141: signal is true;
	signal G27142: std_logic; attribute dont_touch of G27142: signal is true;
	signal G27145: std_logic; attribute dont_touch of G27145: signal is true;
	signal G27146: std_logic; attribute dont_touch of G27146: signal is true;
	signal G27147: std_logic; attribute dont_touch of G27147: signal is true;
	signal G27148: std_logic; attribute dont_touch of G27148: signal is true;
	signal G27149: std_logic; attribute dont_touch of G27149: signal is true;
	signal G27150: std_logic; attribute dont_touch of G27150: signal is true;
	signal G27151: std_logic; attribute dont_touch of G27151: signal is true;
	signal G27152: std_logic; attribute dont_touch of G27152: signal is true;
	signal G27153: std_logic; attribute dont_touch of G27153: signal is true;
	signal G27154: std_logic; attribute dont_touch of G27154: signal is true;
	signal G27155: std_logic; attribute dont_touch of G27155: signal is true;
	signal G27158: std_logic; attribute dont_touch of G27158: signal is true;
	signal G27159: std_logic; attribute dont_touch of G27159: signal is true;
	signal G27160: std_logic; attribute dont_touch of G27160: signal is true;
	signal G27161: std_logic; attribute dont_touch of G27161: signal is true;
	signal G27162: std_logic; attribute dont_touch of G27162: signal is true;
	signal G27163: std_logic; attribute dont_touch of G27163: signal is true;
	signal G27177: std_logic; attribute dont_touch of G27177: signal is true;
	signal G27178: std_logic; attribute dont_touch of G27178: signal is true;
	signal G27179: std_logic; attribute dont_touch of G27179: signal is true;
	signal G27180: std_logic; attribute dont_touch of G27180: signal is true;
	signal G27181: std_logic; attribute dont_touch of G27181: signal is true;
	signal G27182: std_logic; attribute dont_touch of G27182: signal is true;
	signal G27183: std_logic; attribute dont_touch of G27183: signal is true;
	signal G27184: std_logic; attribute dont_touch of G27184: signal is true;
	signal G27185: std_logic; attribute dont_touch of G27185: signal is true;
	signal G27186: std_logic; attribute dont_touch of G27186: signal is true;
	signal G27187: std_logic; attribute dont_touch of G27187: signal is true;
	signal G27201: std_logic; attribute dont_touch of G27201: signal is true;
	signal G27202: std_logic; attribute dont_touch of G27202: signal is true;
	signal G27203: std_logic; attribute dont_touch of G27203: signal is true;
	signal G27204: std_logic; attribute dont_touch of G27204: signal is true;
	signal G27205: std_logic; attribute dont_touch of G27205: signal is true;
	signal G27206: std_logic; attribute dont_touch of G27206: signal is true;
	signal G27207: std_logic; attribute dont_touch of G27207: signal is true;
	signal G27208: std_logic; attribute dont_touch of G27208: signal is true;
	signal G27209: std_logic; attribute dont_touch of G27209: signal is true;
	signal G27210: std_logic; attribute dont_touch of G27210: signal is true;
	signal G27211: std_logic; attribute dont_touch of G27211: signal is true;
	signal G27212: std_logic; attribute dont_touch of G27212: signal is true;
	signal G27213: std_logic; attribute dont_touch of G27213: signal is true;
	signal G27214: std_logic; attribute dont_touch of G27214: signal is true;
	signal G27215: std_logic; attribute dont_touch of G27215: signal is true;
	signal G27216: std_logic; attribute dont_touch of G27216: signal is true;
	signal G27217: std_logic; attribute dont_touch of G27217: signal is true;
	signal G27218: std_logic; attribute dont_touch of G27218: signal is true;
	signal G27219: std_logic; attribute dont_touch of G27219: signal is true;
	signal G27220: std_logic; attribute dont_touch of G27220: signal is true;
	signal G27221: std_logic; attribute dont_touch of G27221: signal is true;
	signal G27222: std_logic; attribute dont_touch of G27222: signal is true;
	signal G27223: std_logic; attribute dont_touch of G27223: signal is true;
	signal G27224: std_logic; attribute dont_touch of G27224: signal is true;
	signal G27225: std_logic; attribute dont_touch of G27225: signal is true;
	signal G27226: std_logic; attribute dont_touch of G27226: signal is true;
	signal G27227: std_logic; attribute dont_touch of G27227: signal is true;
	signal G27228: std_logic; attribute dont_touch of G27228: signal is true;
	signal G27229: std_logic; attribute dont_touch of G27229: signal is true;
	signal G27230: std_logic; attribute dont_touch of G27230: signal is true;
	signal G27231: std_logic; attribute dont_touch of G27231: signal is true;
	signal G27232: std_logic; attribute dont_touch of G27232: signal is true;
	signal G27233: std_logic; attribute dont_touch of G27233: signal is true;
	signal G27234: std_logic; attribute dont_touch of G27234: signal is true;
	signal G27235: std_logic; attribute dont_touch of G27235: signal is true;
	signal G27236: std_logic; attribute dont_touch of G27236: signal is true;
	signal G27237: std_logic; attribute dont_touch of G27237: signal is true;
	signal G27238: std_logic; attribute dont_touch of G27238: signal is true;
	signal G27239: std_logic; attribute dont_touch of G27239: signal is true;
	signal G27240: std_logic; attribute dont_touch of G27240: signal is true;
	signal G27241: std_logic; attribute dont_touch of G27241: signal is true;
	signal G27242: std_logic; attribute dont_touch of G27242: signal is true;
	signal G27243: std_logic; attribute dont_touch of G27243: signal is true;
	signal G27244: std_logic; attribute dont_touch of G27244: signal is true;
	signal G27245: std_logic; attribute dont_touch of G27245: signal is true;
	signal G27246: std_logic; attribute dont_touch of G27246: signal is true;
	signal G27247: std_logic; attribute dont_touch of G27247: signal is true;
	signal G27248: std_logic; attribute dont_touch of G27248: signal is true;
	signal G27249: std_logic; attribute dont_touch of G27249: signal is true;
	signal G27250: std_logic; attribute dont_touch of G27250: signal is true;
	signal G27251: std_logic; attribute dont_touch of G27251: signal is true;
	signal G27252: std_logic; attribute dont_touch of G27252: signal is true;
	signal G27253: std_logic; attribute dont_touch of G27253: signal is true;
	signal G27254: std_logic; attribute dont_touch of G27254: signal is true;
	signal G27255: std_logic; attribute dont_touch of G27255: signal is true;
	signal G27256: std_logic; attribute dont_touch of G27256: signal is true;
	signal G27257: std_logic; attribute dont_touch of G27257: signal is true;
	signal G27258: std_logic; attribute dont_touch of G27258: signal is true;
	signal G27259: std_logic; attribute dont_touch of G27259: signal is true;
	signal G27260: std_logic; attribute dont_touch of G27260: signal is true;
	signal G27261: std_logic; attribute dont_touch of G27261: signal is true;
	signal G27262: std_logic; attribute dont_touch of G27262: signal is true;
	signal G27263: std_logic; attribute dont_touch of G27263: signal is true;
	signal G27264: std_logic; attribute dont_touch of G27264: signal is true;
	signal G27265: std_logic; attribute dont_touch of G27265: signal is true;
	signal G27266: std_logic; attribute dont_touch of G27266: signal is true;
	signal G27267: std_logic; attribute dont_touch of G27267: signal is true;
	signal G27268: std_logic; attribute dont_touch of G27268: signal is true;
	signal G27269: std_logic; attribute dont_touch of G27269: signal is true;
	signal G27270: std_logic; attribute dont_touch of G27270: signal is true;
	signal G27271: std_logic; attribute dont_touch of G27271: signal is true;
	signal G27272: std_logic; attribute dont_touch of G27272: signal is true;
	signal G27273: std_logic; attribute dont_touch of G27273: signal is true;
	signal G27274: std_logic; attribute dont_touch of G27274: signal is true;
	signal G27275: std_logic; attribute dont_touch of G27275: signal is true;
	signal G27276: std_logic; attribute dont_touch of G27276: signal is true;
	signal G27277: std_logic; attribute dont_touch of G27277: signal is true;
	signal G27278: std_logic; attribute dont_touch of G27278: signal is true;
	signal G27279: std_logic; attribute dont_touch of G27279: signal is true;
	signal G27280: std_logic; attribute dont_touch of G27280: signal is true;
	signal G27281: std_logic; attribute dont_touch of G27281: signal is true;
	signal G27282: std_logic; attribute dont_touch of G27282: signal is true;
	signal G27283: std_logic; attribute dont_touch of G27283: signal is true;
	signal G27284: std_logic; attribute dont_touch of G27284: signal is true;
	signal G27285: std_logic; attribute dont_touch of G27285: signal is true;
	signal G27286: std_logic; attribute dont_touch of G27286: signal is true;
	signal G27287: std_logic; attribute dont_touch of G27287: signal is true;
	signal G27288: std_logic; attribute dont_touch of G27288: signal is true;
	signal G27289: std_logic; attribute dont_touch of G27289: signal is true;
	signal G27290: std_logic; attribute dont_touch of G27290: signal is true;
	signal G27291: std_logic; attribute dont_touch of G27291: signal is true;
	signal G27292: std_logic; attribute dont_touch of G27292: signal is true;
	signal G27293: std_logic; attribute dont_touch of G27293: signal is true;
	signal G27294: std_logic; attribute dont_touch of G27294: signal is true;
	signal G27295: std_logic; attribute dont_touch of G27295: signal is true;
	signal G27298: std_logic; attribute dont_touch of G27298: signal is true;
	signal G27299: std_logic; attribute dont_touch of G27299: signal is true;
	signal G27300: std_logic; attribute dont_touch of G27300: signal is true;
	signal G27301: std_logic; attribute dont_touch of G27301: signal is true;
	signal G27302: std_logic; attribute dont_touch of G27302: signal is true;
	signal G27303: std_logic; attribute dont_touch of G27303: signal is true;
	signal G27304: std_logic; attribute dont_touch of G27304: signal is true;
	signal G27305: std_logic; attribute dont_touch of G27305: signal is true;
	signal G27306: std_logic; attribute dont_touch of G27306: signal is true;
	signal G27309: std_logic; attribute dont_touch of G27309: signal is true;
	signal G27310: std_logic; attribute dont_touch of G27310: signal is true;
	signal G27311: std_logic; attribute dont_touch of G27311: signal is true;
	signal G27312: std_logic; attribute dont_touch of G27312: signal is true;
	signal G27313: std_logic; attribute dont_touch of G27313: signal is true;
	signal G27314: std_logic; attribute dont_touch of G27314: signal is true;
	signal G27315: std_logic; attribute dont_touch of G27315: signal is true;
	signal G27316: std_logic; attribute dont_touch of G27316: signal is true;
	signal G27317: std_logic; attribute dont_touch of G27317: signal is true;
	signal G27320: std_logic; attribute dont_touch of G27320: signal is true;
	signal G27323: std_logic; attribute dont_touch of G27323: signal is true;
	signal G27324: std_logic; attribute dont_touch of G27324: signal is true;
	signal G27325: std_logic; attribute dont_touch of G27325: signal is true;
	signal G27326: std_logic; attribute dont_touch of G27326: signal is true;
	signal G27327: std_logic; attribute dont_touch of G27327: signal is true;
	signal G27328: std_logic; attribute dont_touch of G27328: signal is true;
	signal G27329: std_logic; attribute dont_touch of G27329: signal is true;
	signal G27330: std_logic; attribute dont_touch of G27330: signal is true;
	signal G27331: std_logic; attribute dont_touch of G27331: signal is true;
	signal G27332: std_logic; attribute dont_touch of G27332: signal is true;
	signal G27333: std_logic; attribute dont_touch of G27333: signal is true;
	signal G27334: std_logic; attribute dont_touch of G27334: signal is true;
	signal G27335: std_logic; attribute dont_touch of G27335: signal is true;
	signal G27336: std_logic; attribute dont_touch of G27336: signal is true;
	signal G27337: std_logic; attribute dont_touch of G27337: signal is true;
	signal G27338: std_logic; attribute dont_touch of G27338: signal is true;
	signal G27339: std_logic; attribute dont_touch of G27339: signal is true;
	signal G27340: std_logic; attribute dont_touch of G27340: signal is true;
	signal G27341: std_logic; attribute dont_touch of G27341: signal is true;
	signal G27342: std_logic; attribute dont_touch of G27342: signal is true;
	signal G27343: std_logic; attribute dont_touch of G27343: signal is true;
	signal G27344: std_logic; attribute dont_touch of G27344: signal is true;
	signal G27345: std_logic; attribute dont_touch of G27345: signal is true;
	signal G27346: std_logic; attribute dont_touch of G27346: signal is true;
	signal G27347: std_logic; attribute dont_touch of G27347: signal is true;
	signal G27348: std_logic; attribute dont_touch of G27348: signal is true;
	signal G27349: std_logic; attribute dont_touch of G27349: signal is true;
	signal G27350: std_logic; attribute dont_touch of G27350: signal is true;
	signal G27351: std_logic; attribute dont_touch of G27351: signal is true;
	signal G27352: std_logic; attribute dont_touch of G27352: signal is true;
	signal G27353: std_logic; attribute dont_touch of G27353: signal is true;
	signal G27354: std_logic; attribute dont_touch of G27354: signal is true;
	signal G27355: std_logic; attribute dont_touch of G27355: signal is true;
	signal G27356: std_logic; attribute dont_touch of G27356: signal is true;
	signal G27357: std_logic; attribute dont_touch of G27357: signal is true;
	signal G27358: std_logic; attribute dont_touch of G27358: signal is true;
	signal G27359: std_logic; attribute dont_touch of G27359: signal is true;
	signal G27360: std_logic; attribute dont_touch of G27360: signal is true;
	signal G27361: std_logic; attribute dont_touch of G27361: signal is true;
	signal G27362: std_logic; attribute dont_touch of G27362: signal is true;
	signal G27363: std_logic; attribute dont_touch of G27363: signal is true;
	signal G27364: std_logic; attribute dont_touch of G27364: signal is true;
	signal G27365: std_logic; attribute dont_touch of G27365: signal is true;
	signal G27366: std_logic; attribute dont_touch of G27366: signal is true;
	signal G27367: std_logic; attribute dont_touch of G27367: signal is true;
	signal G27368: std_logic; attribute dont_touch of G27368: signal is true;
	signal G27369: std_logic; attribute dont_touch of G27369: signal is true;
	signal G27370: std_logic; attribute dont_touch of G27370: signal is true;
	signal G27371: std_logic; attribute dont_touch of G27371: signal is true;
	signal G27372: std_logic; attribute dont_touch of G27372: signal is true;
	signal G27373: std_logic; attribute dont_touch of G27373: signal is true;
	signal G27374: std_logic; attribute dont_touch of G27374: signal is true;
	signal G27375: std_logic; attribute dont_touch of G27375: signal is true;
	signal G27376: std_logic; attribute dont_touch of G27376: signal is true;
	signal G27377: std_logic; attribute dont_touch of G27377: signal is true;
	signal G27378: std_logic; attribute dont_touch of G27378: signal is true;
	signal G27379: std_logic; attribute dont_touch of G27379: signal is true;
	signal G27380: std_logic; attribute dont_touch of G27380: signal is true;
	signal G27381: std_logic; attribute dont_touch of G27381: signal is true;
	signal G27382: std_logic; attribute dont_touch of G27382: signal is true;
	signal G27383: std_logic; attribute dont_touch of G27383: signal is true;
	signal G27384: std_logic; attribute dont_touch of G27384: signal is true;
	signal G27385: std_logic; attribute dont_touch of G27385: signal is true;
	signal G27386: std_logic; attribute dont_touch of G27386: signal is true;
	signal G27387: std_logic; attribute dont_touch of G27387: signal is true;
	signal G27388: std_logic; attribute dont_touch of G27388: signal is true;
	signal G27389: std_logic; attribute dont_touch of G27389: signal is true;
	signal G27390: std_logic; attribute dont_touch of G27390: signal is true;
	signal G27391: std_logic; attribute dont_touch of G27391: signal is true;
	signal G27392: std_logic; attribute dont_touch of G27392: signal is true;
	signal G27393: std_logic; attribute dont_touch of G27393: signal is true;
	signal G27394: std_logic; attribute dont_touch of G27394: signal is true;
	signal G27395: std_logic; attribute dont_touch of G27395: signal is true;
	signal G27400: std_logic; attribute dont_touch of G27400: signal is true;
	signal G27401: std_logic; attribute dont_touch of G27401: signal is true;
	signal G27402: std_logic; attribute dont_touch of G27402: signal is true;
	signal G27403: std_logic; attribute dont_touch of G27403: signal is true;
	signal G27404: std_logic; attribute dont_touch of G27404: signal is true;
	signal G27405: std_logic; attribute dont_touch of G27405: signal is true;
	signal G27406: std_logic; attribute dont_touch of G27406: signal is true;
	signal G27407: std_logic; attribute dont_touch of G27407: signal is true;
	signal G27408: std_logic; attribute dont_touch of G27408: signal is true;
	signal G27409: std_logic; attribute dont_touch of G27409: signal is true;
	signal G27410: std_logic; attribute dont_touch of G27410: signal is true;
	signal G27411: std_logic; attribute dont_touch of G27411: signal is true;
	signal G27412: std_logic; attribute dont_touch of G27412: signal is true;
	signal G27413: std_logic; attribute dont_touch of G27413: signal is true;
	signal G27414: std_logic; attribute dont_touch of G27414: signal is true;
	signal G27415: std_logic; attribute dont_touch of G27415: signal is true;
	signal G27416: std_logic; attribute dont_touch of G27416: signal is true;
	signal G27421: std_logic; attribute dont_touch of G27421: signal is true;
	signal G27426: std_logic; attribute dont_touch of G27426: signal is true;
	signal G27427: std_logic; attribute dont_touch of G27427: signal is true;
	signal G27428: std_logic; attribute dont_touch of G27428: signal is true;
	signal G27429: std_logic; attribute dont_touch of G27429: signal is true;
	signal G27430: std_logic; attribute dont_touch of G27430: signal is true;
	signal G27431: std_logic; attribute dont_touch of G27431: signal is true;
	signal G27432: std_logic; attribute dont_touch of G27432: signal is true;
	signal G27433: std_logic; attribute dont_touch of G27433: signal is true;
	signal G27434: std_logic; attribute dont_touch of G27434: signal is true;
	signal G27435: std_logic; attribute dont_touch of G27435: signal is true;
	signal G27436: std_logic; attribute dont_touch of G27436: signal is true;
	signal G27437: std_logic; attribute dont_touch of G27437: signal is true;
	signal G27438: std_logic; attribute dont_touch of G27438: signal is true;
	signal G27439: std_logic; attribute dont_touch of G27439: signal is true;
	signal G27440: std_logic; attribute dont_touch of G27440: signal is true;
	signal G27445: std_logic; attribute dont_touch of G27445: signal is true;
	signal G27450: std_logic; attribute dont_touch of G27450: signal is true;
	signal G27451: std_logic; attribute dont_touch of G27451: signal is true;
	signal G27452: std_logic; attribute dont_touch of G27452: signal is true;
	signal G27453: std_logic; attribute dont_touch of G27453: signal is true;
	signal G27454: std_logic; attribute dont_touch of G27454: signal is true;
	signal G27455: std_logic; attribute dont_touch of G27455: signal is true;
	signal G27456: std_logic; attribute dont_touch of G27456: signal is true;
	signal G27457: std_logic; attribute dont_touch of G27457: signal is true;
	signal G27458: std_logic; attribute dont_touch of G27458: signal is true;
	signal G27459: std_logic; attribute dont_touch of G27459: signal is true;
	signal G27460: std_logic; attribute dont_touch of G27460: signal is true;
	signal G27461: std_logic; attribute dont_touch of G27461: signal is true;
	signal G27462: std_logic; attribute dont_touch of G27462: signal is true;
	signal G27463: std_logic; attribute dont_touch of G27463: signal is true;
	signal G27467: std_logic; attribute dont_touch of G27467: signal is true;
	signal G27468: std_logic; attribute dont_touch of G27468: signal is true;
	signal G27469: std_logic; attribute dont_touch of G27469: signal is true;
	signal G27474: std_logic; attribute dont_touch of G27474: signal is true;
	signal G27479: std_logic; attribute dont_touch of G27479: signal is true;
	signal G27480: std_logic; attribute dont_touch of G27480: signal is true;
	signal G27481: std_logic; attribute dont_touch of G27481: signal is true;
	signal G27482: std_logic; attribute dont_touch of G27482: signal is true;
	signal G27483: std_logic; attribute dont_touch of G27483: signal is true;
	signal G27484: std_logic; attribute dont_touch of G27484: signal is true;
	signal G27485: std_logic; attribute dont_touch of G27485: signal is true;
	signal G27486: std_logic; attribute dont_touch of G27486: signal is true;
	signal G27487: std_logic; attribute dont_touch of G27487: signal is true;
	signal G27488: std_logic; attribute dont_touch of G27488: signal is true;
	signal G27489: std_logic; attribute dont_touch of G27489: signal is true;
	signal G27490: std_logic; attribute dont_touch of G27490: signal is true;
	signal G27491: std_logic; attribute dont_touch of G27491: signal is true;
	signal G27492: std_logic; attribute dont_touch of G27492: signal is true;
	signal G27493: std_logic; attribute dont_touch of G27493: signal is true;
	signal G27494: std_logic; attribute dont_touch of G27494: signal is true;
	signal G27499: std_logic; attribute dont_touch of G27499: signal is true;
	signal G27500: std_logic; attribute dont_touch of G27500: signal is true;
	signal G27501: std_logic; attribute dont_touch of G27501: signal is true;
	signal G27502: std_logic; attribute dont_touch of G27502: signal is true;
	signal G27503: std_logic; attribute dont_touch of G27503: signal is true;
	signal G27504: std_logic; attribute dont_touch of G27504: signal is true;
	signal G27505: std_logic; attribute dont_touch of G27505: signal is true;
	signal G27506: std_logic; attribute dont_touch of G27506: signal is true;
	signal G27507: std_logic; attribute dont_touch of G27507: signal is true;
	signal G27508: std_logic; attribute dont_touch of G27508: signal is true;
	signal G27509: std_logic; attribute dont_touch of G27509: signal is true;
	signal G27510: std_logic; attribute dont_touch of G27510: signal is true;
	signal G27511: std_logic; attribute dont_touch of G27511: signal is true;
	signal G27515: std_logic; attribute dont_touch of G27515: signal is true;
	signal G27516: std_logic; attribute dont_touch of G27516: signal is true;
	signal G27517: std_logic; attribute dont_touch of G27517: signal is true;
	signal G27518: std_logic; attribute dont_touch of G27518: signal is true;
	signal G27519: std_logic; attribute dont_touch of G27519: signal is true;
	signal G27520: std_logic; attribute dont_touch of G27520: signal is true;
	signal G27521: std_logic; attribute dont_touch of G27521: signal is true;
	signal G27522: std_logic; attribute dont_touch of G27522: signal is true;
	signal G27523: std_logic; attribute dont_touch of G27523: signal is true;
	signal G27524: std_logic; attribute dont_touch of G27524: signal is true;
	signal G27525: std_logic; attribute dont_touch of G27525: signal is true;
	signal G27526: std_logic; attribute dont_touch of G27526: signal is true;
	signal G27527: std_logic; attribute dont_touch of G27527: signal is true;
	signal G27528: std_logic; attribute dont_touch of G27528: signal is true;
	signal G27532: std_logic; attribute dont_touch of G27532: signal is true;
	signal G27533: std_logic; attribute dont_touch of G27533: signal is true;
	signal G27534: std_logic; attribute dont_touch of G27534: signal is true;
	signal G27535: std_logic; attribute dont_touch of G27535: signal is true;
	signal G27536: std_logic; attribute dont_touch of G27536: signal is true;
	signal G27537: std_logic; attribute dont_touch of G27537: signal is true;
	signal G27538: std_logic; attribute dont_touch of G27538: signal is true;
	signal G27539: std_logic; attribute dont_touch of G27539: signal is true;
	signal G27540: std_logic; attribute dont_touch of G27540: signal is true;
	signal G27541: std_logic; attribute dont_touch of G27541: signal is true;
	signal G27542: std_logic; attribute dont_touch of G27542: signal is true;
	signal G27543: std_logic; attribute dont_touch of G27543: signal is true;
	signal G27544: std_logic; attribute dont_touch of G27544: signal is true;
	signal G27545: std_logic; attribute dont_touch of G27545: signal is true;
	signal G27546: std_logic; attribute dont_touch of G27546: signal is true;
	signal G27547: std_logic; attribute dont_touch of G27547: signal is true;
	signal G27548: std_logic; attribute dont_touch of G27548: signal is true;
	signal G27549: std_logic; attribute dont_touch of G27549: signal is true;
	signal G27550: std_logic; attribute dont_touch of G27550: signal is true;
	signal G27551: std_logic; attribute dont_touch of G27551: signal is true;
	signal G27552: std_logic; attribute dont_touch of G27552: signal is true;
	signal G27553: std_logic; attribute dont_touch of G27553: signal is true;
	signal G27554: std_logic; attribute dont_touch of G27554: signal is true;
	signal G27555: std_logic; attribute dont_touch of G27555: signal is true;
	signal G27556: std_logic; attribute dont_touch of G27556: signal is true;
	signal G27557: std_logic; attribute dont_touch of G27557: signal is true;
	signal G27558: std_logic; attribute dont_touch of G27558: signal is true;
	signal G27559: std_logic; attribute dont_touch of G27559: signal is true;
	signal G27560: std_logic; attribute dont_touch of G27560: signal is true;
	signal G27561: std_logic; attribute dont_touch of G27561: signal is true;
	signal G27562: std_logic; attribute dont_touch of G27562: signal is true;
	signal G27563: std_logic; attribute dont_touch of G27563: signal is true;
	signal G27564: std_logic; attribute dont_touch of G27564: signal is true;
	signal G27565: std_logic; attribute dont_touch of G27565: signal is true;
	signal G27566: std_logic; attribute dont_touch of G27566: signal is true;
	signal G27567: std_logic; attribute dont_touch of G27567: signal is true;
	signal G27568: std_logic; attribute dont_touch of G27568: signal is true;
	signal G27569: std_logic; attribute dont_touch of G27569: signal is true;
	signal G27570: std_logic; attribute dont_touch of G27570: signal is true;
	signal G27571: std_logic; attribute dont_touch of G27571: signal is true;
	signal G27572: std_logic; attribute dont_touch of G27572: signal is true;
	signal G27573: std_logic; attribute dont_touch of G27573: signal is true;
	signal G27574: std_logic; attribute dont_touch of G27574: signal is true;
	signal G27575: std_logic; attribute dont_touch of G27575: signal is true;
	signal G27576: std_logic; attribute dont_touch of G27576: signal is true;
	signal G27577: std_logic; attribute dont_touch of G27577: signal is true;
	signal G27578: std_logic; attribute dont_touch of G27578: signal is true;
	signal G27579: std_logic; attribute dont_touch of G27579: signal is true;
	signal G27580: std_logic; attribute dont_touch of G27580: signal is true;
	signal G27581: std_logic; attribute dont_touch of G27581: signal is true;
	signal G27582: std_logic; attribute dont_touch of G27582: signal is true;
	signal G27583: std_logic; attribute dont_touch of G27583: signal is true;
	signal G27584: std_logic; attribute dont_touch of G27584: signal is true;
	signal G27585: std_logic; attribute dont_touch of G27585: signal is true;
	signal G27586: std_logic; attribute dont_touch of G27586: signal is true;
	signal G27587: std_logic; attribute dont_touch of G27587: signal is true;
	signal G27588: std_logic; attribute dont_touch of G27588: signal is true;
	signal G27589: std_logic; attribute dont_touch of G27589: signal is true;
	signal G27590: std_logic; attribute dont_touch of G27590: signal is true;
	signal G27591: std_logic; attribute dont_touch of G27591: signal is true;
	signal G27592: std_logic; attribute dont_touch of G27592: signal is true;
	signal G27593: std_logic; attribute dont_touch of G27593: signal is true;
	signal G27594: std_logic; attribute dont_touch of G27594: signal is true;
	signal G27595: std_logic; attribute dont_touch of G27595: signal is true;
	signal G27596: std_logic; attribute dont_touch of G27596: signal is true;
	signal G27597: std_logic; attribute dont_touch of G27597: signal is true;
	signal G27598: std_logic; attribute dont_touch of G27598: signal is true;
	signal G27599: std_logic; attribute dont_touch of G27599: signal is true;
	signal G27600: std_logic; attribute dont_touch of G27600: signal is true;
	signal G27601: std_logic; attribute dont_touch of G27601: signal is true;
	signal G27602: std_logic; attribute dont_touch of G27602: signal is true;
	signal G27612: std_logic; attribute dont_touch of G27612: signal is true;
	signal G27613: std_logic; attribute dont_touch of G27613: signal is true;
	signal G27614: std_logic; attribute dont_touch of G27614: signal is true;
	signal G27615: std_logic; attribute dont_touch of G27615: signal is true;
	signal G27616: std_logic; attribute dont_touch of G27616: signal is true;
	signal G27617: std_logic; attribute dont_touch of G27617: signal is true;
	signal G27627: std_logic; attribute dont_touch of G27627: signal is true;
	signal G27628: std_logic; attribute dont_touch of G27628: signal is true;
	signal G27629: std_logic; attribute dont_touch of G27629: signal is true;
	signal G27633: std_logic; attribute dont_touch of G27633: signal is true;
	signal G27634: std_logic; attribute dont_touch of G27634: signal is true;
	signal G27635: std_logic; attribute dont_touch of G27635: signal is true;
	signal G27645: std_logic; attribute dont_touch of G27645: signal is true;
	signal G27646: std_logic; attribute dont_touch of G27646: signal is true;
	signal G27647: std_logic; attribute dont_touch of G27647: signal is true;
	signal G27648: std_logic; attribute dont_touch of G27648: signal is true;
	signal G27649: std_logic; attribute dont_touch of G27649: signal is true;
	signal G27650: std_logic; attribute dont_touch of G27650: signal is true;
	signal G27651: std_logic; attribute dont_touch of G27651: signal is true;
	signal G27652: std_logic; attribute dont_touch of G27652: signal is true;
	signal G27653: std_logic; attribute dont_touch of G27653: signal is true;
	signal G27654: std_logic; attribute dont_touch of G27654: signal is true;
	signal G27658: std_logic; attribute dont_touch of G27658: signal is true;
	signal G27659: std_logic; attribute dont_touch of G27659: signal is true;
	signal G27660: std_logic; attribute dont_touch of G27660: signal is true;
	signal G27661: std_logic; attribute dont_touch of G27661: signal is true;
	signal G27662: std_logic; attribute dont_touch of G27662: signal is true;
	signal G27663: std_logic; attribute dont_touch of G27663: signal is true;
	signal G27664: std_logic; attribute dont_touch of G27664: signal is true;
	signal G27665: std_logic; attribute dont_touch of G27665: signal is true;
	signal G27666: std_logic; attribute dont_touch of G27666: signal is true;
	signal G27667: std_logic; attribute dont_touch of G27667: signal is true;
	signal G27668: std_logic; attribute dont_touch of G27668: signal is true;
	signal G27669: std_logic; attribute dont_touch of G27669: signal is true;
	signal G27670: std_logic; attribute dont_touch of G27670: signal is true;
	signal G27673: std_logic; attribute dont_touch of G27673: signal is true;
	signal G27674: std_logic; attribute dont_touch of G27674: signal is true;
	signal G27675: std_logic; attribute dont_touch of G27675: signal is true;
	signal G27676: std_logic; attribute dont_touch of G27676: signal is true;
	signal G27677: std_logic; attribute dont_touch of G27677: signal is true;
	signal G27678: std_logic; attribute dont_touch of G27678: signal is true;
	signal G27679: std_logic; attribute dont_touch of G27679: signal is true;
	signal G27682: std_logic; attribute dont_touch of G27682: signal is true;
	signal G27683: std_logic; attribute dont_touch of G27683: signal is true;
	signal G27684: std_logic; attribute dont_touch of G27684: signal is true;
	signal G27685: std_logic; attribute dont_touch of G27685: signal is true;
	signal G27686: std_logic; attribute dont_touch of G27686: signal is true;
	signal G27687: std_logic; attribute dont_touch of G27687: signal is true;
	signal G27690: std_logic; attribute dont_touch of G27690: signal is true;
	signal G27691: std_logic; attribute dont_touch of G27691: signal is true;
	signal G27692: std_logic; attribute dont_touch of G27692: signal is true;
	signal G27693: std_logic; attribute dont_touch of G27693: signal is true;
	signal G27696: std_logic; attribute dont_touch of G27696: signal is true;
	signal G27697: std_logic; attribute dont_touch of G27697: signal is true;
	signal G27698: std_logic; attribute dont_touch of G27698: signal is true;
	signal G27699: std_logic; attribute dont_touch of G27699: signal is true;
	signal G27700: std_logic; attribute dont_touch of G27700: signal is true;
	signal G27703: std_logic; attribute dont_touch of G27703: signal is true;
	signal G27704: std_logic; attribute dont_touch of G27704: signal is true;
	signal G27705: std_logic; attribute dont_touch of G27705: signal is true;
	signal G27708: std_logic; attribute dont_touch of G27708: signal is true;
	signal G27709: std_logic; attribute dont_touch of G27709: signal is true;
	signal G27710: std_logic; attribute dont_touch of G27710: signal is true;
	signal G27711: std_logic; attribute dont_touch of G27711: signal is true;
	signal G27714: std_logic; attribute dont_touch of G27714: signal is true;
	signal G27717: std_logic; attribute dont_touch of G27717: signal is true;
	signal G27720: std_logic; attribute dont_touch of G27720: signal is true;
	signal G27721: std_logic; attribute dont_touch of G27721: signal is true;
	signal G27722: std_logic; attribute dont_touch of G27722: signal is true;
	signal G27723: std_logic; attribute dont_touch of G27723: signal is true;
	signal G27724: std_logic; attribute dont_touch of G27724: signal is true;
	signal G27727: std_logic; attribute dont_touch of G27727: signal is true;
	signal G27730: std_logic; attribute dont_touch of G27730: signal is true;
	signal G27731: std_logic; attribute dont_touch of G27731: signal is true;
	signal G27732: std_logic; attribute dont_touch of G27732: signal is true;
	signal G27733: std_logic; attribute dont_touch of G27733: signal is true;
	signal G27734: std_logic; attribute dont_touch of G27734: signal is true;
	signal G27735: std_logic; attribute dont_touch of G27735: signal is true;
	signal G27736: std_logic; attribute dont_touch of G27736: signal is true;
	signal G27737: std_logic; attribute dont_touch of G27737: signal is true;
	signal G27738: std_logic; attribute dont_touch of G27738: signal is true;
	signal G27742: std_logic; attribute dont_touch of G27742: signal is true;
	signal G27759: std_logic; attribute dont_touch of G27759: signal is true;
	signal G27762: std_logic; attribute dont_touch of G27762: signal is true;
	signal G27765: std_logic; attribute dont_touch of G27765: signal is true;
	signal G27766: std_logic; attribute dont_touch of G27766: signal is true;
	signal G27767: std_logic; attribute dont_touch of G27767: signal is true;
	signal G27768: std_logic; attribute dont_touch of G27768: signal is true;
	signal G27769: std_logic; attribute dont_touch of G27769: signal is true;
	signal G27770: std_logic; attribute dont_touch of G27770: signal is true;
	signal G27771: std_logic; attribute dont_touch of G27771: signal is true;
	signal G27772: std_logic; attribute dont_touch of G27772: signal is true;
	signal G27773: std_logic; attribute dont_touch of G27773: signal is true;
	signal G27774: std_logic; attribute dont_touch of G27774: signal is true;
	signal G27775: std_logic; attribute dont_touch of G27775: signal is true;
	signal G27779: std_logic; attribute dont_touch of G27779: signal is true;
	signal G27796: std_logic; attribute dont_touch of G27796: signal is true;
	signal G27800: std_logic; attribute dont_touch of G27800: signal is true;
	signal G27817: std_logic; attribute dont_touch of G27817: signal is true;
	signal G27820: std_logic; attribute dont_touch of G27820: signal is true;
	signal G27821: std_logic; attribute dont_touch of G27821: signal is true;
	signal G27822: std_logic; attribute dont_touch of G27822: signal is true;
	signal G27823: std_logic; attribute dont_touch of G27823: signal is true;
	signal G27824: std_logic; attribute dont_touch of G27824: signal is true;
	signal G27825: std_logic; attribute dont_touch of G27825: signal is true;
	signal G27826: std_logic; attribute dont_touch of G27826: signal is true;
	signal G27827: std_logic; attribute dont_touch of G27827: signal is true;
	signal G27828: std_logic; attribute dont_touch of G27828: signal is true;
	signal G27829: std_logic; attribute dont_touch of G27829: signal is true;
	signal G27830: std_logic; attribute dont_touch of G27830: signal is true;
	signal G27832: std_logic; attribute dont_touch of G27832: signal is true;
	signal G27833: std_logic; attribute dont_touch of G27833: signal is true;
	signal G27837: std_logic; attribute dont_touch of G27837: signal is true;
	signal G27854: std_logic; attribute dont_touch of G27854: signal is true;
	signal G27858: std_logic; attribute dont_touch of G27858: signal is true;
	signal G27875: std_logic; attribute dont_touch of G27875: signal is true;
	signal G27876: std_logic; attribute dont_touch of G27876: signal is true;
	signal G27877: std_logic; attribute dont_touch of G27877: signal is true;
	signal G27878: std_logic; attribute dont_touch of G27878: signal is true;
	signal G27879: std_logic; attribute dont_touch of G27879: signal is true;
	signal G27880: std_logic; attribute dont_touch of G27880: signal is true;
	signal G27881: std_logic; attribute dont_touch of G27881: signal is true;
	signal G27882: std_logic; attribute dont_touch of G27882: signal is true;
	signal G27886: std_logic; attribute dont_touch of G27886: signal is true;
	signal G27903: std_logic; attribute dont_touch of G27903: signal is true;
	signal G27907: std_logic; attribute dont_touch of G27907: signal is true;
	signal G27924: std_logic; attribute dont_touch of G27924: signal is true;
	signal G27925: std_logic; attribute dont_touch of G27925: signal is true;
	signal G27926: std_logic; attribute dont_touch of G27926: signal is true;
	signal G27927: std_logic; attribute dont_touch of G27927: signal is true;
	signal G27928: std_logic; attribute dont_touch of G27928: signal is true;
	signal G27929: std_logic; attribute dont_touch of G27929: signal is true;
	signal G27930: std_logic; attribute dont_touch of G27930: signal is true;
	signal G27931: std_logic; attribute dont_touch of G27931: signal is true;
	signal G27932: std_logic; attribute dont_touch of G27932: signal is true;
	signal G27933: std_logic; attribute dont_touch of G27933: signal is true;
	signal G27937: std_logic; attribute dont_touch of G27937: signal is true;
	signal G27954: std_logic; attribute dont_touch of G27954: signal is true;
	signal G27955: std_logic; attribute dont_touch of G27955: signal is true;
	signal G27956: std_logic; attribute dont_touch of G27956: signal is true;
	signal G27957: std_logic; attribute dont_touch of G27957: signal is true;
	signal G27958: std_logic; attribute dont_touch of G27958: signal is true;
	signal G27959: std_logic; attribute dont_touch of G27959: signal is true;
	signal G27960: std_logic; attribute dont_touch of G27960: signal is true;
	signal G27961: std_logic; attribute dont_touch of G27961: signal is true;
	signal G27962: std_logic; attribute dont_touch of G27962: signal is true;
	signal G27963: std_logic; attribute dont_touch of G27963: signal is true;
	signal G27964: std_logic; attribute dont_touch of G27964: signal is true;
	signal G27965: std_logic; attribute dont_touch of G27965: signal is true;
	signal G27966: std_logic; attribute dont_touch of G27966: signal is true;
	signal G27967: std_logic; attribute dont_touch of G27967: signal is true;
	signal G27968: std_logic; attribute dont_touch of G27968: signal is true;
	signal G27969: std_logic; attribute dont_touch of G27969: signal is true;
	signal G27970: std_logic; attribute dont_touch of G27970: signal is true;
	signal G27971: std_logic; attribute dont_touch of G27971: signal is true;
	signal G27972: std_logic; attribute dont_touch of G27972: signal is true;
	signal G27973: std_logic; attribute dont_touch of G27973: signal is true;
	signal G27974: std_logic; attribute dont_touch of G27974: signal is true;
	signal G27975: std_logic; attribute dont_touch of G27975: signal is true;
	signal G27976: std_logic; attribute dont_touch of G27976: signal is true;
	signal G27977: std_logic; attribute dont_touch of G27977: signal is true;
	signal G27980: std_logic; attribute dont_touch of G27980: signal is true;
	signal G27981: std_logic; attribute dont_touch of G27981: signal is true;
	signal G27982: std_logic; attribute dont_touch of G27982: signal is true;
	signal G27983: std_logic; attribute dont_touch of G27983: signal is true;
	signal G27984: std_logic; attribute dont_touch of G27984: signal is true;
	signal G27985: std_logic; attribute dont_touch of G27985: signal is true;
	signal G27988: std_logic; attribute dont_touch of G27988: signal is true;
	signal G27989: std_logic; attribute dont_touch of G27989: signal is true;
	signal G27990: std_logic; attribute dont_touch of G27990: signal is true;
	signal G27991: std_logic; attribute dont_touch of G27991: signal is true;
	signal G27992: std_logic; attribute dont_touch of G27992: signal is true;
	signal G27993: std_logic; attribute dont_touch of G27993: signal is true;
	signal G27994: std_logic; attribute dont_touch of G27994: signal is true;
	signal G27995: std_logic; attribute dont_touch of G27995: signal is true;
	signal G27996: std_logic; attribute dont_touch of G27996: signal is true;
	signal G27997: std_logic; attribute dont_touch of G27997: signal is true;
	signal G27998: std_logic; attribute dont_touch of G27998: signal is true;
	signal G27999: std_logic; attribute dont_touch of G27999: signal is true;
	signal G28009: std_logic; attribute dont_touch of G28009: signal is true;
	signal G28010: std_logic; attribute dont_touch of G28010: signal is true;
	signal G28020: std_logic; attribute dont_touch of G28020: signal is true;
	signal G28031: std_logic; attribute dont_touch of G28031: signal is true;
	signal G28032: std_logic; attribute dont_touch of G28032: signal is true;
	signal G28033: std_logic; attribute dont_touch of G28033: signal is true;
	signal G28034: std_logic; attribute dont_touch of G28034: signal is true;
	signal G28035: std_logic; attribute dont_touch of G28035: signal is true;
	signal G28036: std_logic; attribute dont_touch of G28036: signal is true;
	signal G28037: std_logic; attribute dont_touch of G28037: signal is true;
	signal G28038: std_logic; attribute dont_touch of G28038: signal is true;
	signal G28039: std_logic; attribute dont_touch of G28039: signal is true;
	signal G28040: std_logic; attribute dont_touch of G28040: signal is true;
	signal G28043: std_logic; attribute dont_touch of G28043: signal is true;
	signal G28044: std_logic; attribute dont_touch of G28044: signal is true;
	signal G28045: std_logic; attribute dont_touch of G28045: signal is true;
	signal G28046: std_logic; attribute dont_touch of G28046: signal is true;
	signal G28047: std_logic; attribute dont_touch of G28047: signal is true;
	signal G28048: std_logic; attribute dont_touch of G28048: signal is true;
	signal G28049: std_logic; attribute dont_touch of G28049: signal is true;
	signal G28050: std_logic; attribute dont_touch of G28050: signal is true;
	signal G28051: std_logic; attribute dont_touch of G28051: signal is true;
	signal G28052: std_logic; attribute dont_touch of G28052: signal is true;
	signal G28053: std_logic; attribute dont_touch of G28053: signal is true;
	signal G28054: std_logic; attribute dont_touch of G28054: signal is true;
	signal G28055: std_logic; attribute dont_touch of G28055: signal is true;
	signal G28056: std_logic; attribute dont_touch of G28056: signal is true;
	signal G28057: std_logic; attribute dont_touch of G28057: signal is true;
	signal G28058: std_logic; attribute dont_touch of G28058: signal is true;
	signal G28059: std_logic; attribute dont_touch of G28059: signal is true;
	signal G28060: std_logic; attribute dont_touch of G28060: signal is true;
	signal G28061: std_logic; attribute dont_touch of G28061: signal is true;
	signal G28062: std_logic; attribute dont_touch of G28062: signal is true;
	signal G28063: std_logic; attribute dont_touch of G28063: signal is true;
	signal G28064: std_logic; attribute dont_touch of G28064: signal is true;
	signal G28065: std_logic; attribute dont_touch of G28065: signal is true;
	signal G28066: std_logic; attribute dont_touch of G28066: signal is true;
	signal G28067: std_logic; attribute dont_touch of G28067: signal is true;
	signal G28068: std_logic; attribute dont_touch of G28068: signal is true;
	signal G28069: std_logic; attribute dont_touch of G28069: signal is true;
	signal G28070: std_logic; attribute dont_touch of G28070: signal is true;
	signal G28071: std_logic; attribute dont_touch of G28071: signal is true;
	signal G28072: std_logic; attribute dont_touch of G28072: signal is true;
	signal G28073: std_logic; attribute dont_touch of G28073: signal is true;
	signal G28074: std_logic; attribute dont_touch of G28074: signal is true;
	signal G28075: std_logic; attribute dont_touch of G28075: signal is true;
	signal G28076: std_logic; attribute dont_touch of G28076: signal is true;
	signal G28077: std_logic; attribute dont_touch of G28077: signal is true;
	signal G28078: std_logic; attribute dont_touch of G28078: signal is true;
	signal G28079: std_logic; attribute dont_touch of G28079: signal is true;
	signal G28080: std_logic; attribute dont_touch of G28080: signal is true;
	signal G28081: std_logic; attribute dont_touch of G28081: signal is true;
	signal G28082: std_logic; attribute dont_touch of G28082: signal is true;
	signal G28083: std_logic; attribute dont_touch of G28083: signal is true;
	signal G28084: std_logic; attribute dont_touch of G28084: signal is true;
	signal G28085: std_logic; attribute dont_touch of G28085: signal is true;
	signal G28086: std_logic; attribute dont_touch of G28086: signal is true;
	signal G28087: std_logic; attribute dont_touch of G28087: signal is true;
	signal G28088: std_logic; attribute dont_touch of G28088: signal is true;
	signal G28089: std_logic; attribute dont_touch of G28089: signal is true;
	signal G28090: std_logic; attribute dont_touch of G28090: signal is true;
	signal G28091: std_logic; attribute dont_touch of G28091: signal is true;
	signal G28092: std_logic; attribute dont_touch of G28092: signal is true;
	signal G28093: std_logic; attribute dont_touch of G28093: signal is true;
	signal G28094: std_logic; attribute dont_touch of G28094: signal is true;
	signal G28095: std_logic; attribute dont_touch of G28095: signal is true;
	signal G28096: std_logic; attribute dont_touch of G28096: signal is true;
	signal G28097: std_logic; attribute dont_touch of G28097: signal is true;
	signal G28098: std_logic; attribute dont_touch of G28098: signal is true;
	signal G28099: std_logic; attribute dont_touch of G28099: signal is true;
	signal G28100: std_logic; attribute dont_touch of G28100: signal is true;
	signal G28101: std_logic; attribute dont_touch of G28101: signal is true;
	signal G28102: std_logic; attribute dont_touch of G28102: signal is true;
	signal G28103: std_logic; attribute dont_touch of G28103: signal is true;
	signal G28104: std_logic; attribute dont_touch of G28104: signal is true;
	signal G28105: std_logic; attribute dont_touch of G28105: signal is true;
	signal G28106: std_logic; attribute dont_touch of G28106: signal is true;
	signal G28107: std_logic; attribute dont_touch of G28107: signal is true;
	signal G28108: std_logic; attribute dont_touch of G28108: signal is true;
	signal G28109: std_logic; attribute dont_touch of G28109: signal is true;
	signal G28110: std_logic; attribute dont_touch of G28110: signal is true;
	signal G28111: std_logic; attribute dont_touch of G28111: signal is true;
	signal G28112: std_logic; attribute dont_touch of G28112: signal is true;
	signal G28113: std_logic; attribute dont_touch of G28113: signal is true;
	signal G28114: std_logic; attribute dont_touch of G28114: signal is true;
	signal G28115: std_logic; attribute dont_touch of G28115: signal is true;
	signal G28116: std_logic; attribute dont_touch of G28116: signal is true;
	signal G28117: std_logic; attribute dont_touch of G28117: signal is true;
	signal G28118: std_logic; attribute dont_touch of G28118: signal is true;
	signal G28119: std_logic; attribute dont_touch of G28119: signal is true;
	signal G28120: std_logic; attribute dont_touch of G28120: signal is true;
	signal G28121: std_logic; attribute dont_touch of G28121: signal is true;
	signal G28124: std_logic; attribute dont_touch of G28124: signal is true;
	signal G28125: std_logic; attribute dont_touch of G28125: signal is true;
	signal G28126: std_logic; attribute dont_touch of G28126: signal is true;
	signal G28127: std_logic; attribute dont_touch of G28127: signal is true;
	signal G28130: std_logic; attribute dont_touch of G28130: signal is true;
	signal G28131: std_logic; attribute dont_touch of G28131: signal is true;
	signal G28132: std_logic; attribute dont_touch of G28132: signal is true;
	signal G28133: std_logic; attribute dont_touch of G28133: signal is true;
	signal G28134: std_logic; attribute dont_touch of G28134: signal is true;
	signal G28135: std_logic; attribute dont_touch of G28135: signal is true;
	signal G28136: std_logic; attribute dont_touch of G28136: signal is true;
	signal G28137: std_logic; attribute dont_touch of G28137: signal is true;
	signal G28138: std_logic; attribute dont_touch of G28138: signal is true;
	signal G28139: std_logic; attribute dont_touch of G28139: signal is true;
	signal G28140: std_logic; attribute dont_touch of G28140: signal is true;
	signal G28141: std_logic; attribute dont_touch of G28141: signal is true;
	signal G28142: std_logic; attribute dont_touch of G28142: signal is true;
	signal G28143: std_logic; attribute dont_touch of G28143: signal is true;
	signal G28144: std_logic; attribute dont_touch of G28144: signal is true;
	signal G28147: std_logic; attribute dont_touch of G28147: signal is true;
	signal G28148: std_logic; attribute dont_touch of G28148: signal is true;
	signal G28149: std_logic; attribute dont_touch of G28149: signal is true;
	signal G28150: std_logic; attribute dont_touch of G28150: signal is true;
	signal G28151: std_logic; attribute dont_touch of G28151: signal is true;
	signal G28152: std_logic; attribute dont_touch of G28152: signal is true;
	signal G28153: std_logic; attribute dont_touch of G28153: signal is true;
	signal G28154: std_logic; attribute dont_touch of G28154: signal is true;
	signal G28155: std_logic; attribute dont_touch of G28155: signal is true;
	signal G28156: std_logic; attribute dont_touch of G28156: signal is true;
	signal G28157: std_logic; attribute dont_touch of G28157: signal is true;
	signal G28158: std_logic; attribute dont_touch of G28158: signal is true;
	signal G28159: std_logic; attribute dont_touch of G28159: signal is true;
	signal G28160: std_logic; attribute dont_touch of G28160: signal is true;
	signal G28161: std_logic; attribute dont_touch of G28161: signal is true;
	signal G28162: std_logic; attribute dont_touch of G28162: signal is true;
	signal G28163: std_logic; attribute dont_touch of G28163: signal is true;
	signal G28164: std_logic; attribute dont_touch of G28164: signal is true;
	signal G28165: std_logic; attribute dont_touch of G28165: signal is true;
	signal G28166: std_logic; attribute dont_touch of G28166: signal is true;
	signal G28167: std_logic; attribute dont_touch of G28167: signal is true;
	signal G28171: std_logic; attribute dont_touch of G28171: signal is true;
	signal G28172: std_logic; attribute dont_touch of G28172: signal is true;
	signal G28173: std_logic; attribute dont_touch of G28173: signal is true;
	signal G28174: std_logic; attribute dont_touch of G28174: signal is true;
	signal G28178: std_logic; attribute dont_touch of G28178: signal is true;
	signal G28179: std_logic; attribute dont_touch of G28179: signal is true;
	signal G28180: std_logic; attribute dont_touch of G28180: signal is true;
	signal G28181: std_logic; attribute dont_touch of G28181: signal is true;
	signal G28182: std_logic; attribute dont_touch of G28182: signal is true;
	signal G28183: std_logic; attribute dont_touch of G28183: signal is true;
	signal G28184: std_logic; attribute dont_touch of G28184: signal is true;
	signal G28185: std_logic; attribute dont_touch of G28185: signal is true;
	signal G28186: std_logic; attribute dont_touch of G28186: signal is true;
	signal G28187: std_logic; attribute dont_touch of G28187: signal is true;
	signal G28188: std_logic; attribute dont_touch of G28188: signal is true;
	signal G28191: std_logic; attribute dont_touch of G28191: signal is true;
	signal G28192: std_logic; attribute dont_touch of G28192: signal is true;
	signal G28193: std_logic; attribute dont_touch of G28193: signal is true;
	signal G28194: std_logic; attribute dont_touch of G28194: signal is true;
	signal G28197: std_logic; attribute dont_touch of G28197: signal is true;
	signal G28198: std_logic; attribute dont_touch of G28198: signal is true;
	signal G28199: std_logic; attribute dont_touch of G28199: signal is true;
	signal G28200: std_logic; attribute dont_touch of G28200: signal is true;
	signal G28201: std_logic; attribute dont_touch of G28201: signal is true;
	signal G28202: std_logic; attribute dont_touch of G28202: signal is true;
	signal G28203: std_logic; attribute dont_touch of G28203: signal is true;
	signal G28204: std_logic; attribute dont_touch of G28204: signal is true;
	signal G28205: std_logic; attribute dont_touch of G28205: signal is true;
	signal G28206: std_logic; attribute dont_touch of G28206: signal is true;
	signal G28207: std_logic; attribute dont_touch of G28207: signal is true;
	signal G28208: std_logic; attribute dont_touch of G28208: signal is true;
	signal G28209: std_logic; attribute dont_touch of G28209: signal is true;
	signal G28210: std_logic; attribute dont_touch of G28210: signal is true;
	signal G28211: std_logic; attribute dont_touch of G28211: signal is true;
	signal G28212: std_logic; attribute dont_touch of G28212: signal is true;
	signal G28213: std_logic; attribute dont_touch of G28213: signal is true;
	signal G28214: std_logic; attribute dont_touch of G28214: signal is true;
	signal G28215: std_logic; attribute dont_touch of G28215: signal is true;
	signal G28216: std_logic; attribute dont_touch of G28216: signal is true;
	signal G28217: std_logic; attribute dont_touch of G28217: signal is true;
	signal G28218: std_logic; attribute dont_touch of G28218: signal is true;
	signal G28219: std_logic; attribute dont_touch of G28219: signal is true;
	signal G28220: std_logic; attribute dont_touch of G28220: signal is true;
	signal G28223: std_logic; attribute dont_touch of G28223: signal is true;
	signal G28224: std_logic; attribute dont_touch of G28224: signal is true;
	signal G28225: std_logic; attribute dont_touch of G28225: signal is true;
	signal G28226: std_logic; attribute dont_touch of G28226: signal is true;
	signal G28227: std_logic; attribute dont_touch of G28227: signal is true;
	signal G28228: std_logic; attribute dont_touch of G28228: signal is true;
	signal G28229: std_logic; attribute dont_touch of G28229: signal is true;
	signal G28230: std_logic; attribute dont_touch of G28230: signal is true;
	signal G28231: std_logic; attribute dont_touch of G28231: signal is true;
	signal G28232: std_logic; attribute dont_touch of G28232: signal is true;
	signal G28233: std_logic; attribute dont_touch of G28233: signal is true;
	signal G28234: std_logic; attribute dont_touch of G28234: signal is true;
	signal G28235: std_logic; attribute dont_touch of G28235: signal is true;
	signal G28236: std_logic; attribute dont_touch of G28236: signal is true;
	signal G28237: std_logic; attribute dont_touch of G28237: signal is true;
	signal G28238: std_logic; attribute dont_touch of G28238: signal is true;
	signal G28239: std_logic; attribute dont_touch of G28239: signal is true;
	signal G28240: std_logic; attribute dont_touch of G28240: signal is true;
	signal G28241: std_logic; attribute dont_touch of G28241: signal is true;
	signal G28242: std_logic; attribute dont_touch of G28242: signal is true;
	signal G28243: std_logic; attribute dont_touch of G28243: signal is true;
	signal G28244: std_logic; attribute dont_touch of G28244: signal is true;
	signal G28245: std_logic; attribute dont_touch of G28245: signal is true;
	signal G28246: std_logic; attribute dont_touch of G28246: signal is true;
	signal G28247: std_logic; attribute dont_touch of G28247: signal is true;
	signal G28248: std_logic; attribute dont_touch of G28248: signal is true;
	signal G28249: std_logic; attribute dont_touch of G28249: signal is true;
	signal G28250: std_logic; attribute dont_touch of G28250: signal is true;
	signal G28251: std_logic; attribute dont_touch of G28251: signal is true;
	signal G28252: std_logic; attribute dont_touch of G28252: signal is true;
	signal G28253: std_logic; attribute dont_touch of G28253: signal is true;
	signal G28254: std_logic; attribute dont_touch of G28254: signal is true;
	signal G28255: std_logic; attribute dont_touch of G28255: signal is true;
	signal G28256: std_logic; attribute dont_touch of G28256: signal is true;
	signal G28257: std_logic; attribute dont_touch of G28257: signal is true;
	signal G28258: std_logic; attribute dont_touch of G28258: signal is true;
	signal G28259: std_logic; attribute dont_touch of G28259: signal is true;
	signal G28260: std_logic; attribute dont_touch of G28260: signal is true;
	signal G28261: std_logic; attribute dont_touch of G28261: signal is true;
	signal G28262: std_logic; attribute dont_touch of G28262: signal is true;
	signal G28263: std_logic; attribute dont_touch of G28263: signal is true;
	signal G28264: std_logic; attribute dont_touch of G28264: signal is true;
	signal G28265: std_logic; attribute dont_touch of G28265: signal is true;
	signal G28266: std_logic; attribute dont_touch of G28266: signal is true;
	signal G28267: std_logic; attribute dont_touch of G28267: signal is true;
	signal G28268: std_logic; attribute dont_touch of G28268: signal is true;
	signal G28269: std_logic; attribute dont_touch of G28269: signal is true;
	signal G28270: std_logic; attribute dont_touch of G28270: signal is true;
	signal G28271: std_logic; attribute dont_touch of G28271: signal is true;
	signal G28272: std_logic; attribute dont_touch of G28272: signal is true;
	signal G28273: std_logic; attribute dont_touch of G28273: signal is true;
	signal G28274: std_logic; attribute dont_touch of G28274: signal is true;
	signal G28279: std_logic; attribute dont_touch of G28279: signal is true;
	signal G28280: std_logic; attribute dont_touch of G28280: signal is true;
	signal G28281: std_logic; attribute dont_touch of G28281: signal is true;
	signal G28282: std_logic; attribute dont_touch of G28282: signal is true;
	signal G28283: std_logic; attribute dont_touch of G28283: signal is true;
	signal G28284: std_logic; attribute dont_touch of G28284: signal is true;
	signal G28285: std_logic; attribute dont_touch of G28285: signal is true;
	signal G28286: std_logic; attribute dont_touch of G28286: signal is true;
	signal G28287: std_logic; attribute dont_touch of G28287: signal is true;
	signal G28288: std_logic; attribute dont_touch of G28288: signal is true;
	signal G28289: std_logic; attribute dont_touch of G28289: signal is true;
	signal G28290: std_logic; attribute dont_touch of G28290: signal is true;
	signal G28291: std_logic; attribute dont_touch of G28291: signal is true;
	signal G28292: std_logic; attribute dont_touch of G28292: signal is true;
	signal G28293: std_logic; attribute dont_touch of G28293: signal is true;
	signal G28294: std_logic; attribute dont_touch of G28294: signal is true;
	signal G28295: std_logic; attribute dont_touch of G28295: signal is true;
	signal G28296: std_logic; attribute dont_touch of G28296: signal is true;
	signal G28297: std_logic; attribute dont_touch of G28297: signal is true;
	signal G28298: std_logic; attribute dont_touch of G28298: signal is true;
	signal G28299: std_logic; attribute dont_touch of G28299: signal is true;
	signal G28300: std_logic; attribute dont_touch of G28300: signal is true;
	signal G28301: std_logic; attribute dont_touch of G28301: signal is true;
	signal G28302: std_logic; attribute dont_touch of G28302: signal is true;
	signal G28303: std_logic; attribute dont_touch of G28303: signal is true;
	signal G28304: std_logic; attribute dont_touch of G28304: signal is true;
	signal G28305: std_logic; attribute dont_touch of G28305: signal is true;
	signal G28306: std_logic; attribute dont_touch of G28306: signal is true;
	signal G28307: std_logic; attribute dont_touch of G28307: signal is true;
	signal G28308: std_logic; attribute dont_touch of G28308: signal is true;
	signal G28309: std_logic; attribute dont_touch of G28309: signal is true;
	signal G28310: std_logic; attribute dont_touch of G28310: signal is true;
	signal G28311: std_logic; attribute dont_touch of G28311: signal is true;
	signal G28312: std_logic; attribute dont_touch of G28312: signal is true;
	signal G28313: std_logic; attribute dont_touch of G28313: signal is true;
	signal G28314: std_logic; attribute dont_touch of G28314: signal is true;
	signal G28315: std_logic; attribute dont_touch of G28315: signal is true;
	signal G28316: std_logic; attribute dont_touch of G28316: signal is true;
	signal G28317: std_logic; attribute dont_touch of G28317: signal is true;
	signal G28318: std_logic; attribute dont_touch of G28318: signal is true;
	signal G28319: std_logic; attribute dont_touch of G28319: signal is true;
	signal G28320: std_logic; attribute dont_touch of G28320: signal is true;
	signal G28321: std_logic; attribute dont_touch of G28321: signal is true;
	signal G28322: std_logic; attribute dont_touch of G28322: signal is true;
	signal G28323: std_logic; attribute dont_touch of G28323: signal is true;
	signal G28324: std_logic; attribute dont_touch of G28324: signal is true;
	signal G28325: std_logic; attribute dont_touch of G28325: signal is true;
	signal G28326: std_logic; attribute dont_touch of G28326: signal is true;
	signal G28327: std_logic; attribute dont_touch of G28327: signal is true;
	signal G28328: std_logic; attribute dont_touch of G28328: signal is true;
	signal G28329: std_logic; attribute dont_touch of G28329: signal is true;
	signal G28330: std_logic; attribute dont_touch of G28330: signal is true;
	signal G28331: std_logic; attribute dont_touch of G28331: signal is true;
	signal G28332: std_logic; attribute dont_touch of G28332: signal is true;
	signal G28333: std_logic; attribute dont_touch of G28333: signal is true;
	signal G28334: std_logic; attribute dont_touch of G28334: signal is true;
	signal G28335: std_logic; attribute dont_touch of G28335: signal is true;
	signal G28336: std_logic; attribute dont_touch of G28336: signal is true;
	signal G28339: std_logic; attribute dont_touch of G28339: signal is true;
	signal G28340: std_logic; attribute dont_touch of G28340: signal is true;
	signal G28341: std_logic; attribute dont_touch of G28341: signal is true;
	signal G28342: std_logic; attribute dont_touch of G28342: signal is true;
	signal G28343: std_logic; attribute dont_touch of G28343: signal is true;
	signal G28344: std_logic; attribute dont_touch of G28344: signal is true;
	signal G28345: std_logic; attribute dont_touch of G28345: signal is true;
	signal G28346: std_logic; attribute dont_touch of G28346: signal is true;
	signal G28347: std_logic; attribute dont_touch of G28347: signal is true;
	signal G28348: std_logic; attribute dont_touch of G28348: signal is true;
	signal G28349: std_logic; attribute dont_touch of G28349: signal is true;
	signal G28352: std_logic; attribute dont_touch of G28352: signal is true;
	signal G28353: std_logic; attribute dont_touch of G28353: signal is true;
	signal G28357: std_logic; attribute dont_touch of G28357: signal is true;
	signal G28358: std_logic; attribute dont_touch of G28358: signal is true;
	signal G28359: std_logic; attribute dont_touch of G28359: signal is true;
	signal G28360: std_logic; attribute dont_touch of G28360: signal is true;
	signal G28361: std_logic; attribute dont_touch of G28361: signal is true;
	signal G28362: std_logic; attribute dont_touch of G28362: signal is true;
	signal G28363: std_logic; attribute dont_touch of G28363: signal is true;
	signal G28367: std_logic; attribute dont_touch of G28367: signal is true;
	signal G28368: std_logic; attribute dont_touch of G28368: signal is true;
	signal G28369: std_logic; attribute dont_touch of G28369: signal is true;
	signal G28370: std_logic; attribute dont_touch of G28370: signal is true;
	signal G28371: std_logic; attribute dont_touch of G28371: signal is true;
	signal G28372: std_logic; attribute dont_touch of G28372: signal is true;
	signal G28373: std_logic; attribute dont_touch of G28373: signal is true;
	signal G28374: std_logic; attribute dont_touch of G28374: signal is true;
	signal G28375: std_logic; attribute dont_touch of G28375: signal is true;
	signal G28376: std_logic; attribute dont_touch of G28376: signal is true;
	signal G28380: std_logic; attribute dont_touch of G28380: signal is true;
	signal G28381: std_logic; attribute dont_touch of G28381: signal is true;
	signal G28385: std_logic; attribute dont_touch of G28385: signal is true;
	signal G28386: std_logic; attribute dont_touch of G28386: signal is true;
	signal G28387: std_logic; attribute dont_touch of G28387: signal is true;
	signal G28388: std_logic; attribute dont_touch of G28388: signal is true;
	signal G28389: std_logic; attribute dont_touch of G28389: signal is true;
	signal G28390: std_logic; attribute dont_touch of G28390: signal is true;
	signal G28391: std_logic; attribute dont_touch of G28391: signal is true;
	signal G28395: std_logic; attribute dont_touch of G28395: signal is true;
	signal G28399: std_logic; attribute dont_touch of G28399: signal is true;
	signal G28400: std_logic; attribute dont_touch of G28400: signal is true;
	signal G28401: std_logic; attribute dont_touch of G28401: signal is true;
	signal G28402: std_logic; attribute dont_touch of G28402: signal is true;
	signal G28403: std_logic; attribute dont_touch of G28403: signal is true;
	signal G28404: std_logic; attribute dont_touch of G28404: signal is true;
	signal G28405: std_logic; attribute dont_touch of G28405: signal is true;
	signal G28406: std_logic; attribute dont_touch of G28406: signal is true;
	signal G28410: std_logic; attribute dont_touch of G28410: signal is true;
	signal G28414: std_logic; attribute dont_touch of G28414: signal is true;
	signal G28415: std_logic; attribute dont_touch of G28415: signal is true;
	signal G28416: std_logic; attribute dont_touch of G28416: signal is true;
	signal G28417: std_logic; attribute dont_touch of G28417: signal is true;
	signal G28418: std_logic; attribute dont_touch of G28418: signal is true;
	signal G28419: std_logic; attribute dont_touch of G28419: signal is true;
	signal G28420: std_logic; attribute dont_touch of G28420: signal is true;
	signal G28421: std_logic; attribute dont_touch of G28421: signal is true;
	signal G28425: std_logic; attribute dont_touch of G28425: signal is true;
	signal G28426: std_logic; attribute dont_touch of G28426: signal is true;
	signal G28427: std_logic; attribute dont_touch of G28427: signal is true;
	signal G28428: std_logic; attribute dont_touch of G28428: signal is true;
	signal G28429: std_logic; attribute dont_touch of G28429: signal is true;
	signal G28430: std_logic; attribute dont_touch of G28430: signal is true;
	signal G28431: std_logic; attribute dont_touch of G28431: signal is true;
	signal G28435: std_logic; attribute dont_touch of G28435: signal is true;
	signal G28436: std_logic; attribute dont_touch of G28436: signal is true;
	signal G28439: std_logic; attribute dont_touch of G28439: signal is true;
	signal G28440: std_logic; attribute dont_touch of G28440: signal is true;
	signal G28441: std_logic; attribute dont_touch of G28441: signal is true;
	signal G28442: std_logic; attribute dont_touch of G28442: signal is true;
	signal G28443: std_logic; attribute dont_touch of G28443: signal is true;
	signal G28444: std_logic; attribute dont_touch of G28444: signal is true;
	signal G28448: std_logic; attribute dont_touch of G28448: signal is true;
	signal G28451: std_logic; attribute dont_touch of G28451: signal is true;
	signal G28452: std_logic; attribute dont_touch of G28452: signal is true;
	signal G28453: std_logic; attribute dont_touch of G28453: signal is true;
	signal G28454: std_logic; attribute dont_touch of G28454: signal is true;
	signal G28455: std_logic; attribute dont_touch of G28455: signal is true;
	signal G28456: std_logic; attribute dont_touch of G28456: signal is true;
	signal G28457: std_logic; attribute dont_touch of G28457: signal is true;
	signal G28458: std_logic; attribute dont_touch of G28458: signal is true;
	signal G28462: std_logic; attribute dont_touch of G28462: signal is true;
	signal G28463: std_logic; attribute dont_touch of G28463: signal is true;
	signal G28466: std_logic; attribute dont_touch of G28466: signal is true;
	signal G28467: std_logic; attribute dont_touch of G28467: signal is true;
	signal G28468: std_logic; attribute dont_touch of G28468: signal is true;
	signal G28469: std_logic; attribute dont_touch of G28469: signal is true;
	signal G28470: std_logic; attribute dont_touch of G28470: signal is true;
	signal G28471: std_logic; attribute dont_touch of G28471: signal is true;
	signal G28475: std_logic; attribute dont_touch of G28475: signal is true;
	signal G28476: std_logic; attribute dont_touch of G28476: signal is true;
	signal G28477: std_logic; attribute dont_touch of G28477: signal is true;
	signal G28478: std_logic; attribute dont_touch of G28478: signal is true;
	signal G28479: std_logic; attribute dont_touch of G28479: signal is true;
	signal G28480: std_logic; attribute dont_touch of G28480: signal is true;
	signal G28481: std_logic; attribute dont_touch of G28481: signal is true;
	signal G28482: std_logic; attribute dont_touch of G28482: signal is true;
	signal G28483: std_logic; attribute dont_touch of G28483: signal is true;
	signal G28484: std_logic; attribute dont_touch of G28484: signal is true;
	signal G28488: std_logic; attribute dont_touch of G28488: signal is true;
	signal G28489: std_logic; attribute dont_touch of G28489: signal is true;
	signal G28490: std_logic; attribute dont_touch of G28490: signal is true;
	signal G28491: std_logic; attribute dont_touch of G28491: signal is true;
	signal G28492: std_logic; attribute dont_touch of G28492: signal is true;
	signal G28493: std_logic; attribute dont_touch of G28493: signal is true;
	signal G28494: std_logic; attribute dont_touch of G28494: signal is true;
	signal G28495: std_logic; attribute dont_touch of G28495: signal is true;
	signal G28496: std_logic; attribute dont_touch of G28496: signal is true;
	signal G28497: std_logic; attribute dont_touch of G28497: signal is true;
	signal G28498: std_logic; attribute dont_touch of G28498: signal is true;
	signal G28499: std_logic; attribute dont_touch of G28499: signal is true;
	signal G28500: std_logic; attribute dont_touch of G28500: signal is true;
	signal G28504: std_logic; attribute dont_touch of G28504: signal is true;
	signal G28508: std_logic; attribute dont_touch of G28508: signal is true;
	signal G28509: std_logic; attribute dont_touch of G28509: signal is true;
	signal G28510: std_logic; attribute dont_touch of G28510: signal is true;
	signal G28511: std_logic; attribute dont_touch of G28511: signal is true;
	signal G28512: std_logic; attribute dont_touch of G28512: signal is true;
	signal G28513: std_logic; attribute dont_touch of G28513: signal is true;
	signal G28514: std_logic; attribute dont_touch of G28514: signal is true;
	signal G28515: std_logic; attribute dont_touch of G28515: signal is true;
	signal G28516: std_logic; attribute dont_touch of G28516: signal is true;
	signal G28517: std_logic; attribute dont_touch of G28517: signal is true;
	signal G28518: std_logic; attribute dont_touch of G28518: signal is true;
	signal G28519: std_logic; attribute dont_touch of G28519: signal is true;
	signal G28520: std_logic; attribute dont_touch of G28520: signal is true;
	signal G28521: std_logic; attribute dont_touch of G28521: signal is true;
	signal G28522: std_logic; attribute dont_touch of G28522: signal is true;
	signal G28523: std_logic; attribute dont_touch of G28523: signal is true;
	signal G28524: std_logic; attribute dont_touch of G28524: signal is true;
	signal G28525: std_logic; attribute dont_touch of G28525: signal is true;
	signal G28526: std_logic; attribute dont_touch of G28526: signal is true;
	signal G28527: std_logic; attribute dont_touch of G28527: signal is true;
	signal G28528: std_logic; attribute dont_touch of G28528: signal is true;
	signal G28529: std_logic; attribute dont_touch of G28529: signal is true;
	signal G28530: std_logic; attribute dont_touch of G28530: signal is true;
	signal G28531: std_logic; attribute dont_touch of G28531: signal is true;
	signal G28532: std_logic; attribute dont_touch of G28532: signal is true;
	signal G28533: std_logic; attribute dont_touch of G28533: signal is true;
	signal G28534: std_logic; attribute dont_touch of G28534: signal is true;
	signal G28535: std_logic; attribute dont_touch of G28535: signal is true;
	signal G28536: std_logic; attribute dont_touch of G28536: signal is true;
	signal G28537: std_logic; attribute dont_touch of G28537: signal is true;
	signal G28538: std_logic; attribute dont_touch of G28538: signal is true;
	signal G28539: std_logic; attribute dont_touch of G28539: signal is true;
	signal G28540: std_logic; attribute dont_touch of G28540: signal is true;
	signal G28541: std_logic; attribute dont_touch of G28541: signal is true;
	signal G28542: std_logic; attribute dont_touch of G28542: signal is true;
	signal G28543: std_logic; attribute dont_touch of G28543: signal is true;
	signal G28544: std_logic; attribute dont_touch of G28544: signal is true;
	signal G28545: std_logic; attribute dont_touch of G28545: signal is true;
	signal G28546: std_logic; attribute dont_touch of G28546: signal is true;
	signal G28547: std_logic; attribute dont_touch of G28547: signal is true;
	signal G28548: std_logic; attribute dont_touch of G28548: signal is true;
	signal G28549: std_logic; attribute dont_touch of G28549: signal is true;
	signal G28550: std_logic; attribute dont_touch of G28550: signal is true;
	signal G28551: std_logic; attribute dont_touch of G28551: signal is true;
	signal G28552: std_logic; attribute dont_touch of G28552: signal is true;
	signal G28553: std_logic; attribute dont_touch of G28553: signal is true;
	signal G28554: std_logic; attribute dont_touch of G28554: signal is true;
	signal G28555: std_logic; attribute dont_touch of G28555: signal is true;
	signal G28556: std_logic; attribute dont_touch of G28556: signal is true;
	signal G28557: std_logic; attribute dont_touch of G28557: signal is true;
	signal G28558: std_logic; attribute dont_touch of G28558: signal is true;
	signal G28559: std_logic; attribute dont_touch of G28559: signal is true;
	signal G28560: std_logic; attribute dont_touch of G28560: signal is true;
	signal G28561: std_logic; attribute dont_touch of G28561: signal is true;
	signal G28562: std_logic; attribute dont_touch of G28562: signal is true;
	signal G28563: std_logic; attribute dont_touch of G28563: signal is true;
	signal G28564: std_logic; attribute dont_touch of G28564: signal is true;
	signal G28565: std_logic; attribute dont_touch of G28565: signal is true;
	signal G28566: std_logic; attribute dont_touch of G28566: signal is true;
	signal G28567: std_logic; attribute dont_touch of G28567: signal is true;
	signal G28568: std_logic; attribute dont_touch of G28568: signal is true;
	signal G28569: std_logic; attribute dont_touch of G28569: signal is true;
	signal G28570: std_logic; attribute dont_touch of G28570: signal is true;
	signal G28571: std_logic; attribute dont_touch of G28571: signal is true;
	signal G28572: std_logic; attribute dont_touch of G28572: signal is true;
	signal G28573: std_logic; attribute dont_touch of G28573: signal is true;
	signal G28574: std_logic; attribute dont_touch of G28574: signal is true;
	signal G28575: std_logic; attribute dont_touch of G28575: signal is true;
	signal G28576: std_logic; attribute dont_touch of G28576: signal is true;
	signal G28577: std_logic; attribute dont_touch of G28577: signal is true;
	signal G28578: std_logic; attribute dont_touch of G28578: signal is true;
	signal G28579: std_logic; attribute dont_touch of G28579: signal is true;
	signal G28580: std_logic; attribute dont_touch of G28580: signal is true;
	signal G28581: std_logic; attribute dont_touch of G28581: signal is true;
	signal G28582: std_logic; attribute dont_touch of G28582: signal is true;
	signal G28583: std_logic; attribute dont_touch of G28583: signal is true;
	signal G28584: std_logic; attribute dont_touch of G28584: signal is true;
	signal G28585: std_logic; attribute dont_touch of G28585: signal is true;
	signal G28586: std_logic; attribute dont_touch of G28586: signal is true;
	signal G28587: std_logic; attribute dont_touch of G28587: signal is true;
	signal G28588: std_logic; attribute dont_touch of G28588: signal is true;
	signal G28589: std_logic; attribute dont_touch of G28589: signal is true;
	signal G28590: std_logic; attribute dont_touch of G28590: signal is true;
	signal G28591: std_logic; attribute dont_touch of G28591: signal is true;
	signal G28592: std_logic; attribute dont_touch of G28592: signal is true;
	signal G28593: std_logic; attribute dont_touch of G28593: signal is true;
	signal G28594: std_logic; attribute dont_touch of G28594: signal is true;
	signal G28595: std_logic; attribute dont_touch of G28595: signal is true;
	signal G28596: std_logic; attribute dont_touch of G28596: signal is true;
	signal G28597: std_logic; attribute dont_touch of G28597: signal is true;
	signal G28598: std_logic; attribute dont_touch of G28598: signal is true;
	signal G28599: std_logic; attribute dont_touch of G28599: signal is true;
	signal G28600: std_logic; attribute dont_touch of G28600: signal is true;
	signal G28601: std_logic; attribute dont_touch of G28601: signal is true;
	signal G28602: std_logic; attribute dont_touch of G28602: signal is true;
	signal G28603: std_logic; attribute dont_touch of G28603: signal is true;
	signal G28604: std_logic; attribute dont_touch of G28604: signal is true;
	signal G28605: std_logic; attribute dont_touch of G28605: signal is true;
	signal G28606: std_logic; attribute dont_touch of G28606: signal is true;
	signal G28607: std_logic; attribute dont_touch of G28607: signal is true;
	signal G28608: std_logic; attribute dont_touch of G28608: signal is true;
	signal G28609: std_logic; attribute dont_touch of G28609: signal is true;
	signal G28610: std_logic; attribute dont_touch of G28610: signal is true;
	signal G28611: std_logic; attribute dont_touch of G28611: signal is true;
	signal G28612: std_logic; attribute dont_touch of G28612: signal is true;
	signal G28613: std_logic; attribute dont_touch of G28613: signal is true;
	signal G28614: std_logic; attribute dont_touch of G28614: signal is true;
	signal G28615: std_logic; attribute dont_touch of G28615: signal is true;
	signal G28616: std_logic; attribute dont_touch of G28616: signal is true;
	signal G28617: std_logic; attribute dont_touch of G28617: signal is true;
	signal G28618: std_logic; attribute dont_touch of G28618: signal is true;
	signal G28619: std_logic; attribute dont_touch of G28619: signal is true;
	signal G28620: std_logic; attribute dont_touch of G28620: signal is true;
	signal G28621: std_logic; attribute dont_touch of G28621: signal is true;
	signal G28622: std_logic; attribute dont_touch of G28622: signal is true;
	signal G28623: std_logic; attribute dont_touch of G28623: signal is true;
	signal G28624: std_logic; attribute dont_touch of G28624: signal is true;
	signal G28625: std_logic; attribute dont_touch of G28625: signal is true;
	signal G28626: std_logic; attribute dont_touch of G28626: signal is true;
	signal G28627: std_logic; attribute dont_touch of G28627: signal is true;
	signal G28628: std_logic; attribute dont_touch of G28628: signal is true;
	signal G28629: std_logic; attribute dont_touch of G28629: signal is true;
	signal G28630: std_logic; attribute dont_touch of G28630: signal is true;
	signal G28631: std_logic; attribute dont_touch of G28631: signal is true;
	signal G28632: std_logic; attribute dont_touch of G28632: signal is true;
	signal G28633: std_logic; attribute dont_touch of G28633: signal is true;
	signal G28634: std_logic; attribute dont_touch of G28634: signal is true;
	signal G28635: std_logic; attribute dont_touch of G28635: signal is true;
	signal G28636: std_logic; attribute dont_touch of G28636: signal is true;
	signal G28637: std_logic; attribute dont_touch of G28637: signal is true;
	signal G28638: std_logic; attribute dont_touch of G28638: signal is true;
	signal G28639: std_logic; attribute dont_touch of G28639: signal is true;
	signal G28640: std_logic; attribute dont_touch of G28640: signal is true;
	signal G28641: std_logic; attribute dont_touch of G28641: signal is true;
	signal G28642: std_logic; attribute dont_touch of G28642: signal is true;
	signal G28643: std_logic; attribute dont_touch of G28643: signal is true;
	signal G28644: std_logic; attribute dont_touch of G28644: signal is true;
	signal G28645: std_logic; attribute dont_touch of G28645: signal is true;
	signal G28646: std_logic; attribute dont_touch of G28646: signal is true;
	signal G28647: std_logic; attribute dont_touch of G28647: signal is true;
	signal G28648: std_logic; attribute dont_touch of G28648: signal is true;
	signal G28649: std_logic; attribute dont_touch of G28649: signal is true;
	signal G28650: std_logic; attribute dont_touch of G28650: signal is true;
	signal G28651: std_logic; attribute dont_touch of G28651: signal is true;
	signal G28652: std_logic; attribute dont_touch of G28652: signal is true;
	signal G28653: std_logic; attribute dont_touch of G28653: signal is true;
	signal G28654: std_logic; attribute dont_touch of G28654: signal is true;
	signal G28655: std_logic; attribute dont_touch of G28655: signal is true;
	signal G28656: std_logic; attribute dont_touch of G28656: signal is true;
	signal G28657: std_logic; attribute dont_touch of G28657: signal is true;
	signal G28658: std_logic; attribute dont_touch of G28658: signal is true;
	signal G28659: std_logic; attribute dont_touch of G28659: signal is true;
	signal G28660: std_logic; attribute dont_touch of G28660: signal is true;
	signal G28661: std_logic; attribute dont_touch of G28661: signal is true;
	signal G28662: std_logic; attribute dont_touch of G28662: signal is true;
	signal G28663: std_logic; attribute dont_touch of G28663: signal is true;
	signal G28664: std_logic; attribute dont_touch of G28664: signal is true;
	signal G28665: std_logic; attribute dont_touch of G28665: signal is true;
	signal G28666: std_logic; attribute dont_touch of G28666: signal is true;
	signal G28667: std_logic; attribute dont_touch of G28667: signal is true;
	signal G28668: std_logic; attribute dont_touch of G28668: signal is true;
	signal G28669: std_logic; attribute dont_touch of G28669: signal is true;
	signal G28670: std_logic; attribute dont_touch of G28670: signal is true;
	signal G28671: std_logic; attribute dont_touch of G28671: signal is true;
	signal G28672: std_logic; attribute dont_touch of G28672: signal is true;
	signal G28673: std_logic; attribute dont_touch of G28673: signal is true;
	signal G28674: std_logic; attribute dont_touch of G28674: signal is true;
	signal G28675: std_logic; attribute dont_touch of G28675: signal is true;
	signal G28676: std_logic; attribute dont_touch of G28676: signal is true;
	signal G28677: std_logic; attribute dont_touch of G28677: signal is true;
	signal G28678: std_logic; attribute dont_touch of G28678: signal is true;
	signal G28679: std_logic; attribute dont_touch of G28679: signal is true;
	signal G28680: std_logic; attribute dont_touch of G28680: signal is true;
	signal G28681: std_logic; attribute dont_touch of G28681: signal is true;
	signal G28682: std_logic; attribute dont_touch of G28682: signal is true;
	signal G28683: std_logic; attribute dont_touch of G28683: signal is true;
	signal G28684: std_logic; attribute dont_touch of G28684: signal is true;
	signal G28685: std_logic; attribute dont_touch of G28685: signal is true;
	signal G28686: std_logic; attribute dont_touch of G28686: signal is true;
	signal G28687: std_logic; attribute dont_touch of G28687: signal is true;
	signal G28688: std_logic; attribute dont_touch of G28688: signal is true;
	signal G28689: std_logic; attribute dont_touch of G28689: signal is true;
	signal G28690: std_logic; attribute dont_touch of G28690: signal is true;
	signal G28691: std_logic; attribute dont_touch of G28691: signal is true;
	signal G28692: std_logic; attribute dont_touch of G28692: signal is true;
	signal G28693: std_logic; attribute dont_touch of G28693: signal is true;
	signal G28694: std_logic; attribute dont_touch of G28694: signal is true;
	signal G28695: std_logic; attribute dont_touch of G28695: signal is true;
	signal G28696: std_logic; attribute dont_touch of G28696: signal is true;
	signal G28697: std_logic; attribute dont_touch of G28697: signal is true;
	signal G28698: std_logic; attribute dont_touch of G28698: signal is true;
	signal G28699: std_logic; attribute dont_touch of G28699: signal is true;
	signal G28700: std_logic; attribute dont_touch of G28700: signal is true;
	signal G28701: std_logic; attribute dont_touch of G28701: signal is true;
	signal G28702: std_logic; attribute dont_touch of G28702: signal is true;
	signal G28703: std_logic; attribute dont_touch of G28703: signal is true;
	signal G28704: std_logic; attribute dont_touch of G28704: signal is true;
	signal G28705: std_logic; attribute dont_touch of G28705: signal is true;
	signal G28706: std_logic; attribute dont_touch of G28706: signal is true;
	signal G28707: std_logic; attribute dont_touch of G28707: signal is true;
	signal G28708: std_logic; attribute dont_touch of G28708: signal is true;
	signal G28709: std_logic; attribute dont_touch of G28709: signal is true;
	signal G28710: std_logic; attribute dont_touch of G28710: signal is true;
	signal G28711: std_logic; attribute dont_touch of G28711: signal is true;
	signal G28712: std_logic; attribute dont_touch of G28712: signal is true;
	signal G28713: std_logic; attribute dont_touch of G28713: signal is true;
	signal G28714: std_logic; attribute dont_touch of G28714: signal is true;
	signal G28715: std_logic; attribute dont_touch of G28715: signal is true;
	signal G28716: std_logic; attribute dont_touch of G28716: signal is true;
	signal G28717: std_logic; attribute dont_touch of G28717: signal is true;
	signal G28718: std_logic; attribute dont_touch of G28718: signal is true;
	signal G28719: std_logic; attribute dont_touch of G28719: signal is true;
	signal G28720: std_logic; attribute dont_touch of G28720: signal is true;
	signal G28721: std_logic; attribute dont_touch of G28721: signal is true;
	signal G28722: std_logic; attribute dont_touch of G28722: signal is true;
	signal G28723: std_logic; attribute dont_touch of G28723: signal is true;
	signal G28724: std_logic; attribute dont_touch of G28724: signal is true;
	signal G28725: std_logic; attribute dont_touch of G28725: signal is true;
	signal G28726: std_logic; attribute dont_touch of G28726: signal is true;
	signal G28727: std_logic; attribute dont_touch of G28727: signal is true;
	signal G28728: std_logic; attribute dont_touch of G28728: signal is true;
	signal G28729: std_logic; attribute dont_touch of G28729: signal is true;
	signal G28730: std_logic; attribute dont_touch of G28730: signal is true;
	signal G28731: std_logic; attribute dont_touch of G28731: signal is true;
	signal G28732: std_logic; attribute dont_touch of G28732: signal is true;
	signal G28733: std_logic; attribute dont_touch of G28733: signal is true;
	signal G28734: std_logic; attribute dont_touch of G28734: signal is true;
	signal G28735: std_logic; attribute dont_touch of G28735: signal is true;
	signal G28736: std_logic; attribute dont_touch of G28736: signal is true;
	signal G28739: std_logic; attribute dont_touch of G28739: signal is true;
	signal G28743: std_logic; attribute dont_touch of G28743: signal is true;
	signal G28744: std_logic; attribute dont_touch of G28744: signal is true;
	signal G28745: std_logic; attribute dont_touch of G28745: signal is true;
	signal G28746: std_logic; attribute dont_touch of G28746: signal is true;
	signal G28747: std_logic; attribute dont_touch of G28747: signal is true;
	signal G28748: std_logic; attribute dont_touch of G28748: signal is true;
	signal G28749: std_logic; attribute dont_touch of G28749: signal is true;
	signal G28750: std_logic; attribute dont_touch of G28750: signal is true;
	signal G28751: std_logic; attribute dont_touch of G28751: signal is true;
	signal G28752: std_logic; attribute dont_touch of G28752: signal is true;
	signal G28754: std_logic; attribute dont_touch of G28754: signal is true;
	signal G28755: std_logic; attribute dont_touch of G28755: signal is true;
	signal G28758: std_logic; attribute dont_touch of G28758: signal is true;
	signal G28761: std_logic; attribute dont_touch of G28761: signal is true;
	signal G28765: std_logic; attribute dont_touch of G28765: signal is true;
	signal G28768: std_logic; attribute dont_touch of G28768: signal is true;
	signal G28772: std_logic; attribute dont_touch of G28772: signal is true;
	signal G28773: std_logic; attribute dont_touch of G28773: signal is true;
	signal G28774: std_logic; attribute dont_touch of G28774: signal is true;
	signal G28775: std_logic; attribute dont_touch of G28775: signal is true;
	signal G28776: std_logic; attribute dont_touch of G28776: signal is true;
	signal G28777: std_logic; attribute dont_touch of G28777: signal is true;
	signal G28778: std_logic; attribute dont_touch of G28778: signal is true;
	signal G28779: std_logic; attribute dont_touch of G28779: signal is true;
	signal G28780: std_logic; attribute dont_touch of G28780: signal is true;
	signal G28783: std_logic; attribute dont_touch of G28783: signal is true;
	signal G28786: std_logic; attribute dont_touch of G28786: signal is true;
	signal G28789: std_logic; attribute dont_touch of G28789: signal is true;
	signal G28793: std_logic; attribute dont_touch of G28793: signal is true;
	signal G28796: std_logic; attribute dont_touch of G28796: signal is true;
	signal G28799: std_logic; attribute dont_touch of G28799: signal is true;
	signal G28803: std_logic; attribute dont_touch of G28803: signal is true;
	signal G28812: std_logic; attribute dont_touch of G28812: signal is true;
	signal G28813: std_logic; attribute dont_touch of G28813: signal is true;
	signal G28814: std_logic; attribute dont_touch of G28814: signal is true;
	signal G28815: std_logic; attribute dont_touch of G28815: signal is true;
	signal G28816: std_logic; attribute dont_touch of G28816: signal is true;
	signal G28817: std_logic; attribute dont_touch of G28817: signal is true;
	signal G28818: std_logic; attribute dont_touch of G28818: signal is true;
	signal G28819: std_logic; attribute dont_touch of G28819: signal is true;
	signal G28820: std_logic; attribute dont_touch of G28820: signal is true;
	signal G28823: std_logic; attribute dont_touch of G28823: signal is true;
	signal G28824: std_logic; attribute dont_touch of G28824: signal is true;
	signal G28827: std_logic; attribute dont_touch of G28827: signal is true;
	signal G28830: std_logic; attribute dont_touch of G28830: signal is true;
	signal G28833: std_logic; attribute dont_touch of G28833: signal is true;
	signal G28837: std_logic; attribute dont_touch of G28837: signal is true;
	signal G28840: std_logic; attribute dont_touch of G28840: signal is true;
	signal G28843: std_logic; attribute dont_touch of G28843: signal is true;
	signal G28846: std_logic; attribute dont_touch of G28846: signal is true;
	signal G28850: std_logic; attribute dont_touch of G28850: signal is true;
	signal G28851: std_logic; attribute dont_touch of G28851: signal is true;
	signal G28852: std_logic; attribute dont_touch of G28852: signal is true;
	signal G28853: std_logic; attribute dont_touch of G28853: signal is true;
	signal G28856: std_logic; attribute dont_touch of G28856: signal is true;
	signal G28857: std_logic; attribute dont_touch of G28857: signal is true;
	signal G28860: std_logic; attribute dont_touch of G28860: signal is true;
	signal G28861: std_logic; attribute dont_touch of G28861: signal is true;
	signal G28864: std_logic; attribute dont_touch of G28864: signal is true;
	signal G28867: std_logic; attribute dont_touch of G28867: signal is true;
	signal G28870: std_logic; attribute dont_touch of G28870: signal is true;
	signal G28871: std_logic; attribute dont_touch of G28871: signal is true;
	signal G28874: std_logic; attribute dont_touch of G28874: signal is true;
	signal G28877: std_logic; attribute dont_touch of G28877: signal is true;
	signal G28880: std_logic; attribute dont_touch of G28880: signal is true;
	signal G28884: std_logic; attribute dont_touch of G28884: signal is true;
	signal G28885: std_logic; attribute dont_touch of G28885: signal is true;
	signal G28888: std_logic; attribute dont_touch of G28888: signal is true;
	signal G28889: std_logic; attribute dont_touch of G28889: signal is true;
	signal G28892: std_logic; attribute dont_touch of G28892: signal is true;
	signal G28895: std_logic; attribute dont_touch of G28895: signal is true;
	signal G28896: std_logic; attribute dont_touch of G28896: signal is true;
	signal G28899: std_logic; attribute dont_touch of G28899: signal is true;
	signal G28900: std_logic; attribute dont_touch of G28900: signal is true;
	signal G28903: std_logic; attribute dont_touch of G28903: signal is true;
	signal G28906: std_logic; attribute dont_touch of G28906: signal is true;
	signal G28907: std_logic; attribute dont_touch of G28907: signal is true;
	signal G28910: std_logic; attribute dont_touch of G28910: signal is true;
	signal G28911: std_logic; attribute dont_touch of G28911: signal is true;
	signal G28914: std_logic; attribute dont_touch of G28914: signal is true;
	signal G28917: std_logic; attribute dont_touch of G28917: signal is true;
	signal G28918: std_logic; attribute dont_touch of G28918: signal is true;
	signal G28919: std_logic; attribute dont_touch of G28919: signal is true;
	signal G28920: std_logic; attribute dont_touch of G28920: signal is true;
	signal G28923: std_logic; attribute dont_touch of G28923: signal is true;
	signal G28924: std_logic; attribute dont_touch of G28924: signal is true;
	signal G28927: std_logic; attribute dont_touch of G28927: signal is true;
	signal G28930: std_logic; attribute dont_touch of G28930: signal is true;
	signal G28931: std_logic; attribute dont_touch of G28931: signal is true;
	signal G28934: std_logic; attribute dont_touch of G28934: signal is true;
	signal G28935: std_logic; attribute dont_touch of G28935: signal is true;
	signal G28938: std_logic; attribute dont_touch of G28938: signal is true;
	signal G28939: std_logic; attribute dont_touch of G28939: signal is true;
	signal G28942: std_logic; attribute dont_touch of G28942: signal is true;
	signal G28945: std_logic; attribute dont_touch of G28945: signal is true;
	signal G28946: std_logic; attribute dont_touch of G28946: signal is true;
	signal G28949: std_logic; attribute dont_touch of G28949: signal is true;
	signal G28950: std_logic; attribute dont_touch of G28950: signal is true;
	signal G28953: std_logic; attribute dont_touch of G28953: signal is true;
	signal G28954: std_logic; attribute dont_touch of G28954: signal is true;
	signal G28955: std_logic; attribute dont_touch of G28955: signal is true;
	signal G28958: std_logic; attribute dont_touch of G28958: signal is true;
	signal G28959: std_logic; attribute dont_touch of G28959: signal is true;
	signal G28962: std_logic; attribute dont_touch of G28962: signal is true;
	signal G28965: std_logic; attribute dont_touch of G28965: signal is true;
	signal G28966: std_logic; attribute dont_touch of G28966: signal is true;
	signal G28969: std_logic; attribute dont_touch of G28969: signal is true;
	signal G28970: std_logic; attribute dont_touch of G28970: signal is true;
	signal G28973: std_logic; attribute dont_touch of G28973: signal is true;
	signal G28976: std_logic; attribute dont_touch of G28976: signal is true;
	signal G28977: std_logic; attribute dont_touch of G28977: signal is true;
	signal G28980: std_logic; attribute dont_touch of G28980: signal is true;
	signal G28981: std_logic; attribute dont_touch of G28981: signal is true;
	signal G28982: std_logic; attribute dont_touch of G28982: signal is true;
	signal G28986: std_logic; attribute dont_touch of G28986: signal is true;
	signal G28987: std_logic; attribute dont_touch of G28987: signal is true;
	signal G28990: std_logic; attribute dont_touch of G28990: signal is true;
	signal G28991: std_logic; attribute dont_touch of G28991: signal is true;
	signal G28994: std_logic; attribute dont_touch of G28994: signal is true;
	signal G28997: std_logic; attribute dont_touch of G28997: signal is true;
	signal G28998: std_logic; attribute dont_touch of G28998: signal is true;
	signal G29001: std_logic; attribute dont_touch of G29001: signal is true;
	signal G29004: std_logic; attribute dont_touch of G29004: signal is true;
	signal G29005: std_logic; attribute dont_touch of G29005: signal is true;
	signal G29006: std_logic; attribute dont_touch of G29006: signal is true;
	signal G29007: std_logic; attribute dont_touch of G29007: signal is true;
	signal G29008: std_logic; attribute dont_touch of G29008: signal is true;
	signal G29012: std_logic; attribute dont_touch of G29012: signal is true;
	signal G29013: std_logic; attribute dont_touch of G29013: signal is true;
	signal G29014: std_logic; attribute dont_touch of G29014: signal is true;
	signal G29015: std_logic; attribute dont_touch of G29015: signal is true;
	signal G29018: std_logic; attribute dont_touch of G29018: signal is true;
	signal G29025: std_logic; attribute dont_touch of G29025: signal is true;
	signal G29028: std_logic; attribute dont_touch of G29028: signal is true;
	signal G29029: std_logic; attribute dont_touch of G29029: signal is true;
	signal G29032: std_logic; attribute dont_touch of G29032: signal is true;
	signal G29033: std_logic; attribute dont_touch of G29033: signal is true;
	signal G29034: std_logic; attribute dont_touch of G29034: signal is true;
	signal G29035: std_logic; attribute dont_touch of G29035: signal is true;
	signal G29036: std_logic; attribute dont_touch of G29036: signal is true;
	signal G29040: std_logic; attribute dont_touch of G29040: signal is true;
	signal G29041: std_logic; attribute dont_touch of G29041: signal is true;
	signal G29042: std_logic; attribute dont_touch of G29042: signal is true;
	signal G29043: std_logic; attribute dont_touch of G29043: signal is true;
	signal G29044: std_logic; attribute dont_touch of G29044: signal is true;
	signal G29045: std_logic; attribute dont_touch of G29045: signal is true;
	signal G29046: std_logic; attribute dont_touch of G29046: signal is true;
	signal G29049: std_logic; attribute dont_touch of G29049: signal is true;
	signal G29056: std_logic; attribute dont_touch of G29056: signal is true;
	signal G29057: std_logic; attribute dont_touch of G29057: signal is true;
	signal G29060: std_logic; attribute dont_touch of G29060: signal is true;
	signal G29067: std_logic; attribute dont_touch of G29067: signal is true;
	signal G29068: std_logic; attribute dont_touch of G29068: signal is true;
	signal G29069: std_logic; attribute dont_touch of G29069: signal is true;
	signal G29070: std_logic; attribute dont_touch of G29070: signal is true;
	signal G29071: std_logic; attribute dont_touch of G29071: signal is true;
	signal G29072: std_logic; attribute dont_touch of G29072: signal is true;
	signal G29073: std_logic; attribute dont_touch of G29073: signal is true;
	signal G29077: std_logic; attribute dont_touch of G29077: signal is true;
	signal G29078: std_logic; attribute dont_touch of G29078: signal is true;
	signal G29079: std_logic; attribute dont_touch of G29079: signal is true;
	signal G29080: std_logic; attribute dont_touch of G29080: signal is true;
	signal G29081: std_logic; attribute dont_touch of G29081: signal is true;
	signal G29082: std_logic; attribute dont_touch of G29082: signal is true;
	signal G29085: std_logic; attribute dont_touch of G29085: signal is true;
	signal G29092: std_logic; attribute dont_touch of G29092: signal is true;
	signal G29093: std_logic; attribute dont_touch of G29093: signal is true;
	signal G29094: std_logic; attribute dont_touch of G29094: signal is true;
	signal G29097: std_logic; attribute dont_touch of G29097: signal is true;
	signal G29104: std_logic; attribute dont_touch of G29104: signal is true;
	signal G29105: std_logic; attribute dont_touch of G29105: signal is true;
	signal G29106: std_logic; attribute dont_touch of G29106: signal is true;
	signal G29107: std_logic; attribute dont_touch of G29107: signal is true;
	signal G29108: std_logic; attribute dont_touch of G29108: signal is true;
	signal G29109: std_logic; attribute dont_touch of G29109: signal is true;
	signal G29110: std_logic; attribute dont_touch of G29110: signal is true;
	signal G29114: std_logic; attribute dont_touch of G29114: signal is true;
	signal G29115: std_logic; attribute dont_touch of G29115: signal is true;
	signal G29116: std_logic; attribute dont_touch of G29116: signal is true;
	signal G29117: std_logic; attribute dont_touch of G29117: signal is true;
	signal G29118: std_logic; attribute dont_touch of G29118: signal is true;
	signal G29121: std_logic; attribute dont_touch of G29121: signal is true;
	signal G29128: std_logic; attribute dont_touch of G29128: signal is true;
	signal G29129: std_logic; attribute dont_touch of G29129: signal is true;
	signal G29130: std_logic; attribute dont_touch of G29130: signal is true;
	signal G29131: std_logic; attribute dont_touch of G29131: signal is true;
	signal G29134: std_logic; attribute dont_touch of G29134: signal is true;
	signal G29141: std_logic; attribute dont_touch of G29141: signal is true;
	signal G29142: std_logic; attribute dont_touch of G29142: signal is true;
	signal G29143: std_logic; attribute dont_touch of G29143: signal is true;
	signal G29144: std_logic; attribute dont_touch of G29144: signal is true;
	signal G29145: std_logic; attribute dont_touch of G29145: signal is true;
	signal G29146: std_logic; attribute dont_touch of G29146: signal is true;
	signal G29147: std_logic; attribute dont_touch of G29147: signal is true;
	signal G29148: std_logic; attribute dont_touch of G29148: signal is true;
	signal G29149: std_logic; attribute dont_touch of G29149: signal is true;
	signal G29150: std_logic; attribute dont_touch of G29150: signal is true;
	signal G29151: std_logic; attribute dont_touch of G29151: signal is true;
	signal G29152: std_logic; attribute dont_touch of G29152: signal is true;
	signal G29153: std_logic; attribute dont_touch of G29153: signal is true;
	signal G29154: std_logic; attribute dont_touch of G29154: signal is true;
	signal G29157: std_logic; attribute dont_touch of G29157: signal is true;
	signal G29164: std_logic; attribute dont_touch of G29164: signal is true;
	signal G29165: std_logic; attribute dont_touch of G29165: signal is true;
	signal G29166: std_logic; attribute dont_touch of G29166: signal is true;
	signal G29167: std_logic; attribute dont_touch of G29167: signal is true;
	signal G29168: std_logic; attribute dont_touch of G29168: signal is true;
	signal G29169: std_logic; attribute dont_touch of G29169: signal is true;
	signal G29170: std_logic; attribute dont_touch of G29170: signal is true;
	signal G29171: std_logic; attribute dont_touch of G29171: signal is true;
	signal G29172: std_logic; attribute dont_touch of G29172: signal is true;
	signal G29173: std_logic; attribute dont_touch of G29173: signal is true;
	signal G29174: std_logic; attribute dont_touch of G29174: signal is true;
	signal G29175: std_logic; attribute dont_touch of G29175: signal is true;
	signal G29176: std_logic; attribute dont_touch of G29176: signal is true;
	signal G29177: std_logic; attribute dont_touch of G29177: signal is true;
	signal G29178: std_logic; attribute dont_touch of G29178: signal is true;
	signal G29179: std_logic; attribute dont_touch of G29179: signal is true;
	signal G29180: std_logic; attribute dont_touch of G29180: signal is true;
	signal G29181: std_logic; attribute dont_touch of G29181: signal is true;
	signal G29182: std_logic; attribute dont_touch of G29182: signal is true;
	signal G29183: std_logic; attribute dont_touch of G29183: signal is true;
	signal G29184: std_logic; attribute dont_touch of G29184: signal is true;
	signal G29185: std_logic; attribute dont_touch of G29185: signal is true;
	signal G29186: std_logic; attribute dont_touch of G29186: signal is true;
	signal G29187: std_logic; attribute dont_touch of G29187: signal is true;
	signal G29188: std_logic; attribute dont_touch of G29188: signal is true;
	signal G29189: std_logic; attribute dont_touch of G29189: signal is true;
	signal G29190: std_logic; attribute dont_touch of G29190: signal is true;
	signal G29191: std_logic; attribute dont_touch of G29191: signal is true;
	signal G29192: std_logic; attribute dont_touch of G29192: signal is true;
	signal G29193: std_logic; attribute dont_touch of G29193: signal is true;
	signal G29194: std_logic; attribute dont_touch of G29194: signal is true;
	signal G29195: std_logic; attribute dont_touch of G29195: signal is true;
	signal G29196: std_logic; attribute dont_touch of G29196: signal is true;
	signal G29197: std_logic; attribute dont_touch of G29197: signal is true;
	signal G29198: std_logic; attribute dont_touch of G29198: signal is true;
	signal G29199: std_logic; attribute dont_touch of G29199: signal is true;
	signal G29200: std_logic; attribute dont_touch of G29200: signal is true;
	signal G29201: std_logic; attribute dont_touch of G29201: signal is true;
	signal G29202: std_logic; attribute dont_touch of G29202: signal is true;
	signal G29203: std_logic; attribute dont_touch of G29203: signal is true;
	signal G29204: std_logic; attribute dont_touch of G29204: signal is true;
	signal G29205: std_logic; attribute dont_touch of G29205: signal is true;
	signal G29206: std_logic; attribute dont_touch of G29206: signal is true;
	signal G29207: std_logic; attribute dont_touch of G29207: signal is true;
	signal G29208: std_logic; attribute dont_touch of G29208: signal is true;
	signal G29209: std_logic; attribute dont_touch of G29209: signal is true;
	signal G29222: std_logic; attribute dont_touch of G29222: signal is true;
	signal G29223: std_logic; attribute dont_touch of G29223: signal is true;
	signal G29224: std_logic; attribute dont_touch of G29224: signal is true;
	signal G29225: std_logic; attribute dont_touch of G29225: signal is true;
	signal G29226: std_logic; attribute dont_touch of G29226: signal is true;
	signal G29227: std_logic; attribute dont_touch of G29227: signal is true;
	signal G29228: std_logic; attribute dont_touch of G29228: signal is true;
	signal G29229: std_logic; attribute dont_touch of G29229: signal is true;
	signal G29230: std_logic; attribute dont_touch of G29230: signal is true;
	signal G29231: std_logic; attribute dont_touch of G29231: signal is true;
	signal G29232: std_logic; attribute dont_touch of G29232: signal is true;
	signal G29233: std_logic; attribute dont_touch of G29233: signal is true;
	signal G29234: std_logic; attribute dont_touch of G29234: signal is true;
	signal G29235: std_logic; attribute dont_touch of G29235: signal is true;
	signal G29236: std_logic; attribute dont_touch of G29236: signal is true;
	signal G29237: std_logic; attribute dont_touch of G29237: signal is true;
	signal G29238: std_logic; attribute dont_touch of G29238: signal is true;
	signal G29239: std_logic; attribute dont_touch of G29239: signal is true;
	signal G29240: std_logic; attribute dont_touch of G29240: signal is true;
	signal G29241: std_logic; attribute dont_touch of G29241: signal is true;
	signal G29242: std_logic; attribute dont_touch of G29242: signal is true;
	signal G29243: std_logic; attribute dont_touch of G29243: signal is true;
	signal G29244: std_logic; attribute dont_touch of G29244: signal is true;
	signal G29245: std_logic; attribute dont_touch of G29245: signal is true;
	signal G29246: std_logic; attribute dont_touch of G29246: signal is true;
	signal G29247: std_logic; attribute dont_touch of G29247: signal is true;
	signal G29248: std_logic; attribute dont_touch of G29248: signal is true;
	signal G29249: std_logic; attribute dont_touch of G29249: signal is true;
	signal G29250: std_logic; attribute dont_touch of G29250: signal is true;
	signal G29251: std_logic; attribute dont_touch of G29251: signal is true;
	signal G29252: std_logic; attribute dont_touch of G29252: signal is true;
	signal G29253: std_logic; attribute dont_touch of G29253: signal is true;
	signal G29254: std_logic; attribute dont_touch of G29254: signal is true;
	signal G29255: std_logic; attribute dont_touch of G29255: signal is true;
	signal G29256: std_logic; attribute dont_touch of G29256: signal is true;
	signal G29257: std_logic; attribute dont_touch of G29257: signal is true;
	signal G29258: std_logic; attribute dont_touch of G29258: signal is true;
	signal G29259: std_logic; attribute dont_touch of G29259: signal is true;
	signal G29260: std_logic; attribute dont_touch of G29260: signal is true;
	signal G29261: std_logic; attribute dont_touch of G29261: signal is true;
	signal G29262: std_logic; attribute dont_touch of G29262: signal is true;
	signal G29263: std_logic; attribute dont_touch of G29263: signal is true;
	signal G29264: std_logic; attribute dont_touch of G29264: signal is true;
	signal G29265: std_logic; attribute dont_touch of G29265: signal is true;
	signal G29266: std_logic; attribute dont_touch of G29266: signal is true;
	signal G29267: std_logic; attribute dont_touch of G29267: signal is true;
	signal G29268: std_logic; attribute dont_touch of G29268: signal is true;
	signal G29269: std_logic; attribute dont_touch of G29269: signal is true;
	signal G29270: std_logic; attribute dont_touch of G29270: signal is true;
	signal G29271: std_logic; attribute dont_touch of G29271: signal is true;
	signal G29272: std_logic; attribute dont_touch of G29272: signal is true;
	signal G29273: std_logic; attribute dont_touch of G29273: signal is true;
	signal G29274: std_logic; attribute dont_touch of G29274: signal is true;
	signal G29275: std_logic; attribute dont_touch of G29275: signal is true;
	signal G29276: std_logic; attribute dont_touch of G29276: signal is true;
	signal G29277: std_logic; attribute dont_touch of G29277: signal is true;
	signal G29278: std_logic; attribute dont_touch of G29278: signal is true;
	signal G29279: std_logic; attribute dont_touch of G29279: signal is true;
	signal G29280: std_logic; attribute dont_touch of G29280: signal is true;
	signal G29281: std_logic; attribute dont_touch of G29281: signal is true;
	signal G29282: std_logic; attribute dont_touch of G29282: signal is true;
	signal G29283: std_logic; attribute dont_touch of G29283: signal is true;
	signal G29284: std_logic; attribute dont_touch of G29284: signal is true;
	signal G29285: std_logic; attribute dont_touch of G29285: signal is true;
	signal G29286: std_logic; attribute dont_touch of G29286: signal is true;
	signal G29287: std_logic; attribute dont_touch of G29287: signal is true;
	signal G29288: std_logic; attribute dont_touch of G29288: signal is true;
	signal G29289: std_logic; attribute dont_touch of G29289: signal is true;
	signal G29290: std_logic; attribute dont_touch of G29290: signal is true;
	signal G29291: std_logic; attribute dont_touch of G29291: signal is true;
	signal G29292: std_logic; attribute dont_touch of G29292: signal is true;
	signal G29293: std_logic; attribute dont_touch of G29293: signal is true;
	signal G29294: std_logic; attribute dont_touch of G29294: signal is true;
	signal G29295: std_logic; attribute dont_touch of G29295: signal is true;
	signal G29296: std_logic; attribute dont_touch of G29296: signal is true;
	signal G29297: std_logic; attribute dont_touch of G29297: signal is true;
	signal G29298: std_logic; attribute dont_touch of G29298: signal is true;
	signal G29299: std_logic; attribute dont_touch of G29299: signal is true;
	signal G29300: std_logic; attribute dont_touch of G29300: signal is true;
	signal G29301: std_logic; attribute dont_touch of G29301: signal is true;
	signal G29302: std_logic; attribute dont_touch of G29302: signal is true;
	signal G29303: std_logic; attribute dont_touch of G29303: signal is true;
	signal G29304: std_logic; attribute dont_touch of G29304: signal is true;
	signal G29305: std_logic; attribute dont_touch of G29305: signal is true;
	signal G29306: std_logic; attribute dont_touch of G29306: signal is true;
	signal G29307: std_logic; attribute dont_touch of G29307: signal is true;
	signal G29308: std_logic; attribute dont_touch of G29308: signal is true;
	signal G29309: std_logic; attribute dont_touch of G29309: signal is true;
	signal G29310: std_logic; attribute dont_touch of G29310: signal is true;
	signal G29311: std_logic; attribute dont_touch of G29311: signal is true;
	signal G29312: std_logic; attribute dont_touch of G29312: signal is true;
	signal G29313: std_logic; attribute dont_touch of G29313: signal is true;
	signal G29314: std_logic; attribute dont_touch of G29314: signal is true;
	signal G29315: std_logic; attribute dont_touch of G29315: signal is true;
	signal G29316: std_logic; attribute dont_touch of G29316: signal is true;
	signal G29317: std_logic; attribute dont_touch of G29317: signal is true;
	signal G29318: std_logic; attribute dont_touch of G29318: signal is true;
	signal G29319: std_logic; attribute dont_touch of G29319: signal is true;
	signal G29320: std_logic; attribute dont_touch of G29320: signal is true;
	signal G29321: std_logic; attribute dont_touch of G29321: signal is true;
	signal G29322: std_logic; attribute dont_touch of G29322: signal is true;
	signal G29323: std_logic; attribute dont_touch of G29323: signal is true;
	signal G29324: std_logic; attribute dont_touch of G29324: signal is true;
	signal G29325: std_logic; attribute dont_touch of G29325: signal is true;
	signal G29326: std_logic; attribute dont_touch of G29326: signal is true;
	signal G29327: std_logic; attribute dont_touch of G29327: signal is true;
	signal G29328: std_logic; attribute dont_touch of G29328: signal is true;
	signal G29329: std_logic; attribute dont_touch of G29329: signal is true;
	signal G29330: std_logic; attribute dont_touch of G29330: signal is true;
	signal G29331: std_logic; attribute dont_touch of G29331: signal is true;
	signal G29332: std_logic; attribute dont_touch of G29332: signal is true;
	signal G29333: std_logic; attribute dont_touch of G29333: signal is true;
	signal G29334: std_logic; attribute dont_touch of G29334: signal is true;
	signal G29335: std_logic; attribute dont_touch of G29335: signal is true;
	signal G29336: std_logic; attribute dont_touch of G29336: signal is true;
	signal G29337: std_logic; attribute dont_touch of G29337: signal is true;
	signal G29338: std_logic; attribute dont_touch of G29338: signal is true;
	signal G29339: std_logic; attribute dont_touch of G29339: signal is true;
	signal G29342: std_logic; attribute dont_touch of G29342: signal is true;
	signal G29343: std_logic; attribute dont_touch of G29343: signal is true;
	signal G29344: std_logic; attribute dont_touch of G29344: signal is true;
	signal G29345: std_logic; attribute dont_touch of G29345: signal is true;
	signal G29346: std_logic; attribute dont_touch of G29346: signal is true;
	signal G29347: std_logic; attribute dont_touch of G29347: signal is true;
	signal G29348: std_logic; attribute dont_touch of G29348: signal is true;
	signal G29349: std_logic; attribute dont_touch of G29349: signal is true;
	signal G29350: std_logic; attribute dont_touch of G29350: signal is true;
	signal G29351: std_logic; attribute dont_touch of G29351: signal is true;
	signal G29352: std_logic; attribute dont_touch of G29352: signal is true;
	signal G29353: std_logic; attribute dont_touch of G29353: signal is true;
	signal G29354: std_logic; attribute dont_touch of G29354: signal is true;
	signal G29355: std_logic; attribute dont_touch of G29355: signal is true;
	signal G29358: std_logic; attribute dont_touch of G29358: signal is true;
	signal G29359: std_logic; attribute dont_touch of G29359: signal is true;
	signal G29360: std_logic; attribute dont_touch of G29360: signal is true;
	signal G29361: std_logic; attribute dont_touch of G29361: signal is true;
	signal G29362: std_logic; attribute dont_touch of G29362: signal is true;
	signal G29363: std_logic; attribute dont_touch of G29363: signal is true;
	signal G29364: std_logic; attribute dont_touch of G29364: signal is true;
	signal G29365: std_logic; attribute dont_touch of G29365: signal is true;
	signal G29366: std_logic; attribute dont_touch of G29366: signal is true;
	signal G29367: std_logic; attribute dont_touch of G29367: signal is true;
	signal G29368: std_logic; attribute dont_touch of G29368: signal is true;
	signal G29369: std_logic; attribute dont_touch of G29369: signal is true;
	signal G29370: std_logic; attribute dont_touch of G29370: signal is true;
	signal G29371: std_logic; attribute dont_touch of G29371: signal is true;
	signal G29372: std_logic; attribute dont_touch of G29372: signal is true;
	signal G29373: std_logic; attribute dont_touch of G29373: signal is true;
	signal G29374: std_logic; attribute dont_touch of G29374: signal is true;
	signal G29375: std_logic; attribute dont_touch of G29375: signal is true;
	signal G29376: std_logic; attribute dont_touch of G29376: signal is true;
	signal G29377: std_logic; attribute dont_touch of G29377: signal is true;
	signal G29378: std_logic; attribute dont_touch of G29378: signal is true;
	signal G29379: std_logic; attribute dont_touch of G29379: signal is true;
	signal G29380: std_logic; attribute dont_touch of G29380: signal is true;
	signal G29381: std_logic; attribute dont_touch of G29381: signal is true;
	signal G29382: std_logic; attribute dont_touch of G29382: signal is true;
	signal G29383: std_logic; attribute dont_touch of G29383: signal is true;
	signal G29384: std_logic; attribute dont_touch of G29384: signal is true;
	signal G29385: std_logic; attribute dont_touch of G29385: signal is true;
	signal G29474: std_logic; attribute dont_touch of G29474: signal is true;
	signal G29475: std_logic; attribute dont_touch of G29475: signal is true;
	signal G29476: std_logic; attribute dont_touch of G29476: signal is true;
	signal G29477: std_logic; attribute dont_touch of G29477: signal is true;
	signal G29478: std_logic; attribute dont_touch of G29478: signal is true;
	signal G29479: std_logic; attribute dont_touch of G29479: signal is true;
	signal G29480: std_logic; attribute dont_touch of G29480: signal is true;
	signal G29481: std_logic; attribute dont_touch of G29481: signal is true;
	signal G29482: std_logic; attribute dont_touch of G29482: signal is true;
	signal G29483: std_logic; attribute dont_touch of G29483: signal is true;
	signal G29484: std_logic; attribute dont_touch of G29484: signal is true;
	signal G29485: std_logic; attribute dont_touch of G29485: signal is true;
	signal G29486: std_logic; attribute dont_touch of G29486: signal is true;
	signal G29487: std_logic; attribute dont_touch of G29487: signal is true;
	signal G29488: std_logic; attribute dont_touch of G29488: signal is true;
	signal G29489: std_logic; attribute dont_touch of G29489: signal is true;
	signal G29490: std_logic; attribute dont_touch of G29490: signal is true;
	signal G29491: std_logic; attribute dont_touch of G29491: signal is true;
	signal G29494: std_logic; attribute dont_touch of G29494: signal is true;
	signal G29495: std_logic; attribute dont_touch of G29495: signal is true;
	signal G29496: std_logic; attribute dont_touch of G29496: signal is true;
	signal G29497: std_logic; attribute dont_touch of G29497: signal is true;
	signal G29498: std_logic; attribute dont_touch of G29498: signal is true;
	signal G29501: std_logic; attribute dont_touch of G29501: signal is true;
	signal G29502: std_logic; attribute dont_touch of G29502: signal is true;
	signal G29503: std_logic; attribute dont_touch of G29503: signal is true;
	signal G29504: std_logic; attribute dont_touch of G29504: signal is true;
	signal G29505: std_logic; attribute dont_touch of G29505: signal is true;
	signal G29506: std_logic; attribute dont_touch of G29506: signal is true;
	signal G29507: std_logic; attribute dont_touch of G29507: signal is true;
	signal G29508: std_logic; attribute dont_touch of G29508: signal is true;
	signal G29509: std_logic; attribute dont_touch of G29509: signal is true;
	signal G29510: std_logic; attribute dont_touch of G29510: signal is true;
	signal G29511: std_logic; attribute dont_touch of G29511: signal is true;
	signal G29512: std_logic; attribute dont_touch of G29512: signal is true;
	signal G29513: std_logic; attribute dont_touch of G29513: signal is true;
	signal G29514: std_logic; attribute dont_touch of G29514: signal is true;
	signal G29515: std_logic; attribute dont_touch of G29515: signal is true;
	signal G29516: std_logic; attribute dont_touch of G29516: signal is true;
	signal G29517: std_logic; attribute dont_touch of G29517: signal is true;
	signal G29518: std_logic; attribute dont_touch of G29518: signal is true;
	signal G29519: std_logic; attribute dont_touch of G29519: signal is true;
	signal G29520: std_logic; attribute dont_touch of G29520: signal is true;
	signal G29521: std_logic; attribute dont_touch of G29521: signal is true;
	signal G29522: std_logic; attribute dont_touch of G29522: signal is true;
	signal G29523: std_logic; attribute dont_touch of G29523: signal is true;
	signal G29524: std_logic; attribute dont_touch of G29524: signal is true;
	signal G29525: std_logic; attribute dont_touch of G29525: signal is true;
	signal G29526: std_logic; attribute dont_touch of G29526: signal is true;
	signal G29527: std_logic; attribute dont_touch of G29527: signal is true;
	signal G29528: std_logic; attribute dont_touch of G29528: signal is true;
	signal G29529: std_logic; attribute dont_touch of G29529: signal is true;
	signal G29530: std_logic; attribute dont_touch of G29530: signal is true;
	signal G29531: std_logic; attribute dont_touch of G29531: signal is true;
	signal G29532: std_logic; attribute dont_touch of G29532: signal is true;
	signal G29533: std_logic; attribute dont_touch of G29533: signal is true;
	signal G29534: std_logic; attribute dont_touch of G29534: signal is true;
	signal G29535: std_logic; attribute dont_touch of G29535: signal is true;
	signal G29536: std_logic; attribute dont_touch of G29536: signal is true;
	signal G29537: std_logic; attribute dont_touch of G29537: signal is true;
	signal G29538: std_logic; attribute dont_touch of G29538: signal is true;
	signal G29539: std_logic; attribute dont_touch of G29539: signal is true;
	signal G29540: std_logic; attribute dont_touch of G29540: signal is true;
	signal G29547: std_logic; attribute dont_touch of G29547: signal is true;
	signal G29548: std_logic; attribute dont_touch of G29548: signal is true;
	signal G29549: std_logic; attribute dont_touch of G29549: signal is true;
	signal G29550: std_logic; attribute dont_touch of G29550: signal is true;
	signal G29551: std_logic; attribute dont_touch of G29551: signal is true;
	signal G29552: std_logic; attribute dont_touch of G29552: signal is true;
	signal G29553: std_logic; attribute dont_touch of G29553: signal is true;
	signal G29554: std_logic; attribute dont_touch of G29554: signal is true;
	signal G29555: std_logic; attribute dont_touch of G29555: signal is true;
	signal G29556: std_logic; attribute dont_touch of G29556: signal is true;
	signal G29563: std_logic; attribute dont_touch of G29563: signal is true;
	signal G29564: std_logic; attribute dont_touch of G29564: signal is true;
	signal G29565: std_logic; attribute dont_touch of G29565: signal is true;
	signal G29566: std_logic; attribute dont_touch of G29566: signal is true;
	signal G29567: std_logic; attribute dont_touch of G29567: signal is true;
	signal G29568: std_logic; attribute dont_touch of G29568: signal is true;
	signal G29569: std_logic; attribute dont_touch of G29569: signal is true;
	signal G29570: std_logic; attribute dont_touch of G29570: signal is true;
	signal G29571: std_logic; attribute dont_touch of G29571: signal is true;
	signal G29572: std_logic; attribute dont_touch of G29572: signal is true;
	signal G29573: std_logic; attribute dont_touch of G29573: signal is true;
	signal G29574: std_logic; attribute dont_touch of G29574: signal is true;
	signal G29575: std_logic; attribute dont_touch of G29575: signal is true;
	signal G29576: std_logic; attribute dont_touch of G29576: signal is true;
	signal G29577: std_logic; attribute dont_touch of G29577: signal is true;
	signal G29578: std_logic; attribute dont_touch of G29578: signal is true;
	signal G29579: std_logic; attribute dont_touch of G29579: signal is true;
	signal G29580: std_logic; attribute dont_touch of G29580: signal is true;
	signal G29581: std_logic; attribute dont_touch of G29581: signal is true;
	signal G29582: std_logic; attribute dont_touch of G29582: signal is true;
	signal G29583: std_logic; attribute dont_touch of G29583: signal is true;
	signal G29584: std_logic; attribute dont_touch of G29584: signal is true;
	signal G29585: std_logic; attribute dont_touch of G29585: signal is true;
	signal G29586: std_logic; attribute dont_touch of G29586: signal is true;
	signal G29587: std_logic; attribute dont_touch of G29587: signal is true;
	signal G29588: std_logic; attribute dont_touch of G29588: signal is true;
	signal G29589: std_logic; attribute dont_touch of G29589: signal is true;
	signal G29590: std_logic; attribute dont_touch of G29590: signal is true;
	signal G29591: std_logic; attribute dont_touch of G29591: signal is true;
	signal G29592: std_logic; attribute dont_touch of G29592: signal is true;
	signal G29593: std_logic; attribute dont_touch of G29593: signal is true;
	signal G29594: std_logic; attribute dont_touch of G29594: signal is true;
	signal G29595: std_logic; attribute dont_touch of G29595: signal is true;
	signal G29596: std_logic; attribute dont_touch of G29596: signal is true;
	signal G29597: std_logic; attribute dont_touch of G29597: signal is true;
	signal G29598: std_logic; attribute dont_touch of G29598: signal is true;
	signal G29599: std_logic; attribute dont_touch of G29599: signal is true;
	signal G29600: std_logic; attribute dont_touch of G29600: signal is true;
	signal G29601: std_logic; attribute dont_touch of G29601: signal is true;
	signal G29602: std_logic; attribute dont_touch of G29602: signal is true;
	signal G29603: std_logic; attribute dont_touch of G29603: signal is true;
	signal G29604: std_logic; attribute dont_touch of G29604: signal is true;
	signal G29605: std_logic; attribute dont_touch of G29605: signal is true;
	signal G29606: std_logic; attribute dont_touch of G29606: signal is true;
	signal G29607: std_logic; attribute dont_touch of G29607: signal is true;
	signal G29608: std_logic; attribute dont_touch of G29608: signal is true;
	signal G29609: std_logic; attribute dont_touch of G29609: signal is true;
	signal G29610: std_logic; attribute dont_touch of G29610: signal is true;
	signal G29611: std_logic; attribute dont_touch of G29611: signal is true;
	signal G29612: std_logic; attribute dont_touch of G29612: signal is true;
	signal G29613: std_logic; attribute dont_touch of G29613: signal is true;
	signal G29614: std_logic; attribute dont_touch of G29614: signal is true;
	signal G29615: std_logic; attribute dont_touch of G29615: signal is true;
	signal G29616: std_logic; attribute dont_touch of G29616: signal is true;
	signal G29617: std_logic; attribute dont_touch of G29617: signal is true;
	signal G29618: std_logic; attribute dont_touch of G29618: signal is true;
	signal G29619: std_logic; attribute dont_touch of G29619: signal is true;
	signal G29620: std_logic; attribute dont_touch of G29620: signal is true;
	signal G29621: std_logic; attribute dont_touch of G29621: signal is true;
	signal G29622: std_logic; attribute dont_touch of G29622: signal is true;
	signal G29623: std_logic; attribute dont_touch of G29623: signal is true;
	signal G29624: std_logic; attribute dont_touch of G29624: signal is true;
	signal G29625: std_logic; attribute dont_touch of G29625: signal is true;
	signal G29626: std_logic; attribute dont_touch of G29626: signal is true;
	signal G29627: std_logic; attribute dont_touch of G29627: signal is true;
	signal G29628: std_logic; attribute dont_touch of G29628: signal is true;
	signal G29629: std_logic; attribute dont_touch of G29629: signal is true;
	signal G29630: std_logic; attribute dont_touch of G29630: signal is true;
	signal G29631: std_logic; attribute dont_touch of G29631: signal is true;
	signal G29632: std_logic; attribute dont_touch of G29632: signal is true;
	signal G29633: std_logic; attribute dont_touch of G29633: signal is true;
	signal G29634: std_logic; attribute dont_touch of G29634: signal is true;
	signal G29635: std_logic; attribute dont_touch of G29635: signal is true;
	signal G29636: std_logic; attribute dont_touch of G29636: signal is true;
	signal G29637: std_logic; attribute dont_touch of G29637: signal is true;
	signal G29638: std_logic; attribute dont_touch of G29638: signal is true;
	signal G29639: std_logic; attribute dont_touch of G29639: signal is true;
	signal G29640: std_logic; attribute dont_touch of G29640: signal is true;
	signal G29641: std_logic; attribute dont_touch of G29641: signal is true;
	signal G29642: std_logic; attribute dont_touch of G29642: signal is true;
	signal G29643: std_logic; attribute dont_touch of G29643: signal is true;
	signal G29644: std_logic; attribute dont_touch of G29644: signal is true;
	signal G29645: std_logic; attribute dont_touch of G29645: signal is true;
	signal G29646: std_logic; attribute dont_touch of G29646: signal is true;
	signal G29647: std_logic; attribute dont_touch of G29647: signal is true;
	signal G29648: std_logic; attribute dont_touch of G29648: signal is true;
	signal G29649: std_logic; attribute dont_touch of G29649: signal is true;
	signal G29650: std_logic; attribute dont_touch of G29650: signal is true;
	signal G29651: std_logic; attribute dont_touch of G29651: signal is true;
	signal G29652: std_logic; attribute dont_touch of G29652: signal is true;
	signal G29653: std_logic; attribute dont_touch of G29653: signal is true;
	signal G29656: std_logic; attribute dont_touch of G29656: signal is true;
	signal G29657: std_logic; attribute dont_touch of G29657: signal is true;
	signal G29660: std_logic; attribute dont_touch of G29660: signal is true;
	signal G29661: std_logic; attribute dont_touch of G29661: signal is true;
	signal G29662: std_logic; attribute dont_touch of G29662: signal is true;
	signal G29663: std_logic; attribute dont_touch of G29663: signal is true;
	signal G29664: std_logic; attribute dont_touch of G29664: signal is true;
	signal G29665: std_logic; attribute dont_touch of G29665: signal is true;
	signal G29666: std_logic; attribute dont_touch of G29666: signal is true;
	signal G29667: std_logic; attribute dont_touch of G29667: signal is true;
	signal G29668: std_logic; attribute dont_touch of G29668: signal is true;
	signal G29669: std_logic; attribute dont_touch of G29669: signal is true;
	signal G29672: std_logic; attribute dont_touch of G29672: signal is true;
	signal G29675: std_logic; attribute dont_touch of G29675: signal is true;
	signal G29676: std_logic; attribute dont_touch of G29676: signal is true;
	signal G29679: std_logic; attribute dont_touch of G29679: signal is true;
	signal G29683: std_logic; attribute dont_touch of G29683: signal is true;
	signal G29684: std_logic; attribute dont_touch of G29684: signal is true;
	signal G29685: std_logic; attribute dont_touch of G29685: signal is true;
	signal G29686: std_logic; attribute dont_touch of G29686: signal is true;
	signal G29687: std_logic; attribute dont_touch of G29687: signal is true;
	signal G29688: std_logic; attribute dont_touch of G29688: signal is true;
	signal G29689: std_logic; attribute dont_touch of G29689: signal is true;
	signal G29692: std_logic; attribute dont_touch of G29692: signal is true;
	signal G29693: std_logic; attribute dont_touch of G29693: signal is true;
	signal G29694: std_logic; attribute dont_touch of G29694: signal is true;
	signal G29697: std_logic; attribute dont_touch of G29697: signal is true;
	signal G29702: std_logic; attribute dont_touch of G29702: signal is true;
	signal G29705: std_logic; attribute dont_touch of G29705: signal is true;
	signal G29706: std_logic; attribute dont_touch of G29706: signal is true;
	signal G29707: std_logic; attribute dont_touch of G29707: signal is true;
	signal G29708: std_logic; attribute dont_touch of G29708: signal is true;
	signal G29709: std_logic; attribute dont_touch of G29709: signal is true;
	signal G29710: std_logic; attribute dont_touch of G29710: signal is true;
	signal G29711: std_logic; attribute dont_touch of G29711: signal is true;
	signal G29712: std_logic; attribute dont_touch of G29712: signal is true;
	signal G29713: std_logic; attribute dont_touch of G29713: signal is true;
	signal G29716: std_logic; attribute dont_touch of G29716: signal is true;
	signal G29717: std_logic; attribute dont_touch of G29717: signal is true;
	signal G29718: std_logic; attribute dont_touch of G29718: signal is true;
	signal G29719: std_logic; attribute dont_touch of G29719: signal is true;
	signal G29722: std_logic; attribute dont_touch of G29722: signal is true;
	signal G29725: std_logic; attribute dont_touch of G29725: signal is true;
	signal G29730: std_logic; attribute dont_touch of G29730: signal is true;
	signal G29731: std_logic; attribute dont_touch of G29731: signal is true;
	signal G29732: std_logic; attribute dont_touch of G29732: signal is true;
	signal G29733: std_logic; attribute dont_touch of G29733: signal is true;
	signal G29734: std_logic; attribute dont_touch of G29734: signal is true;
	signal G29735: std_logic; attribute dont_touch of G29735: signal is true;
	signal G29736: std_logic; attribute dont_touch of G29736: signal is true;
	signal G29737: std_logic; attribute dont_touch of G29737: signal is true;
	signal G29740: std_logic; attribute dont_touch of G29740: signal is true;
	signal G29741: std_logic; attribute dont_touch of G29741: signal is true;
	signal G29742: std_logic; attribute dont_touch of G29742: signal is true;
	signal G29743: std_logic; attribute dont_touch of G29743: signal is true;
	signal G29744: std_logic; attribute dont_touch of G29744: signal is true;
	signal G29745: std_logic; attribute dont_touch of G29745: signal is true;
	signal G29746: std_logic; attribute dont_touch of G29746: signal is true;
	signal G29747: std_logic; attribute dont_touch of G29747: signal is true;
	signal G29748: std_logic; attribute dont_touch of G29748: signal is true;
	signal G29749: std_logic; attribute dont_touch of G29749: signal is true;
	signal G29750: std_logic; attribute dont_touch of G29750: signal is true;
	signal G29751: std_logic; attribute dont_touch of G29751: signal is true;
	signal G29752: std_logic; attribute dont_touch of G29752: signal is true;
	signal G29753: std_logic; attribute dont_touch of G29753: signal is true;
	signal G29754: std_logic; attribute dont_touch of G29754: signal is true;
	signal G29755: std_logic; attribute dont_touch of G29755: signal is true;
	signal G29756: std_logic; attribute dont_touch of G29756: signal is true;
	signal G29757: std_logic; attribute dont_touch of G29757: signal is true;
	signal G29758: std_logic; attribute dont_touch of G29758: signal is true;
	signal G29759: std_logic; attribute dont_touch of G29759: signal is true;
	signal G29760: std_logic; attribute dont_touch of G29760: signal is true;
	signal G29761: std_logic; attribute dont_touch of G29761: signal is true;
	signal G29762: std_logic; attribute dont_touch of G29762: signal is true;
	signal G29763: std_logic; attribute dont_touch of G29763: signal is true;
	signal G29764: std_logic; attribute dont_touch of G29764: signal is true;
	signal G29765: std_logic; attribute dont_touch of G29765: signal is true;
	signal G29766: std_logic; attribute dont_touch of G29766: signal is true;
	signal G29767: std_logic; attribute dont_touch of G29767: signal is true;
	signal G29768: std_logic; attribute dont_touch of G29768: signal is true;
	signal G29769: std_logic; attribute dont_touch of G29769: signal is true;
	signal G29770: std_logic; attribute dont_touch of G29770: signal is true;
	signal G29771: std_logic; attribute dont_touch of G29771: signal is true;
	signal G29772: std_logic; attribute dont_touch of G29772: signal is true;
	signal G29773: std_logic; attribute dont_touch of G29773: signal is true;
	signal G29774: std_logic; attribute dont_touch of G29774: signal is true;
	signal G29775: std_logic; attribute dont_touch of G29775: signal is true;
	signal G29776: std_logic; attribute dont_touch of G29776: signal is true;
	signal G29777: std_logic; attribute dont_touch of G29777: signal is true;
	signal G29778: std_logic; attribute dont_touch of G29778: signal is true;
	signal G29782: std_logic; attribute dont_touch of G29782: signal is true;
	signal G29783: std_logic; attribute dont_touch of G29783: signal is true;
	signal G29784: std_logic; attribute dont_touch of G29784: signal is true;
	signal G29785: std_logic; attribute dont_touch of G29785: signal is true;
	signal G29786: std_logic; attribute dont_touch of G29786: signal is true;
	signal G29787: std_logic; attribute dont_touch of G29787: signal is true;
	signal G29788: std_logic; attribute dont_touch of G29788: signal is true;
	signal G29789: std_logic; attribute dont_touch of G29789: signal is true;
	signal G29790: std_logic; attribute dont_touch of G29790: signal is true;
	signal G29791: std_logic; attribute dont_touch of G29791: signal is true;
	signal G29792: std_logic; attribute dont_touch of G29792: signal is true;
	signal G29793: std_logic; attribute dont_touch of G29793: signal is true;
	signal G29794: std_logic; attribute dont_touch of G29794: signal is true;
	signal G29795: std_logic; attribute dont_touch of G29795: signal is true;
	signal G29796: std_logic; attribute dont_touch of G29796: signal is true;
	signal G29797: std_logic; attribute dont_touch of G29797: signal is true;
	signal G29798: std_logic; attribute dont_touch of G29798: signal is true;
	signal G29799: std_logic; attribute dont_touch of G29799: signal is true;
	signal G29800: std_logic; attribute dont_touch of G29800: signal is true;
	signal G29801: std_logic; attribute dont_touch of G29801: signal is true;
	signal G29802: std_logic; attribute dont_touch of G29802: signal is true;
	signal G29803: std_logic; attribute dont_touch of G29803: signal is true;
	signal G29804: std_logic; attribute dont_touch of G29804: signal is true;
	signal G29805: std_logic; attribute dont_touch of G29805: signal is true;
	signal G29806: std_logic; attribute dont_touch of G29806: signal is true;
	signal G29807: std_logic; attribute dont_touch of G29807: signal is true;
	signal G29808: std_logic; attribute dont_touch of G29808: signal is true;
	signal G29809: std_logic; attribute dont_touch of G29809: signal is true;
	signal G29810: std_logic; attribute dont_touch of G29810: signal is true;
	signal G29811: std_logic; attribute dont_touch of G29811: signal is true;
	signal G29812: std_logic; attribute dont_touch of G29812: signal is true;
	signal G29813: std_logic; attribute dont_touch of G29813: signal is true;
	signal G29814: std_logic; attribute dont_touch of G29814: signal is true;
	signal G29834: std_logic; attribute dont_touch of G29834: signal is true;
	signal G29835: std_logic; attribute dont_touch of G29835: signal is true;
	signal G29836: std_logic; attribute dont_touch of G29836: signal is true;
	signal G29837: std_logic; attribute dont_touch of G29837: signal is true;
	signal G29838: std_logic; attribute dont_touch of G29838: signal is true;
	signal G29839: std_logic; attribute dont_touch of G29839: signal is true;
	signal G29840: std_logic; attribute dont_touch of G29840: signal is true;
	signal G29841: std_logic; attribute dont_touch of G29841: signal is true;
	signal G29842: std_logic; attribute dont_touch of G29842: signal is true;
	signal G29843: std_logic; attribute dont_touch of G29843: signal is true;
	signal G29844: std_logic; attribute dont_touch of G29844: signal is true;
	signal G29845: std_logic; attribute dont_touch of G29845: signal is true;
	signal G29846: std_logic; attribute dont_touch of G29846: signal is true;
	signal G29847: std_logic; attribute dont_touch of G29847: signal is true;
	signal G29848: std_logic; attribute dont_touch of G29848: signal is true;
	signal G29849: std_logic; attribute dont_touch of G29849: signal is true;
	signal G29850: std_logic; attribute dont_touch of G29850: signal is true;
	signal G29851: std_logic; attribute dont_touch of G29851: signal is true;
	signal G29852: std_logic; attribute dont_touch of G29852: signal is true;
	signal G29853: std_logic; attribute dont_touch of G29853: signal is true;
	signal G29854: std_logic; attribute dont_touch of G29854: signal is true;
	signal G29855: std_logic; attribute dont_touch of G29855: signal is true;
	signal G29856: std_logic; attribute dont_touch of G29856: signal is true;
	signal G29857: std_logic; attribute dont_touch of G29857: signal is true;
	signal G29858: std_logic; attribute dont_touch of G29858: signal is true;
	signal G29859: std_logic; attribute dont_touch of G29859: signal is true;
	signal G29860: std_logic; attribute dont_touch of G29860: signal is true;
	signal G29861: std_logic; attribute dont_touch of G29861: signal is true;
	signal G29862: std_logic; attribute dont_touch of G29862: signal is true;
	signal G29863: std_logic; attribute dont_touch of G29863: signal is true;
	signal G29864: std_logic; attribute dont_touch of G29864: signal is true;
	signal G29865: std_logic; attribute dont_touch of G29865: signal is true;
	signal G29866: std_logic; attribute dont_touch of G29866: signal is true;
	signal G29867: std_logic; attribute dont_touch of G29867: signal is true;
	signal G29868: std_logic; attribute dont_touch of G29868: signal is true;
	signal G29869: std_logic; attribute dont_touch of G29869: signal is true;
	signal G29870: std_logic; attribute dont_touch of G29870: signal is true;
	signal G29871: std_logic; attribute dont_touch of G29871: signal is true;
	signal G29872: std_logic; attribute dont_touch of G29872: signal is true;
	signal G29873: std_logic; attribute dont_touch of G29873: signal is true;
	signal G29874: std_logic; attribute dont_touch of G29874: signal is true;
	signal G29875: std_logic; attribute dont_touch of G29875: signal is true;
	signal G29876: std_logic; attribute dont_touch of G29876: signal is true;
	signal G29877: std_logic; attribute dont_touch of G29877: signal is true;
	signal G29878: std_logic; attribute dont_touch of G29878: signal is true;
	signal G29879: std_logic; attribute dont_touch of G29879: signal is true;
	signal G29880: std_logic; attribute dont_touch of G29880: signal is true;
	signal G29881: std_logic; attribute dont_touch of G29881: signal is true;
	signal G29882: std_logic; attribute dont_touch of G29882: signal is true;
	signal G29883: std_logic; attribute dont_touch of G29883: signal is true;
	signal G29884: std_logic; attribute dont_touch of G29884: signal is true;
	signal G29885: std_logic; attribute dont_touch of G29885: signal is true;
	signal G29886: std_logic; attribute dont_touch of G29886: signal is true;
	signal G29887: std_logic; attribute dont_touch of G29887: signal is true;
	signal G29888: std_logic; attribute dont_touch of G29888: signal is true;
	signal G29889: std_logic; attribute dont_touch of G29889: signal is true;
	signal G29890: std_logic; attribute dont_touch of G29890: signal is true;
	signal G29891: std_logic; attribute dont_touch of G29891: signal is true;
	signal G29892: std_logic; attribute dont_touch of G29892: signal is true;
	signal G29893: std_logic; attribute dont_touch of G29893: signal is true;
	signal G29894: std_logic; attribute dont_touch of G29894: signal is true;
	signal G29895: std_logic; attribute dont_touch of G29895: signal is true;
	signal G29896: std_logic; attribute dont_touch of G29896: signal is true;
	signal G29897: std_logic; attribute dont_touch of G29897: signal is true;
	signal G29898: std_logic; attribute dont_touch of G29898: signal is true;
	signal G29899: std_logic; attribute dont_touch of G29899: signal is true;
	signal G29900: std_logic; attribute dont_touch of G29900: signal is true;
	signal G29901: std_logic; attribute dont_touch of G29901: signal is true;
	signal G29902: std_logic; attribute dont_touch of G29902: signal is true;
	signal G29903: std_logic; attribute dont_touch of G29903: signal is true;
	signal G29904: std_logic; attribute dont_touch of G29904: signal is true;
	signal G29905: std_logic; attribute dont_touch of G29905: signal is true;
	signal G29906: std_logic; attribute dont_touch of G29906: signal is true;
	signal G29907: std_logic; attribute dont_touch of G29907: signal is true;
	signal G29908: std_logic; attribute dont_touch of G29908: signal is true;
	signal G29909: std_logic; attribute dont_touch of G29909: signal is true;
	signal G29910: std_logic; attribute dont_touch of G29910: signal is true;
	signal G29911: std_logic; attribute dont_touch of G29911: signal is true;
	signal G29912: std_logic; attribute dont_touch of G29912: signal is true;
	signal G29913: std_logic; attribute dont_touch of G29913: signal is true;
	signal G29914: std_logic; attribute dont_touch of G29914: signal is true;
	signal G29915: std_logic; attribute dont_touch of G29915: signal is true;
	signal G29916: std_logic; attribute dont_touch of G29916: signal is true;
	signal G29920: std_logic; attribute dont_touch of G29920: signal is true;
	signal G29921: std_logic; attribute dont_touch of G29921: signal is true;
	signal G29922: std_logic; attribute dont_touch of G29922: signal is true;
	signal G29923: std_logic; attribute dont_touch of G29923: signal is true;
	signal G29924: std_logic; attribute dont_touch of G29924: signal is true;
	signal G29925: std_logic; attribute dont_touch of G29925: signal is true;
	signal G29926: std_logic; attribute dont_touch of G29926: signal is true;
	signal G29927: std_logic; attribute dont_touch of G29927: signal is true;
	signal G29928: std_logic; attribute dont_touch of G29928: signal is true;
	signal G29929: std_logic; attribute dont_touch of G29929: signal is true;
	signal G29930: std_logic; attribute dont_touch of G29930: signal is true;
	signal G29933: std_logic; attribute dont_touch of G29933: signal is true;
	signal G29937: std_logic; attribute dont_touch of G29937: signal is true;
	signal G29938: std_logic; attribute dont_touch of G29938: signal is true;
	signal G29939: std_logic; attribute dont_touch of G29939: signal is true;
	signal G29940: std_logic; attribute dont_touch of G29940: signal is true;
	signal G29941: std_logic; attribute dont_touch of G29941: signal is true;
	signal G29942: std_logic; attribute dont_touch of G29942: signal is true;
	signal G29943: std_logic; attribute dont_touch of G29943: signal is true;
	signal G29944: std_logic; attribute dont_touch of G29944: signal is true;
	signal G29945: std_logic; attribute dont_touch of G29945: signal is true;
	signal G29948: std_logic; attribute dont_touch of G29948: signal is true;
	signal G29949: std_logic; attribute dont_touch of G29949: signal is true;
	signal G29950: std_logic; attribute dont_touch of G29950: signal is true;
	signal G29951: std_logic; attribute dont_touch of G29951: signal is true;
	signal G29952: std_logic; attribute dont_touch of G29952: signal is true;
	signal G29953: std_logic; attribute dont_touch of G29953: signal is true;
	signal G29954: std_logic; attribute dont_touch of G29954: signal is true;
	signal G29955: std_logic; attribute dont_touch of G29955: signal is true;
	signal G29956: std_logic; attribute dont_touch of G29956: signal is true;
	signal G29959: std_logic; attribute dont_touch of G29959: signal is true;
	signal G29960: std_logic; attribute dont_touch of G29960: signal is true;
	signal G29961: std_logic; attribute dont_touch of G29961: signal is true;
	signal G29962: std_logic; attribute dont_touch of G29962: signal is true;
	signal G29963: std_logic; attribute dont_touch of G29963: signal is true;
	signal G29964: std_logic; attribute dont_touch of G29964: signal is true;
	signal G29965: std_logic; attribute dont_touch of G29965: signal is true;
	signal G29966: std_logic; attribute dont_touch of G29966: signal is true;
	signal G29967: std_logic; attribute dont_touch of G29967: signal is true;
	signal G29968: std_logic; attribute dont_touch of G29968: signal is true;
	signal G29969: std_logic; attribute dont_touch of G29969: signal is true;
	signal G29970: std_logic; attribute dont_touch of G29970: signal is true;
	signal G29973: std_logic; attribute dont_touch of G29973: signal is true;
	signal G29974: std_logic; attribute dont_touch of G29974: signal is true;
	signal G29975: std_logic; attribute dont_touch of G29975: signal is true;
	signal G29976: std_logic; attribute dont_touch of G29976: signal is true;
	signal G29977: std_logic; attribute dont_touch of G29977: signal is true;
	signal G29978: std_logic; attribute dont_touch of G29978: signal is true;
	signal G29979: std_logic; attribute dont_touch of G29979: signal is true;
	signal G29980: std_logic; attribute dont_touch of G29980: signal is true;
	signal G29981: std_logic; attribute dont_touch of G29981: signal is true;
	signal G29982: std_logic; attribute dont_touch of G29982: signal is true;
	signal G29983: std_logic; attribute dont_touch of G29983: signal is true;
	signal G29984: std_logic; attribute dont_touch of G29984: signal is true;
	signal G29985: std_logic; attribute dont_touch of G29985: signal is true;
	signal G29986: std_logic; attribute dont_touch of G29986: signal is true;
	signal G29987: std_logic; attribute dont_touch of G29987: signal is true;
	signal G29988: std_logic; attribute dont_touch of G29988: signal is true;
	signal G29989: std_logic; attribute dont_touch of G29989: signal is true;
	signal G29990: std_logic; attribute dont_touch of G29990: signal is true;
	signal G29991: std_logic; attribute dont_touch of G29991: signal is true;
	signal G29992: std_logic; attribute dont_touch of G29992: signal is true;
	signal G29993: std_logic; attribute dont_touch of G29993: signal is true;
	signal G29994: std_logic; attribute dont_touch of G29994: signal is true;
	signal G29995: std_logic; attribute dont_touch of G29995: signal is true;
	signal G29996: std_logic; attribute dont_touch of G29996: signal is true;
	signal G29997: std_logic; attribute dont_touch of G29997: signal is true;
	signal G29998: std_logic; attribute dont_touch of G29998: signal is true;
	signal G29999: std_logic; attribute dont_touch of G29999: signal is true;
	signal G30000: std_logic; attribute dont_touch of G30000: signal is true;
	signal G30001: std_logic; attribute dont_touch of G30001: signal is true;
	signal G30002: std_logic; attribute dont_touch of G30002: signal is true;
	signal G30003: std_logic; attribute dont_touch of G30003: signal is true;
	signal G30004: std_logic; attribute dont_touch of G30004: signal is true;
	signal G30005: std_logic; attribute dont_touch of G30005: signal is true;
	signal G30006: std_logic; attribute dont_touch of G30006: signal is true;
	signal G30007: std_logic; attribute dont_touch of G30007: signal is true;
	signal G30008: std_logic; attribute dont_touch of G30008: signal is true;
	signal G30009: std_logic; attribute dont_touch of G30009: signal is true;
	signal G30010: std_logic; attribute dont_touch of G30010: signal is true;
	signal G30011: std_logic; attribute dont_touch of G30011: signal is true;
	signal G30012: std_logic; attribute dont_touch of G30012: signal is true;
	signal G30015: std_logic; attribute dont_touch of G30015: signal is true;
	signal G30016: std_logic; attribute dont_touch of G30016: signal is true;
	signal G30017: std_logic; attribute dont_touch of G30017: signal is true;
	signal G30018: std_logic; attribute dont_touch of G30018: signal is true;
	signal G30019: std_logic; attribute dont_touch of G30019: signal is true;
	signal G30020: std_logic; attribute dont_touch of G30020: signal is true;
	signal G30021: std_logic; attribute dont_touch of G30021: signal is true;
	signal G30022: std_logic; attribute dont_touch of G30022: signal is true;
	signal G30023: std_logic; attribute dont_touch of G30023: signal is true;
	signal G30024: std_logic; attribute dont_touch of G30024: signal is true;
	signal G30025: std_logic; attribute dont_touch of G30025: signal is true;
	signal G30026: std_logic; attribute dont_touch of G30026: signal is true;
	signal G30027: std_logic; attribute dont_touch of G30027: signal is true;
	signal G30028: std_logic; attribute dont_touch of G30028: signal is true;
	signal G30029: std_logic; attribute dont_touch of G30029: signal is true;
	signal G30030: std_logic; attribute dont_touch of G30030: signal is true;
	signal G30031: std_logic; attribute dont_touch of G30031: signal is true;
	signal G30032: std_logic; attribute dont_touch of G30032: signal is true;
	signal G30033: std_logic; attribute dont_touch of G30033: signal is true;
	signal G30034: std_logic; attribute dont_touch of G30034: signal is true;
	signal G30035: std_logic; attribute dont_touch of G30035: signal is true;
	signal G30036: std_logic; attribute dont_touch of G30036: signal is true;
	signal G30037: std_logic; attribute dont_touch of G30037: signal is true;
	signal G30038: std_logic; attribute dont_touch of G30038: signal is true;
	signal G30039: std_logic; attribute dont_touch of G30039: signal is true;
	signal G30040: std_logic; attribute dont_touch of G30040: signal is true;
	signal G30041: std_logic; attribute dont_touch of G30041: signal is true;
	signal G30042: std_logic; attribute dont_touch of G30042: signal is true;
	signal G30043: std_logic; attribute dont_touch of G30043: signal is true;
	signal G30044: std_logic; attribute dont_touch of G30044: signal is true;
	signal G30045: std_logic; attribute dont_touch of G30045: signal is true;
	signal G30046: std_logic; attribute dont_touch of G30046: signal is true;
	signal G30047: std_logic; attribute dont_touch of G30047: signal is true;
	signal G30048: std_logic; attribute dont_touch of G30048: signal is true;
	signal G30049: std_logic; attribute dont_touch of G30049: signal is true;
	signal G30050: std_logic; attribute dont_touch of G30050: signal is true;
	signal G30051: std_logic; attribute dont_touch of G30051: signal is true;
	signal G30052: std_logic; attribute dont_touch of G30052: signal is true;
	signal G30053: std_logic; attribute dont_touch of G30053: signal is true;
	signal G30054: std_logic; attribute dont_touch of G30054: signal is true;
	signal G30055: std_logic; attribute dont_touch of G30055: signal is true;
	signal G30056: std_logic; attribute dont_touch of G30056: signal is true;
	signal G30057: std_logic; attribute dont_touch of G30057: signal is true;
	signal G30058: std_logic; attribute dont_touch of G30058: signal is true;
	signal G30059: std_logic; attribute dont_touch of G30059: signal is true;
	signal G30060: std_logic; attribute dont_touch of G30060: signal is true;
	signal G30061: std_logic; attribute dont_touch of G30061: signal is true;
	signal G30062: std_logic; attribute dont_touch of G30062: signal is true;
	signal G30063: std_logic; attribute dont_touch of G30063: signal is true;
	signal G30064: std_logic; attribute dont_touch of G30064: signal is true;
	signal G30065: std_logic; attribute dont_touch of G30065: signal is true;
	signal G30066: std_logic; attribute dont_touch of G30066: signal is true;
	signal G30067: std_logic; attribute dont_touch of G30067: signal is true;
	signal G30068: std_logic; attribute dont_touch of G30068: signal is true;
	signal G30069: std_logic; attribute dont_touch of G30069: signal is true;
	signal G30070: std_logic; attribute dont_touch of G30070: signal is true;
	signal G30071: std_logic; attribute dont_touch of G30071: signal is true;
	signal G30072: std_logic; attribute dont_touch of G30072: signal is true;
	signal G30073: std_logic; attribute dont_touch of G30073: signal is true;
	signal G30074: std_logic; attribute dont_touch of G30074: signal is true;
	signal G30075: std_logic; attribute dont_touch of G30075: signal is true;
	signal G30076: std_logic; attribute dont_touch of G30076: signal is true;
	signal G30077: std_logic; attribute dont_touch of G30077: signal is true;
	signal G30078: std_logic; attribute dont_touch of G30078: signal is true;
	signal G30079: std_logic; attribute dont_touch of G30079: signal is true;
	signal G30080: std_logic; attribute dont_touch of G30080: signal is true;
	signal G30081: std_logic; attribute dont_touch of G30081: signal is true;
	signal G30082: std_logic; attribute dont_touch of G30082: signal is true;
	signal G30083: std_logic; attribute dont_touch of G30083: signal is true;
	signal G30084: std_logic; attribute dont_touch of G30084: signal is true;
	signal G30085: std_logic; attribute dont_touch of G30085: signal is true;
	signal G30086: std_logic; attribute dont_touch of G30086: signal is true;
	signal G30087: std_logic; attribute dont_touch of G30087: signal is true;
	signal G30088: std_logic; attribute dont_touch of G30088: signal is true;
	signal G30089: std_logic; attribute dont_touch of G30089: signal is true;
	signal G30090: std_logic; attribute dont_touch of G30090: signal is true;
	signal G30091: std_logic; attribute dont_touch of G30091: signal is true;
	signal G30092: std_logic; attribute dont_touch of G30092: signal is true;
	signal G30093: std_logic; attribute dont_touch of G30093: signal is true;
	signal G30094: std_logic; attribute dont_touch of G30094: signal is true;
	signal G30095: std_logic; attribute dont_touch of G30095: signal is true;
	signal G30096: std_logic; attribute dont_touch of G30096: signal is true;
	signal G30097: std_logic; attribute dont_touch of G30097: signal is true;
	signal G30098: std_logic; attribute dont_touch of G30098: signal is true;
	signal G30099: std_logic; attribute dont_touch of G30099: signal is true;
	signal G30100: std_logic; attribute dont_touch of G30100: signal is true;
	signal G30101: std_logic; attribute dont_touch of G30101: signal is true;
	signal G30102: std_logic; attribute dont_touch of G30102: signal is true;
	signal G30103: std_logic; attribute dont_touch of G30103: signal is true;
	signal G30104: std_logic; attribute dont_touch of G30104: signal is true;
	signal G30105: std_logic; attribute dont_touch of G30105: signal is true;
	signal G30106: std_logic; attribute dont_touch of G30106: signal is true;
	signal G30107: std_logic; attribute dont_touch of G30107: signal is true;
	signal G30108: std_logic; attribute dont_touch of G30108: signal is true;
	signal G30109: std_logic; attribute dont_touch of G30109: signal is true;
	signal G30110: std_logic; attribute dont_touch of G30110: signal is true;
	signal G30111: std_logic; attribute dont_touch of G30111: signal is true;
	signal G30112: std_logic; attribute dont_touch of G30112: signal is true;
	signal G30113: std_logic; attribute dont_touch of G30113: signal is true;
	signal G30114: std_logic; attribute dont_touch of G30114: signal is true;
	signal G30115: std_logic; attribute dont_touch of G30115: signal is true;
	signal G30116: std_logic; attribute dont_touch of G30116: signal is true;
	signal G30117: std_logic; attribute dont_touch of G30117: signal is true;
	signal G30118: std_logic; attribute dont_touch of G30118: signal is true;
	signal G30119: std_logic; attribute dont_touch of G30119: signal is true;
	signal G30120: std_logic; attribute dont_touch of G30120: signal is true;
	signal G30121: std_logic; attribute dont_touch of G30121: signal is true;
	signal G30122: std_logic; attribute dont_touch of G30122: signal is true;
	signal G30123: std_logic; attribute dont_touch of G30123: signal is true;
	signal G30124: std_logic; attribute dont_touch of G30124: signal is true;
	signal G30125: std_logic; attribute dont_touch of G30125: signal is true;
	signal G30126: std_logic; attribute dont_touch of G30126: signal is true;
	signal G30127: std_logic; attribute dont_touch of G30127: signal is true;
	signal G30128: std_logic; attribute dont_touch of G30128: signal is true;
	signal G30129: std_logic; attribute dont_touch of G30129: signal is true;
	signal G30130: std_logic; attribute dont_touch of G30130: signal is true;
	signal G30131: std_logic; attribute dont_touch of G30131: signal is true;
	signal G30132: std_logic; attribute dont_touch of G30132: signal is true;
	signal G30133: std_logic; attribute dont_touch of G30133: signal is true;
	signal G30134: std_logic; attribute dont_touch of G30134: signal is true;
	signal G30135: std_logic; attribute dont_touch of G30135: signal is true;
	signal G30136: std_logic; attribute dont_touch of G30136: signal is true;
	signal G30137: std_logic; attribute dont_touch of G30137: signal is true;
	signal G30138: std_logic; attribute dont_touch of G30138: signal is true;
	signal G30139: std_logic; attribute dont_touch of G30139: signal is true;
	signal G30140: std_logic; attribute dont_touch of G30140: signal is true;
	signal G30141: std_logic; attribute dont_touch of G30141: signal is true;
	signal G30142: std_logic; attribute dont_touch of G30142: signal is true;
	signal G30143: std_logic; attribute dont_touch of G30143: signal is true;
	signal G30144: std_logic; attribute dont_touch of G30144: signal is true;
	signal G30145: std_logic; attribute dont_touch of G30145: signal is true;
	signal G30146: std_logic; attribute dont_touch of G30146: signal is true;
	signal G30147: std_logic; attribute dont_touch of G30147: signal is true;
	signal G30148: std_logic; attribute dont_touch of G30148: signal is true;
	signal G30149: std_logic; attribute dont_touch of G30149: signal is true;
	signal G30150: std_logic; attribute dont_touch of G30150: signal is true;
	signal G30151: std_logic; attribute dont_touch of G30151: signal is true;
	signal G30152: std_logic; attribute dont_touch of G30152: signal is true;
	signal G30153: std_logic; attribute dont_touch of G30153: signal is true;
	signal G30154: std_logic; attribute dont_touch of G30154: signal is true;
	signal G30155: std_logic; attribute dont_touch of G30155: signal is true;
	signal G30156: std_logic; attribute dont_touch of G30156: signal is true;
	signal G30157: std_logic; attribute dont_touch of G30157: signal is true;
	signal G30158: std_logic; attribute dont_touch of G30158: signal is true;
	signal G30159: std_logic; attribute dont_touch of G30159: signal is true;
	signal G30160: std_logic; attribute dont_touch of G30160: signal is true;
	signal G30161: std_logic; attribute dont_touch of G30161: signal is true;
	signal G30162: std_logic; attribute dont_touch of G30162: signal is true;
	signal G30163: std_logic; attribute dont_touch of G30163: signal is true;
	signal G30164: std_logic; attribute dont_touch of G30164: signal is true;
	signal G30165: std_logic; attribute dont_touch of G30165: signal is true;
	signal G30166: std_logic; attribute dont_touch of G30166: signal is true;
	signal G30167: std_logic; attribute dont_touch of G30167: signal is true;
	signal G30168: std_logic; attribute dont_touch of G30168: signal is true;
	signal G30169: std_logic; attribute dont_touch of G30169: signal is true;
	signal G30170: std_logic; attribute dont_touch of G30170: signal is true;
	signal G30171: std_logic; attribute dont_touch of G30171: signal is true;
	signal G30172: std_logic; attribute dont_touch of G30172: signal is true;
	signal G30173: std_logic; attribute dont_touch of G30173: signal is true;
	signal G30174: std_logic; attribute dont_touch of G30174: signal is true;
	signal G30175: std_logic; attribute dont_touch of G30175: signal is true;
	signal G30176: std_logic; attribute dont_touch of G30176: signal is true;
	signal G30177: std_logic; attribute dont_touch of G30177: signal is true;
	signal G30178: std_logic; attribute dont_touch of G30178: signal is true;
	signal G30179: std_logic; attribute dont_touch of G30179: signal is true;
	signal G30180: std_logic; attribute dont_touch of G30180: signal is true;
	signal G30181: std_logic; attribute dont_touch of G30181: signal is true;
	signal G30182: std_logic; attribute dont_touch of G30182: signal is true;
	signal G30183: std_logic; attribute dont_touch of G30183: signal is true;
	signal G30184: std_logic; attribute dont_touch of G30184: signal is true;
	signal G30185: std_logic; attribute dont_touch of G30185: signal is true;
	signal G30186: std_logic; attribute dont_touch of G30186: signal is true;
	signal G30187: std_logic; attribute dont_touch of G30187: signal is true;
	signal G30188: std_logic; attribute dont_touch of G30188: signal is true;
	signal G30189: std_logic; attribute dont_touch of G30189: signal is true;
	signal G30190: std_logic; attribute dont_touch of G30190: signal is true;
	signal G30191: std_logic; attribute dont_touch of G30191: signal is true;
	signal G30192: std_logic; attribute dont_touch of G30192: signal is true;
	signal G30193: std_logic; attribute dont_touch of G30193: signal is true;
	signal G30194: std_logic; attribute dont_touch of G30194: signal is true;
	signal G30195: std_logic; attribute dont_touch of G30195: signal is true;
	signal G30196: std_logic; attribute dont_touch of G30196: signal is true;
	signal G30197: std_logic; attribute dont_touch of G30197: signal is true;
	signal G30198: std_logic; attribute dont_touch of G30198: signal is true;
	signal G30199: std_logic; attribute dont_touch of G30199: signal is true;
	signal G30200: std_logic; attribute dont_touch of G30200: signal is true;
	signal G30201: std_logic; attribute dont_touch of G30201: signal is true;
	signal G30202: std_logic; attribute dont_touch of G30202: signal is true;
	signal G30203: std_logic; attribute dont_touch of G30203: signal is true;
	signal G30204: std_logic; attribute dont_touch of G30204: signal is true;
	signal G30205: std_logic; attribute dont_touch of G30205: signal is true;
	signal G30206: std_logic; attribute dont_touch of G30206: signal is true;
	signal G30207: std_logic; attribute dont_touch of G30207: signal is true;
	signal G30208: std_logic; attribute dont_touch of G30208: signal is true;
	signal G30209: std_logic; attribute dont_touch of G30209: signal is true;
	signal G30210: std_logic; attribute dont_touch of G30210: signal is true;
	signal G30211: std_logic; attribute dont_touch of G30211: signal is true;
	signal G30212: std_logic; attribute dont_touch of G30212: signal is true;
	signal G30213: std_logic; attribute dont_touch of G30213: signal is true;
	signal G30214: std_logic; attribute dont_touch of G30214: signal is true;
	signal G30215: std_logic; attribute dont_touch of G30215: signal is true;
	signal G30216: std_logic; attribute dont_touch of G30216: signal is true;
	signal G30217: std_logic; attribute dont_touch of G30217: signal is true;
	signal G30218: std_logic; attribute dont_touch of G30218: signal is true;
	signal G30219: std_logic; attribute dont_touch of G30219: signal is true;
	signal G30220: std_logic; attribute dont_touch of G30220: signal is true;
	signal G30221: std_logic; attribute dont_touch of G30221: signal is true;
	signal G30222: std_logic; attribute dont_touch of G30222: signal is true;
	signal G30223: std_logic; attribute dont_touch of G30223: signal is true;
	signal G30224: std_logic; attribute dont_touch of G30224: signal is true;
	signal G30225: std_logic; attribute dont_touch of G30225: signal is true;
	signal G30226: std_logic; attribute dont_touch of G30226: signal is true;
	signal G30227: std_logic; attribute dont_touch of G30227: signal is true;
	signal G30228: std_logic; attribute dont_touch of G30228: signal is true;
	signal G30229: std_logic; attribute dont_touch of G30229: signal is true;
	signal G30230: std_logic; attribute dont_touch of G30230: signal is true;
	signal G30231: std_logic; attribute dont_touch of G30231: signal is true;
	signal G30232: std_logic; attribute dont_touch of G30232: signal is true;
	signal G30233: std_logic; attribute dont_touch of G30233: signal is true;
	signal G30234: std_logic; attribute dont_touch of G30234: signal is true;
	signal G30235: std_logic; attribute dont_touch of G30235: signal is true;
	signal G30236: std_logic; attribute dont_touch of G30236: signal is true;
	signal G30237: std_logic; attribute dont_touch of G30237: signal is true;
	signal G30238: std_logic; attribute dont_touch of G30238: signal is true;
	signal G30239: std_logic; attribute dont_touch of G30239: signal is true;
	signal G30240: std_logic; attribute dont_touch of G30240: signal is true;
	signal G30241: std_logic; attribute dont_touch of G30241: signal is true;
	signal G30242: std_logic; attribute dont_touch of G30242: signal is true;
	signal G30243: std_logic; attribute dont_touch of G30243: signal is true;
	signal G30244: std_logic; attribute dont_touch of G30244: signal is true;
	signal G30245: std_logic; attribute dont_touch of G30245: signal is true;
	signal G30246: std_logic; attribute dont_touch of G30246: signal is true;
	signal G30247: std_logic; attribute dont_touch of G30247: signal is true;
	signal G30248: std_logic; attribute dont_touch of G30248: signal is true;
	signal G30249: std_logic; attribute dont_touch of G30249: signal is true;
	signal G30250: std_logic; attribute dont_touch of G30250: signal is true;
	signal G30251: std_logic; attribute dont_touch of G30251: signal is true;
	signal G30252: std_logic; attribute dont_touch of G30252: signal is true;
	signal G30253: std_logic; attribute dont_touch of G30253: signal is true;
	signal G30254: std_logic; attribute dont_touch of G30254: signal is true;
	signal G30255: std_logic; attribute dont_touch of G30255: signal is true;
	signal G30256: std_logic; attribute dont_touch of G30256: signal is true;
	signal G30257: std_logic; attribute dont_touch of G30257: signal is true;
	signal G30258: std_logic; attribute dont_touch of G30258: signal is true;
	signal G30259: std_logic; attribute dont_touch of G30259: signal is true;
	signal G30260: std_logic; attribute dont_touch of G30260: signal is true;
	signal G30261: std_logic; attribute dont_touch of G30261: signal is true;
	signal G30262: std_logic; attribute dont_touch of G30262: signal is true;
	signal G30263: std_logic; attribute dont_touch of G30263: signal is true;
	signal G30264: std_logic; attribute dont_touch of G30264: signal is true;
	signal G30265: std_logic; attribute dont_touch of G30265: signal is true;
	signal G30266: std_logic; attribute dont_touch of G30266: signal is true;
	signal G30267: std_logic; attribute dont_touch of G30267: signal is true;
	signal G30268: std_logic; attribute dont_touch of G30268: signal is true;
	signal G30269: std_logic; attribute dont_touch of G30269: signal is true;
	signal G30270: std_logic; attribute dont_touch of G30270: signal is true;
	signal G30271: std_logic; attribute dont_touch of G30271: signal is true;
	signal G30272: std_logic; attribute dont_touch of G30272: signal is true;
	signal G30273: std_logic; attribute dont_touch of G30273: signal is true;
	signal G30274: std_logic; attribute dont_touch of G30274: signal is true;
	signal G30275: std_logic; attribute dont_touch of G30275: signal is true;
	signal G30276: std_logic; attribute dont_touch of G30276: signal is true;
	signal G30277: std_logic; attribute dont_touch of G30277: signal is true;
	signal G30278: std_logic; attribute dont_touch of G30278: signal is true;
	signal G30279: std_logic; attribute dont_touch of G30279: signal is true;
	signal G30280: std_logic; attribute dont_touch of G30280: signal is true;
	signal G30281: std_logic; attribute dont_touch of G30281: signal is true;
	signal G30282: std_logic; attribute dont_touch of G30282: signal is true;
	signal G30283: std_logic; attribute dont_touch of G30283: signal is true;
	signal G30284: std_logic; attribute dont_touch of G30284: signal is true;
	signal G30285: std_logic; attribute dont_touch of G30285: signal is true;
	signal G30286: std_logic; attribute dont_touch of G30286: signal is true;
	signal G30287: std_logic; attribute dont_touch of G30287: signal is true;
	signal G30288: std_logic; attribute dont_touch of G30288: signal is true;
	signal G30289: std_logic; attribute dont_touch of G30289: signal is true;
	signal G30290: std_logic; attribute dont_touch of G30290: signal is true;
	signal G30291: std_logic; attribute dont_touch of G30291: signal is true;
	signal G30292: std_logic; attribute dont_touch of G30292: signal is true;
	signal G30293: std_logic; attribute dont_touch of G30293: signal is true;
	signal G30294: std_logic; attribute dont_touch of G30294: signal is true;
	signal G30295: std_logic; attribute dont_touch of G30295: signal is true;
	signal G30296: std_logic; attribute dont_touch of G30296: signal is true;
	signal G30297: std_logic; attribute dont_touch of G30297: signal is true;
	signal G30298: std_logic; attribute dont_touch of G30298: signal is true;
	signal G30299: std_logic; attribute dont_touch of G30299: signal is true;
	signal G30300: std_logic; attribute dont_touch of G30300: signal is true;
	signal G30301: std_logic; attribute dont_touch of G30301: signal is true;
	signal G30302: std_logic; attribute dont_touch of G30302: signal is true;
	signal G30303: std_logic; attribute dont_touch of G30303: signal is true;
	signal G30304: std_logic; attribute dont_touch of G30304: signal is true;
	signal G30305: std_logic; attribute dont_touch of G30305: signal is true;
	signal G30306: std_logic; attribute dont_touch of G30306: signal is true;
	signal G30307: std_logic; attribute dont_touch of G30307: signal is true;
	signal G30308: std_logic; attribute dont_touch of G30308: signal is true;
	signal G30309: std_logic; attribute dont_touch of G30309: signal is true;
	signal G30310: std_logic; attribute dont_touch of G30310: signal is true;
	signal G30311: std_logic; attribute dont_touch of G30311: signal is true;
	signal G30312: std_logic; attribute dont_touch of G30312: signal is true;
	signal G30313: std_logic; attribute dont_touch of G30313: signal is true;
	signal G30314: std_logic; attribute dont_touch of G30314: signal is true;
	signal G30315: std_logic; attribute dont_touch of G30315: signal is true;
	signal G30316: std_logic; attribute dont_touch of G30316: signal is true;
	signal G30317: std_logic; attribute dont_touch of G30317: signal is true;
	signal G30318: std_logic; attribute dont_touch of G30318: signal is true;
	signal G30321: std_logic; attribute dont_touch of G30321: signal is true;
	signal G30322: std_logic; attribute dont_touch of G30322: signal is true;
	signal G30325: std_logic; attribute dont_touch of G30325: signal is true;
	signal G30326: std_logic; attribute dont_touch of G30326: signal is true;
	signal G30328: std_logic; attribute dont_touch of G30328: signal is true;
	signal G30333: std_logic; attribute dont_touch of G30333: signal is true;
	signal G30334: std_logic; attribute dont_touch of G30334: signal is true;
	signal G30335: std_logic; attribute dont_touch of G30335: signal is true;
	signal G30336: std_logic; attribute dont_touch of G30336: signal is true;
	signal G30337: std_logic; attribute dont_touch of G30337: signal is true;
	signal G30338: std_logic; attribute dont_touch of G30338: signal is true;
	signal G30339: std_logic; attribute dont_touch of G30339: signal is true;
	signal G30340: std_logic; attribute dont_touch of G30340: signal is true;
	signal G30341: std_logic; attribute dont_touch of G30341: signal is true;
	signal G30342: std_logic; attribute dont_touch of G30342: signal is true;
	signal G30343: std_logic; attribute dont_touch of G30343: signal is true;
	signal G30344: std_logic; attribute dont_touch of G30344: signal is true;
	signal G30345: std_logic; attribute dont_touch of G30345: signal is true;
	signal G30346: std_logic; attribute dont_touch of G30346: signal is true;
	signal G30347: std_logic; attribute dont_touch of G30347: signal is true;
	signal G30348: std_logic; attribute dont_touch of G30348: signal is true;
	signal G30349: std_logic; attribute dont_touch of G30349: signal is true;
	signal G30350: std_logic; attribute dont_touch of G30350: signal is true;
	signal G30351: std_logic; attribute dont_touch of G30351: signal is true;
	signal G30352: std_logic; attribute dont_touch of G30352: signal is true;
	signal G30353: std_logic; attribute dont_touch of G30353: signal is true;
	signal G30354: std_logic; attribute dont_touch of G30354: signal is true;
	signal G30355: std_logic; attribute dont_touch of G30355: signal is true;
	signal G30356: std_logic; attribute dont_touch of G30356: signal is true;
	signal G30357: std_logic; attribute dont_touch of G30357: signal is true;
	signal G30358: std_logic; attribute dont_touch of G30358: signal is true;
	signal G30359: std_logic; attribute dont_touch of G30359: signal is true;
	signal G30360: std_logic; attribute dont_touch of G30360: signal is true;
	signal G30361: std_logic; attribute dont_touch of G30361: signal is true;
	signal G30362: std_logic; attribute dont_touch of G30362: signal is true;
	signal G30363: std_logic; attribute dont_touch of G30363: signal is true;
	signal G30364: std_logic; attribute dont_touch of G30364: signal is true;
	signal G30365: std_logic; attribute dont_touch of G30365: signal is true;
	signal G30366: std_logic; attribute dont_touch of G30366: signal is true;
	signal G30367: std_logic; attribute dont_touch of G30367: signal is true;
	signal G30368: std_logic; attribute dont_touch of G30368: signal is true;
	signal G30369: std_logic; attribute dont_touch of G30369: signal is true;
	signal G30370: std_logic; attribute dont_touch of G30370: signal is true;
	signal G30371: std_logic; attribute dont_touch of G30371: signal is true;
	signal G30372: std_logic; attribute dont_touch of G30372: signal is true;
	signal G30373: std_logic; attribute dont_touch of G30373: signal is true;
	signal G30374: std_logic; attribute dont_touch of G30374: signal is true;
	signal G30375: std_logic; attribute dont_touch of G30375: signal is true;
	signal G30376: std_logic; attribute dont_touch of G30376: signal is true;
	signal G30377: std_logic; attribute dont_touch of G30377: signal is true;
	signal G30378: std_logic; attribute dont_touch of G30378: signal is true;
	signal G30379: std_logic; attribute dont_touch of G30379: signal is true;
	signal G30380: std_logic; attribute dont_touch of G30380: signal is true;
	signal G30381: std_logic; attribute dont_touch of G30381: signal is true;
	signal G30382: std_logic; attribute dont_touch of G30382: signal is true;
	signal G30383: std_logic; attribute dont_touch of G30383: signal is true;
	signal G30384: std_logic; attribute dont_touch of G30384: signal is true;
	signal G30385: std_logic; attribute dont_touch of G30385: signal is true;
	signal G30386: std_logic; attribute dont_touch of G30386: signal is true;
	signal G30387: std_logic; attribute dont_touch of G30387: signal is true;
	signal G30388: std_logic; attribute dont_touch of G30388: signal is true;
	signal G30389: std_logic; attribute dont_touch of G30389: signal is true;
	signal G30390: std_logic; attribute dont_touch of G30390: signal is true;
	signal G30391: std_logic; attribute dont_touch of G30391: signal is true;
	signal G30392: std_logic; attribute dont_touch of G30392: signal is true;
	signal G30393: std_logic; attribute dont_touch of G30393: signal is true;
	signal G30394: std_logic; attribute dont_touch of G30394: signal is true;
	signal G30395: std_logic; attribute dont_touch of G30395: signal is true;
	signal G30396: std_logic; attribute dont_touch of G30396: signal is true;
	signal G30397: std_logic; attribute dont_touch of G30397: signal is true;
	signal G30398: std_logic; attribute dont_touch of G30398: signal is true;
	signal G30399: std_logic; attribute dont_touch of G30399: signal is true;
	signal G30400: std_logic; attribute dont_touch of G30400: signal is true;
	signal G30401: std_logic; attribute dont_touch of G30401: signal is true;
	signal G30402: std_logic; attribute dont_touch of G30402: signal is true;
	signal G30403: std_logic; attribute dont_touch of G30403: signal is true;
	signal G30404: std_logic; attribute dont_touch of G30404: signal is true;
	signal G30405: std_logic; attribute dont_touch of G30405: signal is true;
	signal G30406: std_logic; attribute dont_touch of G30406: signal is true;
	signal G30407: std_logic; attribute dont_touch of G30407: signal is true;
	signal G30408: std_logic; attribute dont_touch of G30408: signal is true;
	signal G30409: std_logic; attribute dont_touch of G30409: signal is true;
	signal G30410: std_logic; attribute dont_touch of G30410: signal is true;
	signal G30411: std_logic; attribute dont_touch of G30411: signal is true;
	signal G30412: std_logic; attribute dont_touch of G30412: signal is true;
	signal G30413: std_logic; attribute dont_touch of G30413: signal is true;
	signal G30414: std_logic; attribute dont_touch of G30414: signal is true;
	signal G30415: std_logic; attribute dont_touch of G30415: signal is true;
	signal G30416: std_logic; attribute dont_touch of G30416: signal is true;
	signal G30417: std_logic; attribute dont_touch of G30417: signal is true;
	signal G30418: std_logic; attribute dont_touch of G30418: signal is true;
	signal G30419: std_logic; attribute dont_touch of G30419: signal is true;
	signal G30420: std_logic; attribute dont_touch of G30420: signal is true;
	signal G30421: std_logic; attribute dont_touch of G30421: signal is true;
	signal G30422: std_logic; attribute dont_touch of G30422: signal is true;
	signal G30423: std_logic; attribute dont_touch of G30423: signal is true;
	signal G30424: std_logic; attribute dont_touch of G30424: signal is true;
	signal G30425: std_logic; attribute dont_touch of G30425: signal is true;
	signal G30426: std_logic; attribute dont_touch of G30426: signal is true;
	signal G30427: std_logic; attribute dont_touch of G30427: signal is true;
	signal G30428: std_logic; attribute dont_touch of G30428: signal is true;
	signal G30429: std_logic; attribute dont_touch of G30429: signal is true;
	signal G30430: std_logic; attribute dont_touch of G30430: signal is true;
	signal G30431: std_logic; attribute dont_touch of G30431: signal is true;
	signal G30432: std_logic; attribute dont_touch of G30432: signal is true;
	signal G30433: std_logic; attribute dont_touch of G30433: signal is true;
	signal G30434: std_logic; attribute dont_touch of G30434: signal is true;
	signal G30435: std_logic; attribute dont_touch of G30435: signal is true;
	signal G30436: std_logic; attribute dont_touch of G30436: signal is true;
	signal G30437: std_logic; attribute dont_touch of G30437: signal is true;
	signal G30438: std_logic; attribute dont_touch of G30438: signal is true;
	signal G30439: std_logic; attribute dont_touch of G30439: signal is true;
	signal G30440: std_logic; attribute dont_touch of G30440: signal is true;
	signal G30441: std_logic; attribute dont_touch of G30441: signal is true;
	signal G30442: std_logic; attribute dont_touch of G30442: signal is true;
	signal G30443: std_logic; attribute dont_touch of G30443: signal is true;
	signal G30444: std_logic; attribute dont_touch of G30444: signal is true;
	signal G30445: std_logic; attribute dont_touch of G30445: signal is true;
	signal G30446: std_logic; attribute dont_touch of G30446: signal is true;
	signal G30447: std_logic; attribute dont_touch of G30447: signal is true;
	signal G30448: std_logic; attribute dont_touch of G30448: signal is true;
	signal G30449: std_logic; attribute dont_touch of G30449: signal is true;
	signal G30450: std_logic; attribute dont_touch of G30450: signal is true;
	signal G30451: std_logic; attribute dont_touch of G30451: signal is true;
	signal G30452: std_logic; attribute dont_touch of G30452: signal is true;
	signal G30453: std_logic; attribute dont_touch of G30453: signal is true;
	signal G30454: std_logic; attribute dont_touch of G30454: signal is true;
	signal G30455: std_logic; attribute dont_touch of G30455: signal is true;
	signal G30456: std_logic; attribute dont_touch of G30456: signal is true;
	signal G30457: std_logic; attribute dont_touch of G30457: signal is true;
	signal G30458: std_logic; attribute dont_touch of G30458: signal is true;
	signal G30459: std_logic; attribute dont_touch of G30459: signal is true;
	signal G30460: std_logic; attribute dont_touch of G30460: signal is true;
	signal G30461: std_logic; attribute dont_touch of G30461: signal is true;
	signal G30462: std_logic; attribute dont_touch of G30462: signal is true;
	signal G30463: std_logic; attribute dont_touch of G30463: signal is true;
	signal G30464: std_logic; attribute dont_touch of G30464: signal is true;
	signal G30465: std_logic; attribute dont_touch of G30465: signal is true;
	signal G30466: std_logic; attribute dont_touch of G30466: signal is true;
	signal G30467: std_logic; attribute dont_touch of G30467: signal is true;
	signal G30468: std_logic; attribute dont_touch of G30468: signal is true;
	signal G30469: std_logic; attribute dont_touch of G30469: signal is true;
	signal G30470: std_logic; attribute dont_touch of G30470: signal is true;
	signal G30471: std_logic; attribute dont_touch of G30471: signal is true;
	signal G30472: std_logic; attribute dont_touch of G30472: signal is true;
	signal G30473: std_logic; attribute dont_touch of G30473: signal is true;
	signal G30474: std_logic; attribute dont_touch of G30474: signal is true;
	signal G30475: std_logic; attribute dont_touch of G30475: signal is true;
	signal G30476: std_logic; attribute dont_touch of G30476: signal is true;
	signal G30477: std_logic; attribute dont_touch of G30477: signal is true;
	signal G30478: std_logic; attribute dont_touch of G30478: signal is true;
	signal G30479: std_logic; attribute dont_touch of G30479: signal is true;
	signal G30480: std_logic; attribute dont_touch of G30480: signal is true;
	signal G30481: std_logic; attribute dont_touch of G30481: signal is true;
	signal G30482: std_logic; attribute dont_touch of G30482: signal is true;
	signal G30483: std_logic; attribute dont_touch of G30483: signal is true;
	signal G30484: std_logic; attribute dont_touch of G30484: signal is true;
	signal G30485: std_logic; attribute dont_touch of G30485: signal is true;
	signal G30486: std_logic; attribute dont_touch of G30486: signal is true;
	signal G30487: std_logic; attribute dont_touch of G30487: signal is true;
	signal G30488: std_logic; attribute dont_touch of G30488: signal is true;
	signal G30489: std_logic; attribute dont_touch of G30489: signal is true;
	signal G30490: std_logic; attribute dont_touch of G30490: signal is true;
	signal G30491: std_logic; attribute dont_touch of G30491: signal is true;
	signal G30492: std_logic; attribute dont_touch of G30492: signal is true;
	signal G30493: std_logic; attribute dont_touch of G30493: signal is true;
	signal G30494: std_logic; attribute dont_touch of G30494: signal is true;
	signal G30495: std_logic; attribute dont_touch of G30495: signal is true;
	signal G30496: std_logic; attribute dont_touch of G30496: signal is true;
	signal G30497: std_logic; attribute dont_touch of G30497: signal is true;
	signal G30498: std_logic; attribute dont_touch of G30498: signal is true;
	signal G30499: std_logic; attribute dont_touch of G30499: signal is true;
	signal G30500: std_logic; attribute dont_touch of G30500: signal is true;
	signal G30501: std_logic; attribute dont_touch of G30501: signal is true;
	signal G30502: std_logic; attribute dont_touch of G30502: signal is true;
	signal G30503: std_logic; attribute dont_touch of G30503: signal is true;
	signal G30504: std_logic; attribute dont_touch of G30504: signal is true;
	signal G30505: std_logic; attribute dont_touch of G30505: signal is true;
	signal G30506: std_logic; attribute dont_touch of G30506: signal is true;
	signal G30507: std_logic; attribute dont_touch of G30507: signal is true;
	signal G30508: std_logic; attribute dont_touch of G30508: signal is true;
	signal G30509: std_logic; attribute dont_touch of G30509: signal is true;
	signal G30510: std_logic; attribute dont_touch of G30510: signal is true;
	signal G30511: std_logic; attribute dont_touch of G30511: signal is true;
	signal G30512: std_logic; attribute dont_touch of G30512: signal is true;
	signal G30513: std_logic; attribute dont_touch of G30513: signal is true;
	signal G30514: std_logic; attribute dont_touch of G30514: signal is true;
	signal G30515: std_logic; attribute dont_touch of G30515: signal is true;
	signal G30516: std_logic; attribute dont_touch of G30516: signal is true;
	signal G30517: std_logic; attribute dont_touch of G30517: signal is true;
	signal G30518: std_logic; attribute dont_touch of G30518: signal is true;
	signal G30519: std_logic; attribute dont_touch of G30519: signal is true;
	signal G30520: std_logic; attribute dont_touch of G30520: signal is true;
	signal G30521: std_logic; attribute dont_touch of G30521: signal is true;
	signal G30522: std_logic; attribute dont_touch of G30522: signal is true;
	signal G30523: std_logic; attribute dont_touch of G30523: signal is true;
	signal G30524: std_logic; attribute dont_touch of G30524: signal is true;
	signal G30525: std_logic; attribute dont_touch of G30525: signal is true;
	signal G30526: std_logic; attribute dont_touch of G30526: signal is true;
	signal G30527: std_logic; attribute dont_touch of G30527: signal is true;
	signal G30528: std_logic; attribute dont_touch of G30528: signal is true;
	signal G30529: std_logic; attribute dont_touch of G30529: signal is true;
	signal G30530: std_logic; attribute dont_touch of G30530: signal is true;
	signal G30531: std_logic; attribute dont_touch of G30531: signal is true;
	signal G30532: std_logic; attribute dont_touch of G30532: signal is true;
	signal G30533: std_logic; attribute dont_touch of G30533: signal is true;
	signal G30534: std_logic; attribute dont_touch of G30534: signal is true;
	signal G30535: std_logic; attribute dont_touch of G30535: signal is true;
	signal G30536: std_logic; attribute dont_touch of G30536: signal is true;
	signal G30537: std_logic; attribute dont_touch of G30537: signal is true;
	signal G30538: std_logic; attribute dont_touch of G30538: signal is true;
	signal G30539: std_logic; attribute dont_touch of G30539: signal is true;
	signal G30540: std_logic; attribute dont_touch of G30540: signal is true;
	signal G30541: std_logic; attribute dont_touch of G30541: signal is true;
	signal G30542: std_logic; attribute dont_touch of G30542: signal is true;
	signal G30543: std_logic; attribute dont_touch of G30543: signal is true;
	signal G30544: std_logic; attribute dont_touch of G30544: signal is true;
	signal G30545: std_logic; attribute dont_touch of G30545: signal is true;
	signal G30546: std_logic; attribute dont_touch of G30546: signal is true;
	signal G30547: std_logic; attribute dont_touch of G30547: signal is true;
	signal G30548: std_logic; attribute dont_touch of G30548: signal is true;
	signal G30549: std_logic; attribute dont_touch of G30549: signal is true;
	signal G30550: std_logic; attribute dont_touch of G30550: signal is true;
	signal G30551: std_logic; attribute dont_touch of G30551: signal is true;
	signal G30552: std_logic; attribute dont_touch of G30552: signal is true;
	signal G30553: std_logic; attribute dont_touch of G30553: signal is true;
	signal G30554: std_logic; attribute dont_touch of G30554: signal is true;
	signal G30555: std_logic; attribute dont_touch of G30555: signal is true;
	signal G30556: std_logic; attribute dont_touch of G30556: signal is true;
	signal G30557: std_logic; attribute dont_touch of G30557: signal is true;
	signal G30558: std_logic; attribute dont_touch of G30558: signal is true;
	signal G30559: std_logic; attribute dont_touch of G30559: signal is true;
	signal G30560: std_logic; attribute dont_touch of G30560: signal is true;
	signal G30561: std_logic; attribute dont_touch of G30561: signal is true;
	signal G30562: std_logic; attribute dont_touch of G30562: signal is true;
	signal G30563: std_logic; attribute dont_touch of G30563: signal is true;
	signal G30564: std_logic; attribute dont_touch of G30564: signal is true;
	signal G30565: std_logic; attribute dont_touch of G30565: signal is true;
	signal G30566: std_logic; attribute dont_touch of G30566: signal is true;
	signal G30567: std_logic; attribute dont_touch of G30567: signal is true;
	signal G30568: std_logic; attribute dont_touch of G30568: signal is true;
	signal G30569: std_logic; attribute dont_touch of G30569: signal is true;
	signal G30572: std_logic; attribute dont_touch of G30572: signal is true;
	signal G30573: std_logic; attribute dont_touch of G30573: signal is true;
	signal G30576: std_logic; attribute dont_touch of G30576: signal is true;
	signal G30577: std_logic; attribute dont_touch of G30577: signal is true;
	signal G30578: std_logic; attribute dont_touch of G30578: signal is true;
	signal G30579: std_logic; attribute dont_touch of G30579: signal is true;
	signal G30580: std_logic; attribute dont_touch of G30580: signal is true;
	signal G30583: std_logic; attribute dont_touch of G30583: signal is true;
	signal G30589: std_logic; attribute dont_touch of G30589: signal is true;
	signal G30590: std_logic; attribute dont_touch of G30590: signal is true;
	signal G30591: std_logic; attribute dont_touch of G30591: signal is true;
	signal G30592: std_logic; attribute dont_touch of G30592: signal is true;
	signal G30593: std_logic; attribute dont_touch of G30593: signal is true;
	signal G30594: std_logic; attribute dont_touch of G30594: signal is true;
	signal G30595: std_logic; attribute dont_touch of G30595: signal is true;
	signal G30596: std_logic; attribute dont_touch of G30596: signal is true;
	signal G30597: std_logic; attribute dont_touch of G30597: signal is true;
	signal G30598: std_logic; attribute dont_touch of G30598: signal is true;
	signal G30599: std_logic; attribute dont_touch of G30599: signal is true;
	signal G30600: std_logic; attribute dont_touch of G30600: signal is true;
	signal G30601: std_logic; attribute dont_touch of G30601: signal is true;
	signal G30604: std_logic; attribute dont_touch of G30604: signal is true;
	signal G30605: std_logic; attribute dont_touch of G30605: signal is true;
	signal G30606: std_logic; attribute dont_touch of G30606: signal is true;
	signal G30607: std_logic; attribute dont_touch of G30607: signal is true;
	signal G30608: std_logic; attribute dont_touch of G30608: signal is true;
	signal G30609: std_logic; attribute dont_touch of G30609: signal is true;
	signal G30610: std_logic; attribute dont_touch of G30610: signal is true;
	signal G30611: std_logic; attribute dont_touch of G30611: signal is true;
	signal G30612: std_logic; attribute dont_touch of G30612: signal is true;
	signal G30613: std_logic; attribute dont_touch of G30613: signal is true;
	signal G30614: std_logic; attribute dont_touch of G30614: signal is true;
	signal G30670: std_logic; attribute dont_touch of G30670: signal is true;
	signal G30671: std_logic; attribute dont_touch of G30671: signal is true;
	signal G30672: std_logic; attribute dont_touch of G30672: signal is true;
	signal G30673: std_logic; attribute dont_touch of G30673: signal is true;
	signal G30729: std_logic; attribute dont_touch of G30729: signal is true;
	signal G30730: std_logic; attribute dont_touch of G30730: signal is true;
	signal G30731: std_logic; attribute dont_touch of G30731: signal is true;
	signal G30732: std_logic; attribute dont_touch of G30732: signal is true;
	signal G30733: std_logic; attribute dont_touch of G30733: signal is true;
	signal G30734: std_logic; attribute dont_touch of G30734: signal is true;
	signal G30735: std_logic; attribute dont_touch of G30735: signal is true;
	signal G30824: std_logic; attribute dont_touch of G30824: signal is true;
	signal G30825: std_logic; attribute dont_touch of G30825: signal is true;
	signal G30914: std_logic; attribute dont_touch of G30914: signal is true;
	signal G30915: std_logic; attribute dont_touch of G30915: signal is true;
	signal G30916: std_logic; attribute dont_touch of G30916: signal is true;
	signal G30917: std_logic; attribute dont_touch of G30917: signal is true;
	signal G30918: std_logic; attribute dont_touch of G30918: signal is true;
	signal G30919: std_logic; attribute dont_touch of G30919: signal is true;
	signal G30920: std_logic; attribute dont_touch of G30920: signal is true;
	signal G30921: std_logic; attribute dont_touch of G30921: signal is true;
	signal G30922: std_logic; attribute dont_touch of G30922: signal is true;
	signal G30925: std_logic; attribute dont_touch of G30925: signal is true;
	signal G30926: std_logic; attribute dont_touch of G30926: signal is true;
	signal G30927: std_logic; attribute dont_touch of G30927: signal is true;
	signal G30928: std_logic; attribute dont_touch of G30928: signal is true;
	signal G30929: std_logic; attribute dont_touch of G30929: signal is true;
	signal G30930: std_logic; attribute dont_touch of G30930: signal is true;
	signal G30931: std_logic; attribute dont_touch of G30931: signal is true;
	signal G30934: std_logic; attribute dont_touch of G30934: signal is true;
	signal G30935: std_logic; attribute dont_touch of G30935: signal is true;
	signal G30936: std_logic; attribute dont_touch of G30936: signal is true;
	signal G30937: std_logic; attribute dont_touch of G30937: signal is true;
	signal G30982: std_logic; attribute dont_touch of G30982: signal is true;
	signal G30983: std_logic; attribute dont_touch of G30983: signal is true;
	signal G30984: std_logic; attribute dont_touch of G30984: signal is true;
	signal G30989: std_logic; attribute dont_touch of G30989: signal is true;
	signal G30990: std_logic; attribute dont_touch of G30990: signal is true;
	signal G30991: std_logic; attribute dont_touch of G30991: signal is true;
	signal G30996: std_logic; attribute dont_touch of G30996: signal is true;
	signal G30997: std_logic; attribute dont_touch of G30997: signal is true;
	signal G30998: std_logic; attribute dont_touch of G30998: signal is true;
	signal G30999: std_logic; attribute dont_touch of G30999: signal is true;
	signal G31000: std_logic; attribute dont_touch of G31000: signal is true;
	signal G31001: std_logic; attribute dont_touch of G31001: signal is true;
	signal G31002: std_logic; attribute dont_touch of G31002: signal is true;
	signal G31003: std_logic; attribute dont_touch of G31003: signal is true;
	signal G31007: std_logic; attribute dont_touch of G31007: signal is true;
	signal G31008: std_logic; attribute dont_touch of G31008: signal is true;
	signal G31009: std_logic; attribute dont_touch of G31009: signal is true;
	signal G31013: std_logic; attribute dont_touch of G31013: signal is true;
	signal G31014: std_logic; attribute dont_touch of G31014: signal is true;
	signal G31015: std_logic; attribute dont_touch of G31015: signal is true;
	signal G31016: std_logic; attribute dont_touch of G31016: signal is true;
	signal G31017: std_logic; attribute dont_touch of G31017: signal is true;
	signal G31018: std_logic; attribute dont_touch of G31018: signal is true;
	signal G31019: std_logic; attribute dont_touch of G31019: signal is true;
	signal G31020: std_logic; attribute dont_touch of G31020: signal is true;
	signal G31021: std_logic; attribute dont_touch of G31021: signal is true;
	signal G31066: std_logic; attribute dont_touch of G31066: signal is true;
	signal G31067: std_logic; attribute dont_touch of G31067: signal is true;
	signal G31068: std_logic; attribute dont_touch of G31068: signal is true;
	signal G31069: std_logic; attribute dont_touch of G31069: signal is true;
	signal G31070: std_logic; attribute dont_touch of G31070: signal is true;
	signal G31115: std_logic; attribute dont_touch of G31115: signal is true;
	signal G31116: std_logic; attribute dont_touch of G31116: signal is true;
	signal G31117: std_logic; attribute dont_touch of G31117: signal is true;
	signal G31118: std_logic; attribute dont_touch of G31118: signal is true;
	signal G31119: std_logic; attribute dont_touch of G31119: signal is true;
	signal G31120: std_logic; attribute dont_touch of G31120: signal is true;
	signal G31121: std_logic; attribute dont_touch of G31121: signal is true;
	signal G31122: std_logic; attribute dont_touch of G31122: signal is true;
	signal G31123: std_logic; attribute dont_touch of G31123: signal is true;
	signal G31124: std_logic; attribute dont_touch of G31124: signal is true;
	signal G31125: std_logic; attribute dont_touch of G31125: signal is true;
	signal G31126: std_logic; attribute dont_touch of G31126: signal is true;
	signal G31127: std_logic; attribute dont_touch of G31127: signal is true;
	signal G31128: std_logic; attribute dont_touch of G31128: signal is true;
	signal G31129: std_logic; attribute dont_touch of G31129: signal is true;
	signal G31130: std_logic; attribute dont_touch of G31130: signal is true;
	signal G31131: std_logic; attribute dont_touch of G31131: signal is true;
	signal G31132: std_logic; attribute dont_touch of G31132: signal is true;
	signal G31133: std_logic; attribute dont_touch of G31133: signal is true;
	signal G31134: std_logic; attribute dont_touch of G31134: signal is true;
	signal G31138: std_logic; attribute dont_touch of G31138: signal is true;
	signal G31139: std_logic; attribute dont_touch of G31139: signal is true;
	signal G31140: std_logic; attribute dont_touch of G31140: signal is true;
	signal G31141: std_logic; attribute dont_touch of G31141: signal is true;
	signal G31142: std_logic; attribute dont_touch of G31142: signal is true;
	signal G31143: std_logic; attribute dont_touch of G31143: signal is true;
	signal G31144: std_logic; attribute dont_touch of G31144: signal is true;
	signal G31145: std_logic; attribute dont_touch of G31145: signal is true;
	signal G31146: std_logic; attribute dont_touch of G31146: signal is true;
	signal G31147: std_logic; attribute dont_touch of G31147: signal is true;
	signal G31148: std_logic; attribute dont_touch of G31148: signal is true;
	signal G31149: std_logic; attribute dont_touch of G31149: signal is true;
	signal G31150: std_logic; attribute dont_touch of G31150: signal is true;
	signal G31151: std_logic; attribute dont_touch of G31151: signal is true;
	signal G31152: std_logic; attribute dont_touch of G31152: signal is true;
	signal G31153: std_logic; attribute dont_touch of G31153: signal is true;
	signal G31154: std_logic; attribute dont_touch of G31154: signal is true;
	signal G31166: std_logic; attribute dont_touch of G31166: signal is true;
	signal G31167: std_logic; attribute dont_touch of G31167: signal is true;
	signal G31168: std_logic; attribute dont_touch of G31168: signal is true;
	signal G31169: std_logic; attribute dont_touch of G31169: signal is true;
	signal G31170: std_logic; attribute dont_touch of G31170: signal is true;
	signal G31182: std_logic; attribute dont_touch of G31182: signal is true;
	signal G31183: std_logic; attribute dont_touch of G31183: signal is true;
	signal G31184: std_logic; attribute dont_touch of G31184: signal is true;
	signal G31185: std_logic; attribute dont_touch of G31185: signal is true;
	signal G31186: std_logic; attribute dont_touch of G31186: signal is true;
	signal G31187: std_logic; attribute dont_touch of G31187: signal is true;
	signal G31188: std_logic; attribute dont_touch of G31188: signal is true;
	signal G31189: std_logic; attribute dont_touch of G31189: signal is true;
	signal G31194: std_logic; attribute dont_touch of G31194: signal is true;
	signal G31206: std_logic; attribute dont_touch of G31206: signal is true;
	signal G31207: std_logic; attribute dont_touch of G31207: signal is true;
	signal G31208: std_logic; attribute dont_touch of G31208: signal is true;
	signal G31209: std_logic; attribute dont_touch of G31209: signal is true;
	signal G31210: std_logic; attribute dont_touch of G31210: signal is true;
	signal G31211: std_logic; attribute dont_touch of G31211: signal is true;
	signal G31212: std_logic; attribute dont_touch of G31212: signal is true;
	signal G31213: std_logic; attribute dont_touch of G31213: signal is true;
	signal G31218: std_logic; attribute dont_touch of G31218: signal is true;
	signal G31219: std_logic; attribute dont_touch of G31219: signal is true;
	signal G31220: std_logic; attribute dont_touch of G31220: signal is true;
	signal G31221: std_logic; attribute dont_touch of G31221: signal is true;
	signal G31222: std_logic; attribute dont_touch of G31222: signal is true;
	signal G31223: std_logic; attribute dont_touch of G31223: signal is true;
	signal G31224: std_logic; attribute dont_touch of G31224: signal is true;
	signal G31225: std_logic; attribute dont_touch of G31225: signal is true;
	signal G31226: std_logic; attribute dont_touch of G31226: signal is true;
	signal G31227: std_logic; attribute dont_touch of G31227: signal is true;
	signal G31228: std_logic; attribute dont_touch of G31228: signal is true;
	signal G31229: std_logic; attribute dont_touch of G31229: signal is true;
	signal G31230: std_logic; attribute dont_touch of G31230: signal is true;
	signal G31231: std_logic; attribute dont_touch of G31231: signal is true;
	signal G31232: std_logic; attribute dont_touch of G31232: signal is true;
	signal G31233: std_logic; attribute dont_touch of G31233: signal is true;
	signal G31237: std_logic; attribute dont_touch of G31237: signal is true;
	signal G31238: std_logic; attribute dont_touch of G31238: signal is true;
	signal G31239: std_logic; attribute dont_touch of G31239: signal is true;
	signal G31240: std_logic; attribute dont_touch of G31240: signal is true;
	signal G31241: std_logic; attribute dont_touch of G31241: signal is true;
	signal G31242: std_logic; attribute dont_touch of G31242: signal is true;
	signal G31243: std_logic; attribute dont_touch of G31243: signal is true;
	signal G31244: std_logic; attribute dont_touch of G31244: signal is true;
	signal G31245: std_logic; attribute dont_touch of G31245: signal is true;
	signal G31246: std_logic; attribute dont_touch of G31246: signal is true;
	signal G31247: std_logic; attribute dont_touch of G31247: signal is true;
	signal G31248: std_logic; attribute dont_touch of G31248: signal is true;
	signal G31249: std_logic; attribute dont_touch of G31249: signal is true;
	signal G31250: std_logic; attribute dont_touch of G31250: signal is true;
	signal G31251: std_logic; attribute dont_touch of G31251: signal is true;
	signal G31252: std_logic; attribute dont_touch of G31252: signal is true;
	signal G31253: std_logic; attribute dont_touch of G31253: signal is true;
	signal G31254: std_logic; attribute dont_touch of G31254: signal is true;
	signal G31255: std_logic; attribute dont_touch of G31255: signal is true;
	signal G31256: std_logic; attribute dont_touch of G31256: signal is true;
	signal G31257: std_logic; attribute dont_touch of G31257: signal is true;
	signal G31258: std_logic; attribute dont_touch of G31258: signal is true;
	signal G31259: std_logic; attribute dont_touch of G31259: signal is true;
	signal G31260: std_logic; attribute dont_touch of G31260: signal is true;
	signal G31261: std_logic; attribute dont_touch of G31261: signal is true;
	signal G31262: std_logic; attribute dont_touch of G31262: signal is true;
	signal G31266: std_logic; attribute dont_touch of G31266: signal is true;
	signal G31267: std_logic; attribute dont_touch of G31267: signal is true;
	signal G31268: std_logic; attribute dont_touch of G31268: signal is true;
	signal G31269: std_logic; attribute dont_touch of G31269: signal is true;
	signal G31270: std_logic; attribute dont_touch of G31270: signal is true;
	signal G31271: std_logic; attribute dont_touch of G31271: signal is true;
	signal G31272: std_logic; attribute dont_touch of G31272: signal is true;
	signal G31273: std_logic; attribute dont_touch of G31273: signal is true;
	signal G31274: std_logic; attribute dont_touch of G31274: signal is true;
	signal G31275: std_logic; attribute dont_touch of G31275: signal is true;
	signal G31276: std_logic; attribute dont_touch of G31276: signal is true;
	signal G31277: std_logic; attribute dont_touch of G31277: signal is true;
	signal G31278: std_logic; attribute dont_touch of G31278: signal is true;
	signal G31279: std_logic; attribute dont_touch of G31279: signal is true;
	signal G31280: std_logic; attribute dont_touch of G31280: signal is true;
	signal G31281: std_logic; attribute dont_touch of G31281: signal is true;
	signal G31282: std_logic; attribute dont_touch of G31282: signal is true;
	signal G31283: std_logic; attribute dont_touch of G31283: signal is true;
	signal G31284: std_logic; attribute dont_touch of G31284: signal is true;
	signal G31285: std_logic; attribute dont_touch of G31285: signal is true;
	signal G31286: std_logic; attribute dont_touch of G31286: signal is true;
	signal G31287: std_logic; attribute dont_touch of G31287: signal is true;
	signal G31288: std_logic; attribute dont_touch of G31288: signal is true;
	signal G31289: std_logic; attribute dont_touch of G31289: signal is true;
	signal G31290: std_logic; attribute dont_touch of G31290: signal is true;
	signal G31291: std_logic; attribute dont_touch of G31291: signal is true;
	signal G31292: std_logic; attribute dont_touch of G31292: signal is true;
	signal G31293: std_logic; attribute dont_touch of G31293: signal is true;
	signal G31294: std_logic; attribute dont_touch of G31294: signal is true;
	signal G31295: std_logic; attribute dont_touch of G31295: signal is true;
	signal G31296: std_logic; attribute dont_touch of G31296: signal is true;
	signal G31297: std_logic; attribute dont_touch of G31297: signal is true;
	signal G31298: std_logic; attribute dont_touch of G31298: signal is true;
	signal G31299: std_logic; attribute dont_touch of G31299: signal is true;
	signal G31300: std_logic; attribute dont_touch of G31300: signal is true;
	signal G31301: std_logic; attribute dont_touch of G31301: signal is true;
	signal G31302: std_logic; attribute dont_touch of G31302: signal is true;
	signal G31303: std_logic; attribute dont_touch of G31303: signal is true;
	signal G31304: std_logic; attribute dont_touch of G31304: signal is true;
	signal G31305: std_logic; attribute dont_touch of G31305: signal is true;
	signal G31306: std_logic; attribute dont_touch of G31306: signal is true;
	signal G31307: std_logic; attribute dont_touch of G31307: signal is true;
	signal G31308: std_logic; attribute dont_touch of G31308: signal is true;
	signal G31309: std_logic; attribute dont_touch of G31309: signal is true;
	signal G31310: std_logic; attribute dont_touch of G31310: signal is true;
	signal G31311: std_logic; attribute dont_touch of G31311: signal is true;
	signal G31312: std_logic; attribute dont_touch of G31312: signal is true;
	signal G31313: std_logic; attribute dont_touch of G31313: signal is true;
	signal G31314: std_logic; attribute dont_touch of G31314: signal is true;
	signal G31315: std_logic; attribute dont_touch of G31315: signal is true;
	signal G31316: std_logic; attribute dont_touch of G31316: signal is true;
	signal G31317: std_logic; attribute dont_touch of G31317: signal is true;
	signal G31318: std_logic; attribute dont_touch of G31318: signal is true;
	signal G31319: std_logic; attribute dont_touch of G31319: signal is true;
	signal G31320: std_logic; attribute dont_touch of G31320: signal is true;
	signal G31321: std_logic; attribute dont_touch of G31321: signal is true;
	signal G31322: std_logic; attribute dont_touch of G31322: signal is true;
	signal G31323: std_logic; attribute dont_touch of G31323: signal is true;
	signal G31324: std_logic; attribute dont_touch of G31324: signal is true;
	signal G31325: std_logic; attribute dont_touch of G31325: signal is true;
	signal G31326: std_logic; attribute dont_touch of G31326: signal is true;
	signal G31327: std_logic; attribute dont_touch of G31327: signal is true;
	signal G31372: std_logic; attribute dont_touch of G31372: signal is true;
	signal G31373: std_logic; attribute dont_touch of G31373: signal is true;
	signal G31374: std_logic; attribute dont_touch of G31374: signal is true;
	signal G31375: std_logic; attribute dont_touch of G31375: signal is true;
	signal G31376: std_logic; attribute dont_touch of G31376: signal is true;
	signal G31465: std_logic; attribute dont_touch of G31465: signal is true;
	signal G31466: std_logic; attribute dont_touch of G31466: signal is true;
	signal G31467: std_logic; attribute dont_touch of G31467: signal is true;
	signal G31468: std_logic; attribute dont_touch of G31468: signal is true;
	signal G31469: std_logic; attribute dont_touch of G31469: signal is true;
	signal G31470: std_logic; attribute dont_touch of G31470: signal is true;
	signal G31471: std_logic; attribute dont_touch of G31471: signal is true;
	signal G31472: std_logic; attribute dont_touch of G31472: signal is true;
	signal G31473: std_logic; attribute dont_touch of G31473: signal is true;
	signal G31474: std_logic; attribute dont_touch of G31474: signal is true;
	signal G31475: std_logic; attribute dont_touch of G31475: signal is true;
	signal G31476: std_logic; attribute dont_touch of G31476: signal is true;
	signal G31477: std_logic; attribute dont_touch of G31477: signal is true;
	signal G31478: std_logic; attribute dont_touch of G31478: signal is true;
	signal G31479: std_logic; attribute dont_touch of G31479: signal is true;
	signal G31480: std_logic; attribute dont_touch of G31480: signal is true;
	signal G31481: std_logic; attribute dont_touch of G31481: signal is true;
	signal G31482: std_logic; attribute dont_touch of G31482: signal is true;
	signal G31483: std_logic; attribute dont_touch of G31483: signal is true;
	signal G31484: std_logic; attribute dont_touch of G31484: signal is true;
	signal G31485: std_logic; attribute dont_touch of G31485: signal is true;
	signal G31486: std_logic; attribute dont_touch of G31486: signal is true;
	signal G31487: std_logic; attribute dont_touch of G31487: signal is true;
	signal G31488: std_logic; attribute dont_touch of G31488: signal is true;
	signal G31489: std_logic; attribute dont_touch of G31489: signal is true;
	signal G31490: std_logic; attribute dont_touch of G31490: signal is true;
	signal G31491: std_logic; attribute dont_touch of G31491: signal is true;
	signal G31492: std_logic; attribute dont_touch of G31492: signal is true;
	signal G31493: std_logic; attribute dont_touch of G31493: signal is true;
	signal G31494: std_logic; attribute dont_touch of G31494: signal is true;
	signal G31495: std_logic; attribute dont_touch of G31495: signal is true;
	signal G31496: std_logic; attribute dont_touch of G31496: signal is true;
	signal G31497: std_logic; attribute dont_touch of G31497: signal is true;
	signal G31498: std_logic; attribute dont_touch of G31498: signal is true;
	signal G31499: std_logic; attribute dont_touch of G31499: signal is true;
	signal G31500: std_logic; attribute dont_touch of G31500: signal is true;
	signal G31501: std_logic; attribute dont_touch of G31501: signal is true;
	signal G31502: std_logic; attribute dont_touch of G31502: signal is true;
	signal G31503: std_logic; attribute dont_touch of G31503: signal is true;
	signal G31504: std_logic; attribute dont_touch of G31504: signal is true;
	signal G31505: std_logic; attribute dont_touch of G31505: signal is true;
	signal G31506: std_logic; attribute dont_touch of G31506: signal is true;
	signal G31507: std_logic; attribute dont_touch of G31507: signal is true;
	signal G31508: std_logic; attribute dont_touch of G31508: signal is true;
	signal G31509: std_logic; attribute dont_touch of G31509: signal is true;
	signal G31513: std_logic; attribute dont_touch of G31513: signal is true;
	signal G31514: std_logic; attribute dont_touch of G31514: signal is true;
	signal G31515: std_logic; attribute dont_touch of G31515: signal is true;
	signal G31516: std_logic; attribute dont_touch of G31516: signal is true;
	signal G31517: std_logic; attribute dont_touch of G31517: signal is true;
	signal G31518: std_logic; attribute dont_touch of G31518: signal is true;
	signal G31519: std_logic; attribute dont_touch of G31519: signal is true;
	signal G31520: std_logic; attribute dont_touch of G31520: signal is true;
	signal G31522: std_logic; attribute dont_touch of G31522: signal is true;
	signal G31523: std_logic; attribute dont_touch of G31523: signal is true;
	signal G31524: std_logic; attribute dont_touch of G31524: signal is true;
	signal G31525: std_logic; attribute dont_touch of G31525: signal is true;
	signal G31526: std_logic; attribute dont_touch of G31526: signal is true;
	signal G31527: std_logic; attribute dont_touch of G31527: signal is true;
	signal G31528: std_logic; attribute dont_touch of G31528: signal is true;
	signal G31540: std_logic; attribute dont_touch of G31540: signal is true;
	signal G31541: std_logic; attribute dont_touch of G31541: signal is true;
	signal G31542: std_logic; attribute dont_touch of G31542: signal is true;
	signal G31554: std_logic; attribute dont_touch of G31554: signal is true;
	signal G31566: std_logic; attribute dont_touch of G31566: signal is true;
	signal G31578: std_logic; attribute dont_touch of G31578: signal is true;
	signal G31579: std_logic; attribute dont_touch of G31579: signal is true;
	signal G31591: std_logic; attribute dont_touch of G31591: signal is true;
	signal G31596: std_logic; attribute dont_touch of G31596: signal is true;
	signal G31601: std_logic; attribute dont_touch of G31601: signal is true;
	signal G31608: std_logic; attribute dont_touch of G31608: signal is true;
	signal G31609: std_logic; attribute dont_touch of G31609: signal is true;
	signal G31616: std_logic; attribute dont_touch of G31616: signal is true;
	signal G31623: std_logic; attribute dont_touch of G31623: signal is true;
	signal G31624: std_logic; attribute dont_touch of G31624: signal is true;
	signal G31631: std_logic; attribute dont_touch of G31631: signal is true;
	signal G31638: std_logic; attribute dont_touch of G31638: signal is true;
	signal G31639: std_logic; attribute dont_touch of G31639: signal is true;
	signal G31646: std_logic; attribute dont_touch of G31646: signal is true;
	signal G31653: std_logic; attribute dont_touch of G31653: signal is true;
	signal G31654: std_logic; attribute dont_touch of G31654: signal is true;
	signal G31655: std_logic; attribute dont_touch of G31655: signal is true;
	signal G31657: std_logic; attribute dont_touch of G31657: signal is true;
	signal G31658: std_logic; attribute dont_touch of G31658: signal is true;
	signal G31666: std_logic; attribute dont_touch of G31666: signal is true;
	signal G31667: std_logic; attribute dont_touch of G31667: signal is true;
	signal G31668: std_logic; attribute dont_touch of G31668: signal is true;
	signal G31669: std_logic; attribute dont_touch of G31669: signal is true;
	signal G31670: std_logic; attribute dont_touch of G31670: signal is true;
	signal G31671: std_logic; attribute dont_touch of G31671: signal is true;
	signal G31672: std_logic; attribute dont_touch of G31672: signal is true;
	signal G31706: std_logic; attribute dont_touch of G31706: signal is true;
	signal G31707: std_logic; attribute dont_touch of G31707: signal is true;
	signal G31708: std_logic; attribute dont_touch of G31708: signal is true;
	signal G31709: std_logic; attribute dont_touch of G31709: signal is true;
	signal G31710: std_logic; attribute dont_touch of G31710: signal is true;
	signal G31744: std_logic; attribute dont_touch of G31744: signal is true;
	signal G31745: std_logic; attribute dont_touch of G31745: signal is true;
	signal G31746: std_logic; attribute dont_touch of G31746: signal is true;
	signal G31747: std_logic; attribute dont_touch of G31747: signal is true;
	signal G31748: std_logic; attribute dont_touch of G31748: signal is true;
	signal G31749: std_logic; attribute dont_touch of G31749: signal is true;
	signal G31750: std_logic; attribute dont_touch of G31750: signal is true;
	signal G31751: std_logic; attribute dont_touch of G31751: signal is true;
	signal G31752: std_logic; attribute dont_touch of G31752: signal is true;
	signal G31753: std_logic; attribute dont_touch of G31753: signal is true;
	signal G31754: std_logic; attribute dont_touch of G31754: signal is true;
	signal G31755: std_logic; attribute dont_touch of G31755: signal is true;
	signal G31756: std_logic; attribute dont_touch of G31756: signal is true;
	signal G31757: std_logic; attribute dont_touch of G31757: signal is true;
	signal G31758: std_logic; attribute dont_touch of G31758: signal is true;
	signal G31759: std_logic; attribute dont_touch of G31759: signal is true;
	signal G31760: std_logic; attribute dont_touch of G31760: signal is true;
	signal G31761: std_logic; attribute dont_touch of G31761: signal is true;
	signal G31762: std_logic; attribute dont_touch of G31762: signal is true;
	signal G31763: std_logic; attribute dont_touch of G31763: signal is true;
	signal G31764: std_logic; attribute dont_touch of G31764: signal is true;
	signal G31765: std_logic; attribute dont_touch of G31765: signal is true;
	signal G31766: std_logic; attribute dont_touch of G31766: signal is true;
	signal G31767: std_logic; attribute dont_touch of G31767: signal is true;
	signal G31768: std_logic; attribute dont_touch of G31768: signal is true;
	signal G31769: std_logic; attribute dont_touch of G31769: signal is true;
	signal G31770: std_logic; attribute dont_touch of G31770: signal is true;
	signal G31771: std_logic; attribute dont_touch of G31771: signal is true;
	signal G31772: std_logic; attribute dont_touch of G31772: signal is true;
	signal G31773: std_logic; attribute dont_touch of G31773: signal is true;
	signal G31774: std_logic; attribute dont_touch of G31774: signal is true;
	signal G31775: std_logic; attribute dont_touch of G31775: signal is true;
	signal G31776: std_logic; attribute dont_touch of G31776: signal is true;
	signal G31777: std_logic; attribute dont_touch of G31777: signal is true;
	signal G31778: std_logic; attribute dont_touch of G31778: signal is true;
	signal G31779: std_logic; attribute dont_touch of G31779: signal is true;
	signal G31780: std_logic; attribute dont_touch of G31780: signal is true;
	signal G31781: std_logic; attribute dont_touch of G31781: signal is true;
	signal G31782: std_logic; attribute dont_touch of G31782: signal is true;
	signal G31783: std_logic; attribute dont_touch of G31783: signal is true;
	signal G31784: std_logic; attribute dont_touch of G31784: signal is true;
	signal G31785: std_logic; attribute dont_touch of G31785: signal is true;
	signal G31786: std_logic; attribute dont_touch of G31786: signal is true;
	signal G31787: std_logic; attribute dont_touch of G31787: signal is true;
	signal G31788: std_logic; attribute dont_touch of G31788: signal is true;
	signal G31789: std_logic; attribute dont_touch of G31789: signal is true;
	signal G31790: std_logic; attribute dont_touch of G31790: signal is true;
	signal G31791: std_logic; attribute dont_touch of G31791: signal is true;
	signal G31792: std_logic; attribute dont_touch of G31792: signal is true;
	signal G31794: std_logic; attribute dont_touch of G31794: signal is true;
	signal G31795: std_logic; attribute dont_touch of G31795: signal is true;
	signal G31796: std_logic; attribute dont_touch of G31796: signal is true;
	signal G31797: std_logic; attribute dont_touch of G31797: signal is true;
	signal G31798: std_logic; attribute dont_touch of G31798: signal is true;
	signal G31799: std_logic; attribute dont_touch of G31799: signal is true;
	signal G31800: std_logic; attribute dont_touch of G31800: signal is true;
	signal G31801: std_logic; attribute dont_touch of G31801: signal is true;
	signal G31802: std_logic; attribute dont_touch of G31802: signal is true;
	signal G31803: std_logic; attribute dont_touch of G31803: signal is true;
	signal G31804: std_logic; attribute dont_touch of G31804: signal is true;
	signal G31805: std_logic; attribute dont_touch of G31805: signal is true;
	signal G31806: std_logic; attribute dont_touch of G31806: signal is true;
	signal G31807: std_logic; attribute dont_touch of G31807: signal is true;
	signal G31808: std_logic; attribute dont_touch of G31808: signal is true;
	signal G31809: std_logic; attribute dont_touch of G31809: signal is true;
	signal G31810: std_logic; attribute dont_touch of G31810: signal is true;
	signal G31811: std_logic; attribute dont_touch of G31811: signal is true;
	signal G31812: std_logic; attribute dont_touch of G31812: signal is true;
	signal G31813: std_logic; attribute dont_touch of G31813: signal is true;
	signal G31814: std_logic; attribute dont_touch of G31814: signal is true;
	signal G31815: std_logic; attribute dont_touch of G31815: signal is true;
	signal G31816: std_logic; attribute dont_touch of G31816: signal is true;
	signal G31817: std_logic; attribute dont_touch of G31817: signal is true;
	signal G31818: std_logic; attribute dont_touch of G31818: signal is true;
	signal G31819: std_logic; attribute dont_touch of G31819: signal is true;
	signal G31820: std_logic; attribute dont_touch of G31820: signal is true;
	signal G31821: std_logic; attribute dont_touch of G31821: signal is true;
	signal G31822: std_logic; attribute dont_touch of G31822: signal is true;
	signal G31823: std_logic; attribute dont_touch of G31823: signal is true;
	signal G31824: std_logic; attribute dont_touch of G31824: signal is true;
	signal G31825: std_logic; attribute dont_touch of G31825: signal is true;
	signal G31826: std_logic; attribute dont_touch of G31826: signal is true;
	signal G31827: std_logic; attribute dont_touch of G31827: signal is true;
	signal G31828: std_logic; attribute dont_touch of G31828: signal is true;
	signal G31829: std_logic; attribute dont_touch of G31829: signal is true;
	signal G31830: std_logic; attribute dont_touch of G31830: signal is true;
	signal G31831: std_logic; attribute dont_touch of G31831: signal is true;
	signal G31832: std_logic; attribute dont_touch of G31832: signal is true;
	signal G31833: std_logic; attribute dont_touch of G31833: signal is true;
	signal G31834: std_logic; attribute dont_touch of G31834: signal is true;
	signal G31835: std_logic; attribute dont_touch of G31835: signal is true;
	signal G31836: std_logic; attribute dont_touch of G31836: signal is true;
	signal G31837: std_logic; attribute dont_touch of G31837: signal is true;
	signal G31838: std_logic; attribute dont_touch of G31838: signal is true;
	signal G31839: std_logic; attribute dont_touch of G31839: signal is true;
	signal G31840: std_logic; attribute dont_touch of G31840: signal is true;
	signal G31841: std_logic; attribute dont_touch of G31841: signal is true;
	signal G31842: std_logic; attribute dont_touch of G31842: signal is true;
	signal G31843: std_logic; attribute dont_touch of G31843: signal is true;
	signal G31844: std_logic; attribute dont_touch of G31844: signal is true;
	signal G31845: std_logic; attribute dont_touch of G31845: signal is true;
	signal G31846: std_logic; attribute dont_touch of G31846: signal is true;
	signal G31847: std_logic; attribute dont_touch of G31847: signal is true;
	signal G31848: std_logic; attribute dont_touch of G31848: signal is true;
	signal G31849: std_logic; attribute dont_touch of G31849: signal is true;
	signal G31850: std_logic; attribute dont_touch of G31850: signal is true;
	signal G31851: std_logic; attribute dont_touch of G31851: signal is true;
	signal G31852: std_logic; attribute dont_touch of G31852: signal is true;
	signal G31853: std_logic; attribute dont_touch of G31853: signal is true;
	signal G31854: std_logic; attribute dont_touch of G31854: signal is true;
	signal G31855: std_logic; attribute dont_touch of G31855: signal is true;
	signal G31856: std_logic; attribute dont_touch of G31856: signal is true;
	signal G31857: std_logic; attribute dont_touch of G31857: signal is true;
	signal G31858: std_logic; attribute dont_touch of G31858: signal is true;
	signal G31859: std_logic; attribute dont_touch of G31859: signal is true;
	signal G31864: std_logic; attribute dont_touch of G31864: signal is true;
	signal G31865: std_logic; attribute dont_touch of G31865: signal is true;
	signal G31866: std_logic; attribute dont_touch of G31866: signal is true;
	signal G31867: std_logic; attribute dont_touch of G31867: signal is true;
	signal G31868: std_logic; attribute dont_touch of G31868: signal is true;
	signal G31869: std_logic; attribute dont_touch of G31869: signal is true;
	signal G31870: std_logic; attribute dont_touch of G31870: signal is true;
	signal G31871: std_logic; attribute dont_touch of G31871: signal is true;
	signal G31872: std_logic; attribute dont_touch of G31872: signal is true;
	signal G31873: std_logic; attribute dont_touch of G31873: signal is true;
	signal G31874: std_logic; attribute dont_touch of G31874: signal is true;
	signal G31875: std_logic; attribute dont_touch of G31875: signal is true;
	signal G31876: std_logic; attribute dont_touch of G31876: signal is true;
	signal G31877: std_logic; attribute dont_touch of G31877: signal is true;
	signal G31878: std_logic; attribute dont_touch of G31878: signal is true;
	signal G31879: std_logic; attribute dont_touch of G31879: signal is true;
	signal G31880: std_logic; attribute dont_touch of G31880: signal is true;
	signal G31881: std_logic; attribute dont_touch of G31881: signal is true;
	signal G31882: std_logic; attribute dont_touch of G31882: signal is true;
	signal G31883: std_logic; attribute dont_touch of G31883: signal is true;
	signal G31884: std_logic; attribute dont_touch of G31884: signal is true;
	signal G31885: std_logic; attribute dont_touch of G31885: signal is true;
	signal G31886: std_logic; attribute dont_touch of G31886: signal is true;
	signal G31887: std_logic; attribute dont_touch of G31887: signal is true;
	signal G31888: std_logic; attribute dont_touch of G31888: signal is true;
	signal G31889: std_logic; attribute dont_touch of G31889: signal is true;
	signal G31890: std_logic; attribute dont_touch of G31890: signal is true;
	signal G31891: std_logic; attribute dont_touch of G31891: signal is true;
	signal G31892: std_logic; attribute dont_touch of G31892: signal is true;
	signal G31893: std_logic; attribute dont_touch of G31893: signal is true;
	signal G31894: std_logic; attribute dont_touch of G31894: signal is true;
	signal G31895: std_logic; attribute dont_touch of G31895: signal is true;
	signal G31896: std_logic; attribute dont_touch of G31896: signal is true;
	signal G31897: std_logic; attribute dont_touch of G31897: signal is true;
	signal G31898: std_logic; attribute dont_touch of G31898: signal is true;
	signal G31899: std_logic; attribute dont_touch of G31899: signal is true;
	signal G31900: std_logic; attribute dont_touch of G31900: signal is true;
	signal G31901: std_logic; attribute dont_touch of G31901: signal is true;
	signal G31902: std_logic; attribute dont_touch of G31902: signal is true;
	signal G31903: std_logic; attribute dont_touch of G31903: signal is true;
	signal G31904: std_logic; attribute dont_touch of G31904: signal is true;
	signal G31905: std_logic; attribute dont_touch of G31905: signal is true;
	signal G31906: std_logic; attribute dont_touch of G31906: signal is true;
	signal G31907: std_logic; attribute dont_touch of G31907: signal is true;
	signal G31908: std_logic; attribute dont_touch of G31908: signal is true;
	signal G31909: std_logic; attribute dont_touch of G31909: signal is true;
	signal G31910: std_logic; attribute dont_touch of G31910: signal is true;
	signal G31911: std_logic; attribute dont_touch of G31911: signal is true;
	signal G31912: std_logic; attribute dont_touch of G31912: signal is true;
	signal G31913: std_logic; attribute dont_touch of G31913: signal is true;
	signal G31914: std_logic; attribute dont_touch of G31914: signal is true;
	signal G31915: std_logic; attribute dont_touch of G31915: signal is true;
	signal G31916: std_logic; attribute dont_touch of G31916: signal is true;
	signal G31917: std_logic; attribute dont_touch of G31917: signal is true;
	signal G31918: std_logic; attribute dont_touch of G31918: signal is true;
	signal G31919: std_logic; attribute dont_touch of G31919: signal is true;
	signal G31920: std_logic; attribute dont_touch of G31920: signal is true;
	signal G31921: std_logic; attribute dont_touch of G31921: signal is true;
	signal G31922: std_logic; attribute dont_touch of G31922: signal is true;
	signal G31923: std_logic; attribute dont_touch of G31923: signal is true;
	signal G31924: std_logic; attribute dont_touch of G31924: signal is true;
	signal G31925: std_logic; attribute dont_touch of G31925: signal is true;
	signal G31926: std_logic; attribute dont_touch of G31926: signal is true;
	signal G31927: std_logic; attribute dont_touch of G31927: signal is true;
	signal G31928: std_logic; attribute dont_touch of G31928: signal is true;
	signal G31929: std_logic; attribute dont_touch of G31929: signal is true;
	signal G31930: std_logic; attribute dont_touch of G31930: signal is true;
	signal G31931: std_logic; attribute dont_touch of G31931: signal is true;
	signal G31932: std_logic; attribute dont_touch of G31932: signal is true;
	signal G31933: std_logic; attribute dont_touch of G31933: signal is true;
	signal G31934: std_logic; attribute dont_touch of G31934: signal is true;
	signal G31935: std_logic; attribute dont_touch of G31935: signal is true;
	signal G31936: std_logic; attribute dont_touch of G31936: signal is true;
	signal G31937: std_logic; attribute dont_touch of G31937: signal is true;
	signal G31940: std_logic; attribute dont_touch of G31940: signal is true;
	signal G31941: std_logic; attribute dont_touch of G31941: signal is true;
	signal G31942: std_logic; attribute dont_touch of G31942: signal is true;
	signal G31943: std_logic; attribute dont_touch of G31943: signal is true;
	signal G31944: std_logic; attribute dont_touch of G31944: signal is true;
	signal G31945: std_logic; attribute dont_touch of G31945: signal is true;
	signal G31948: std_logic; attribute dont_touch of G31948: signal is true;
	signal G31949: std_logic; attribute dont_touch of G31949: signal is true;
	signal G31950: std_logic; attribute dont_touch of G31950: signal is true;
	signal G31959: std_logic; attribute dont_touch of G31959: signal is true;
	signal G31960: std_logic; attribute dont_touch of G31960: signal is true;
	signal G31961: std_logic; attribute dont_touch of G31961: signal is true;
	signal G31962: std_logic; attribute dont_touch of G31962: signal is true;
	signal G31963: std_logic; attribute dont_touch of G31963: signal is true;
	signal G31964: std_logic; attribute dont_touch of G31964: signal is true;
	signal G31965: std_logic; attribute dont_touch of G31965: signal is true;
	signal G31966: std_logic; attribute dont_touch of G31966: signal is true;
	signal G31967: std_logic; attribute dont_touch of G31967: signal is true;
	signal G31968: std_logic; attribute dont_touch of G31968: signal is true;
	signal G31969: std_logic; attribute dont_touch of G31969: signal is true;
	signal G31970: std_logic; attribute dont_touch of G31970: signal is true;
	signal G31971: std_logic; attribute dont_touch of G31971: signal is true;
	signal G31974: std_logic; attribute dont_touch of G31974: signal is true;
	signal G31975: std_logic; attribute dont_touch of G31975: signal is true;
	signal G31976: std_logic; attribute dont_touch of G31976: signal is true;
	signal G31977: std_logic; attribute dont_touch of G31977: signal is true;
	signal G31978: std_logic; attribute dont_touch of G31978: signal is true;
	signal G31985: std_logic; attribute dont_touch of G31985: signal is true;
	signal G31986: std_logic; attribute dont_touch of G31986: signal is true;
	signal G31987: std_logic; attribute dont_touch of G31987: signal is true;
	signal G31988: std_logic; attribute dont_touch of G31988: signal is true;
	signal G31989: std_logic; attribute dont_touch of G31989: signal is true;
	signal G31990: std_logic; attribute dont_touch of G31990: signal is true;
	signal G31991: std_logic; attribute dont_touch of G31991: signal is true;
	signal G31992: std_logic; attribute dont_touch of G31992: signal is true;
	signal G31993: std_logic; attribute dont_touch of G31993: signal is true;
	signal G31994: std_logic; attribute dont_touch of G31994: signal is true;
	signal G31995: std_logic; attribute dont_touch of G31995: signal is true;
	signal G31996: std_logic; attribute dont_touch of G31996: signal is true;
	signal G31997: std_logic; attribute dont_touch of G31997: signal is true;
	signal G32008: std_logic; attribute dont_touch of G32008: signal is true;
	signal G32009: std_logic; attribute dont_touch of G32009: signal is true;
	signal G32010: std_logic; attribute dont_touch of G32010: signal is true;
	signal G32011: std_logic; attribute dont_touch of G32011: signal is true;
	signal G32012: std_logic; attribute dont_touch of G32012: signal is true;
	signal G32013: std_logic; attribute dont_touch of G32013: signal is true;
	signal G32014: std_logic; attribute dont_touch of G32014: signal is true;
	signal G32015: std_logic; attribute dont_touch of G32015: signal is true;
	signal G32016: std_logic; attribute dont_touch of G32016: signal is true;
	signal G32017: std_logic; attribute dont_touch of G32017: signal is true;
	signal G32018: std_logic; attribute dont_touch of G32018: signal is true;
	signal G32019: std_logic; attribute dont_touch of G32019: signal is true;
	signal G32020: std_logic; attribute dont_touch of G32020: signal is true;
	signal G32021: std_logic; attribute dont_touch of G32021: signal is true;
	signal G32024: std_logic; attribute dont_touch of G32024: signal is true;
	signal G32027: std_logic; attribute dont_touch of G32027: signal is true;
	signal G32028: std_logic; attribute dont_touch of G32028: signal is true;
	signal G32029: std_logic; attribute dont_touch of G32029: signal is true;
	signal G32030: std_logic; attribute dont_touch of G32030: signal is true;
	signal G32031: std_logic; attribute dont_touch of G32031: signal is true;
	signal G32032: std_logic; attribute dont_touch of G32032: signal is true;
	signal G32033: std_logic; attribute dont_touch of G32033: signal is true;
	signal G32034: std_logic; attribute dont_touch of G32034: signal is true;
	signal G32035: std_logic; attribute dont_touch of G32035: signal is true;
	signal G32036: std_logic; attribute dont_touch of G32036: signal is true;
	signal G32037: std_logic; attribute dont_touch of G32037: signal is true;
	signal G32038: std_logic; attribute dont_touch of G32038: signal is true;
	signal G32039: std_logic; attribute dont_touch of G32039: signal is true;
	signal G32040: std_logic; attribute dont_touch of G32040: signal is true;
	signal G32041: std_logic; attribute dont_touch of G32041: signal is true;
	signal G32042: std_logic; attribute dont_touch of G32042: signal is true;
	signal G32043: std_logic; attribute dont_touch of G32043: signal is true;
	signal G32044: std_logic; attribute dont_touch of G32044: signal is true;
	signal G32045: std_logic; attribute dont_touch of G32045: signal is true;
	signal G32046: std_logic; attribute dont_touch of G32046: signal is true;
	signal G32047: std_logic; attribute dont_touch of G32047: signal is true;
	signal G32048: std_logic; attribute dont_touch of G32048: signal is true;
	signal G32049: std_logic; attribute dont_touch of G32049: signal is true;
	signal G32050: std_logic; attribute dont_touch of G32050: signal is true;
	signal G32051: std_logic; attribute dont_touch of G32051: signal is true;
	signal G32052: std_logic; attribute dont_touch of G32052: signal is true;
	signal G32053: std_logic; attribute dont_touch of G32053: signal is true;
	signal G32054: std_logic; attribute dont_touch of G32054: signal is true;
	signal G32055: std_logic; attribute dont_touch of G32055: signal is true;
	signal G32056: std_logic; attribute dont_touch of G32056: signal is true;
	signal G32057: std_logic; attribute dont_touch of G32057: signal is true;
	signal G32067: std_logic; attribute dont_touch of G32067: signal is true;
	signal G32068: std_logic; attribute dont_touch of G32068: signal is true;
	signal G32069: std_logic; attribute dont_touch of G32069: signal is true;
	signal G32070: std_logic; attribute dont_touch of G32070: signal is true;
	signal G32071: std_logic; attribute dont_touch of G32071: signal is true;
	signal G32072: std_logic; attribute dont_touch of G32072: signal is true;
	signal G32082: std_logic; attribute dont_touch of G32082: signal is true;
	signal G32083: std_logic; attribute dont_touch of G32083: signal is true;
	signal G32084: std_logic; attribute dont_touch of G32084: signal is true;
	signal G32085: std_logic; attribute dont_touch of G32085: signal is true;
	signal G32086: std_logic; attribute dont_touch of G32086: signal is true;
	signal G32087: std_logic; attribute dont_touch of G32087: signal is true;
	signal G32088: std_logic; attribute dont_touch of G32088: signal is true;
	signal G32089: std_logic; attribute dont_touch of G32089: signal is true;
	signal G32090: std_logic; attribute dont_touch of G32090: signal is true;
	signal G32094: std_logic; attribute dont_touch of G32094: signal is true;
	signal G32095: std_logic; attribute dont_touch of G32095: signal is true;
	signal G32096: std_logic; attribute dont_touch of G32096: signal is true;
	signal G32097: std_logic; attribute dont_touch of G32097: signal is true;
	signal G32098: std_logic; attribute dont_touch of G32098: signal is true;
	signal G32099: std_logic; attribute dont_touch of G32099: signal is true;
	signal G32103: std_logic; attribute dont_touch of G32103: signal is true;
	signal G32104: std_logic; attribute dont_touch of G32104: signal is true;
	signal G32105: std_logic; attribute dont_touch of G32105: signal is true;
	signal G32106: std_logic; attribute dont_touch of G32106: signal is true;
	signal G32107: std_logic; attribute dont_touch of G32107: signal is true;
	signal G32108: std_logic; attribute dont_touch of G32108: signal is true;
	signal G32109: std_logic; attribute dont_touch of G32109: signal is true;
	signal G32110: std_logic; attribute dont_touch of G32110: signal is true;
	signal G32111: std_logic; attribute dont_touch of G32111: signal is true;
	signal G32112: std_logic; attribute dont_touch of G32112: signal is true;
	signal G32113: std_logic; attribute dont_touch of G32113: signal is true;
	signal G32114: std_logic; attribute dont_touch of G32114: signal is true;
	signal G32115: std_logic; attribute dont_touch of G32115: signal is true;
	signal G32116: std_logic; attribute dont_touch of G32116: signal is true;
	signal G32117: std_logic; attribute dont_touch of G32117: signal is true;
	signal G32118: std_logic; attribute dont_touch of G32118: signal is true;
	signal G32119: std_logic; attribute dont_touch of G32119: signal is true;
	signal G32120: std_logic; attribute dont_touch of G32120: signal is true;
	signal G32121: std_logic; attribute dont_touch of G32121: signal is true;
	signal G32122: std_logic; attribute dont_touch of G32122: signal is true;
	signal G32123: std_logic; attribute dont_touch of G32123: signal is true;
	signal G32124: std_logic; attribute dont_touch of G32124: signal is true;
	signal G32125: std_logic; attribute dont_touch of G32125: signal is true;
	signal G32126: std_logic; attribute dont_touch of G32126: signal is true;
	signal G32127: std_logic; attribute dont_touch of G32127: signal is true;
	signal G32128: std_logic; attribute dont_touch of G32128: signal is true;
	signal G32129: std_logic; attribute dont_touch of G32129: signal is true;
	signal G32130: std_logic; attribute dont_touch of G32130: signal is true;
	signal G32131: std_logic; attribute dont_touch of G32131: signal is true;
	signal G32132: std_logic; attribute dont_touch of G32132: signal is true;
	signal G32137: std_logic; attribute dont_touch of G32137: signal is true;
	signal G32138: std_logic; attribute dont_touch of G32138: signal is true;
	signal G32139: std_logic; attribute dont_touch of G32139: signal is true;
	signal G32140: std_logic; attribute dont_touch of G32140: signal is true;
	signal G32141: std_logic; attribute dont_touch of G32141: signal is true;
	signal G32142: std_logic; attribute dont_touch of G32142: signal is true;
	signal G32143: std_logic; attribute dont_touch of G32143: signal is true;
	signal G32144: std_logic; attribute dont_touch of G32144: signal is true;
	signal G32145: std_logic; attribute dont_touch of G32145: signal is true;
	signal G32146: std_logic; attribute dont_touch of G32146: signal is true;
	signal G32147: std_logic; attribute dont_touch of G32147: signal is true;
	signal G32148: std_logic; attribute dont_touch of G32148: signal is true;
	signal G32149: std_logic; attribute dont_touch of G32149: signal is true;
	signal G32150: std_logic; attribute dont_touch of G32150: signal is true;
	signal G32151: std_logic; attribute dont_touch of G32151: signal is true;
	signal G32152: std_logic; attribute dont_touch of G32152: signal is true;
	signal G32153: std_logic; attribute dont_touch of G32153: signal is true;
	signal G32154: std_logic; attribute dont_touch of G32154: signal is true;
	signal G32155: std_logic; attribute dont_touch of G32155: signal is true;
	signal G32156: std_logic; attribute dont_touch of G32156: signal is true;
	signal G32157: std_logic; attribute dont_touch of G32157: signal is true;
	signal G32158: std_logic; attribute dont_touch of G32158: signal is true;
	signal G32159: std_logic; attribute dont_touch of G32159: signal is true;
	signal G32160: std_logic; attribute dont_touch of G32160: signal is true;
	signal G32161: std_logic; attribute dont_touch of G32161: signal is true;
	signal G32162: std_logic; attribute dont_touch of G32162: signal is true;
	signal G32163: std_logic; attribute dont_touch of G32163: signal is true;
	signal G32164: std_logic; attribute dont_touch of G32164: signal is true;
	signal G32165: std_logic; attribute dont_touch of G32165: signal is true;
	signal G32166: std_logic; attribute dont_touch of G32166: signal is true;
	signal G32167: std_logic; attribute dont_touch of G32167: signal is true;
	signal G32168: std_logic; attribute dont_touch of G32168: signal is true;
	signal G32169: std_logic; attribute dont_touch of G32169: signal is true;
	signal G32170: std_logic; attribute dont_touch of G32170: signal is true;
	signal G32171: std_logic; attribute dont_touch of G32171: signal is true;
	signal G32172: std_logic; attribute dont_touch of G32172: signal is true;
	signal G32173: std_logic; attribute dont_touch of G32173: signal is true;
	signal G32174: std_logic; attribute dont_touch of G32174: signal is true;
	signal G32175: std_logic; attribute dont_touch of G32175: signal is true;
	signal G32176: std_logic; attribute dont_touch of G32176: signal is true;
	signal G32177: std_logic; attribute dont_touch of G32177: signal is true;
	signal G32178: std_logic; attribute dont_touch of G32178: signal is true;
	signal G32179: std_logic; attribute dont_touch of G32179: signal is true;
	signal G32180: std_logic; attribute dont_touch of G32180: signal is true;
	signal G32181: std_logic; attribute dont_touch of G32181: signal is true;
	signal G32182: std_logic; attribute dont_touch of G32182: signal is true;
	signal G32183: std_logic; attribute dont_touch of G32183: signal is true;
	signal G32184: std_logic; attribute dont_touch of G32184: signal is true;
	signal G32186: std_logic; attribute dont_touch of G32186: signal is true;
	signal G32187: std_logic; attribute dont_touch of G32187: signal is true;
	signal G32188: std_logic; attribute dont_touch of G32188: signal is true;
	signal G32189: std_logic; attribute dont_touch of G32189: signal is true;
	signal G32190: std_logic; attribute dont_touch of G32190: signal is true;
	signal G32191: std_logic; attribute dont_touch of G32191: signal is true;
	signal G32192: std_logic; attribute dont_touch of G32192: signal is true;
	signal G32193: std_logic; attribute dont_touch of G32193: signal is true;
	signal G32194: std_logic; attribute dont_touch of G32194: signal is true;
	signal G32195: std_logic; attribute dont_touch of G32195: signal is true;
	signal G32196: std_logic; attribute dont_touch of G32196: signal is true;
	signal G32197: std_logic; attribute dont_touch of G32197: signal is true;
	signal G32198: std_logic; attribute dont_touch of G32198: signal is true;
	signal G32199: std_logic; attribute dont_touch of G32199: signal is true;
	signal G32200: std_logic; attribute dont_touch of G32200: signal is true;
	signal G32201: std_logic; attribute dont_touch of G32201: signal is true;
	signal G32202: std_logic; attribute dont_touch of G32202: signal is true;
	signal G32203: std_logic; attribute dont_touch of G32203: signal is true;
	signal G32204: std_logic; attribute dont_touch of G32204: signal is true;
	signal G32205: std_logic; attribute dont_touch of G32205: signal is true;
	signal G32206: std_logic; attribute dont_touch of G32206: signal is true;
	signal G32207: std_logic; attribute dont_touch of G32207: signal is true;
	signal G32208: std_logic; attribute dont_touch of G32208: signal is true;
	signal G32209: std_logic; attribute dont_touch of G32209: signal is true;
	signal G32210: std_logic; attribute dont_touch of G32210: signal is true;
	signal G32211: std_logic; attribute dont_touch of G32211: signal is true;
	signal G32212: std_logic; attribute dont_touch of G32212: signal is true;
	signal G32216: std_logic; attribute dont_touch of G32216: signal is true;
	signal G32217: std_logic; attribute dont_touch of G32217: signal is true;
	signal G32218: std_logic; attribute dont_touch of G32218: signal is true;
	signal G32219: std_logic; attribute dont_touch of G32219: signal is true;
	signal G32220: std_logic; attribute dont_touch of G32220: signal is true;
	signal G32221: std_logic; attribute dont_touch of G32221: signal is true;
	signal G32222: std_logic; attribute dont_touch of G32222: signal is true;
	signal G32223: std_logic; attribute dont_touch of G32223: signal is true;
	signal G32224: std_logic; attribute dont_touch of G32224: signal is true;
	signal G32225: std_logic; attribute dont_touch of G32225: signal is true;
	signal G32226: std_logic; attribute dont_touch of G32226: signal is true;
	signal G32227: std_logic; attribute dont_touch of G32227: signal is true;
	signal G32228: std_logic; attribute dont_touch of G32228: signal is true;
	signal G32229: std_logic; attribute dont_touch of G32229: signal is true;
	signal G32230: std_logic; attribute dont_touch of G32230: signal is true;
	signal G32231: std_logic; attribute dont_touch of G32231: signal is true;
	signal G32232: std_logic; attribute dont_touch of G32232: signal is true;
	signal G32233: std_logic; attribute dont_touch of G32233: signal is true;
	signal G32234: std_logic; attribute dont_touch of G32234: signal is true;
	signal G32235: std_logic; attribute dont_touch of G32235: signal is true;
	signal G32236: std_logic; attribute dont_touch of G32236: signal is true;
	signal G32237: std_logic; attribute dont_touch of G32237: signal is true;
	signal G32238: std_logic; attribute dont_touch of G32238: signal is true;
	signal G32239: std_logic; attribute dont_touch of G32239: signal is true;
	signal G32240: std_logic; attribute dont_touch of G32240: signal is true;
	signal G32241: std_logic; attribute dont_touch of G32241: signal is true;
	signal G32242: std_logic; attribute dont_touch of G32242: signal is true;
	signal G32243: std_logic; attribute dont_touch of G32243: signal is true;
	signal G32244: std_logic; attribute dont_touch of G32244: signal is true;
	signal G32245: std_logic; attribute dont_touch of G32245: signal is true;
	signal G32246: std_logic; attribute dont_touch of G32246: signal is true;
	signal G32247: std_logic; attribute dont_touch of G32247: signal is true;
	signal G32248: std_logic; attribute dont_touch of G32248: signal is true;
	signal G32249: std_logic; attribute dont_touch of G32249: signal is true;
	signal G32250: std_logic; attribute dont_touch of G32250: signal is true;
	signal G32251: std_logic; attribute dont_touch of G32251: signal is true;
	signal G32252: std_logic; attribute dont_touch of G32252: signal is true;
	signal G32253: std_logic; attribute dont_touch of G32253: signal is true;
	signal G32254: std_logic; attribute dont_touch of G32254: signal is true;
	signal G32255: std_logic; attribute dont_touch of G32255: signal is true;
	signal G32256: std_logic; attribute dont_touch of G32256: signal is true;
	signal G32257: std_logic; attribute dont_touch of G32257: signal is true;
	signal G32258: std_logic; attribute dont_touch of G32258: signal is true;
	signal G32259: std_logic; attribute dont_touch of G32259: signal is true;
	signal G32260: std_logic; attribute dont_touch of G32260: signal is true;
	signal G32261: std_logic; attribute dont_touch of G32261: signal is true;
	signal G32262: std_logic; attribute dont_touch of G32262: signal is true;
	signal G32263: std_logic; attribute dont_touch of G32263: signal is true;
	signal G32264: std_logic; attribute dont_touch of G32264: signal is true;
	signal G32265: std_logic; attribute dont_touch of G32265: signal is true;
	signal G32266: std_logic; attribute dont_touch of G32266: signal is true;
	signal G32267: std_logic; attribute dont_touch of G32267: signal is true;
	signal G32268: std_logic; attribute dont_touch of G32268: signal is true;
	signal G32269: std_logic; attribute dont_touch of G32269: signal is true;
	signal G32270: std_logic; attribute dont_touch of G32270: signal is true;
	signal G32271: std_logic; attribute dont_touch of G32271: signal is true;
	signal G32272: std_logic; attribute dont_touch of G32272: signal is true;
	signal G32273: std_logic; attribute dont_touch of G32273: signal is true;
	signal G32274: std_logic; attribute dont_touch of G32274: signal is true;
	signal G32275: std_logic; attribute dont_touch of G32275: signal is true;
	signal G32276: std_logic; attribute dont_touch of G32276: signal is true;
	signal G32277: std_logic; attribute dont_touch of G32277: signal is true;
	signal G32278: std_logic; attribute dont_touch of G32278: signal is true;
	signal G32279: std_logic; attribute dont_touch of G32279: signal is true;
	signal G32280: std_logic; attribute dont_touch of G32280: signal is true;
	signal G32281: std_logic; attribute dont_touch of G32281: signal is true;
	signal G32282: std_logic; attribute dont_touch of G32282: signal is true;
	signal G32283: std_logic; attribute dont_touch of G32283: signal is true;
	signal G32284: std_logic; attribute dont_touch of G32284: signal is true;
	signal G32285: std_logic; attribute dont_touch of G32285: signal is true;
	signal G32286: std_logic; attribute dont_touch of G32286: signal is true;
	signal G32287: std_logic; attribute dont_touch of G32287: signal is true;
	signal G32288: std_logic; attribute dont_touch of G32288: signal is true;
	signal G32289: std_logic; attribute dont_touch of G32289: signal is true;
	signal G32290: std_logic; attribute dont_touch of G32290: signal is true;
	signal G32291: std_logic; attribute dont_touch of G32291: signal is true;
	signal G32292: std_logic; attribute dont_touch of G32292: signal is true;
	signal G32293: std_logic; attribute dont_touch of G32293: signal is true;
	signal G32294: std_logic; attribute dont_touch of G32294: signal is true;
	signal G32295: std_logic; attribute dont_touch of G32295: signal is true;
	signal G32296: std_logic; attribute dont_touch of G32296: signal is true;
	signal G32300: std_logic; attribute dont_touch of G32300: signal is true;
	signal G32301: std_logic; attribute dont_touch of G32301: signal is true;
	signal G32302: std_logic; attribute dont_touch of G32302: signal is true;
	signal G32303: std_logic; attribute dont_touch of G32303: signal is true;
	signal G32304: std_logic; attribute dont_touch of G32304: signal is true;
	signal G32305: std_logic; attribute dont_touch of G32305: signal is true;
	signal G32306: std_logic; attribute dont_touch of G32306: signal is true;
	signal G32307: std_logic; attribute dont_touch of G32307: signal is true;
	signal G32308: std_logic; attribute dont_touch of G32308: signal is true;
	signal G32309: std_logic; attribute dont_touch of G32309: signal is true;
	signal G32310: std_logic; attribute dont_touch of G32310: signal is true;
	signal G32311: std_logic; attribute dont_touch of G32311: signal is true;
	signal G32312: std_logic; attribute dont_touch of G32312: signal is true;
	signal G32313: std_logic; attribute dont_touch of G32313: signal is true;
	signal G32314: std_logic; attribute dont_touch of G32314: signal is true;
	signal G32315: std_logic; attribute dont_touch of G32315: signal is true;
	signal G32316: std_logic; attribute dont_touch of G32316: signal is true;
	signal G32317: std_logic; attribute dont_touch of G32317: signal is true;
	signal G32318: std_logic; attribute dont_touch of G32318: signal is true;
	signal G32321: std_logic; attribute dont_touch of G32321: signal is true;
	signal G32322: std_logic; attribute dont_touch of G32322: signal is true;
	signal G32323: std_logic; attribute dont_touch of G32323: signal is true;
	signal G32324: std_logic; attribute dont_touch of G32324: signal is true;
	signal G32325: std_logic; attribute dont_touch of G32325: signal is true;
	signal G32326: std_logic; attribute dont_touch of G32326: signal is true;
	signal G32327: std_logic; attribute dont_touch of G32327: signal is true;
	signal G32328: std_logic; attribute dont_touch of G32328: signal is true;
	signal G32329: std_logic; attribute dont_touch of G32329: signal is true;
	signal G32330: std_logic; attribute dont_touch of G32330: signal is true;
	signal G32331: std_logic; attribute dont_touch of G32331: signal is true;
	signal G32332: std_logic; attribute dont_touch of G32332: signal is true;
	signal G32333: std_logic; attribute dont_touch of G32333: signal is true;
	signal G32334: std_logic; attribute dont_touch of G32334: signal is true;
	signal G32335: std_logic; attribute dont_touch of G32335: signal is true;
	signal G32336: std_logic; attribute dont_touch of G32336: signal is true;
	signal G32337: std_logic; attribute dont_touch of G32337: signal is true;
	signal G32338: std_logic; attribute dont_touch of G32338: signal is true;
	signal G32339: std_logic; attribute dont_touch of G32339: signal is true;
	signal G32340: std_logic; attribute dont_touch of G32340: signal is true;
	signal G32341: std_logic; attribute dont_touch of G32341: signal is true;
	signal G32342: std_logic; attribute dont_touch of G32342: signal is true;
	signal G32343: std_logic; attribute dont_touch of G32343: signal is true;
	signal G32344: std_logic; attribute dont_touch of G32344: signal is true;
	signal G32345: std_logic; attribute dont_touch of G32345: signal is true;
	signal G32346: std_logic; attribute dont_touch of G32346: signal is true;
	signal G32347: std_logic; attribute dont_touch of G32347: signal is true;
	signal G32348: std_logic; attribute dont_touch of G32348: signal is true;
	signal G32349: std_logic; attribute dont_touch of G32349: signal is true;
	signal G32350: std_logic; attribute dont_touch of G32350: signal is true;
	signal G32351: std_logic; attribute dont_touch of G32351: signal is true;
	signal G32352: std_logic; attribute dont_touch of G32352: signal is true;
	signal G32353: std_logic; attribute dont_touch of G32353: signal is true;
	signal G32354: std_logic; attribute dont_touch of G32354: signal is true;
	signal G32355: std_logic; attribute dont_touch of G32355: signal is true;
	signal G32356: std_logic; attribute dont_touch of G32356: signal is true;
	signal G32357: std_logic; attribute dont_touch of G32357: signal is true;
	signal G32358: std_logic; attribute dont_touch of G32358: signal is true;
	signal G32359: std_logic; attribute dont_touch of G32359: signal is true;
	signal G32360: std_logic; attribute dont_touch of G32360: signal is true;
	signal G32361: std_logic; attribute dont_touch of G32361: signal is true;
	signal G32362: std_logic; attribute dont_touch of G32362: signal is true;
	signal G32363: std_logic; attribute dont_touch of G32363: signal is true;
	signal G32364: std_logic; attribute dont_touch of G32364: signal is true;
	signal G32367: std_logic; attribute dont_touch of G32367: signal is true;
	signal G32368: std_logic; attribute dont_touch of G32368: signal is true;
	signal G32369: std_logic; attribute dont_touch of G32369: signal is true;
	signal G32370: std_logic; attribute dont_touch of G32370: signal is true;
	signal G32371: std_logic; attribute dont_touch of G32371: signal is true;
	signal G32372: std_logic; attribute dont_touch of G32372: signal is true;
	signal G32373: std_logic; attribute dont_touch of G32373: signal is true;
	signal G32374: std_logic; attribute dont_touch of G32374: signal is true;
	signal G32375: std_logic; attribute dont_touch of G32375: signal is true;
	signal G32376: std_logic; attribute dont_touch of G32376: signal is true;
	signal G32377: std_logic; attribute dont_touch of G32377: signal is true;
	signal G32380: std_logic; attribute dont_touch of G32380: signal is true;
	signal G32381: std_logic; attribute dont_touch of G32381: signal is true;
	signal G32382: std_logic; attribute dont_touch of G32382: signal is true;
	signal G32383: std_logic; attribute dont_touch of G32383: signal is true;
	signal G32384: std_logic; attribute dont_touch of G32384: signal is true;
	signal G32385: std_logic; attribute dont_touch of G32385: signal is true;
	signal G32386: std_logic; attribute dont_touch of G32386: signal is true;
	signal G32387: std_logic; attribute dont_touch of G32387: signal is true;
	signal G32388: std_logic; attribute dont_touch of G32388: signal is true;
	signal G32389: std_logic; attribute dont_touch of G32389: signal is true;
	signal G32390: std_logic; attribute dont_touch of G32390: signal is true;
	signal G32391: std_logic; attribute dont_touch of G32391: signal is true;
	signal G32392: std_logic; attribute dont_touch of G32392: signal is true;
	signal G32393: std_logic; attribute dont_touch of G32393: signal is true;
	signal G32394: std_logic; attribute dont_touch of G32394: signal is true;
	signal G32395: std_logic; attribute dont_touch of G32395: signal is true;
	signal G32396: std_logic; attribute dont_touch of G32396: signal is true;
	signal G32397: std_logic; attribute dont_touch of G32397: signal is true;
	signal G32398: std_logic; attribute dont_touch of G32398: signal is true;
	signal G32399: std_logic; attribute dont_touch of G32399: signal is true;
	signal G32400: std_logic; attribute dont_touch of G32400: signal is true;
	signal G32401: std_logic; attribute dont_touch of G32401: signal is true;
	signal G32402: std_logic; attribute dont_touch of G32402: signal is true;
	signal G32403: std_logic; attribute dont_touch of G32403: signal is true;
	signal G32404: std_logic; attribute dont_touch of G32404: signal is true;
	signal G32407: std_logic; attribute dont_touch of G32407: signal is true;
	signal G32408: std_logic; attribute dont_touch of G32408: signal is true;
	signal G32409: std_logic; attribute dont_touch of G32409: signal is true;
	signal G32410: std_logic; attribute dont_touch of G32410: signal is true;
	signal G32411: std_logic; attribute dont_touch of G32411: signal is true;
	signal G32412: std_logic; attribute dont_touch of G32412: signal is true;
	signal G32413: std_logic; attribute dont_touch of G32413: signal is true;
	signal G32414: std_logic; attribute dont_touch of G32414: signal is true;
	signal G32415: std_logic; attribute dont_touch of G32415: signal is true;
	signal G32418: std_logic; attribute dont_touch of G32418: signal is true;
	signal G32419: std_logic; attribute dont_touch of G32419: signal is true;
	signal G32420: std_logic; attribute dont_touch of G32420: signal is true;
	signal G32421: std_logic; attribute dont_touch of G32421: signal is true;
	signal G32424: std_logic; attribute dont_touch of G32424: signal is true;
	signal G32425: std_logic; attribute dont_touch of G32425: signal is true;
	signal G32426: std_logic; attribute dont_touch of G32426: signal is true;
	signal G32427: std_logic; attribute dont_touch of G32427: signal is true;
	signal G32428: std_logic; attribute dont_touch of G32428: signal is true;
	signal G32430: std_logic; attribute dont_touch of G32430: signal is true;
	signal G32433: std_logic; attribute dont_touch of G32433: signal is true;
	signal G32434: std_logic; attribute dont_touch of G32434: signal is true;
	signal G32437: std_logic; attribute dont_touch of G32437: signal is true;
	signal G32438: std_logic; attribute dont_touch of G32438: signal is true;
	signal G32441: std_logic; attribute dont_touch of G32441: signal is true;
	signal G32442: std_logic; attribute dont_touch of G32442: signal is true;
	signal G32445: std_logic; attribute dont_touch of G32445: signal is true;
	signal G32446: std_logic; attribute dont_touch of G32446: signal is true;
	signal G32449: std_logic; attribute dont_touch of G32449: signal is true;
	signal G32450: std_logic; attribute dont_touch of G32450: signal is true;
	signal G32453: std_logic; attribute dont_touch of G32453: signal is true;
	signal G32455: std_logic; attribute dont_touch of G32455: signal is true;
	signal G32456: std_logic; attribute dont_touch of G32456: signal is true;
	signal G32457: std_logic; attribute dont_touch of G32457: signal is true;
	signal G32458: std_logic; attribute dont_touch of G32458: signal is true;
	signal G32459: std_logic; attribute dont_touch of G32459: signal is true;
	signal G32460: std_logic; attribute dont_touch of G32460: signal is true;
	signal G32461: std_logic; attribute dont_touch of G32461: signal is true;
	signal G32462: std_logic; attribute dont_touch of G32462: signal is true;
	signal G32463: std_logic; attribute dont_touch of G32463: signal is true;
	signal G32464: std_logic; attribute dont_touch of G32464: signal is true;
	signal G32465: std_logic; attribute dont_touch of G32465: signal is true;
	signal G32466: std_logic; attribute dont_touch of G32466: signal is true;
	signal G32467: std_logic; attribute dont_touch of G32467: signal is true;
	signal G32468: std_logic; attribute dont_touch of G32468: signal is true;
	signal G32469: std_logic; attribute dont_touch of G32469: signal is true;
	signal G32470: std_logic; attribute dont_touch of G32470: signal is true;
	signal G32471: std_logic; attribute dont_touch of G32471: signal is true;
	signal G32472: std_logic; attribute dont_touch of G32472: signal is true;
	signal G32473: std_logic; attribute dont_touch of G32473: signal is true;
	signal G32474: std_logic; attribute dont_touch of G32474: signal is true;
	signal G32475: std_logic; attribute dont_touch of G32475: signal is true;
	signal G32476: std_logic; attribute dont_touch of G32476: signal is true;
	signal G32477: std_logic; attribute dont_touch of G32477: signal is true;
	signal G32478: std_logic; attribute dont_touch of G32478: signal is true;
	signal G32479: std_logic; attribute dont_touch of G32479: signal is true;
	signal G32480: std_logic; attribute dont_touch of G32480: signal is true;
	signal G32481: std_logic; attribute dont_touch of G32481: signal is true;
	signal G32482: std_logic; attribute dont_touch of G32482: signal is true;
	signal G32483: std_logic; attribute dont_touch of G32483: signal is true;
	signal G32484: std_logic; attribute dont_touch of G32484: signal is true;
	signal G32485: std_logic; attribute dont_touch of G32485: signal is true;
	signal G32486: std_logic; attribute dont_touch of G32486: signal is true;
	signal G32487: std_logic; attribute dont_touch of G32487: signal is true;
	signal G32488: std_logic; attribute dont_touch of G32488: signal is true;
	signal G32489: std_logic; attribute dont_touch of G32489: signal is true;
	signal G32490: std_logic; attribute dont_touch of G32490: signal is true;
	signal G32491: std_logic; attribute dont_touch of G32491: signal is true;
	signal G32492: std_logic; attribute dont_touch of G32492: signal is true;
	signal G32493: std_logic; attribute dont_touch of G32493: signal is true;
	signal G32494: std_logic; attribute dont_touch of G32494: signal is true;
	signal G32495: std_logic; attribute dont_touch of G32495: signal is true;
	signal G32496: std_logic; attribute dont_touch of G32496: signal is true;
	signal G32497: std_logic; attribute dont_touch of G32497: signal is true;
	signal G32498: std_logic; attribute dont_touch of G32498: signal is true;
	signal G32499: std_logic; attribute dont_touch of G32499: signal is true;
	signal G32500: std_logic; attribute dont_touch of G32500: signal is true;
	signal G32501: std_logic; attribute dont_touch of G32501: signal is true;
	signal G32502: std_logic; attribute dont_touch of G32502: signal is true;
	signal G32503: std_logic; attribute dont_touch of G32503: signal is true;
	signal G32504: std_logic; attribute dont_touch of G32504: signal is true;
	signal G32505: std_logic; attribute dont_touch of G32505: signal is true;
	signal G32506: std_logic; attribute dont_touch of G32506: signal is true;
	signal G32507: std_logic; attribute dont_touch of G32507: signal is true;
	signal G32508: std_logic; attribute dont_touch of G32508: signal is true;
	signal G32509: std_logic; attribute dont_touch of G32509: signal is true;
	signal G32510: std_logic; attribute dont_touch of G32510: signal is true;
	signal G32511: std_logic; attribute dont_touch of G32511: signal is true;
	signal G32512: std_logic; attribute dont_touch of G32512: signal is true;
	signal G32513: std_logic; attribute dont_touch of G32513: signal is true;
	signal G32514: std_logic; attribute dont_touch of G32514: signal is true;
	signal G32515: std_logic; attribute dont_touch of G32515: signal is true;
	signal G32516: std_logic; attribute dont_touch of G32516: signal is true;
	signal G32517: std_logic; attribute dont_touch of G32517: signal is true;
	signal G32518: std_logic; attribute dont_touch of G32518: signal is true;
	signal G32519: std_logic; attribute dont_touch of G32519: signal is true;
	signal G32520: std_logic; attribute dont_touch of G32520: signal is true;
	signal G32521: std_logic; attribute dont_touch of G32521: signal is true;
	signal G32522: std_logic; attribute dont_touch of G32522: signal is true;
	signal G32523: std_logic; attribute dont_touch of G32523: signal is true;
	signal G32524: std_logic; attribute dont_touch of G32524: signal is true;
	signal G32525: std_logic; attribute dont_touch of G32525: signal is true;
	signal G32526: std_logic; attribute dont_touch of G32526: signal is true;
	signal G32527: std_logic; attribute dont_touch of G32527: signal is true;
	signal G32528: std_logic; attribute dont_touch of G32528: signal is true;
	signal G32529: std_logic; attribute dont_touch of G32529: signal is true;
	signal G32530: std_logic; attribute dont_touch of G32530: signal is true;
	signal G32531: std_logic; attribute dont_touch of G32531: signal is true;
	signal G32532: std_logic; attribute dont_touch of G32532: signal is true;
	signal G32533: std_logic; attribute dont_touch of G32533: signal is true;
	signal G32534: std_logic; attribute dont_touch of G32534: signal is true;
	signal G32535: std_logic; attribute dont_touch of G32535: signal is true;
	signal G32536: std_logic; attribute dont_touch of G32536: signal is true;
	signal G32537: std_logic; attribute dont_touch of G32537: signal is true;
	signal G32538: std_logic; attribute dont_touch of G32538: signal is true;
	signal G32539: std_logic; attribute dont_touch of G32539: signal is true;
	signal G32540: std_logic; attribute dont_touch of G32540: signal is true;
	signal G32541: std_logic; attribute dont_touch of G32541: signal is true;
	signal G32542: std_logic; attribute dont_touch of G32542: signal is true;
	signal G32543: std_logic; attribute dont_touch of G32543: signal is true;
	signal G32544: std_logic; attribute dont_touch of G32544: signal is true;
	signal G32545: std_logic; attribute dont_touch of G32545: signal is true;
	signal G32546: std_logic; attribute dont_touch of G32546: signal is true;
	signal G32547: std_logic; attribute dont_touch of G32547: signal is true;
	signal G32548: std_logic; attribute dont_touch of G32548: signal is true;
	signal G32549: std_logic; attribute dont_touch of G32549: signal is true;
	signal G32550: std_logic; attribute dont_touch of G32550: signal is true;
	signal G32551: std_logic; attribute dont_touch of G32551: signal is true;
	signal G32552: std_logic; attribute dont_touch of G32552: signal is true;
	signal G32553: std_logic; attribute dont_touch of G32553: signal is true;
	signal G32554: std_logic; attribute dont_touch of G32554: signal is true;
	signal G32555: std_logic; attribute dont_touch of G32555: signal is true;
	signal G32556: std_logic; attribute dont_touch of G32556: signal is true;
	signal G32557: std_logic; attribute dont_touch of G32557: signal is true;
	signal G32558: std_logic; attribute dont_touch of G32558: signal is true;
	signal G32559: std_logic; attribute dont_touch of G32559: signal is true;
	signal G32560: std_logic; attribute dont_touch of G32560: signal is true;
	signal G32561: std_logic; attribute dont_touch of G32561: signal is true;
	signal G32562: std_logic; attribute dont_touch of G32562: signal is true;
	signal G32563: std_logic; attribute dont_touch of G32563: signal is true;
	signal G32564: std_logic; attribute dont_touch of G32564: signal is true;
	signal G32565: std_logic; attribute dont_touch of G32565: signal is true;
	signal G32566: std_logic; attribute dont_touch of G32566: signal is true;
	signal G32567: std_logic; attribute dont_touch of G32567: signal is true;
	signal G32568: std_logic; attribute dont_touch of G32568: signal is true;
	signal G32569: std_logic; attribute dont_touch of G32569: signal is true;
	signal G32570: std_logic; attribute dont_touch of G32570: signal is true;
	signal G32571: std_logic; attribute dont_touch of G32571: signal is true;
	signal G32572: std_logic; attribute dont_touch of G32572: signal is true;
	signal G32573: std_logic; attribute dont_touch of G32573: signal is true;
	signal G32574: std_logic; attribute dont_touch of G32574: signal is true;
	signal G32575: std_logic; attribute dont_touch of G32575: signal is true;
	signal G32576: std_logic; attribute dont_touch of G32576: signal is true;
	signal G32577: std_logic; attribute dont_touch of G32577: signal is true;
	signal G32578: std_logic; attribute dont_touch of G32578: signal is true;
	signal G32579: std_logic; attribute dont_touch of G32579: signal is true;
	signal G32580: std_logic; attribute dont_touch of G32580: signal is true;
	signal G32581: std_logic; attribute dont_touch of G32581: signal is true;
	signal G32582: std_logic; attribute dont_touch of G32582: signal is true;
	signal G32583: std_logic; attribute dont_touch of G32583: signal is true;
	signal G32584: std_logic; attribute dont_touch of G32584: signal is true;
	signal G32585: std_logic; attribute dont_touch of G32585: signal is true;
	signal G32586: std_logic; attribute dont_touch of G32586: signal is true;
	signal G32587: std_logic; attribute dont_touch of G32587: signal is true;
	signal G32588: std_logic; attribute dont_touch of G32588: signal is true;
	signal G32589: std_logic; attribute dont_touch of G32589: signal is true;
	signal G32590: std_logic; attribute dont_touch of G32590: signal is true;
	signal G32591: std_logic; attribute dont_touch of G32591: signal is true;
	signal G32592: std_logic; attribute dont_touch of G32592: signal is true;
	signal G32593: std_logic; attribute dont_touch of G32593: signal is true;
	signal G32594: std_logic; attribute dont_touch of G32594: signal is true;
	signal G32595: std_logic; attribute dont_touch of G32595: signal is true;
	signal G32596: std_logic; attribute dont_touch of G32596: signal is true;
	signal G32597: std_logic; attribute dont_touch of G32597: signal is true;
	signal G32598: std_logic; attribute dont_touch of G32598: signal is true;
	signal G32599: std_logic; attribute dont_touch of G32599: signal is true;
	signal G32600: std_logic; attribute dont_touch of G32600: signal is true;
	signal G32601: std_logic; attribute dont_touch of G32601: signal is true;
	signal G32602: std_logic; attribute dont_touch of G32602: signal is true;
	signal G32603: std_logic; attribute dont_touch of G32603: signal is true;
	signal G32604: std_logic; attribute dont_touch of G32604: signal is true;
	signal G32605: std_logic; attribute dont_touch of G32605: signal is true;
	signal G32606: std_logic; attribute dont_touch of G32606: signal is true;
	signal G32607: std_logic; attribute dont_touch of G32607: signal is true;
	signal G32608: std_logic; attribute dont_touch of G32608: signal is true;
	signal G32609: std_logic; attribute dont_touch of G32609: signal is true;
	signal G32610: std_logic; attribute dont_touch of G32610: signal is true;
	signal G32611: std_logic; attribute dont_touch of G32611: signal is true;
	signal G32612: std_logic; attribute dont_touch of G32612: signal is true;
	signal G32613: std_logic; attribute dont_touch of G32613: signal is true;
	signal G32614: std_logic; attribute dont_touch of G32614: signal is true;
	signal G32615: std_logic; attribute dont_touch of G32615: signal is true;
	signal G32616: std_logic; attribute dont_touch of G32616: signal is true;
	signal G32617: std_logic; attribute dont_touch of G32617: signal is true;
	signal G32618: std_logic; attribute dont_touch of G32618: signal is true;
	signal G32619: std_logic; attribute dont_touch of G32619: signal is true;
	signal G32620: std_logic; attribute dont_touch of G32620: signal is true;
	signal G32621: std_logic; attribute dont_touch of G32621: signal is true;
	signal G32622: std_logic; attribute dont_touch of G32622: signal is true;
	signal G32623: std_logic; attribute dont_touch of G32623: signal is true;
	signal G32624: std_logic; attribute dont_touch of G32624: signal is true;
	signal G32625: std_logic; attribute dont_touch of G32625: signal is true;
	signal G32626: std_logic; attribute dont_touch of G32626: signal is true;
	signal G32627: std_logic; attribute dont_touch of G32627: signal is true;
	signal G32628: std_logic; attribute dont_touch of G32628: signal is true;
	signal G32629: std_logic; attribute dont_touch of G32629: signal is true;
	signal G32630: std_logic; attribute dont_touch of G32630: signal is true;
	signal G32631: std_logic; attribute dont_touch of G32631: signal is true;
	signal G32632: std_logic; attribute dont_touch of G32632: signal is true;
	signal G32633: std_logic; attribute dont_touch of G32633: signal is true;
	signal G32634: std_logic; attribute dont_touch of G32634: signal is true;
	signal G32635: std_logic; attribute dont_touch of G32635: signal is true;
	signal G32636: std_logic; attribute dont_touch of G32636: signal is true;
	signal G32637: std_logic; attribute dont_touch of G32637: signal is true;
	signal G32638: std_logic; attribute dont_touch of G32638: signal is true;
	signal G32639: std_logic; attribute dont_touch of G32639: signal is true;
	signal G32640: std_logic; attribute dont_touch of G32640: signal is true;
	signal G32641: std_logic; attribute dont_touch of G32641: signal is true;
	signal G32642: std_logic; attribute dont_touch of G32642: signal is true;
	signal G32643: std_logic; attribute dont_touch of G32643: signal is true;
	signal G32644: std_logic; attribute dont_touch of G32644: signal is true;
	signal G32645: std_logic; attribute dont_touch of G32645: signal is true;
	signal G32646: std_logic; attribute dont_touch of G32646: signal is true;
	signal G32647: std_logic; attribute dont_touch of G32647: signal is true;
	signal G32648: std_logic; attribute dont_touch of G32648: signal is true;
	signal G32649: std_logic; attribute dont_touch of G32649: signal is true;
	signal G32650: std_logic; attribute dont_touch of G32650: signal is true;
	signal G32651: std_logic; attribute dont_touch of G32651: signal is true;
	signal G32652: std_logic; attribute dont_touch of G32652: signal is true;
	signal G32653: std_logic; attribute dont_touch of G32653: signal is true;
	signal G32654: std_logic; attribute dont_touch of G32654: signal is true;
	signal G32655: std_logic; attribute dont_touch of G32655: signal is true;
	signal G32656: std_logic; attribute dont_touch of G32656: signal is true;
	signal G32657: std_logic; attribute dont_touch of G32657: signal is true;
	signal G32658: std_logic; attribute dont_touch of G32658: signal is true;
	signal G32659: std_logic; attribute dont_touch of G32659: signal is true;
	signal G32660: std_logic; attribute dont_touch of G32660: signal is true;
	signal G32661: std_logic; attribute dont_touch of G32661: signal is true;
	signal G32662: std_logic; attribute dont_touch of G32662: signal is true;
	signal G32663: std_logic; attribute dont_touch of G32663: signal is true;
	signal G32664: std_logic; attribute dont_touch of G32664: signal is true;
	signal G32665: std_logic; attribute dont_touch of G32665: signal is true;
	signal G32666: std_logic; attribute dont_touch of G32666: signal is true;
	signal G32667: std_logic; attribute dont_touch of G32667: signal is true;
	signal G32668: std_logic; attribute dont_touch of G32668: signal is true;
	signal G32669: std_logic; attribute dont_touch of G32669: signal is true;
	signal G32670: std_logic; attribute dont_touch of G32670: signal is true;
	signal G32671: std_logic; attribute dont_touch of G32671: signal is true;
	signal G32672: std_logic; attribute dont_touch of G32672: signal is true;
	signal G32673: std_logic; attribute dont_touch of G32673: signal is true;
	signal G32674: std_logic; attribute dont_touch of G32674: signal is true;
	signal G32675: std_logic; attribute dont_touch of G32675: signal is true;
	signal G32676: std_logic; attribute dont_touch of G32676: signal is true;
	signal G32677: std_logic; attribute dont_touch of G32677: signal is true;
	signal G32678: std_logic; attribute dont_touch of G32678: signal is true;
	signal G32679: std_logic; attribute dont_touch of G32679: signal is true;
	signal G32680: std_logic; attribute dont_touch of G32680: signal is true;
	signal G32681: std_logic; attribute dont_touch of G32681: signal is true;
	signal G32682: std_logic; attribute dont_touch of G32682: signal is true;
	signal G32683: std_logic; attribute dont_touch of G32683: signal is true;
	signal G32684: std_logic; attribute dont_touch of G32684: signal is true;
	signal G32685: std_logic; attribute dont_touch of G32685: signal is true;
	signal G32686: std_logic; attribute dont_touch of G32686: signal is true;
	signal G32687: std_logic; attribute dont_touch of G32687: signal is true;
	signal G32688: std_logic; attribute dont_touch of G32688: signal is true;
	signal G32689: std_logic; attribute dont_touch of G32689: signal is true;
	signal G32690: std_logic; attribute dont_touch of G32690: signal is true;
	signal G32691: std_logic; attribute dont_touch of G32691: signal is true;
	signal G32692: std_logic; attribute dont_touch of G32692: signal is true;
	signal G32693: std_logic; attribute dont_touch of G32693: signal is true;
	signal G32694: std_logic; attribute dont_touch of G32694: signal is true;
	signal G32695: std_logic; attribute dont_touch of G32695: signal is true;
	signal G32696: std_logic; attribute dont_touch of G32696: signal is true;
	signal G32697: std_logic; attribute dont_touch of G32697: signal is true;
	signal G32698: std_logic; attribute dont_touch of G32698: signal is true;
	signal G32699: std_logic; attribute dont_touch of G32699: signal is true;
	signal G32700: std_logic; attribute dont_touch of G32700: signal is true;
	signal G32701: std_logic; attribute dont_touch of G32701: signal is true;
	signal G32702: std_logic; attribute dont_touch of G32702: signal is true;
	signal G32703: std_logic; attribute dont_touch of G32703: signal is true;
	signal G32704: std_logic; attribute dont_touch of G32704: signal is true;
	signal G32705: std_logic; attribute dont_touch of G32705: signal is true;
	signal G32706: std_logic; attribute dont_touch of G32706: signal is true;
	signal G32707: std_logic; attribute dont_touch of G32707: signal is true;
	signal G32708: std_logic; attribute dont_touch of G32708: signal is true;
	signal G32709: std_logic; attribute dont_touch of G32709: signal is true;
	signal G32710: std_logic; attribute dont_touch of G32710: signal is true;
	signal G32711: std_logic; attribute dont_touch of G32711: signal is true;
	signal G32712: std_logic; attribute dont_touch of G32712: signal is true;
	signal G32713: std_logic; attribute dont_touch of G32713: signal is true;
	signal G32714: std_logic; attribute dont_touch of G32714: signal is true;
	signal G32715: std_logic; attribute dont_touch of G32715: signal is true;
	signal G32716: std_logic; attribute dont_touch of G32716: signal is true;
	signal G32717: std_logic; attribute dont_touch of G32717: signal is true;
	signal G32718: std_logic; attribute dont_touch of G32718: signal is true;
	signal G32719: std_logic; attribute dont_touch of G32719: signal is true;
	signal G32720: std_logic; attribute dont_touch of G32720: signal is true;
	signal G32721: std_logic; attribute dont_touch of G32721: signal is true;
	signal G32722: std_logic; attribute dont_touch of G32722: signal is true;
	signal G32723: std_logic; attribute dont_touch of G32723: signal is true;
	signal G32724: std_logic; attribute dont_touch of G32724: signal is true;
	signal G32725: std_logic; attribute dont_touch of G32725: signal is true;
	signal G32726: std_logic; attribute dont_touch of G32726: signal is true;
	signal G32727: std_logic; attribute dont_touch of G32727: signal is true;
	signal G32728: std_logic; attribute dont_touch of G32728: signal is true;
	signal G32729: std_logic; attribute dont_touch of G32729: signal is true;
	signal G32730: std_logic; attribute dont_touch of G32730: signal is true;
	signal G32731: std_logic; attribute dont_touch of G32731: signal is true;
	signal G32732: std_logic; attribute dont_touch of G32732: signal is true;
	signal G32733: std_logic; attribute dont_touch of G32733: signal is true;
	signal G32734: std_logic; attribute dont_touch of G32734: signal is true;
	signal G32735: std_logic; attribute dont_touch of G32735: signal is true;
	signal G32736: std_logic; attribute dont_touch of G32736: signal is true;
	signal G32737: std_logic; attribute dont_touch of G32737: signal is true;
	signal G32738: std_logic; attribute dont_touch of G32738: signal is true;
	signal G32739: std_logic; attribute dont_touch of G32739: signal is true;
	signal G32740: std_logic; attribute dont_touch of G32740: signal is true;
	signal G32741: std_logic; attribute dont_touch of G32741: signal is true;
	signal G32742: std_logic; attribute dont_touch of G32742: signal is true;
	signal G32743: std_logic; attribute dont_touch of G32743: signal is true;
	signal G32744: std_logic; attribute dont_touch of G32744: signal is true;
	signal G32745: std_logic; attribute dont_touch of G32745: signal is true;
	signal G32746: std_logic; attribute dont_touch of G32746: signal is true;
	signal G32747: std_logic; attribute dont_touch of G32747: signal is true;
	signal G32748: std_logic; attribute dont_touch of G32748: signal is true;
	signal G32749: std_logic; attribute dont_touch of G32749: signal is true;
	signal G32750: std_logic; attribute dont_touch of G32750: signal is true;
	signal G32751: std_logic; attribute dont_touch of G32751: signal is true;
	signal G32752: std_logic; attribute dont_touch of G32752: signal is true;
	signal G32753: std_logic; attribute dont_touch of G32753: signal is true;
	signal G32754: std_logic; attribute dont_touch of G32754: signal is true;
	signal G32755: std_logic; attribute dont_touch of G32755: signal is true;
	signal G32756: std_logic; attribute dont_touch of G32756: signal is true;
	signal G32757: std_logic; attribute dont_touch of G32757: signal is true;
	signal G32758: std_logic; attribute dont_touch of G32758: signal is true;
	signal G32759: std_logic; attribute dont_touch of G32759: signal is true;
	signal G32760: std_logic; attribute dont_touch of G32760: signal is true;
	signal G32761: std_logic; attribute dont_touch of G32761: signal is true;
	signal G32762: std_logic; attribute dont_touch of G32762: signal is true;
	signal G32763: std_logic; attribute dont_touch of G32763: signal is true;
	signal G32764: std_logic; attribute dont_touch of G32764: signal is true;
	signal G32765: std_logic; attribute dont_touch of G32765: signal is true;
	signal G32766: std_logic; attribute dont_touch of G32766: signal is true;
	signal G32767: std_logic; attribute dont_touch of G32767: signal is true;
	signal G32768: std_logic; attribute dont_touch of G32768: signal is true;
	signal G32769: std_logic; attribute dont_touch of G32769: signal is true;
	signal G32770: std_logic; attribute dont_touch of G32770: signal is true;
	signal G32771: std_logic; attribute dont_touch of G32771: signal is true;
	signal G32772: std_logic; attribute dont_touch of G32772: signal is true;
	signal G32773: std_logic; attribute dont_touch of G32773: signal is true;
	signal G32774: std_logic; attribute dont_touch of G32774: signal is true;
	signal G32775: std_logic; attribute dont_touch of G32775: signal is true;
	signal G32776: std_logic; attribute dont_touch of G32776: signal is true;
	signal G32777: std_logic; attribute dont_touch of G32777: signal is true;
	signal G32778: std_logic; attribute dont_touch of G32778: signal is true;
	signal G32779: std_logic; attribute dont_touch of G32779: signal is true;
	signal G32780: std_logic; attribute dont_touch of G32780: signal is true;
	signal G32781: std_logic; attribute dont_touch of G32781: signal is true;
	signal G32782: std_logic; attribute dont_touch of G32782: signal is true;
	signal G32783: std_logic; attribute dont_touch of G32783: signal is true;
	signal G32784: std_logic; attribute dont_touch of G32784: signal is true;
	signal G32785: std_logic; attribute dont_touch of G32785: signal is true;
	signal G32786: std_logic; attribute dont_touch of G32786: signal is true;
	signal G32787: std_logic; attribute dont_touch of G32787: signal is true;
	signal G32788: std_logic; attribute dont_touch of G32788: signal is true;
	signal G32789: std_logic; attribute dont_touch of G32789: signal is true;
	signal G32790: std_logic; attribute dont_touch of G32790: signal is true;
	signal G32791: std_logic; attribute dont_touch of G32791: signal is true;
	signal G32792: std_logic; attribute dont_touch of G32792: signal is true;
	signal G32793: std_logic; attribute dont_touch of G32793: signal is true;
	signal G32794: std_logic; attribute dont_touch of G32794: signal is true;
	signal G32795: std_logic; attribute dont_touch of G32795: signal is true;
	signal G32796: std_logic; attribute dont_touch of G32796: signal is true;
	signal G32797: std_logic; attribute dont_touch of G32797: signal is true;
	signal G32798: std_logic; attribute dont_touch of G32798: signal is true;
	signal G32799: std_logic; attribute dont_touch of G32799: signal is true;
	signal G32800: std_logic; attribute dont_touch of G32800: signal is true;
	signal G32801: std_logic; attribute dont_touch of G32801: signal is true;
	signal G32802: std_logic; attribute dont_touch of G32802: signal is true;
	signal G32803: std_logic; attribute dont_touch of G32803: signal is true;
	signal G32804: std_logic; attribute dont_touch of G32804: signal is true;
	signal G32805: std_logic; attribute dont_touch of G32805: signal is true;
	signal G32806: std_logic; attribute dont_touch of G32806: signal is true;
	signal G32807: std_logic; attribute dont_touch of G32807: signal is true;
	signal G32808: std_logic; attribute dont_touch of G32808: signal is true;
	signal G32809: std_logic; attribute dont_touch of G32809: signal is true;
	signal G32810: std_logic; attribute dont_touch of G32810: signal is true;
	signal G32811: std_logic; attribute dont_touch of G32811: signal is true;
	signal G32812: std_logic; attribute dont_touch of G32812: signal is true;
	signal G32813: std_logic; attribute dont_touch of G32813: signal is true;
	signal G32814: std_logic; attribute dont_touch of G32814: signal is true;
	signal G32815: std_logic; attribute dont_touch of G32815: signal is true;
	signal G32816: std_logic; attribute dont_touch of G32816: signal is true;
	signal G32817: std_logic; attribute dont_touch of G32817: signal is true;
	signal G32818: std_logic; attribute dont_touch of G32818: signal is true;
	signal G32819: std_logic; attribute dont_touch of G32819: signal is true;
	signal G32820: std_logic; attribute dont_touch of G32820: signal is true;
	signal G32821: std_logic; attribute dont_touch of G32821: signal is true;
	signal G32822: std_logic; attribute dont_touch of G32822: signal is true;
	signal G32823: std_logic; attribute dont_touch of G32823: signal is true;
	signal G32824: std_logic; attribute dont_touch of G32824: signal is true;
	signal G32825: std_logic; attribute dont_touch of G32825: signal is true;
	signal G32826: std_logic; attribute dont_touch of G32826: signal is true;
	signal G32827: std_logic; attribute dont_touch of G32827: signal is true;
	signal G32828: std_logic; attribute dont_touch of G32828: signal is true;
	signal G32829: std_logic; attribute dont_touch of G32829: signal is true;
	signal G32830: std_logic; attribute dont_touch of G32830: signal is true;
	signal G32831: std_logic; attribute dont_touch of G32831: signal is true;
	signal G32832: std_logic; attribute dont_touch of G32832: signal is true;
	signal G32833: std_logic; attribute dont_touch of G32833: signal is true;
	signal G32834: std_logic; attribute dont_touch of G32834: signal is true;
	signal G32835: std_logic; attribute dont_touch of G32835: signal is true;
	signal G32836: std_logic; attribute dont_touch of G32836: signal is true;
	signal G32837: std_logic; attribute dont_touch of G32837: signal is true;
	signal G32838: std_logic; attribute dont_touch of G32838: signal is true;
	signal G32839: std_logic; attribute dont_touch of G32839: signal is true;
	signal G32840: std_logic; attribute dont_touch of G32840: signal is true;
	signal G32841: std_logic; attribute dont_touch of G32841: signal is true;
	signal G32842: std_logic; attribute dont_touch of G32842: signal is true;
	signal G32843: std_logic; attribute dont_touch of G32843: signal is true;
	signal G32844: std_logic; attribute dont_touch of G32844: signal is true;
	signal G32845: std_logic; attribute dont_touch of G32845: signal is true;
	signal G32846: std_logic; attribute dont_touch of G32846: signal is true;
	signal G32847: std_logic; attribute dont_touch of G32847: signal is true;
	signal G32848: std_logic; attribute dont_touch of G32848: signal is true;
	signal G32849: std_logic; attribute dont_touch of G32849: signal is true;
	signal G32850: std_logic; attribute dont_touch of G32850: signal is true;
	signal G32851: std_logic; attribute dont_touch of G32851: signal is true;
	signal G32852: std_logic; attribute dont_touch of G32852: signal is true;
	signal G32853: std_logic; attribute dont_touch of G32853: signal is true;
	signal G32854: std_logic; attribute dont_touch of G32854: signal is true;
	signal G32855: std_logic; attribute dont_touch of G32855: signal is true;
	signal G32856: std_logic; attribute dont_touch of G32856: signal is true;
	signal G32857: std_logic; attribute dont_touch of G32857: signal is true;
	signal G32858: std_logic; attribute dont_touch of G32858: signal is true;
	signal G32859: std_logic; attribute dont_touch of G32859: signal is true;
	signal G32860: std_logic; attribute dont_touch of G32860: signal is true;
	signal G32861: std_logic; attribute dont_touch of G32861: signal is true;
	signal G32862: std_logic; attribute dont_touch of G32862: signal is true;
	signal G32863: std_logic; attribute dont_touch of G32863: signal is true;
	signal G32864: std_logic; attribute dont_touch of G32864: signal is true;
	signal G32865: std_logic; attribute dont_touch of G32865: signal is true;
	signal G32866: std_logic; attribute dont_touch of G32866: signal is true;
	signal G32867: std_logic; attribute dont_touch of G32867: signal is true;
	signal G32868: std_logic; attribute dont_touch of G32868: signal is true;
	signal G32869: std_logic; attribute dont_touch of G32869: signal is true;
	signal G32870: std_logic; attribute dont_touch of G32870: signal is true;
	signal G32871: std_logic; attribute dont_touch of G32871: signal is true;
	signal G32872: std_logic; attribute dont_touch of G32872: signal is true;
	signal G32873: std_logic; attribute dont_touch of G32873: signal is true;
	signal G32874: std_logic; attribute dont_touch of G32874: signal is true;
	signal G32875: std_logic; attribute dont_touch of G32875: signal is true;
	signal G32876: std_logic; attribute dont_touch of G32876: signal is true;
	signal G32877: std_logic; attribute dont_touch of G32877: signal is true;
	signal G32878: std_logic; attribute dont_touch of G32878: signal is true;
	signal G32879: std_logic; attribute dont_touch of G32879: signal is true;
	signal G32880: std_logic; attribute dont_touch of G32880: signal is true;
	signal G32881: std_logic; attribute dont_touch of G32881: signal is true;
	signal G32882: std_logic; attribute dont_touch of G32882: signal is true;
	signal G32883: std_logic; attribute dont_touch of G32883: signal is true;
	signal G32884: std_logic; attribute dont_touch of G32884: signal is true;
	signal G32885: std_logic; attribute dont_touch of G32885: signal is true;
	signal G32886: std_logic; attribute dont_touch of G32886: signal is true;
	signal G32887: std_logic; attribute dont_touch of G32887: signal is true;
	signal G32888: std_logic; attribute dont_touch of G32888: signal is true;
	signal G32889: std_logic; attribute dont_touch of G32889: signal is true;
	signal G32890: std_logic; attribute dont_touch of G32890: signal is true;
	signal G32891: std_logic; attribute dont_touch of G32891: signal is true;
	signal G32892: std_logic; attribute dont_touch of G32892: signal is true;
	signal G32893: std_logic; attribute dont_touch of G32893: signal is true;
	signal G32894: std_logic; attribute dont_touch of G32894: signal is true;
	signal G32895: std_logic; attribute dont_touch of G32895: signal is true;
	signal G32896: std_logic; attribute dont_touch of G32896: signal is true;
	signal G32897: std_logic; attribute dont_touch of G32897: signal is true;
	signal G32898: std_logic; attribute dont_touch of G32898: signal is true;
	signal G32899: std_logic; attribute dont_touch of G32899: signal is true;
	signal G32900: std_logic; attribute dont_touch of G32900: signal is true;
	signal G32901: std_logic; attribute dont_touch of G32901: signal is true;
	signal G32902: std_logic; attribute dont_touch of G32902: signal is true;
	signal G32903: std_logic; attribute dont_touch of G32903: signal is true;
	signal G32904: std_logic; attribute dont_touch of G32904: signal is true;
	signal G32905: std_logic; attribute dont_touch of G32905: signal is true;
	signal G32906: std_logic; attribute dont_touch of G32906: signal is true;
	signal G32907: std_logic; attribute dont_touch of G32907: signal is true;
	signal G32908: std_logic; attribute dont_touch of G32908: signal is true;
	signal G32909: std_logic; attribute dont_touch of G32909: signal is true;
	signal G32910: std_logic; attribute dont_touch of G32910: signal is true;
	signal G32911: std_logic; attribute dont_touch of G32911: signal is true;
	signal G32912: std_logic; attribute dont_touch of G32912: signal is true;
	signal G32913: std_logic; attribute dont_touch of G32913: signal is true;
	signal G32914: std_logic; attribute dont_touch of G32914: signal is true;
	signal G32915: std_logic; attribute dont_touch of G32915: signal is true;
	signal G32916: std_logic; attribute dont_touch of G32916: signal is true;
	signal G32917: std_logic; attribute dont_touch of G32917: signal is true;
	signal G32918: std_logic; attribute dont_touch of G32918: signal is true;
	signal G32919: std_logic; attribute dont_touch of G32919: signal is true;
	signal G32920: std_logic; attribute dont_touch of G32920: signal is true;
	signal G32921: std_logic; attribute dont_touch of G32921: signal is true;
	signal G32922: std_logic; attribute dont_touch of G32922: signal is true;
	signal G32923: std_logic; attribute dont_touch of G32923: signal is true;
	signal G32924: std_logic; attribute dont_touch of G32924: signal is true;
	signal G32925: std_logic; attribute dont_touch of G32925: signal is true;
	signal G32926: std_logic; attribute dont_touch of G32926: signal is true;
	signal G32927: std_logic; attribute dont_touch of G32927: signal is true;
	signal G32928: std_logic; attribute dont_touch of G32928: signal is true;
	signal G32929: std_logic; attribute dont_touch of G32929: signal is true;
	signal G32930: std_logic; attribute dont_touch of G32930: signal is true;
	signal G32931: std_logic; attribute dont_touch of G32931: signal is true;
	signal G32932: std_logic; attribute dont_touch of G32932: signal is true;
	signal G32933: std_logic; attribute dont_touch of G32933: signal is true;
	signal G32934: std_logic; attribute dont_touch of G32934: signal is true;
	signal G32935: std_logic; attribute dont_touch of G32935: signal is true;
	signal G32936: std_logic; attribute dont_touch of G32936: signal is true;
	signal G32937: std_logic; attribute dont_touch of G32937: signal is true;
	signal G32938: std_logic; attribute dont_touch of G32938: signal is true;
	signal G32939: std_logic; attribute dont_touch of G32939: signal is true;
	signal G32940: std_logic; attribute dont_touch of G32940: signal is true;
	signal G32941: std_logic; attribute dont_touch of G32941: signal is true;
	signal G32942: std_logic; attribute dont_touch of G32942: signal is true;
	signal G32943: std_logic; attribute dont_touch of G32943: signal is true;
	signal G32944: std_logic; attribute dont_touch of G32944: signal is true;
	signal G32945: std_logic; attribute dont_touch of G32945: signal is true;
	signal G32946: std_logic; attribute dont_touch of G32946: signal is true;
	signal G32947: std_logic; attribute dont_touch of G32947: signal is true;
	signal G32948: std_logic; attribute dont_touch of G32948: signal is true;
	signal G32949: std_logic; attribute dont_touch of G32949: signal is true;
	signal G32950: std_logic; attribute dont_touch of G32950: signal is true;
	signal G32951: std_logic; attribute dont_touch of G32951: signal is true;
	signal G32952: std_logic; attribute dont_touch of G32952: signal is true;
	signal G32953: std_logic; attribute dont_touch of G32953: signal is true;
	signal G32954: std_logic; attribute dont_touch of G32954: signal is true;
	signal G32955: std_logic; attribute dont_touch of G32955: signal is true;
	signal G32956: std_logic; attribute dont_touch of G32956: signal is true;
	signal G32957: std_logic; attribute dont_touch of G32957: signal is true;
	signal G32958: std_logic; attribute dont_touch of G32958: signal is true;
	signal G32959: std_logic; attribute dont_touch of G32959: signal is true;
	signal G32960: std_logic; attribute dont_touch of G32960: signal is true;
	signal G32961: std_logic; attribute dont_touch of G32961: signal is true;
	signal G32962: std_logic; attribute dont_touch of G32962: signal is true;
	signal G32963: std_logic; attribute dont_touch of G32963: signal is true;
	signal G32964: std_logic; attribute dont_touch of G32964: signal is true;
	signal G32965: std_logic; attribute dont_touch of G32965: signal is true;
	signal G32966: std_logic; attribute dont_touch of G32966: signal is true;
	signal G32967: std_logic; attribute dont_touch of G32967: signal is true;
	signal G32968: std_logic; attribute dont_touch of G32968: signal is true;
	signal G32969: std_logic; attribute dont_touch of G32969: signal is true;
	signal G32970: std_logic; attribute dont_touch of G32970: signal is true;
	signal G32971: std_logic; attribute dont_touch of G32971: signal is true;
	signal G32972: std_logic; attribute dont_touch of G32972: signal is true;
	signal G32973: std_logic; attribute dont_touch of G32973: signal is true;
	signal G32974: std_logic; attribute dont_touch of G32974: signal is true;
	signal G32976: std_logic; attribute dont_touch of G32976: signal is true;
	signal G32977: std_logic; attribute dont_touch of G32977: signal is true;
	signal G32978: std_logic; attribute dont_touch of G32978: signal is true;
	signal G32979: std_logic; attribute dont_touch of G32979: signal is true;
	signal G32980: std_logic; attribute dont_touch of G32980: signal is true;
	signal G32981: std_logic; attribute dont_touch of G32981: signal is true;
	signal G32982: std_logic; attribute dont_touch of G32982: signal is true;
	signal G32983: std_logic; attribute dont_touch of G32983: signal is true;
	signal G32984: std_logic; attribute dont_touch of G32984: signal is true;
	signal G32985: std_logic; attribute dont_touch of G32985: signal is true;
	signal G32986: std_logic; attribute dont_touch of G32986: signal is true;
	signal G32987: std_logic; attribute dont_touch of G32987: signal is true;
	signal G32988: std_logic; attribute dont_touch of G32988: signal is true;
	signal G32989: std_logic; attribute dont_touch of G32989: signal is true;
	signal G32990: std_logic; attribute dont_touch of G32990: signal is true;
	signal G32991: std_logic; attribute dont_touch of G32991: signal is true;
	signal G32992: std_logic; attribute dont_touch of G32992: signal is true;
	signal G32993: std_logic; attribute dont_touch of G32993: signal is true;
	signal G32994: std_logic; attribute dont_touch of G32994: signal is true;
	signal G32995: std_logic; attribute dont_touch of G32995: signal is true;
	signal G32996: std_logic; attribute dont_touch of G32996: signal is true;
	signal G32997: std_logic; attribute dont_touch of G32997: signal is true;
	signal G32998: std_logic; attribute dont_touch of G32998: signal is true;
	signal G32999: std_logic; attribute dont_touch of G32999: signal is true;
	signal G33000: std_logic; attribute dont_touch of G33000: signal is true;
	signal G33001: std_logic; attribute dont_touch of G33001: signal is true;
	signal G33002: std_logic; attribute dont_touch of G33002: signal is true;
	signal G33003: std_logic; attribute dont_touch of G33003: signal is true;
	signal G33004: std_logic; attribute dont_touch of G33004: signal is true;
	signal G33005: std_logic; attribute dont_touch of G33005: signal is true;
	signal G33006: std_logic; attribute dont_touch of G33006: signal is true;
	signal G33007: std_logic; attribute dont_touch of G33007: signal is true;
	signal G33008: std_logic; attribute dont_touch of G33008: signal is true;
	signal G33009: std_logic; attribute dont_touch of G33009: signal is true;
	signal G33010: std_logic; attribute dont_touch of G33010: signal is true;
	signal G33011: std_logic; attribute dont_touch of G33011: signal is true;
	signal G33012: std_logic; attribute dont_touch of G33012: signal is true;
	signal G33013: std_logic; attribute dont_touch of G33013: signal is true;
	signal G33014: std_logic; attribute dont_touch of G33014: signal is true;
	signal G33015: std_logic; attribute dont_touch of G33015: signal is true;
	signal G33016: std_logic; attribute dont_touch of G33016: signal is true;
	signal G33017: std_logic; attribute dont_touch of G33017: signal is true;
	signal G33018: std_logic; attribute dont_touch of G33018: signal is true;
	signal G33019: std_logic; attribute dont_touch of G33019: signal is true;
	signal G33020: std_logic; attribute dont_touch of G33020: signal is true;
	signal G33021: std_logic; attribute dont_touch of G33021: signal is true;
	signal G33022: std_logic; attribute dont_touch of G33022: signal is true;
	signal G33023: std_logic; attribute dont_touch of G33023: signal is true;
	signal G33024: std_logic; attribute dont_touch of G33024: signal is true;
	signal G33025: std_logic; attribute dont_touch of G33025: signal is true;
	signal G33026: std_logic; attribute dont_touch of G33026: signal is true;
	signal G33027: std_logic; attribute dont_touch of G33027: signal is true;
	signal G33028: std_logic; attribute dont_touch of G33028: signal is true;
	signal G33029: std_logic; attribute dont_touch of G33029: signal is true;
	signal G33030: std_logic; attribute dont_touch of G33030: signal is true;
	signal G33031: std_logic; attribute dont_touch of G33031: signal is true;
	signal G33032: std_logic; attribute dont_touch of G33032: signal is true;
	signal G33033: std_logic; attribute dont_touch of G33033: signal is true;
	signal G33034: std_logic; attribute dont_touch of G33034: signal is true;
	signal G33035: std_logic; attribute dont_touch of G33035: signal is true;
	signal G33036: std_logic; attribute dont_touch of G33036: signal is true;
	signal G33037: std_logic; attribute dont_touch of G33037: signal is true;
	signal G33038: std_logic; attribute dont_touch of G33038: signal is true;
	signal G33039: std_logic; attribute dont_touch of G33039: signal is true;
	signal G33040: std_logic; attribute dont_touch of G33040: signal is true;
	signal G33041: std_logic; attribute dont_touch of G33041: signal is true;
	signal G33042: std_logic; attribute dont_touch of G33042: signal is true;
	signal G33043: std_logic; attribute dont_touch of G33043: signal is true;
	signal G33044: std_logic; attribute dont_touch of G33044: signal is true;
	signal G33045: std_logic; attribute dont_touch of G33045: signal is true;
	signal G33046: std_logic; attribute dont_touch of G33046: signal is true;
	signal G33047: std_logic; attribute dont_touch of G33047: signal is true;
	signal G33048: std_logic; attribute dont_touch of G33048: signal is true;
	signal G33049: std_logic; attribute dont_touch of G33049: signal is true;
	signal G33050: std_logic; attribute dont_touch of G33050: signal is true;
	signal G33051: std_logic; attribute dont_touch of G33051: signal is true;
	signal G33052: std_logic; attribute dont_touch of G33052: signal is true;
	signal G33053: std_logic; attribute dont_touch of G33053: signal is true;
	signal G33054: std_logic; attribute dont_touch of G33054: signal is true;
	signal G33055: std_logic; attribute dont_touch of G33055: signal is true;
	signal G33056: std_logic; attribute dont_touch of G33056: signal is true;
	signal G33057: std_logic; attribute dont_touch of G33057: signal is true;
	signal G33058: std_logic; attribute dont_touch of G33058: signal is true;
	signal G33059: std_logic; attribute dont_touch of G33059: signal is true;
	signal G33060: std_logic; attribute dont_touch of G33060: signal is true;
	signal G33061: std_logic; attribute dont_touch of G33061: signal is true;
	signal G33062: std_logic; attribute dont_touch of G33062: signal is true;
	signal G33063: std_logic; attribute dont_touch of G33063: signal is true;
	signal G33064: std_logic; attribute dont_touch of G33064: signal is true;
	signal G33065: std_logic; attribute dont_touch of G33065: signal is true;
	signal G33066: std_logic; attribute dont_touch of G33066: signal is true;
	signal G33067: std_logic; attribute dont_touch of G33067: signal is true;
	signal G33068: std_logic; attribute dont_touch of G33068: signal is true;
	signal G33069: std_logic; attribute dont_touch of G33069: signal is true;
	signal G33070: std_logic; attribute dont_touch of G33070: signal is true;
	signal G33071: std_logic; attribute dont_touch of G33071: signal is true;
	signal G33072: std_logic; attribute dont_touch of G33072: signal is true;
	signal G33073: std_logic; attribute dont_touch of G33073: signal is true;
	signal G33074: std_logic; attribute dont_touch of G33074: signal is true;
	signal G33075: std_logic; attribute dont_touch of G33075: signal is true;
	signal G33076: std_logic; attribute dont_touch of G33076: signal is true;
	signal G33080: std_logic; attribute dont_touch of G33080: signal is true;
	signal G33081: std_logic; attribute dont_touch of G33081: signal is true;
	signal G33082: std_logic; attribute dont_touch of G33082: signal is true;
	signal G33083: std_logic; attribute dont_touch of G33083: signal is true;
	signal G33084: std_logic; attribute dont_touch of G33084: signal is true;
	signal G33085: std_logic; attribute dont_touch of G33085: signal is true;
	signal G33086: std_logic; attribute dont_touch of G33086: signal is true;
	signal G33087: std_logic; attribute dont_touch of G33087: signal is true;
	signal G33088: std_logic; attribute dont_touch of G33088: signal is true;
	signal G33089: std_logic; attribute dont_touch of G33089: signal is true;
	signal G33090: std_logic; attribute dont_touch of G33090: signal is true;
	signal G33091: std_logic; attribute dont_touch of G33091: signal is true;
	signal G33092: std_logic; attribute dont_touch of G33092: signal is true;
	signal G33093: std_logic; attribute dont_touch of G33093: signal is true;
	signal G33094: std_logic; attribute dont_touch of G33094: signal is true;
	signal G33095: std_logic; attribute dont_touch of G33095: signal is true;
	signal G33096: std_logic; attribute dont_touch of G33096: signal is true;
	signal G33097: std_logic; attribute dont_touch of G33097: signal is true;
	signal G33098: std_logic; attribute dont_touch of G33098: signal is true;
	signal G33099: std_logic; attribute dont_touch of G33099: signal is true;
	signal G33100: std_logic; attribute dont_touch of G33100: signal is true;
	signal G33101: std_logic; attribute dont_touch of G33101: signal is true;
	signal G33102: std_logic; attribute dont_touch of G33102: signal is true;
	signal G33103: std_logic; attribute dont_touch of G33103: signal is true;
	signal G33104: std_logic; attribute dont_touch of G33104: signal is true;
	signal G33105: std_logic; attribute dont_touch of G33105: signal is true;
	signal G33106: std_logic; attribute dont_touch of G33106: signal is true;
	signal G33107: std_logic; attribute dont_touch of G33107: signal is true;
	signal G33108: std_logic; attribute dont_touch of G33108: signal is true;
	signal G33109: std_logic; attribute dont_touch of G33109: signal is true;
	signal G33110: std_logic; attribute dont_touch of G33110: signal is true;
	signal G33111: std_logic; attribute dont_touch of G33111: signal is true;
	signal G33112: std_logic; attribute dont_touch of G33112: signal is true;
	signal G33113: std_logic; attribute dont_touch of G33113: signal is true;
	signal G33114: std_logic; attribute dont_touch of G33114: signal is true;
	signal G33115: std_logic; attribute dont_touch of G33115: signal is true;
	signal G33116: std_logic; attribute dont_touch of G33116: signal is true;
	signal G33117: std_logic; attribute dont_touch of G33117: signal is true;
	signal G33118: std_logic; attribute dont_touch of G33118: signal is true;
	signal G33119: std_logic; attribute dont_touch of G33119: signal is true;
	signal G33120: std_logic; attribute dont_touch of G33120: signal is true;
	signal G33121: std_logic; attribute dont_touch of G33121: signal is true;
	signal G33122: std_logic; attribute dont_touch of G33122: signal is true;
	signal G33123: std_logic; attribute dont_touch of G33123: signal is true;
	signal G33124: std_logic; attribute dont_touch of G33124: signal is true;
	signal G33125: std_logic; attribute dont_touch of G33125: signal is true;
	signal G33126: std_logic; attribute dont_touch of G33126: signal is true;
	signal G33127: std_logic; attribute dont_touch of G33127: signal is true;
	signal G33128: std_logic; attribute dont_touch of G33128: signal is true;
	signal G33129: std_logic; attribute dont_touch of G33129: signal is true;
	signal G33130: std_logic; attribute dont_touch of G33130: signal is true;
	signal G33131: std_logic; attribute dont_touch of G33131: signal is true;
	signal G33132: std_logic; attribute dont_touch of G33132: signal is true;
	signal G33133: std_logic; attribute dont_touch of G33133: signal is true;
	signal G33134: std_logic; attribute dont_touch of G33134: signal is true;
	signal G33135: std_logic; attribute dont_touch of G33135: signal is true;
	signal G33136: std_logic; attribute dont_touch of G33136: signal is true;
	signal G33137: std_logic; attribute dont_touch of G33137: signal is true;
	signal G33138: std_logic; attribute dont_touch of G33138: signal is true;
	signal G33139: std_logic; attribute dont_touch of G33139: signal is true;
	signal G33140: std_logic; attribute dont_touch of G33140: signal is true;
	signal G33141: std_logic; attribute dont_touch of G33141: signal is true;
	signal G33142: std_logic; attribute dont_touch of G33142: signal is true;
	signal G33143: std_logic; attribute dont_touch of G33143: signal is true;
	signal G33144: std_logic; attribute dont_touch of G33144: signal is true;
	signal G33145: std_logic; attribute dont_touch of G33145: signal is true;
	signal G33146: std_logic; attribute dont_touch of G33146: signal is true;
	signal G33147: std_logic; attribute dont_touch of G33147: signal is true;
	signal G33148: std_logic; attribute dont_touch of G33148: signal is true;
	signal G33149: std_logic; attribute dont_touch of G33149: signal is true;
	signal G33159: std_logic; attribute dont_touch of G33159: signal is true;
	signal G33160: std_logic; attribute dont_touch of G33160: signal is true;
	signal G33161: std_logic; attribute dont_touch of G33161: signal is true;
	signal G33162: std_logic; attribute dont_touch of G33162: signal is true;
	signal G33163: std_logic; attribute dont_touch of G33163: signal is true;
	signal G33164: std_logic; attribute dont_touch of G33164: signal is true;
	signal G33174: std_logic; attribute dont_touch of G33174: signal is true;
	signal G33175: std_logic; attribute dont_touch of G33175: signal is true;
	signal G33176: std_logic; attribute dont_touch of G33176: signal is true;
	signal G33186: std_logic; attribute dont_touch of G33186: signal is true;
	signal G33187: std_logic; attribute dont_touch of G33187: signal is true;
	signal G33197: std_logic; attribute dont_touch of G33197: signal is true;
	signal G33204: std_logic; attribute dont_touch of G33204: signal is true;
	signal G33212: std_logic; attribute dont_touch of G33212: signal is true;
	signal G33219: std_logic; attribute dont_touch of G33219: signal is true;
	signal G33227: std_logic; attribute dont_touch of G33227: signal is true;
	signal G33228: std_logic; attribute dont_touch of G33228: signal is true;
	signal G33231: std_logic; attribute dont_touch of G33231: signal is true;
	signal G33232: std_logic; attribute dont_touch of G33232: signal is true;
	signal G33233: std_logic; attribute dont_touch of G33233: signal is true;
	signal G33234: std_logic; attribute dont_touch of G33234: signal is true;
	signal G33235: std_logic; attribute dont_touch of G33235: signal is true;
	signal G33236: std_logic; attribute dont_touch of G33236: signal is true;
	signal G33237: std_logic; attribute dont_touch of G33237: signal is true;
	signal G33238: std_logic; attribute dont_touch of G33238: signal is true;
	signal G33239: std_logic; attribute dont_touch of G33239: signal is true;
	signal G33240: std_logic; attribute dont_touch of G33240: signal is true;
	signal G33241: std_logic; attribute dont_touch of G33241: signal is true;
	signal G33242: std_logic; attribute dont_touch of G33242: signal is true;
	signal G33243: std_logic; attribute dont_touch of G33243: signal is true;
	signal G33244: std_logic; attribute dont_touch of G33244: signal is true;
	signal G33245: std_logic; attribute dont_touch of G33245: signal is true;
	signal G33246: std_logic; attribute dont_touch of G33246: signal is true;
	signal G33247: std_logic; attribute dont_touch of G33247: signal is true;
	signal G33248: std_logic; attribute dont_touch of G33248: signal is true;
	signal G33249: std_logic; attribute dont_touch of G33249: signal is true;
	signal G33250: std_logic; attribute dont_touch of G33250: signal is true;
	signal G33251: std_logic; attribute dont_touch of G33251: signal is true;
	signal G33252: std_logic; attribute dont_touch of G33252: signal is true;
	signal G33253: std_logic; attribute dont_touch of G33253: signal is true;
	signal G33254: std_logic; attribute dont_touch of G33254: signal is true;
	signal G33255: std_logic; attribute dont_touch of G33255: signal is true;
	signal G33256: std_logic; attribute dont_touch of G33256: signal is true;
	signal G33257: std_logic; attribute dont_touch of G33257: signal is true;
	signal G33258: std_logic; attribute dont_touch of G33258: signal is true;
	signal G33259: std_logic; attribute dont_touch of G33259: signal is true;
	signal G33260: std_logic; attribute dont_touch of G33260: signal is true;
	signal G33261: std_logic; attribute dont_touch of G33261: signal is true;
	signal G33262: std_logic; attribute dont_touch of G33262: signal is true;
	signal G33263: std_logic; attribute dont_touch of G33263: signal is true;
	signal G33264: std_logic; attribute dont_touch of G33264: signal is true;
	signal G33265: std_logic; attribute dont_touch of G33265: signal is true;
	signal G33266: std_logic; attribute dont_touch of G33266: signal is true;
	signal G33267: std_logic; attribute dont_touch of G33267: signal is true;
	signal G33268: std_logic; attribute dont_touch of G33268: signal is true;
	signal G33269: std_logic; attribute dont_touch of G33269: signal is true;
	signal G33270: std_logic; attribute dont_touch of G33270: signal is true;
	signal G33271: std_logic; attribute dont_touch of G33271: signal is true;
	signal G33272: std_logic; attribute dont_touch of G33272: signal is true;
	signal G33273: std_logic; attribute dont_touch of G33273: signal is true;
	signal G33274: std_logic; attribute dont_touch of G33274: signal is true;
	signal G33275: std_logic; attribute dont_touch of G33275: signal is true;
	signal G33276: std_logic; attribute dont_touch of G33276: signal is true;
	signal G33277: std_logic; attribute dont_touch of G33277: signal is true;
	signal G33278: std_logic; attribute dont_touch of G33278: signal is true;
	signal G33279: std_logic; attribute dont_touch of G33279: signal is true;
	signal G33280: std_logic; attribute dont_touch of G33280: signal is true;
	signal G33281: std_logic; attribute dont_touch of G33281: signal is true;
	signal G33282: std_logic; attribute dont_touch of G33282: signal is true;
	signal G33283: std_logic; attribute dont_touch of G33283: signal is true;
	signal G33286: std_logic; attribute dont_touch of G33286: signal is true;
	signal G33287: std_logic; attribute dont_touch of G33287: signal is true;
	signal G33288: std_logic; attribute dont_touch of G33288: signal is true;
	signal G33289: std_logic; attribute dont_touch of G33289: signal is true;
	signal G33290: std_logic; attribute dont_touch of G33290: signal is true;
	signal G33291: std_logic; attribute dont_touch of G33291: signal is true;
	signal G33292: std_logic; attribute dont_touch of G33292: signal is true;
	signal G33293: std_logic; attribute dont_touch of G33293: signal is true;
	signal G33294: std_logic; attribute dont_touch of G33294: signal is true;
	signal G33295: std_logic; attribute dont_touch of G33295: signal is true;
	signal G33296: std_logic; attribute dont_touch of G33296: signal is true;
	signal G33297: std_logic; attribute dont_touch of G33297: signal is true;
	signal G33298: std_logic; attribute dont_touch of G33298: signal is true;
	signal G33299: std_logic; attribute dont_touch of G33299: signal is true;
	signal G33303: std_logic; attribute dont_touch of G33303: signal is true;
	signal G33304: std_logic; attribute dont_touch of G33304: signal is true;
	signal G33305: std_logic; attribute dont_touch of G33305: signal is true;
	signal G33306: std_logic; attribute dont_touch of G33306: signal is true;
	signal G33310: std_logic; attribute dont_touch of G33310: signal is true;
	signal G33311: std_logic; attribute dont_touch of G33311: signal is true;
	signal G33312: std_logic; attribute dont_touch of G33312: signal is true;
	signal G33313: std_logic; attribute dont_touch of G33313: signal is true;
	signal G33314: std_logic; attribute dont_touch of G33314: signal is true;
	signal G33315: std_logic; attribute dont_touch of G33315: signal is true;
	signal G33316: std_logic; attribute dont_touch of G33316: signal is true;
	signal G33317: std_logic; attribute dont_touch of G33317: signal is true;
	signal G33318: std_logic; attribute dont_touch of G33318: signal is true;
	signal G33321: std_logic; attribute dont_touch of G33321: signal is true;
	signal G33322: std_logic; attribute dont_touch of G33322: signal is true;
	signal G33323: std_logic; attribute dont_touch of G33323: signal is true;
	signal G33326: std_logic; attribute dont_touch of G33326: signal is true;
	signal G33327: std_logic; attribute dont_touch of G33327: signal is true;
	signal G33328: std_logic; attribute dont_touch of G33328: signal is true;
	signal G33329: std_logic; attribute dont_touch of G33329: signal is true;
	signal G33330: std_logic; attribute dont_touch of G33330: signal is true;
	signal G33331: std_logic; attribute dont_touch of G33331: signal is true;
	signal G33332: std_logic; attribute dont_touch of G33332: signal is true;
	signal G33333: std_logic; attribute dont_touch of G33333: signal is true;
	signal G33334: std_logic; attribute dont_touch of G33334: signal is true;
	signal G33335: std_logic; attribute dont_touch of G33335: signal is true;
	signal G33338: std_logic; attribute dont_touch of G33338: signal is true;
	signal G33339: std_logic; attribute dont_touch of G33339: signal is true;
	signal G33340: std_logic; attribute dont_touch of G33340: signal is true;
	signal G33341: std_logic; attribute dont_touch of G33341: signal is true;
	signal G33342: std_logic; attribute dont_touch of G33342: signal is true;
	signal G33343: std_logic; attribute dont_touch of G33343: signal is true;
	signal G33344: std_logic; attribute dont_touch of G33344: signal is true;
	signal G33345: std_logic; attribute dont_touch of G33345: signal is true;
	signal G33346: std_logic; attribute dont_touch of G33346: signal is true;
	signal G33349: std_logic; attribute dont_touch of G33349: signal is true;
	signal G33350: std_logic; attribute dont_touch of G33350: signal is true;
	signal G33351: std_logic; attribute dont_touch of G33351: signal is true;
	signal G33352: std_logic; attribute dont_touch of G33352: signal is true;
	signal G33353: std_logic; attribute dont_touch of G33353: signal is true;
	signal G33354: std_logic; attribute dont_touch of G33354: signal is true;
	signal G33355: std_logic; attribute dont_touch of G33355: signal is true;
	signal G33356: std_logic; attribute dont_touch of G33356: signal is true;
	signal G33357: std_logic; attribute dont_touch of G33357: signal is true;
	signal G33358: std_logic; attribute dont_touch of G33358: signal is true;
	signal G33359: std_logic; attribute dont_touch of G33359: signal is true;
	signal G33360: std_logic; attribute dont_touch of G33360: signal is true;
	signal G33361: std_logic; attribute dont_touch of G33361: signal is true;
	signal G33362: std_logic; attribute dont_touch of G33362: signal is true;
	signal G33363: std_logic; attribute dont_touch of G33363: signal is true;
	signal G33364: std_logic; attribute dont_touch of G33364: signal is true;
	signal G33365: std_logic; attribute dont_touch of G33365: signal is true;
	signal G33366: std_logic; attribute dont_touch of G33366: signal is true;
	signal G33367: std_logic; attribute dont_touch of G33367: signal is true;
	signal G33368: std_logic; attribute dont_touch of G33368: signal is true;
	signal G33369: std_logic; attribute dont_touch of G33369: signal is true;
	signal G33370: std_logic; attribute dont_touch of G33370: signal is true;
	signal G33371: std_logic; attribute dont_touch of G33371: signal is true;
	signal G33372: std_logic; attribute dont_touch of G33372: signal is true;
	signal G33373: std_logic; attribute dont_touch of G33373: signal is true;
	signal G33374: std_logic; attribute dont_touch of G33374: signal is true;
	signal G33375: std_logic; attribute dont_touch of G33375: signal is true;
	signal G33376: std_logic; attribute dont_touch of G33376: signal is true;
	signal G33377: std_logic; attribute dont_touch of G33377: signal is true;
	signal G33378: std_logic; attribute dont_touch of G33378: signal is true;
	signal G33379: std_logic; attribute dont_touch of G33379: signal is true;
	signal G33380: std_logic; attribute dont_touch of G33380: signal is true;
	signal G33381: std_logic; attribute dont_touch of G33381: signal is true;
	signal G33382: std_logic; attribute dont_touch of G33382: signal is true;
	signal G33383: std_logic; attribute dont_touch of G33383: signal is true;
	signal G33384: std_logic; attribute dont_touch of G33384: signal is true;
	signal G33385: std_logic; attribute dont_touch of G33385: signal is true;
	signal G33386: std_logic; attribute dont_touch of G33386: signal is true;
	signal G33387: std_logic; attribute dont_touch of G33387: signal is true;
	signal G33388: std_logic; attribute dont_touch of G33388: signal is true;
	signal G33389: std_logic; attribute dont_touch of G33389: signal is true;
	signal G33390: std_logic; attribute dont_touch of G33390: signal is true;
	signal G33391: std_logic; attribute dont_touch of G33391: signal is true;
	signal G33392: std_logic; attribute dont_touch of G33392: signal is true;
	signal G33393: std_logic; attribute dont_touch of G33393: signal is true;
	signal G33394: std_logic; attribute dont_touch of G33394: signal is true;
	signal G33399: std_logic; attribute dont_touch of G33399: signal is true;
	signal G33400: std_logic; attribute dont_touch of G33400: signal is true;
	signal G33401: std_logic; attribute dont_touch of G33401: signal is true;
	signal G33402: std_logic; attribute dont_touch of G33402: signal is true;
	signal G33403: std_logic; attribute dont_touch of G33403: signal is true;
	signal G33404: std_logic; attribute dont_touch of G33404: signal is true;
	signal G33405: std_logic; attribute dont_touch of G33405: signal is true;
	signal G33406: std_logic; attribute dont_touch of G33406: signal is true;
	signal G33407: std_logic; attribute dont_touch of G33407: signal is true;
	signal G33408: std_logic; attribute dont_touch of G33408: signal is true;
	signal G33409: std_logic; attribute dont_touch of G33409: signal is true;
	signal G33410: std_logic; attribute dont_touch of G33410: signal is true;
	signal G33411: std_logic; attribute dont_touch of G33411: signal is true;
	signal G33412: std_logic; attribute dont_touch of G33412: signal is true;
	signal G33413: std_logic; attribute dont_touch of G33413: signal is true;
	signal G33414: std_logic; attribute dont_touch of G33414: signal is true;
	signal G33415: std_logic; attribute dont_touch of G33415: signal is true;
	signal G33416: std_logic; attribute dont_touch of G33416: signal is true;
	signal G33417: std_logic; attribute dont_touch of G33417: signal is true;
	signal G33418: std_logic; attribute dont_touch of G33418: signal is true;
	signal G33419: std_logic; attribute dont_touch of G33419: signal is true;
	signal G33420: std_logic; attribute dont_touch of G33420: signal is true;
	signal G33421: std_logic; attribute dont_touch of G33421: signal is true;
	signal G33422: std_logic; attribute dont_touch of G33422: signal is true;
	signal G33423: std_logic; attribute dont_touch of G33423: signal is true;
	signal G33424: std_logic; attribute dont_touch of G33424: signal is true;
	signal G33425: std_logic; attribute dont_touch of G33425: signal is true;
	signal G33426: std_logic; attribute dont_touch of G33426: signal is true;
	signal G33427: std_logic; attribute dont_touch of G33427: signal is true;
	signal G33428: std_logic; attribute dont_touch of G33428: signal is true;
	signal G33429: std_logic; attribute dont_touch of G33429: signal is true;
	signal G33430: std_logic; attribute dont_touch of G33430: signal is true;
	signal G33431: std_logic; attribute dont_touch of G33431: signal is true;
	signal G33432: std_logic; attribute dont_touch of G33432: signal is true;
	signal G33433: std_logic; attribute dont_touch of G33433: signal is true;
	signal G33434: std_logic; attribute dont_touch of G33434: signal is true;
	signal G33436: std_logic; attribute dont_touch of G33436: signal is true;
	signal G33437: std_logic; attribute dont_touch of G33437: signal is true;
	signal G33438: std_logic; attribute dont_touch of G33438: signal is true;
	signal G33439: std_logic; attribute dont_touch of G33439: signal is true;
	signal G33440: std_logic; attribute dont_touch of G33440: signal is true;
	signal G33441: std_logic; attribute dont_touch of G33441: signal is true;
	signal G33442: std_logic; attribute dont_touch of G33442: signal is true;
	signal G33443: std_logic; attribute dont_touch of G33443: signal is true;
	signal G33446: std_logic; attribute dont_touch of G33446: signal is true;
	signal G33447: std_logic; attribute dont_touch of G33447: signal is true;
	signal G33448: std_logic; attribute dont_touch of G33448: signal is true;
	signal G33449: std_logic; attribute dont_touch of G33449: signal is true;
	signal G33450: std_logic; attribute dont_touch of G33450: signal is true;
	signal G33451: std_logic; attribute dont_touch of G33451: signal is true;
	signal G33454: std_logic; attribute dont_touch of G33454: signal is true;
	signal G33455: std_logic; attribute dont_touch of G33455: signal is true;
	signal G33456: std_logic; attribute dont_touch of G33456: signal is true;
	signal G33457: std_logic; attribute dont_touch of G33457: signal is true;
	signal G33458: std_logic; attribute dont_touch of G33458: signal is true;
	signal G33459: std_logic; attribute dont_touch of G33459: signal is true;
	signal G33460: std_logic; attribute dont_touch of G33460: signal is true;
	signal G33461: std_logic; attribute dont_touch of G33461: signal is true;
	signal G33462: std_logic; attribute dont_touch of G33462: signal is true;
	signal G33463: std_logic; attribute dont_touch of G33463: signal is true;
	signal G33464: std_logic; attribute dont_touch of G33464: signal is true;
	signal G33465: std_logic; attribute dont_touch of G33465: signal is true;
	signal G33466: std_logic; attribute dont_touch of G33466: signal is true;
	signal G33467: std_logic; attribute dont_touch of G33467: signal is true;
	signal G33468: std_logic; attribute dont_touch of G33468: signal is true;
	signal G33469: std_logic; attribute dont_touch of G33469: signal is true;
	signal G33470: std_logic; attribute dont_touch of G33470: signal is true;
	signal G33471: std_logic; attribute dont_touch of G33471: signal is true;
	signal G33472: std_logic; attribute dont_touch of G33472: signal is true;
	signal G33473: std_logic; attribute dont_touch of G33473: signal is true;
	signal G33474: std_logic; attribute dont_touch of G33474: signal is true;
	signal G33475: std_logic; attribute dont_touch of G33475: signal is true;
	signal G33476: std_logic; attribute dont_touch of G33476: signal is true;
	signal G33477: std_logic; attribute dont_touch of G33477: signal is true;
	signal G33478: std_logic; attribute dont_touch of G33478: signal is true;
	signal G33479: std_logic; attribute dont_touch of G33479: signal is true;
	signal G33480: std_logic; attribute dont_touch of G33480: signal is true;
	signal G33481: std_logic; attribute dont_touch of G33481: signal is true;
	signal G33482: std_logic; attribute dont_touch of G33482: signal is true;
	signal G33483: std_logic; attribute dont_touch of G33483: signal is true;
	signal G33484: std_logic; attribute dont_touch of G33484: signal is true;
	signal G33485: std_logic; attribute dont_touch of G33485: signal is true;
	signal G33486: std_logic; attribute dont_touch of G33486: signal is true;
	signal G33487: std_logic; attribute dont_touch of G33487: signal is true;
	signal G33488: std_logic; attribute dont_touch of G33488: signal is true;
	signal G33489: std_logic; attribute dont_touch of G33489: signal is true;
	signal G33490: std_logic; attribute dont_touch of G33490: signal is true;
	signal G33491: std_logic; attribute dont_touch of G33491: signal is true;
	signal G33492: std_logic; attribute dont_touch of G33492: signal is true;
	signal G33493: std_logic; attribute dont_touch of G33493: signal is true;
	signal G33494: std_logic; attribute dont_touch of G33494: signal is true;
	signal G33495: std_logic; attribute dont_touch of G33495: signal is true;
	signal G33496: std_logic; attribute dont_touch of G33496: signal is true;
	signal G33497: std_logic; attribute dont_touch of G33497: signal is true;
	signal G33498: std_logic; attribute dont_touch of G33498: signal is true;
	signal G33499: std_logic; attribute dont_touch of G33499: signal is true;
	signal G33500: std_logic; attribute dont_touch of G33500: signal is true;
	signal G33501: std_logic; attribute dont_touch of G33501: signal is true;
	signal G33502: std_logic; attribute dont_touch of G33502: signal is true;
	signal G33503: std_logic; attribute dont_touch of G33503: signal is true;
	signal G33504: std_logic; attribute dont_touch of G33504: signal is true;
	signal G33505: std_logic; attribute dont_touch of G33505: signal is true;
	signal G33506: std_logic; attribute dont_touch of G33506: signal is true;
	signal G33507: std_logic; attribute dont_touch of G33507: signal is true;
	signal G33508: std_logic; attribute dont_touch of G33508: signal is true;
	signal G33509: std_logic; attribute dont_touch of G33509: signal is true;
	signal G33510: std_logic; attribute dont_touch of G33510: signal is true;
	signal G33511: std_logic; attribute dont_touch of G33511: signal is true;
	signal G33512: std_logic; attribute dont_touch of G33512: signal is true;
	signal G33513: std_logic; attribute dont_touch of G33513: signal is true;
	signal G33514: std_logic; attribute dont_touch of G33514: signal is true;
	signal G33515: std_logic; attribute dont_touch of G33515: signal is true;
	signal G33516: std_logic; attribute dont_touch of G33516: signal is true;
	signal G33517: std_logic; attribute dont_touch of G33517: signal is true;
	signal G33518: std_logic; attribute dont_touch of G33518: signal is true;
	signal G33519: std_logic; attribute dont_touch of G33519: signal is true;
	signal G33520: std_logic; attribute dont_touch of G33520: signal is true;
	signal G33521: std_logic; attribute dont_touch of G33521: signal is true;
	signal G33522: std_logic; attribute dont_touch of G33522: signal is true;
	signal G33523: std_logic; attribute dont_touch of G33523: signal is true;
	signal G33524: std_logic; attribute dont_touch of G33524: signal is true;
	signal G33525: std_logic; attribute dont_touch of G33525: signal is true;
	signal G33526: std_logic; attribute dont_touch of G33526: signal is true;
	signal G33527: std_logic; attribute dont_touch of G33527: signal is true;
	signal G33528: std_logic; attribute dont_touch of G33528: signal is true;
	signal G33529: std_logic; attribute dont_touch of G33529: signal is true;
	signal G33530: std_logic; attribute dont_touch of G33530: signal is true;
	signal G33531: std_logic; attribute dont_touch of G33531: signal is true;
	signal G33532: std_logic; attribute dont_touch of G33532: signal is true;
	signal G33534: std_logic; attribute dont_touch of G33534: signal is true;
	signal G33535: std_logic; attribute dont_touch of G33535: signal is true;
	signal G33536: std_logic; attribute dont_touch of G33536: signal is true;
	signal G33537: std_logic; attribute dont_touch of G33537: signal is true;
	signal G33538: std_logic; attribute dont_touch of G33538: signal is true;
	signal G33539: std_logic; attribute dont_touch of G33539: signal is true;
	signal G33540: std_logic; attribute dont_touch of G33540: signal is true;
	signal G33541: std_logic; attribute dont_touch of G33541: signal is true;
	signal G33542: std_logic; attribute dont_touch of G33542: signal is true;
	signal G33543: std_logic; attribute dont_touch of G33543: signal is true;
	signal G33544: std_logic; attribute dont_touch of G33544: signal is true;
	signal G33545: std_logic; attribute dont_touch of G33545: signal is true;
	signal G33546: std_logic; attribute dont_touch of G33546: signal is true;
	signal G33547: std_logic; attribute dont_touch of G33547: signal is true;
	signal G33548: std_logic; attribute dont_touch of G33548: signal is true;
	signal G33549: std_logic; attribute dont_touch of G33549: signal is true;
	signal G33550: std_logic; attribute dont_touch of G33550: signal is true;
	signal G33551: std_logic; attribute dont_touch of G33551: signal is true;
	signal G33552: std_logic; attribute dont_touch of G33552: signal is true;
	signal G33553: std_logic; attribute dont_touch of G33553: signal is true;
	signal G33554: std_logic; attribute dont_touch of G33554: signal is true;
	signal G33555: std_logic; attribute dont_touch of G33555: signal is true;
	signal G33556: std_logic; attribute dont_touch of G33556: signal is true;
	signal G33557: std_logic; attribute dont_touch of G33557: signal is true;
	signal G33558: std_logic; attribute dont_touch of G33558: signal is true;
	signal G33559: std_logic; attribute dont_touch of G33559: signal is true;
	signal G33560: std_logic; attribute dont_touch of G33560: signal is true;
	signal G33561: std_logic; attribute dont_touch of G33561: signal is true;
	signal G33562: std_logic; attribute dont_touch of G33562: signal is true;
	signal G33563: std_logic; attribute dont_touch of G33563: signal is true;
	signal G33564: std_logic; attribute dont_touch of G33564: signal is true;
	signal G33565: std_logic; attribute dont_touch of G33565: signal is true;
	signal G33566: std_logic; attribute dont_touch of G33566: signal is true;
	signal G33567: std_logic; attribute dont_touch of G33567: signal is true;
	signal G33568: std_logic; attribute dont_touch of G33568: signal is true;
	signal G33569: std_logic; attribute dont_touch of G33569: signal is true;
	signal G33570: std_logic; attribute dont_touch of G33570: signal is true;
	signal G33571: std_logic; attribute dont_touch of G33571: signal is true;
	signal G33572: std_logic; attribute dont_touch of G33572: signal is true;
	signal G33573: std_logic; attribute dont_touch of G33573: signal is true;
	signal G33574: std_logic; attribute dont_touch of G33574: signal is true;
	signal G33575: std_logic; attribute dont_touch of G33575: signal is true;
	signal G33576: std_logic; attribute dont_touch of G33576: signal is true;
	signal G33577: std_logic; attribute dont_touch of G33577: signal is true;
	signal G33578: std_logic; attribute dont_touch of G33578: signal is true;
	signal G33579: std_logic; attribute dont_touch of G33579: signal is true;
	signal G33580: std_logic; attribute dont_touch of G33580: signal is true;
	signal G33581: std_logic; attribute dont_touch of G33581: signal is true;
	signal G33582: std_logic; attribute dont_touch of G33582: signal is true;
	signal G33583: std_logic; attribute dont_touch of G33583: signal is true;
	signal G33584: std_logic; attribute dont_touch of G33584: signal is true;
	signal G33585: std_logic; attribute dont_touch of G33585: signal is true;
	signal G33586: std_logic; attribute dont_touch of G33586: signal is true;
	signal G33587: std_logic; attribute dont_touch of G33587: signal is true;
	signal G33588: std_logic; attribute dont_touch of G33588: signal is true;
	signal G33589: std_logic; attribute dont_touch of G33589: signal is true;
	signal G33590: std_logic; attribute dont_touch of G33590: signal is true;
	signal G33591: std_logic; attribute dont_touch of G33591: signal is true;
	signal G33592: std_logic; attribute dont_touch of G33592: signal is true;
	signal G33593: std_logic; attribute dont_touch of G33593: signal is true;
	signal G33594: std_logic; attribute dont_touch of G33594: signal is true;
	signal G33595: std_logic; attribute dont_touch of G33595: signal is true;
	signal G33596: std_logic; attribute dont_touch of G33596: signal is true;
	signal G33597: std_logic; attribute dont_touch of G33597: signal is true;
	signal G33598: std_logic; attribute dont_touch of G33598: signal is true;
	signal G33599: std_logic; attribute dont_touch of G33599: signal is true;
	signal G33600: std_logic; attribute dont_touch of G33600: signal is true;
	signal G33601: std_logic; attribute dont_touch of G33601: signal is true;
	signal G33602: std_logic; attribute dont_touch of G33602: signal is true;
	signal G33603: std_logic; attribute dont_touch of G33603: signal is true;
	signal G33604: std_logic; attribute dont_touch of G33604: signal is true;
	signal G33605: std_logic; attribute dont_touch of G33605: signal is true;
	signal G33606: std_logic; attribute dont_touch of G33606: signal is true;
	signal G33607: std_logic; attribute dont_touch of G33607: signal is true;
	signal G33608: std_logic; attribute dont_touch of G33608: signal is true;
	signal G33609: std_logic; attribute dont_touch of G33609: signal is true;
	signal G33610: std_logic; attribute dont_touch of G33610: signal is true;
	signal G33611: std_logic; attribute dont_touch of G33611: signal is true;
	signal G33612: std_logic; attribute dont_touch of G33612: signal is true;
	signal G33613: std_logic; attribute dont_touch of G33613: signal is true;
	signal G33614: std_logic; attribute dont_touch of G33614: signal is true;
	signal G33615: std_logic; attribute dont_touch of G33615: signal is true;
	signal G33616: std_logic; attribute dont_touch of G33616: signal is true;
	signal G33617: std_logic; attribute dont_touch of G33617: signal is true;
	signal G33618: std_logic; attribute dont_touch of G33618: signal is true;
	signal G33619: std_logic; attribute dont_touch of G33619: signal is true;
	signal G33620: std_logic; attribute dont_touch of G33620: signal is true;
	signal G33621: std_logic; attribute dont_touch of G33621: signal is true;
	signal G33622: std_logic; attribute dont_touch of G33622: signal is true;
	signal G33623: std_logic; attribute dont_touch of G33623: signal is true;
	signal G33624: std_logic; attribute dont_touch of G33624: signal is true;
	signal G33625: std_logic; attribute dont_touch of G33625: signal is true;
	signal G33626: std_logic; attribute dont_touch of G33626: signal is true;
	signal G33627: std_logic; attribute dont_touch of G33627: signal is true;
	signal G33628: std_logic; attribute dont_touch of G33628: signal is true;
	signal G33631: std_logic; attribute dont_touch of G33631: signal is true;
	signal G33635: std_logic; attribute dont_touch of G33635: signal is true;
	signal G33637: std_logic; attribute dont_touch of G33637: signal is true;
	signal G33638: std_logic; attribute dont_touch of G33638: signal is true;
	signal G33639: std_logic; attribute dont_touch of G33639: signal is true;
	signal G33640: std_logic; attribute dont_touch of G33640: signal is true;
	signal G33641: std_logic; attribute dont_touch of G33641: signal is true;
	signal G33645: std_logic; attribute dont_touch of G33645: signal is true;
	signal G33646: std_logic; attribute dont_touch of G33646: signal is true;
	signal G33647: std_logic; attribute dont_touch of G33647: signal is true;
	signal G33648: std_logic; attribute dont_touch of G33648: signal is true;
	signal G33652: std_logic; attribute dont_touch of G33652: signal is true;
	signal G33653: std_logic; attribute dont_touch of G33653: signal is true;
	signal G33657: std_logic; attribute dont_touch of G33657: signal is true;
	signal G33658: std_logic; attribute dont_touch of G33658: signal is true;
	signal G33660: std_logic; attribute dont_touch of G33660: signal is true;
	signal G33661: std_logic; attribute dont_touch of G33661: signal is true;
	signal G33665: std_logic; attribute dont_touch of G33665: signal is true;
	signal G33669: std_logic; attribute dont_touch of G33669: signal is true;
	signal G33670: std_logic; attribute dont_touch of G33670: signal is true;
	signal G33674: std_logic; attribute dont_touch of G33674: signal is true;
	signal G33675: std_logic; attribute dont_touch of G33675: signal is true;
	signal G33676: std_logic; attribute dont_touch of G33676: signal is true;
	signal G33677: std_logic; attribute dont_touch of G33677: signal is true;
	signal G33678: std_logic; attribute dont_touch of G33678: signal is true;
	signal G33679: std_logic; attribute dont_touch of G33679: signal is true;
	signal G33680: std_logic; attribute dont_touch of G33680: signal is true;
	signal G33681: std_logic; attribute dont_touch of G33681: signal is true;
	signal G33682: std_logic; attribute dont_touch of G33682: signal is true;
	signal G33683: std_logic; attribute dont_touch of G33683: signal is true;
	signal G33684: std_logic; attribute dont_touch of G33684: signal is true;
	signal G33685: std_logic; attribute dont_touch of G33685: signal is true;
	signal G33686: std_logic; attribute dont_touch of G33686: signal is true;
	signal G33687: std_logic; attribute dont_touch of G33687: signal is true;
	signal G33688: std_logic; attribute dont_touch of G33688: signal is true;
	signal G33689: std_logic; attribute dont_touch of G33689: signal is true;
	signal G33690: std_logic; attribute dont_touch of G33690: signal is true;
	signal G33691: std_logic; attribute dont_touch of G33691: signal is true;
	signal G33692: std_logic; attribute dont_touch of G33692: signal is true;
	signal G33693: std_logic; attribute dont_touch of G33693: signal is true;
	signal G33694: std_logic; attribute dont_touch of G33694: signal is true;
	signal G33695: std_logic; attribute dont_touch of G33695: signal is true;
	signal G33696: std_logic; attribute dont_touch of G33696: signal is true;
	signal G33697: std_logic; attribute dont_touch of G33697: signal is true;
	signal G33698: std_logic; attribute dont_touch of G33698: signal is true;
	signal G33699: std_logic; attribute dont_touch of G33699: signal is true;
	signal G33700: std_logic; attribute dont_touch of G33700: signal is true;
	signal G33701: std_logic; attribute dont_touch of G33701: signal is true;
	signal G33702: std_logic; attribute dont_touch of G33702: signal is true;
	signal G33703: std_logic; attribute dont_touch of G33703: signal is true;
	signal G33704: std_logic; attribute dont_touch of G33704: signal is true;
	signal G33705: std_logic; attribute dont_touch of G33705: signal is true;
	signal G33706: std_logic; attribute dont_touch of G33706: signal is true;
	signal G33707: std_logic; attribute dont_touch of G33707: signal is true;
	signal G33708: std_logic; attribute dont_touch of G33708: signal is true;
	signal G33709: std_logic; attribute dont_touch of G33709: signal is true;
	signal G33710: std_logic; attribute dont_touch of G33710: signal is true;
	signal G33711: std_logic; attribute dont_touch of G33711: signal is true;
	signal G33712: std_logic; attribute dont_touch of G33712: signal is true;
	signal G33713: std_logic; attribute dont_touch of G33713: signal is true;
	signal G33714: std_logic; attribute dont_touch of G33714: signal is true;
	signal G33715: std_logic; attribute dont_touch of G33715: signal is true;
	signal G33716: std_logic; attribute dont_touch of G33716: signal is true;
	signal G33717: std_logic; attribute dont_touch of G33717: signal is true;
	signal G33718: std_logic; attribute dont_touch of G33718: signal is true;
	signal G33719: std_logic; attribute dont_touch of G33719: signal is true;
	signal G33720: std_logic; attribute dont_touch of G33720: signal is true;
	signal G33721: std_logic; attribute dont_touch of G33721: signal is true;
	signal G33722: std_logic; attribute dont_touch of G33722: signal is true;
	signal G33723: std_logic; attribute dont_touch of G33723: signal is true;
	signal G33724: std_logic; attribute dont_touch of G33724: signal is true;
	signal G33725: std_logic; attribute dont_touch of G33725: signal is true;
	signal G33726: std_logic; attribute dont_touch of G33726: signal is true;
	signal G33727: std_logic; attribute dont_touch of G33727: signal is true;
	signal G33728: std_logic; attribute dont_touch of G33728: signal is true;
	signal G33729: std_logic; attribute dont_touch of G33729: signal is true;
	signal G33730: std_logic; attribute dont_touch of G33730: signal is true;
	signal G33731: std_logic; attribute dont_touch of G33731: signal is true;
	signal G33732: std_logic; attribute dont_touch of G33732: signal is true;
	signal G33733: std_logic; attribute dont_touch of G33733: signal is true;
	signal G33734: std_logic; attribute dont_touch of G33734: signal is true;
	signal G33735: std_logic; attribute dont_touch of G33735: signal is true;
	signal G33736: std_logic; attribute dont_touch of G33736: signal is true;
	signal G33742: std_logic; attribute dont_touch of G33742: signal is true;
	signal G33743: std_logic; attribute dont_touch of G33743: signal is true;
	signal G33744: std_logic; attribute dont_touch of G33744: signal is true;
	signal G33750: std_logic; attribute dont_touch of G33750: signal is true;
	signal G33755: std_logic; attribute dont_touch of G33755: signal is true;
	signal G33758: std_logic; attribute dont_touch of G33758: signal is true;
	signal G33759: std_logic; attribute dont_touch of G33759: signal is true;
	signal G33760: std_logic; attribute dont_touch of G33760: signal is true;
	signal G33761: std_logic; attribute dont_touch of G33761: signal is true;
	signal G33766: std_logic; attribute dont_touch of G33766: signal is true;
	signal G33772: std_logic; attribute dont_touch of G33772: signal is true;
	signal G33778: std_logic; attribute dont_touch of G33778: signal is true;
	signal G33784: std_logic; attribute dont_touch of G33784: signal is true;
	signal G33785: std_logic; attribute dont_touch of G33785: signal is true;
	signal G33786: std_logic; attribute dont_touch of G33786: signal is true;
	signal G33787: std_logic; attribute dont_touch of G33787: signal is true;
	signal G33788: std_logic; attribute dont_touch of G33788: signal is true;
	signal G33789: std_logic; attribute dont_touch of G33789: signal is true;
	signal G33790: std_logic; attribute dont_touch of G33790: signal is true;
	signal G33791: std_logic; attribute dont_touch of G33791: signal is true;
	signal G33794: std_logic; attribute dont_touch of G33794: signal is true;
	signal G33795: std_logic; attribute dont_touch of G33795: signal is true;
	signal G33796: std_logic; attribute dont_touch of G33796: signal is true;
	signal G33797: std_logic; attribute dont_touch of G33797: signal is true;
	signal G33798: std_logic; attribute dont_touch of G33798: signal is true;
	signal G33799: std_logic; attribute dont_touch of G33799: signal is true;
	signal G33800: std_logic; attribute dont_touch of G33800: signal is true;
	signal G33801: std_logic; attribute dont_touch of G33801: signal is true;
	signal G33802: std_logic; attribute dont_touch of G33802: signal is true;
	signal G33803: std_logic; attribute dont_touch of G33803: signal is true;
	signal G33804: std_logic; attribute dont_touch of G33804: signal is true;
	signal G33805: std_logic; attribute dont_touch of G33805: signal is true;
	signal G33806: std_logic; attribute dont_touch of G33806: signal is true;
	signal G33807: std_logic; attribute dont_touch of G33807: signal is true;
	signal G33808: std_logic; attribute dont_touch of G33808: signal is true;
	signal G33809: std_logic; attribute dont_touch of G33809: signal is true;
	signal G33810: std_logic; attribute dont_touch of G33810: signal is true;
	signal G33811: std_logic; attribute dont_touch of G33811: signal is true;
	signal G33812: std_logic; attribute dont_touch of G33812: signal is true;
	signal G33813: std_logic; attribute dont_touch of G33813: signal is true;
	signal G33814: std_logic; attribute dont_touch of G33814: signal is true;
	signal G33815: std_logic; attribute dont_touch of G33815: signal is true;
	signal G33816: std_logic; attribute dont_touch of G33816: signal is true;
	signal G33817: std_logic; attribute dont_touch of G33817: signal is true;
	signal G33818: std_logic; attribute dont_touch of G33818: signal is true;
	signal G33819: std_logic; attribute dont_touch of G33819: signal is true;
	signal G33820: std_logic; attribute dont_touch of G33820: signal is true;
	signal G33821: std_logic; attribute dont_touch of G33821: signal is true;
	signal G33822: std_logic; attribute dont_touch of G33822: signal is true;
	signal G33823: std_logic; attribute dont_touch of G33823: signal is true;
	signal G33827: std_logic; attribute dont_touch of G33827: signal is true;
	signal G33828: std_logic; attribute dont_touch of G33828: signal is true;
	signal G33829: std_logic; attribute dont_touch of G33829: signal is true;
	signal G33830: std_logic; attribute dont_touch of G33830: signal is true;
	signal G33831: std_logic; attribute dont_touch of G33831: signal is true;
	signal G33832: std_logic; attribute dont_touch of G33832: signal is true;
	signal G33833: std_logic; attribute dont_touch of G33833: signal is true;
	signal G33834: std_logic; attribute dont_touch of G33834: signal is true;
	signal G33835: std_logic; attribute dont_touch of G33835: signal is true;
	signal G33836: std_logic; attribute dont_touch of G33836: signal is true;
	signal G33837: std_logic; attribute dont_touch of G33837: signal is true;
	signal G33838: std_logic; attribute dont_touch of G33838: signal is true;
	signal G33839: std_logic; attribute dont_touch of G33839: signal is true;
	signal G33840: std_logic; attribute dont_touch of G33840: signal is true;
	signal G33841: std_logic; attribute dont_touch of G33841: signal is true;
	signal G33842: std_logic; attribute dont_touch of G33842: signal is true;
	signal G33843: std_logic; attribute dont_touch of G33843: signal is true;
	signal G33844: std_logic; attribute dont_touch of G33844: signal is true;
	signal G33845: std_logic; attribute dont_touch of G33845: signal is true;
	signal G33846: std_logic; attribute dont_touch of G33846: signal is true;
	signal G33847: std_logic; attribute dont_touch of G33847: signal is true;
	signal G33848: std_logic; attribute dont_touch of G33848: signal is true;
	signal G33849: std_logic; attribute dont_touch of G33849: signal is true;
	signal G33850: std_logic; attribute dont_touch of G33850: signal is true;
	signal G33851: std_logic; attribute dont_touch of G33851: signal is true;
	signal G33855: std_logic; attribute dont_touch of G33855: signal is true;
	signal G33856: std_logic; attribute dont_touch of G33856: signal is true;
	signal G33857: std_logic; attribute dont_touch of G33857: signal is true;
	signal G33858: std_logic; attribute dont_touch of G33858: signal is true;
	signal G33859: std_logic; attribute dont_touch of G33859: signal is true;
	signal G33860: std_logic; attribute dont_touch of G33860: signal is true;
	signal G33861: std_logic; attribute dont_touch of G33861: signal is true;
	signal G33862: std_logic; attribute dont_touch of G33862: signal is true;
	signal G33863: std_logic; attribute dont_touch of G33863: signal is true;
	signal G33864: std_logic; attribute dont_touch of G33864: signal is true;
	signal G33865: std_logic; attribute dont_touch of G33865: signal is true;
	signal G33866: std_logic; attribute dont_touch of G33866: signal is true;
	signal G33867: std_logic; attribute dont_touch of G33867: signal is true;
	signal G33868: std_logic; attribute dont_touch of G33868: signal is true;
	signal G33869: std_logic; attribute dont_touch of G33869: signal is true;
	signal G33870: std_logic; attribute dont_touch of G33870: signal is true;
	signal G33871: std_logic; attribute dont_touch of G33871: signal is true;
	signal G33872: std_logic; attribute dont_touch of G33872: signal is true;
	signal G33873: std_logic; attribute dont_touch of G33873: signal is true;
	signal G33875: std_logic; attribute dont_touch of G33875: signal is true;
	signal G33876: std_logic; attribute dont_touch of G33876: signal is true;
	signal G33877: std_logic; attribute dont_touch of G33877: signal is true;
	signal G33878: std_logic; attribute dont_touch of G33878: signal is true;
	signal G33879: std_logic; attribute dont_touch of G33879: signal is true;
	signal G33880: std_logic; attribute dont_touch of G33880: signal is true;
	signal G33881: std_logic; attribute dont_touch of G33881: signal is true;
	signal G33882: std_logic; attribute dont_touch of G33882: signal is true;
	signal G33883: std_logic; attribute dont_touch of G33883: signal is true;
	signal G33884: std_logic; attribute dont_touch of G33884: signal is true;
	signal G33885: std_logic; attribute dont_touch of G33885: signal is true;
	signal G33886: std_logic; attribute dont_touch of G33886: signal is true;
	signal G33887: std_logic; attribute dont_touch of G33887: signal is true;
	signal G33888: std_logic; attribute dont_touch of G33888: signal is true;
	signal G33889: std_logic; attribute dont_touch of G33889: signal is true;
	signal G33890: std_logic; attribute dont_touch of G33890: signal is true;
	signal G33891: std_logic; attribute dont_touch of G33891: signal is true;
	signal G33892: std_logic; attribute dont_touch of G33892: signal is true;
	signal G33893: std_logic; attribute dont_touch of G33893: signal is true;
	signal G33895: std_logic; attribute dont_touch of G33895: signal is true;
	signal G33896: std_logic; attribute dont_touch of G33896: signal is true;
	signal G33897: std_logic; attribute dont_touch of G33897: signal is true;
	signal G33898: std_logic; attribute dont_touch of G33898: signal is true;
	signal G33899: std_logic; attribute dont_touch of G33899: signal is true;
	signal G33900: std_logic; attribute dont_touch of G33900: signal is true;
	signal G33901: std_logic; attribute dont_touch of G33901: signal is true;
	signal G33902: std_logic; attribute dont_touch of G33902: signal is true;
	signal G33903: std_logic; attribute dont_touch of G33903: signal is true;
	signal G33904: std_logic; attribute dont_touch of G33904: signal is true;
	signal G33905: std_logic; attribute dont_touch of G33905: signal is true;
	signal G33906: std_logic; attribute dont_touch of G33906: signal is true;
	signal G33907: std_logic; attribute dont_touch of G33907: signal is true;
	signal G33908: std_logic; attribute dont_touch of G33908: signal is true;
	signal G33909: std_logic; attribute dont_touch of G33909: signal is true;
	signal G33910: std_logic; attribute dont_touch of G33910: signal is true;
	signal G33911: std_logic; attribute dont_touch of G33911: signal is true;
	signal G33912: std_logic; attribute dont_touch of G33912: signal is true;
	signal G33913: std_logic; attribute dont_touch of G33913: signal is true;
	signal G33914: std_logic; attribute dont_touch of G33914: signal is true;
	signal G33915: std_logic; attribute dont_touch of G33915: signal is true;
	signal G33916: std_logic; attribute dont_touch of G33916: signal is true;
	signal G33917: std_logic; attribute dont_touch of G33917: signal is true;
	signal G33918: std_logic; attribute dont_touch of G33918: signal is true;
	signal G33919: std_logic; attribute dont_touch of G33919: signal is true;
	signal G33920: std_logic; attribute dont_touch of G33920: signal is true;
	signal G33921: std_logic; attribute dont_touch of G33921: signal is true;
	signal G33922: std_logic; attribute dont_touch of G33922: signal is true;
	signal G33923: std_logic; attribute dont_touch of G33923: signal is true;
	signal G33924: std_logic; attribute dont_touch of G33924: signal is true;
	signal G33925: std_logic; attribute dont_touch of G33925: signal is true;
	signal G33926: std_logic; attribute dont_touch of G33926: signal is true;
	signal G33927: std_logic; attribute dont_touch of G33927: signal is true;
	signal G33928: std_logic; attribute dont_touch of G33928: signal is true;
	signal G33929: std_logic; attribute dont_touch of G33929: signal is true;
	signal G33930: std_logic; attribute dont_touch of G33930: signal is true;
	signal G33931: std_logic; attribute dont_touch of G33931: signal is true;
	signal G33932: std_logic; attribute dont_touch of G33932: signal is true;
	signal G33933: std_logic; attribute dont_touch of G33933: signal is true;
	signal G33934: std_logic; attribute dont_touch of G33934: signal is true;
	signal G33936: std_logic; attribute dont_touch of G33936: signal is true;
	signal G33937: std_logic; attribute dont_touch of G33937: signal is true;
	signal G33941: std_logic; attribute dont_touch of G33941: signal is true;
	signal G33942: std_logic; attribute dont_touch of G33942: signal is true;
	signal G33943: std_logic; attribute dont_touch of G33943: signal is true;
	signal G33944: std_logic; attribute dont_touch of G33944: signal is true;
	signal G33951: std_logic; attribute dont_touch of G33951: signal is true;
	signal G33952: std_logic; attribute dont_touch of G33952: signal is true;
	signal G33953: std_logic; attribute dont_touch of G33953: signal is true;
	signal G33954: std_logic; attribute dont_touch of G33954: signal is true;
	signal G33955: std_logic; attribute dont_touch of G33955: signal is true;
	signal G33956: std_logic; attribute dont_touch of G33956: signal is true;
	signal G33957: std_logic; attribute dont_touch of G33957: signal is true;
	signal G33958: std_logic; attribute dont_touch of G33958: signal is true;
	signal G33960: std_logic; attribute dont_touch of G33960: signal is true;
	signal G33961: std_logic; attribute dont_touch of G33961: signal is true;
	signal G33962: std_logic; attribute dont_touch of G33962: signal is true;
	signal G33963: std_logic; attribute dont_touch of G33963: signal is true;
	signal G33964: std_logic; attribute dont_touch of G33964: signal is true;
	signal G33965: std_logic; attribute dont_touch of G33965: signal is true;
	signal G33966: std_logic; attribute dont_touch of G33966: signal is true;
	signal G33967: std_logic; attribute dont_touch of G33967: signal is true;
	signal G33968: std_logic; attribute dont_touch of G33968: signal is true;
	signal G33969: std_logic; attribute dont_touch of G33969: signal is true;
	signal G33970: std_logic; attribute dont_touch of G33970: signal is true;
	signal G33971: std_logic; attribute dont_touch of G33971: signal is true;
	signal G33972: std_logic; attribute dont_touch of G33972: signal is true;
	signal G33973: std_logic; attribute dont_touch of G33973: signal is true;
	signal G33974: std_logic; attribute dont_touch of G33974: signal is true;
	signal G33975: std_logic; attribute dont_touch of G33975: signal is true;
	signal G33976: std_logic; attribute dont_touch of G33976: signal is true;
	signal G33977: std_logic; attribute dont_touch of G33977: signal is true;
	signal G33978: std_logic; attribute dont_touch of G33978: signal is true;
	signal G33979: std_logic; attribute dont_touch of G33979: signal is true;
	signal G33980: std_logic; attribute dont_touch of G33980: signal is true;
	signal G33981: std_logic; attribute dont_touch of G33981: signal is true;
	signal G33982: std_logic; attribute dont_touch of G33982: signal is true;
	signal G33983: std_logic; attribute dont_touch of G33983: signal is true;
	signal G33984: std_logic; attribute dont_touch of G33984: signal is true;
	signal G33985: std_logic; attribute dont_touch of G33985: signal is true;
	signal G33986: std_logic; attribute dont_touch of G33986: signal is true;
	signal G33987: std_logic; attribute dont_touch of G33987: signal is true;
	signal G33988: std_logic; attribute dont_touch of G33988: signal is true;
	signal G33989: std_logic; attribute dont_touch of G33989: signal is true;
	signal G33990: std_logic; attribute dont_touch of G33990: signal is true;
	signal G33991: std_logic; attribute dont_touch of G33991: signal is true;
	signal G33992: std_logic; attribute dont_touch of G33992: signal is true;
	signal G33993: std_logic; attribute dont_touch of G33993: signal is true;
	signal G33994: std_logic; attribute dont_touch of G33994: signal is true;
	signal G33995: std_logic; attribute dont_touch of G33995: signal is true;
	signal G33996: std_logic; attribute dont_touch of G33996: signal is true;
	signal G33997: std_logic; attribute dont_touch of G33997: signal is true;
	signal G33998: std_logic; attribute dont_touch of G33998: signal is true;
	signal G33999: std_logic; attribute dont_touch of G33999: signal is true;
	signal G34000: std_logic; attribute dont_touch of G34000: signal is true;
	signal G34001: std_logic; attribute dont_touch of G34001: signal is true;
	signal G34002: std_logic; attribute dont_touch of G34002: signal is true;
	signal G34003: std_logic; attribute dont_touch of G34003: signal is true;
	signal G34004: std_logic; attribute dont_touch of G34004: signal is true;
	signal G34005: std_logic; attribute dont_touch of G34005: signal is true;
	signal G34006: std_logic; attribute dont_touch of G34006: signal is true;
	signal G34007: std_logic; attribute dont_touch of G34007: signal is true;
	signal G34008: std_logic; attribute dont_touch of G34008: signal is true;
	signal G34009: std_logic; attribute dont_touch of G34009: signal is true;
	signal G34010: std_logic; attribute dont_touch of G34010: signal is true;
	signal G34011: std_logic; attribute dont_touch of G34011: signal is true;
	signal G34012: std_logic; attribute dont_touch of G34012: signal is true;
	signal G34013: std_logic; attribute dont_touch of G34013: signal is true;
	signal G34014: std_logic; attribute dont_touch of G34014: signal is true;
	signal G34015: std_logic; attribute dont_touch of G34015: signal is true;
	signal G34016: std_logic; attribute dont_touch of G34016: signal is true;
	signal G34017: std_logic; attribute dont_touch of G34017: signal is true;
	signal G34018: std_logic; attribute dont_touch of G34018: signal is true;
	signal G34019: std_logic; attribute dont_touch of G34019: signal is true;
	signal G34020: std_logic; attribute dont_touch of G34020: signal is true;
	signal G34021: std_logic; attribute dont_touch of G34021: signal is true;
	signal G34022: std_logic; attribute dont_touch of G34022: signal is true;
	signal G34023: std_logic; attribute dont_touch of G34023: signal is true;
	signal G34024: std_logic; attribute dont_touch of G34024: signal is true;
	signal G34025: std_logic; attribute dont_touch of G34025: signal is true;
	signal G34026: std_logic; attribute dont_touch of G34026: signal is true;
	signal G34027: std_logic; attribute dont_touch of G34027: signal is true;
	signal G34028: std_logic; attribute dont_touch of G34028: signal is true;
	signal G34029: std_logic; attribute dont_touch of G34029: signal is true;
	signal G34030: std_logic; attribute dont_touch of G34030: signal is true;
	signal G34031: std_logic; attribute dont_touch of G34031: signal is true;
	signal G34032: std_logic; attribute dont_touch of G34032: signal is true;
	signal G34033: std_logic; attribute dont_touch of G34033: signal is true;
	signal G34034: std_logic; attribute dont_touch of G34034: signal is true;
	signal G34035: std_logic; attribute dont_touch of G34035: signal is true;
	signal G34036: std_logic; attribute dont_touch of G34036: signal is true;
	signal G34037: std_logic; attribute dont_touch of G34037: signal is true;
	signal G34038: std_logic; attribute dont_touch of G34038: signal is true;
	signal G34039: std_logic; attribute dont_touch of G34039: signal is true;
	signal G34040: std_logic; attribute dont_touch of G34040: signal is true;
	signal G34041: std_logic; attribute dont_touch of G34041: signal is true;
	signal G34042: std_logic; attribute dont_touch of G34042: signal is true;
	signal G34043: std_logic; attribute dont_touch of G34043: signal is true;
	signal G34044: std_logic; attribute dont_touch of G34044: signal is true;
	signal G34045: std_logic; attribute dont_touch of G34045: signal is true;
	signal G34046: std_logic; attribute dont_touch of G34046: signal is true;
	signal G34047: std_logic; attribute dont_touch of G34047: signal is true;
	signal G34048: std_logic; attribute dont_touch of G34048: signal is true;
	signal G34049: std_logic; attribute dont_touch of G34049: signal is true;
	signal G34050: std_logic; attribute dont_touch of G34050: signal is true;
	signal G34051: std_logic; attribute dont_touch of G34051: signal is true;
	signal G34052: std_logic; attribute dont_touch of G34052: signal is true;
	signal G34053: std_logic; attribute dont_touch of G34053: signal is true;
	signal G34054: std_logic; attribute dont_touch of G34054: signal is true;
	signal G34055: std_logic; attribute dont_touch of G34055: signal is true;
	signal G34056: std_logic; attribute dont_touch of G34056: signal is true;
	signal G34057: std_logic; attribute dont_touch of G34057: signal is true;
	signal G34058: std_logic; attribute dont_touch of G34058: signal is true;
	signal G34059: std_logic; attribute dont_touch of G34059: signal is true;
	signal G34060: std_logic; attribute dont_touch of G34060: signal is true;
	signal G34061: std_logic; attribute dont_touch of G34061: signal is true;
	signal G34062: std_logic; attribute dont_touch of G34062: signal is true;
	signal G34063: std_logic; attribute dont_touch of G34063: signal is true;
	signal G34064: std_logic; attribute dont_touch of G34064: signal is true;
	signal G34065: std_logic; attribute dont_touch of G34065: signal is true;
	signal G34066: std_logic; attribute dont_touch of G34066: signal is true;
	signal G34067: std_logic; attribute dont_touch of G34067: signal is true;
	signal G34068: std_logic; attribute dont_touch of G34068: signal is true;
	signal G34069: std_logic; attribute dont_touch of G34069: signal is true;
	signal G34070: std_logic; attribute dont_touch of G34070: signal is true;
	signal G34071: std_logic; attribute dont_touch of G34071: signal is true;
	signal G34072: std_logic; attribute dont_touch of G34072: signal is true;
	signal G34073: std_logic; attribute dont_touch of G34073: signal is true;
	signal G34074: std_logic; attribute dont_touch of G34074: signal is true;
	signal G34075: std_logic; attribute dont_touch of G34075: signal is true;
	signal G34076: std_logic; attribute dont_touch of G34076: signal is true;
	signal G34077: std_logic; attribute dont_touch of G34077: signal is true;
	signal G34078: std_logic; attribute dont_touch of G34078: signal is true;
	signal G34079: std_logic; attribute dont_touch of G34079: signal is true;
	signal G34080: std_logic; attribute dont_touch of G34080: signal is true;
	signal G34081: std_logic; attribute dont_touch of G34081: signal is true;
	signal G34082: std_logic; attribute dont_touch of G34082: signal is true;
	signal G34083: std_logic; attribute dont_touch of G34083: signal is true;
	signal G34084: std_logic; attribute dont_touch of G34084: signal is true;
	signal G34085: std_logic; attribute dont_touch of G34085: signal is true;
	signal G34086: std_logic; attribute dont_touch of G34086: signal is true;
	signal G34087: std_logic; attribute dont_touch of G34087: signal is true;
	signal G34088: std_logic; attribute dont_touch of G34088: signal is true;
	signal G34089: std_logic; attribute dont_touch of G34089: signal is true;
	signal G34090: std_logic; attribute dont_touch of G34090: signal is true;
	signal G34091: std_logic; attribute dont_touch of G34091: signal is true;
	signal G34092: std_logic; attribute dont_touch of G34092: signal is true;
	signal G34093: std_logic; attribute dont_touch of G34093: signal is true;
	signal G34094: std_logic; attribute dont_touch of G34094: signal is true;
	signal G34095: std_logic; attribute dont_touch of G34095: signal is true;
	signal G34096: std_logic; attribute dont_touch of G34096: signal is true;
	signal G34097: std_logic; attribute dont_touch of G34097: signal is true;
	signal G34098: std_logic; attribute dont_touch of G34098: signal is true;
	signal G34099: std_logic; attribute dont_touch of G34099: signal is true;
	signal G34100: std_logic; attribute dont_touch of G34100: signal is true;
	signal G34101: std_logic; attribute dont_touch of G34101: signal is true;
	signal G34102: std_logic; attribute dont_touch of G34102: signal is true;
	signal G34103: std_logic; attribute dont_touch of G34103: signal is true;
	signal G34104: std_logic; attribute dont_touch of G34104: signal is true;
	signal G34105: std_logic; attribute dont_touch of G34105: signal is true;
	signal G34106: std_logic; attribute dont_touch of G34106: signal is true;
	signal G34107: std_logic; attribute dont_touch of G34107: signal is true;
	signal G34108: std_logic; attribute dont_touch of G34108: signal is true;
	signal G34109: std_logic; attribute dont_touch of G34109: signal is true;
	signal G34110: std_logic; attribute dont_touch of G34110: signal is true;
	signal G34111: std_logic; attribute dont_touch of G34111: signal is true;
	signal G34112: std_logic; attribute dont_touch of G34112: signal is true;
	signal G34113: std_logic; attribute dont_touch of G34113: signal is true;
	signal G34114: std_logic; attribute dont_touch of G34114: signal is true;
	signal G34115: std_logic; attribute dont_touch of G34115: signal is true;
	signal G34116: std_logic; attribute dont_touch of G34116: signal is true;
	signal G34117: std_logic; attribute dont_touch of G34117: signal is true;
	signal G34118: std_logic; attribute dont_touch of G34118: signal is true;
	signal G34119: std_logic; attribute dont_touch of G34119: signal is true;
	signal G34120: std_logic; attribute dont_touch of G34120: signal is true;
	signal G34121: std_logic; attribute dont_touch of G34121: signal is true;
	signal G34122: std_logic; attribute dont_touch of G34122: signal is true;
	signal G34123: std_logic; attribute dont_touch of G34123: signal is true;
	signal G34124: std_logic; attribute dont_touch of G34124: signal is true;
	signal G34125: std_logic; attribute dont_touch of G34125: signal is true;
	signal G34126: std_logic; attribute dont_touch of G34126: signal is true;
	signal G34127: std_logic; attribute dont_touch of G34127: signal is true;
	signal G34130: std_logic; attribute dont_touch of G34130: signal is true;
	signal G34131: std_logic; attribute dont_touch of G34131: signal is true;
	signal G34132: std_logic; attribute dont_touch of G34132: signal is true;
	signal G34133: std_logic; attribute dont_touch of G34133: signal is true;
	signal G34134: std_logic; attribute dont_touch of G34134: signal is true;
	signal G34135: std_logic; attribute dont_touch of G34135: signal is true;
	signal G34136: std_logic; attribute dont_touch of G34136: signal is true;
	signal G34137: std_logic; attribute dont_touch of G34137: signal is true;
	signal G34138: std_logic; attribute dont_touch of G34138: signal is true;
	signal G34139: std_logic; attribute dont_touch of G34139: signal is true;
	signal G34140: std_logic; attribute dont_touch of G34140: signal is true;
	signal G34141: std_logic; attribute dont_touch of G34141: signal is true;
	signal G34142: std_logic; attribute dont_touch of G34142: signal is true;
	signal G34143: std_logic; attribute dont_touch of G34143: signal is true;
	signal G34144: std_logic; attribute dont_touch of G34144: signal is true;
	signal G34145: std_logic; attribute dont_touch of G34145: signal is true;
	signal G34146: std_logic; attribute dont_touch of G34146: signal is true;
	signal G34147: std_logic; attribute dont_touch of G34147: signal is true;
	signal G34148: std_logic; attribute dont_touch of G34148: signal is true;
	signal G34149: std_logic; attribute dont_touch of G34149: signal is true;
	signal G34150: std_logic; attribute dont_touch of G34150: signal is true;
	signal G34151: std_logic; attribute dont_touch of G34151: signal is true;
	signal G34152: std_logic; attribute dont_touch of G34152: signal is true;
	signal G34153: std_logic; attribute dont_touch of G34153: signal is true;
	signal G34156: std_logic; attribute dont_touch of G34156: signal is true;
	signal G34157: std_logic; attribute dont_touch of G34157: signal is true;
	signal G34158: std_logic; attribute dont_touch of G34158: signal is true;
	signal G34159: std_logic; attribute dont_touch of G34159: signal is true;
	signal G34160: std_logic; attribute dont_touch of G34160: signal is true;
	signal G34161: std_logic; attribute dont_touch of G34161: signal is true;
	signal G34162: std_logic; attribute dont_touch of G34162: signal is true;
	signal G34166: std_logic; attribute dont_touch of G34166: signal is true;
	signal G34167: std_logic; attribute dont_touch of G34167: signal is true;
	signal G34168: std_logic; attribute dont_touch of G34168: signal is true;
	signal G34169: std_logic; attribute dont_touch of G34169: signal is true;
	signal G34170: std_logic; attribute dont_touch of G34170: signal is true;
	signal G34171: std_logic; attribute dont_touch of G34171: signal is true;
	signal G34172: std_logic; attribute dont_touch of G34172: signal is true;
	signal G34173: std_logic; attribute dont_touch of G34173: signal is true;
	signal G34174: std_logic; attribute dont_touch of G34174: signal is true;
	signal G34178: std_logic; attribute dont_touch of G34178: signal is true;
	signal G34179: std_logic; attribute dont_touch of G34179: signal is true;
	signal G34180: std_logic; attribute dont_touch of G34180: signal is true;
	signal G34181: std_logic; attribute dont_touch of G34181: signal is true;
	signal G34182: std_logic; attribute dont_touch of G34182: signal is true;
	signal G34183: std_logic; attribute dont_touch of G34183: signal is true;
	signal G34184: std_logic; attribute dont_touch of G34184: signal is true;
	signal G34185: std_logic; attribute dont_touch of G34185: signal is true;
	signal G34186: std_logic; attribute dont_touch of G34186: signal is true;
	signal G34187: std_logic; attribute dont_touch of G34187: signal is true;
	signal G34188: std_logic; attribute dont_touch of G34188: signal is true;
	signal G34189: std_logic; attribute dont_touch of G34189: signal is true;
	signal G34190: std_logic; attribute dont_touch of G34190: signal is true;
	signal G34191: std_logic; attribute dont_touch of G34191: signal is true;
	signal G34192: std_logic; attribute dont_touch of G34192: signal is true;
	signal G34193: std_logic; attribute dont_touch of G34193: signal is true;
	signal G34194: std_logic; attribute dont_touch of G34194: signal is true;
	signal G34195: std_logic; attribute dont_touch of G34195: signal is true;
	signal G34196: std_logic; attribute dont_touch of G34196: signal is true;
	signal G34197: std_logic; attribute dont_touch of G34197: signal is true;
	signal G34198: std_logic; attribute dont_touch of G34198: signal is true;
	signal G34199: std_logic; attribute dont_touch of G34199: signal is true;
	signal G34200: std_logic; attribute dont_touch of G34200: signal is true;
	signal G34202: std_logic; attribute dont_touch of G34202: signal is true;
	signal G34203: std_logic; attribute dont_touch of G34203: signal is true;
	signal G34204: std_logic; attribute dont_touch of G34204: signal is true;
	signal G34205: std_logic; attribute dont_touch of G34205: signal is true;
	signal G34206: std_logic; attribute dont_touch of G34206: signal is true;
	signal G34207: std_logic; attribute dont_touch of G34207: signal is true;
	signal G34208: std_logic; attribute dont_touch of G34208: signal is true;
	signal G34209: std_logic; attribute dont_touch of G34209: signal is true;
	signal G34210: std_logic; attribute dont_touch of G34210: signal is true;
	signal G34211: std_logic; attribute dont_touch of G34211: signal is true;
	signal G34212: std_logic; attribute dont_touch of G34212: signal is true;
	signal G34213: std_logic; attribute dont_touch of G34213: signal is true;
	signal G34214: std_logic; attribute dont_touch of G34214: signal is true;
	signal G34215: std_logic; attribute dont_touch of G34215: signal is true;
	signal G34216: std_logic; attribute dont_touch of G34216: signal is true;
	signal G34217: std_logic; attribute dont_touch of G34217: signal is true;
	signal G34218: std_logic; attribute dont_touch of G34218: signal is true;
	signal G34219: std_logic; attribute dont_touch of G34219: signal is true;
	signal G34220: std_logic; attribute dont_touch of G34220: signal is true;
	signal G34222: std_logic; attribute dont_touch of G34222: signal is true;
	signal G34223: std_logic; attribute dont_touch of G34223: signal is true;
	signal G34224: std_logic; attribute dont_touch of G34224: signal is true;
	signal G34225: std_logic; attribute dont_touch of G34225: signal is true;
	signal G34226: std_logic; attribute dont_touch of G34226: signal is true;
	signal G34227: std_logic; attribute dont_touch of G34227: signal is true;
	signal G34228: std_logic; attribute dont_touch of G34228: signal is true;
	signal G34229: std_logic; attribute dont_touch of G34229: signal is true;
	signal G34230: std_logic; attribute dont_touch of G34230: signal is true;
	signal G34231: std_logic; attribute dont_touch of G34231: signal is true;
	signal G34241: std_logic; attribute dont_touch of G34241: signal is true;
	signal G34242: std_logic; attribute dont_touch of G34242: signal is true;
	signal G34243: std_logic; attribute dont_touch of G34243: signal is true;
	signal G34244: std_logic; attribute dont_touch of G34244: signal is true;
	signal G34245: std_logic; attribute dont_touch of G34245: signal is true;
	signal G34246: std_logic; attribute dont_touch of G34246: signal is true;
	signal G34247: std_logic; attribute dont_touch of G34247: signal is true;
	signal G34248: std_logic; attribute dont_touch of G34248: signal is true;
	signal G34249: std_logic; attribute dont_touch of G34249: signal is true;
	signal G34250: std_logic; attribute dont_touch of G34250: signal is true;
	signal G34251: std_logic; attribute dont_touch of G34251: signal is true;
	signal G34252: std_logic; attribute dont_touch of G34252: signal is true;
	signal G34253: std_logic; attribute dont_touch of G34253: signal is true;
	signal G34254: std_logic; attribute dont_touch of G34254: signal is true;
	signal G34255: std_logic; attribute dont_touch of G34255: signal is true;
	signal G34256: std_logic; attribute dont_touch of G34256: signal is true;
	signal G34257: std_logic; attribute dont_touch of G34257: signal is true;
	signal G34258: std_logic; attribute dont_touch of G34258: signal is true;
	signal G34259: std_logic; attribute dont_touch of G34259: signal is true;
	signal G34260: std_logic; attribute dont_touch of G34260: signal is true;
	signal G34261: std_logic; attribute dont_touch of G34261: signal is true;
	signal G34262: std_logic; attribute dont_touch of G34262: signal is true;
	signal G34263: std_logic; attribute dont_touch of G34263: signal is true;
	signal G34264: std_logic; attribute dont_touch of G34264: signal is true;
	signal G34265: std_logic; attribute dont_touch of G34265: signal is true;
	signal G34266: std_logic; attribute dont_touch of G34266: signal is true;
	signal G34267: std_logic; attribute dont_touch of G34267: signal is true;
	signal G34268: std_logic; attribute dont_touch of G34268: signal is true;
	signal G34269: std_logic; attribute dont_touch of G34269: signal is true;
	signal G34270: std_logic; attribute dont_touch of G34270: signal is true;
	signal G34271: std_logic; attribute dont_touch of G34271: signal is true;
	signal G34272: std_logic; attribute dont_touch of G34272: signal is true;
	signal G34273: std_logic; attribute dont_touch of G34273: signal is true;
	signal G34274: std_logic; attribute dont_touch of G34274: signal is true;
	signal G34275: std_logic; attribute dont_touch of G34275: signal is true;
	signal G34276: std_logic; attribute dont_touch of G34276: signal is true;
	signal G34277: std_logic; attribute dont_touch of G34277: signal is true;
	signal G34278: std_logic; attribute dont_touch of G34278: signal is true;
	signal G34279: std_logic; attribute dont_touch of G34279: signal is true;
	signal G34280: std_logic; attribute dont_touch of G34280: signal is true;
	signal G34281: std_logic; attribute dont_touch of G34281: signal is true;
	signal G34282: std_logic; attribute dont_touch of G34282: signal is true;
	signal G34283: std_logic; attribute dont_touch of G34283: signal is true;
	signal G34284: std_logic; attribute dont_touch of G34284: signal is true;
	signal G34285: std_logic; attribute dont_touch of G34285: signal is true;
	signal G34286: std_logic; attribute dont_touch of G34286: signal is true;
	signal G34287: std_logic; attribute dont_touch of G34287: signal is true;
	signal G34288: std_logic; attribute dont_touch of G34288: signal is true;
	signal G34289: std_logic; attribute dont_touch of G34289: signal is true;
	signal G34290: std_logic; attribute dont_touch of G34290: signal is true;
	signal G34291: std_logic; attribute dont_touch of G34291: signal is true;
	signal G34292: std_logic; attribute dont_touch of G34292: signal is true;
	signal G34293: std_logic; attribute dont_touch of G34293: signal is true;
	signal G34294: std_logic; attribute dont_touch of G34294: signal is true;
	signal G34295: std_logic; attribute dont_touch of G34295: signal is true;
	signal G34296: std_logic; attribute dont_touch of G34296: signal is true;
	signal G34297: std_logic; attribute dont_touch of G34297: signal is true;
	signal G34298: std_logic; attribute dont_touch of G34298: signal is true;
	signal G34299: std_logic; attribute dont_touch of G34299: signal is true;
	signal G34300: std_logic; attribute dont_touch of G34300: signal is true;
	signal G34301: std_logic; attribute dont_touch of G34301: signal is true;
	signal G34302: std_logic; attribute dont_touch of G34302: signal is true;
	signal G34303: std_logic; attribute dont_touch of G34303: signal is true;
	signal G34304: std_logic; attribute dont_touch of G34304: signal is true;
	signal G34305: std_logic; attribute dont_touch of G34305: signal is true;
	signal G34306: std_logic; attribute dont_touch of G34306: signal is true;
	signal G34307: std_logic; attribute dont_touch of G34307: signal is true;
	signal G34308: std_logic; attribute dont_touch of G34308: signal is true;
	signal G34309: std_logic; attribute dont_touch of G34309: signal is true;
	signal G34310: std_logic; attribute dont_touch of G34310: signal is true;
	signal G34311: std_logic; attribute dont_touch of G34311: signal is true;
	signal G34312: std_logic; attribute dont_touch of G34312: signal is true;
	signal G34313: std_logic; attribute dont_touch of G34313: signal is true;
	signal G34314: std_logic; attribute dont_touch of G34314: signal is true;
	signal G34315: std_logic; attribute dont_touch of G34315: signal is true;
	signal G34316: std_logic; attribute dont_touch of G34316: signal is true;
	signal G34317: std_logic; attribute dont_touch of G34317: signal is true;
	signal G34318: std_logic; attribute dont_touch of G34318: signal is true;
	signal G34319: std_logic; attribute dont_touch of G34319: signal is true;
	signal G34320: std_logic; attribute dont_touch of G34320: signal is true;
	signal G34321: std_logic; attribute dont_touch of G34321: signal is true;
	signal G34322: std_logic; attribute dont_touch of G34322: signal is true;
	signal G34323: std_logic; attribute dont_touch of G34323: signal is true;
	signal G34324: std_logic; attribute dont_touch of G34324: signal is true;
	signal G34325: std_logic; attribute dont_touch of G34325: signal is true;
	signal G34326: std_logic; attribute dont_touch of G34326: signal is true;
	signal G34327: std_logic; attribute dont_touch of G34327: signal is true;
	signal G34328: std_logic; attribute dont_touch of G34328: signal is true;
	signal G34329: std_logic; attribute dont_touch of G34329: signal is true;
	signal G34330: std_logic; attribute dont_touch of G34330: signal is true;
	signal G34331: std_logic; attribute dont_touch of G34331: signal is true;
	signal G34332: std_logic; attribute dont_touch of G34332: signal is true;
	signal G34333: std_logic; attribute dont_touch of G34333: signal is true;
	signal G34334: std_logic; attribute dont_touch of G34334: signal is true;
	signal G34335: std_logic; attribute dont_touch of G34335: signal is true;
	signal G34336: std_logic; attribute dont_touch of G34336: signal is true;
	signal G34337: std_logic; attribute dont_touch of G34337: signal is true;
	signal G34338: std_logic; attribute dont_touch of G34338: signal is true;
	signal G34339: std_logic; attribute dont_touch of G34339: signal is true;
	signal G34340: std_logic; attribute dont_touch of G34340: signal is true;
	signal G34341: std_logic; attribute dont_touch of G34341: signal is true;
	signal G34342: std_logic; attribute dont_touch of G34342: signal is true;
	signal G34343: std_logic; attribute dont_touch of G34343: signal is true;
	signal G34344: std_logic; attribute dont_touch of G34344: signal is true;
	signal G34345: std_logic; attribute dont_touch of G34345: signal is true;
	signal G34346: std_logic; attribute dont_touch of G34346: signal is true;
	signal G34347: std_logic; attribute dont_touch of G34347: signal is true;
	signal G34348: std_logic; attribute dont_touch of G34348: signal is true;
	signal G34349: std_logic; attribute dont_touch of G34349: signal is true;
	signal G34350: std_logic; attribute dont_touch of G34350: signal is true;
	signal G34351: std_logic; attribute dont_touch of G34351: signal is true;
	signal G34352: std_logic; attribute dont_touch of G34352: signal is true;
	signal G34353: std_logic; attribute dont_touch of G34353: signal is true;
	signal G34354: std_logic; attribute dont_touch of G34354: signal is true;
	signal G34358: std_logic; attribute dont_touch of G34358: signal is true;
	signal G34359: std_logic; attribute dont_touch of G34359: signal is true;
	signal G34363: std_logic; attribute dont_touch of G34363: signal is true;
	signal G34364: std_logic; attribute dont_touch of G34364: signal is true;
	signal G34365: std_logic; attribute dont_touch of G34365: signal is true;
	signal G34366: std_logic; attribute dont_touch of G34366: signal is true;
	signal G34367: std_logic; attribute dont_touch of G34367: signal is true;
	signal G34368: std_logic; attribute dont_touch of G34368: signal is true;
	signal G34369: std_logic; attribute dont_touch of G34369: signal is true;
	signal G34370: std_logic; attribute dont_touch of G34370: signal is true;
	signal G34371: std_logic; attribute dont_touch of G34371: signal is true;
	signal G34372: std_logic; attribute dont_touch of G34372: signal is true;
	signal G34373: std_logic; attribute dont_touch of G34373: signal is true;
	signal G34374: std_logic; attribute dont_touch of G34374: signal is true;
	signal G34375: std_logic; attribute dont_touch of G34375: signal is true;
	signal G34376: std_logic; attribute dont_touch of G34376: signal is true;
	signal G34377: std_logic; attribute dont_touch of G34377: signal is true;
	signal G34378: std_logic; attribute dont_touch of G34378: signal is true;
	signal G34379: std_logic; attribute dont_touch of G34379: signal is true;
	signal G34380: std_logic; attribute dont_touch of G34380: signal is true;
	signal G34381: std_logic; attribute dont_touch of G34381: signal is true;
	signal G34382: std_logic; attribute dont_touch of G34382: signal is true;
	signal G34384: std_logic; attribute dont_touch of G34384: signal is true;
	signal G34385: std_logic; attribute dont_touch of G34385: signal is true;
	signal G34386: std_logic; attribute dont_touch of G34386: signal is true;
	signal G34387: std_logic; attribute dont_touch of G34387: signal is true;
	signal G34388: std_logic; attribute dont_touch of G34388: signal is true;
	signal G34389: std_logic; attribute dont_touch of G34389: signal is true;
	signal G34390: std_logic; attribute dont_touch of G34390: signal is true;
	signal G34391: std_logic; attribute dont_touch of G34391: signal is true;
	signal G34392: std_logic; attribute dont_touch of G34392: signal is true;
	signal G34393: std_logic; attribute dont_touch of G34393: signal is true;
	signal G34394: std_logic; attribute dont_touch of G34394: signal is true;
	signal G34395: std_logic; attribute dont_touch of G34395: signal is true;
	signal G34396: std_logic; attribute dont_touch of G34396: signal is true;
	signal G34397: std_logic; attribute dont_touch of G34397: signal is true;
	signal G34398: std_logic; attribute dont_touch of G34398: signal is true;
	signal G34399: std_logic; attribute dont_touch of G34399: signal is true;
	signal G34400: std_logic; attribute dont_touch of G34400: signal is true;
	signal G34401: std_logic; attribute dont_touch of G34401: signal is true;
	signal G34402: std_logic; attribute dont_touch of G34402: signal is true;
	signal G34403: std_logic; attribute dont_touch of G34403: signal is true;
	signal G34404: std_logic; attribute dont_touch of G34404: signal is true;
	signal G34405: std_logic; attribute dont_touch of G34405: signal is true;
	signal G34406: std_logic; attribute dont_touch of G34406: signal is true;
	signal G34407: std_logic; attribute dont_touch of G34407: signal is true;
	signal G34408: std_logic; attribute dont_touch of G34408: signal is true;
	signal G34409: std_logic; attribute dont_touch of G34409: signal is true;
	signal G34410: std_logic; attribute dont_touch of G34410: signal is true;
	signal G34411: std_logic; attribute dont_touch of G34411: signal is true;
	signal G34412: std_logic; attribute dont_touch of G34412: signal is true;
	signal G34413: std_logic; attribute dont_touch of G34413: signal is true;
	signal G34414: std_logic; attribute dont_touch of G34414: signal is true;
	signal G34415: std_logic; attribute dont_touch of G34415: signal is true;
	signal G34416: std_logic; attribute dont_touch of G34416: signal is true;
	signal G34417: std_logic; attribute dont_touch of G34417: signal is true;
	signal G34418: std_logic; attribute dont_touch of G34418: signal is true;
	signal G34419: std_logic; attribute dont_touch of G34419: signal is true;
	signal G34420: std_logic; attribute dont_touch of G34420: signal is true;
	signal G34421: std_logic; attribute dont_touch of G34421: signal is true;
	signal G34422: std_logic; attribute dont_touch of G34422: signal is true;
	signal G34423: std_logic; attribute dont_touch of G34423: signal is true;
	signal G34424: std_logic; attribute dont_touch of G34424: signal is true;
	signal G34426: std_logic; attribute dont_touch of G34426: signal is true;
	signal G34427: std_logic; attribute dont_touch of G34427: signal is true;
	signal G34428: std_logic; attribute dont_touch of G34428: signal is true;
	signal G34429: std_logic; attribute dont_touch of G34429: signal is true;
	signal G34430: std_logic; attribute dont_touch of G34430: signal is true;
	signal G34431: std_logic; attribute dont_touch of G34431: signal is true;
	signal G34432: std_logic; attribute dont_touch of G34432: signal is true;
	signal G34433: std_logic; attribute dont_touch of G34433: signal is true;
	signal G34434: std_logic; attribute dont_touch of G34434: signal is true;
	signal G34438: std_logic; attribute dont_touch of G34438: signal is true;
	signal G34439: std_logic; attribute dont_touch of G34439: signal is true;
	signal G34440: std_logic; attribute dont_touch of G34440: signal is true;
	signal G34441: std_logic; attribute dont_touch of G34441: signal is true;
	signal G34442: std_logic; attribute dont_touch of G34442: signal is true;
	signal G34443: std_logic; attribute dont_touch of G34443: signal is true;
	signal G34444: std_logic; attribute dont_touch of G34444: signal is true;
	signal G34445: std_logic; attribute dont_touch of G34445: signal is true;
	signal G34446: std_logic; attribute dont_touch of G34446: signal is true;
	signal G34447: std_logic; attribute dont_touch of G34447: signal is true;
	signal G34448: std_logic; attribute dont_touch of G34448: signal is true;
	signal G34449: std_logic; attribute dont_touch of G34449: signal is true;
	signal G34450: std_logic; attribute dont_touch of G34450: signal is true;
	signal G34451: std_logic; attribute dont_touch of G34451: signal is true;
	signal G34452: std_logic; attribute dont_touch of G34452: signal is true;
	signal G34453: std_logic; attribute dont_touch of G34453: signal is true;
	signal G34454: std_logic; attribute dont_touch of G34454: signal is true;
	signal G34455: std_logic; attribute dont_touch of G34455: signal is true;
	signal G34456: std_logic; attribute dont_touch of G34456: signal is true;
	signal G34457: std_logic; attribute dont_touch of G34457: signal is true;
	signal G34458: std_logic; attribute dont_touch of G34458: signal is true;
	signal G34459: std_logic; attribute dont_touch of G34459: signal is true;
	signal G34460: std_logic; attribute dont_touch of G34460: signal is true;
	signal G34461: std_logic; attribute dont_touch of G34461: signal is true;
	signal G34462: std_logic; attribute dont_touch of G34462: signal is true;
	signal G34463: std_logic; attribute dont_touch of G34463: signal is true;
	signal G34464: std_logic; attribute dont_touch of G34464: signal is true;
	signal G34465: std_logic; attribute dont_touch of G34465: signal is true;
	signal G34466: std_logic; attribute dont_touch of G34466: signal is true;
	signal G34467: std_logic; attribute dont_touch of G34467: signal is true;
	signal G34468: std_logic; attribute dont_touch of G34468: signal is true;
	signal G34469: std_logic; attribute dont_touch of G34469: signal is true;
	signal G34470: std_logic; attribute dont_touch of G34470: signal is true;
	signal G34471: std_logic; attribute dont_touch of G34471: signal is true;
	signal G34472: std_logic; attribute dont_touch of G34472: signal is true;
	signal G34473: std_logic; attribute dont_touch of G34473: signal is true;
	signal G34474: std_logic; attribute dont_touch of G34474: signal is true;
	signal G34475: std_logic; attribute dont_touch of G34475: signal is true;
	signal G34476: std_logic; attribute dont_touch of G34476: signal is true;
	signal G34477: std_logic; attribute dont_touch of G34477: signal is true;
	signal G34478: std_logic; attribute dont_touch of G34478: signal is true;
	signal G34479: std_logic; attribute dont_touch of G34479: signal is true;
	signal G34480: std_logic; attribute dont_touch of G34480: signal is true;
	signal G34481: std_logic; attribute dont_touch of G34481: signal is true;
	signal G34482: std_logic; attribute dont_touch of G34482: signal is true;
	signal G34483: std_logic; attribute dont_touch of G34483: signal is true;
	signal G34484: std_logic; attribute dont_touch of G34484: signal is true;
	signal G34485: std_logic; attribute dont_touch of G34485: signal is true;
	signal G34486: std_logic; attribute dont_touch of G34486: signal is true;
	signal G34487: std_logic; attribute dont_touch of G34487: signal is true;
	signal G34488: std_logic; attribute dont_touch of G34488: signal is true;
	signal G34489: std_logic; attribute dont_touch of G34489: signal is true;
	signal G34490: std_logic; attribute dont_touch of G34490: signal is true;
	signal G34491: std_logic; attribute dont_touch of G34491: signal is true;
	signal G34492: std_logic; attribute dont_touch of G34492: signal is true;
	signal G34493: std_logic; attribute dont_touch of G34493: signal is true;
	signal G34494: std_logic; attribute dont_touch of G34494: signal is true;
	signal G34495: std_logic; attribute dont_touch of G34495: signal is true;
	signal G34496: std_logic; attribute dont_touch of G34496: signal is true;
	signal G34497: std_logic; attribute dont_touch of G34497: signal is true;
	signal G34498: std_logic; attribute dont_touch of G34498: signal is true;
	signal G34499: std_logic; attribute dont_touch of G34499: signal is true;
	signal G34500: std_logic; attribute dont_touch of G34500: signal is true;
	signal G34501: std_logic; attribute dont_touch of G34501: signal is true;
	signal G34502: std_logic; attribute dont_touch of G34502: signal is true;
	signal G34503: std_logic; attribute dont_touch of G34503: signal is true;
	signal G34504: std_logic; attribute dont_touch of G34504: signal is true;
	signal G34505: std_logic; attribute dont_touch of G34505: signal is true;
	signal G34506: std_logic; attribute dont_touch of G34506: signal is true;
	signal G34507: std_logic; attribute dont_touch of G34507: signal is true;
	signal G34508: std_logic; attribute dont_touch of G34508: signal is true;
	signal G34509: std_logic; attribute dont_touch of G34509: signal is true;
	signal G34510: std_logic; attribute dont_touch of G34510: signal is true;
	signal G34511: std_logic; attribute dont_touch of G34511: signal is true;
	signal G34512: std_logic; attribute dont_touch of G34512: signal is true;
	signal G34513: std_logic; attribute dont_touch of G34513: signal is true;
	signal G34514: std_logic; attribute dont_touch of G34514: signal is true;
	signal G34515: std_logic; attribute dont_touch of G34515: signal is true;
	signal G34516: std_logic; attribute dont_touch of G34516: signal is true;
	signal G34517: std_logic; attribute dont_touch of G34517: signal is true;
	signal G34518: std_logic; attribute dont_touch of G34518: signal is true;
	signal G34519: std_logic; attribute dont_touch of G34519: signal is true;
	signal G34520: std_logic; attribute dont_touch of G34520: signal is true;
	signal G34521: std_logic; attribute dont_touch of G34521: signal is true;
	signal G34522: std_logic; attribute dont_touch of G34522: signal is true;
	signal G34523: std_logic; attribute dont_touch of G34523: signal is true;
	signal G34524: std_logic; attribute dont_touch of G34524: signal is true;
	signal G34525: std_logic; attribute dont_touch of G34525: signal is true;
	signal G34526: std_logic; attribute dont_touch of G34526: signal is true;
	signal G34527: std_logic; attribute dont_touch of G34527: signal is true;
	signal G34528: std_logic; attribute dont_touch of G34528: signal is true;
	signal G34529: std_logic; attribute dont_touch of G34529: signal is true;
	signal G34530: std_logic; attribute dont_touch of G34530: signal is true;
	signal G34531: std_logic; attribute dont_touch of G34531: signal is true;
	signal G34532: std_logic; attribute dont_touch of G34532: signal is true;
	signal G34533: std_logic; attribute dont_touch of G34533: signal is true;
	signal G34534: std_logic; attribute dont_touch of G34534: signal is true;
	signal G34535: std_logic; attribute dont_touch of G34535: signal is true;
	signal G34536: std_logic; attribute dont_touch of G34536: signal is true;
	signal G34537: std_logic; attribute dont_touch of G34537: signal is true;
	signal G34538: std_logic; attribute dont_touch of G34538: signal is true;
	signal G34539: std_logic; attribute dont_touch of G34539: signal is true;
	signal G34540: std_logic; attribute dont_touch of G34540: signal is true;
	signal G34541: std_logic; attribute dont_touch of G34541: signal is true;
	signal G34542: std_logic; attribute dont_touch of G34542: signal is true;
	signal G34543: std_logic; attribute dont_touch of G34543: signal is true;
	signal G34544: std_logic; attribute dont_touch of G34544: signal is true;
	signal G34545: std_logic; attribute dont_touch of G34545: signal is true;
	signal G34549: std_logic; attribute dont_touch of G34549: signal is true;
	signal G34550: std_logic; attribute dont_touch of G34550: signal is true;
	signal G34553: std_logic; attribute dont_touch of G34553: signal is true;
	signal G34554: std_logic; attribute dont_touch of G34554: signal is true;
	signal G34555: std_logic; attribute dont_touch of G34555: signal is true;
	signal G34556: std_logic; attribute dont_touch of G34556: signal is true;
	signal G34557: std_logic; attribute dont_touch of G34557: signal is true;
	signal G34558: std_logic; attribute dont_touch of G34558: signal is true;
	signal G34559: std_logic; attribute dont_touch of G34559: signal is true;
	signal G34560: std_logic; attribute dont_touch of G34560: signal is true;
	signal G34561: std_logic; attribute dont_touch of G34561: signal is true;
	signal G34562: std_logic; attribute dont_touch of G34562: signal is true;
	signal G34563: std_logic; attribute dont_touch of G34563: signal is true;
	signal G34564: std_logic; attribute dont_touch of G34564: signal is true;
	signal G34565: std_logic; attribute dont_touch of G34565: signal is true;
	signal G34566: std_logic; attribute dont_touch of G34566: signal is true;
	signal G34567: std_logic; attribute dont_touch of G34567: signal is true;
	signal G34568: std_logic; attribute dont_touch of G34568: signal is true;
	signal G34569: std_logic; attribute dont_touch of G34569: signal is true;
	signal G34570: std_logic; attribute dont_touch of G34570: signal is true;
	signal G34571: std_logic; attribute dont_touch of G34571: signal is true;
	signal G34572: std_logic; attribute dont_touch of G34572: signal is true;
	signal G34573: std_logic; attribute dont_touch of G34573: signal is true;
	signal G34574: std_logic; attribute dont_touch of G34574: signal is true;
	signal G34575: std_logic; attribute dont_touch of G34575: signal is true;
	signal G34576: std_logic; attribute dont_touch of G34576: signal is true;
	signal G34577: std_logic; attribute dont_touch of G34577: signal is true;
	signal G34578: std_logic; attribute dont_touch of G34578: signal is true;
	signal G34579: std_logic; attribute dont_touch of G34579: signal is true;
	signal G34580: std_logic; attribute dont_touch of G34580: signal is true;
	signal G34581: std_logic; attribute dont_touch of G34581: signal is true;
	signal G34582: std_logic; attribute dont_touch of G34582: signal is true;
	signal G34583: std_logic; attribute dont_touch of G34583: signal is true;
	signal G34584: std_logic; attribute dont_touch of G34584: signal is true;
	signal G34585: std_logic; attribute dont_touch of G34585: signal is true;
	signal G34586: std_logic; attribute dont_touch of G34586: signal is true;
	signal G34587: std_logic; attribute dont_touch of G34587: signal is true;
	signal G34588: std_logic; attribute dont_touch of G34588: signal is true;
	signal G34589: std_logic; attribute dont_touch of G34589: signal is true;
	signal G34590: std_logic; attribute dont_touch of G34590: signal is true;
	signal G34591: std_logic; attribute dont_touch of G34591: signal is true;
	signal G34592: std_logic; attribute dont_touch of G34592: signal is true;
	signal G34593: std_logic; attribute dont_touch of G34593: signal is true;
	signal G34594: std_logic; attribute dont_touch of G34594: signal is true;
	signal G34595: std_logic; attribute dont_touch of G34595: signal is true;
	signal G34596: std_logic; attribute dont_touch of G34596: signal is true;
	signal G34598: std_logic; attribute dont_touch of G34598: signal is true;
	signal G34599: std_logic; attribute dont_touch of G34599: signal is true;
	signal G34600: std_logic; attribute dont_touch of G34600: signal is true;
	signal G34601: std_logic; attribute dont_touch of G34601: signal is true;
	signal G34602: std_logic; attribute dont_touch of G34602: signal is true;
	signal G34603: std_logic; attribute dont_touch of G34603: signal is true;
	signal G34604: std_logic; attribute dont_touch of G34604: signal is true;
	signal G34605: std_logic; attribute dont_touch of G34605: signal is true;
	signal G34606: std_logic; attribute dont_touch of G34606: signal is true;
	signal G34607: std_logic; attribute dont_touch of G34607: signal is true;
	signal G34608: std_logic; attribute dont_touch of G34608: signal is true;
	signal G34609: std_logic; attribute dont_touch of G34609: signal is true;
	signal G34610: std_logic; attribute dont_touch of G34610: signal is true;
	signal G34611: std_logic; attribute dont_touch of G34611: signal is true;
	signal G34612: std_logic; attribute dont_touch of G34612: signal is true;
	signal G34613: std_logic; attribute dont_touch of G34613: signal is true;
	signal G34614: std_logic; attribute dont_touch of G34614: signal is true;
	signal G34615: std_logic; attribute dont_touch of G34615: signal is true;
	signal G34616: std_logic; attribute dont_touch of G34616: signal is true;
	signal G34617: std_logic; attribute dont_touch of G34617: signal is true;
	signal G34618: std_logic; attribute dont_touch of G34618: signal is true;
	signal G34619: std_logic; attribute dont_touch of G34619: signal is true;
	signal G34620: std_logic; attribute dont_touch of G34620: signal is true;
	signal G34621: std_logic; attribute dont_touch of G34621: signal is true;
	signal G34622: std_logic; attribute dont_touch of G34622: signal is true;
	signal G34623: std_logic; attribute dont_touch of G34623: signal is true;
	signal G34624: std_logic; attribute dont_touch of G34624: signal is true;
	signal G34625: std_logic; attribute dont_touch of G34625: signal is true;
	signal G34626: std_logic; attribute dont_touch of G34626: signal is true;
	signal G34627: std_logic; attribute dont_touch of G34627: signal is true;
	signal G34628: std_logic; attribute dont_touch of G34628: signal is true;
	signal G34629: std_logic; attribute dont_touch of G34629: signal is true;
	signal G34630: std_logic; attribute dont_touch of G34630: signal is true;
	signal G34631: std_logic; attribute dont_touch of G34631: signal is true;
	signal G34632: std_logic; attribute dont_touch of G34632: signal is true;
	signal G34633: std_logic; attribute dont_touch of G34633: signal is true;
	signal G34634: std_logic; attribute dont_touch of G34634: signal is true;
	signal G34635: std_logic; attribute dont_touch of G34635: signal is true;
	signal G34636: std_logic; attribute dont_touch of G34636: signal is true;
	signal G34637: std_logic; attribute dont_touch of G34637: signal is true;
	signal G34638: std_logic; attribute dont_touch of G34638: signal is true;
	signal G34639: std_logic; attribute dont_touch of G34639: signal is true;
	signal G34640: std_logic; attribute dont_touch of G34640: signal is true;
	signal G34641: std_logic; attribute dont_touch of G34641: signal is true;
	signal G34642: std_logic; attribute dont_touch of G34642: signal is true;
	signal G34643: std_logic; attribute dont_touch of G34643: signal is true;
	signal G34644: std_logic; attribute dont_touch of G34644: signal is true;
	signal G34645: std_logic; attribute dont_touch of G34645: signal is true;
	signal G34646: std_logic; attribute dont_touch of G34646: signal is true;
	signal G34647: std_logic; attribute dont_touch of G34647: signal is true;
	signal G34648: std_logic; attribute dont_touch of G34648: signal is true;
	signal G34649: std_logic; attribute dont_touch of G34649: signal is true;
	signal G34650: std_logic; attribute dont_touch of G34650: signal is true;
	signal G34653: std_logic; attribute dont_touch of G34653: signal is true;
	signal G34654: std_logic; attribute dont_touch of G34654: signal is true;
	signal G34655: std_logic; attribute dont_touch of G34655: signal is true;
	signal G34656: std_logic; attribute dont_touch of G34656: signal is true;
	signal G34657: std_logic; attribute dont_touch of G34657: signal is true;
	signal G34658: std_logic; attribute dont_touch of G34658: signal is true;
	signal G34659: std_logic; attribute dont_touch of G34659: signal is true;
	signal G34660: std_logic; attribute dont_touch of G34660: signal is true;
	signal G34661: std_logic; attribute dont_touch of G34661: signal is true;
	signal G34662: std_logic; attribute dont_touch of G34662: signal is true;
	signal G34663: std_logic; attribute dont_touch of G34663: signal is true;
	signal G34664: std_logic; attribute dont_touch of G34664: signal is true;
	signal G34665: std_logic; attribute dont_touch of G34665: signal is true;
	signal G34666: std_logic; attribute dont_touch of G34666: signal is true;
	signal G34667: std_logic; attribute dont_touch of G34667: signal is true;
	signal G34668: std_logic; attribute dont_touch of G34668: signal is true;
	signal G34669: std_logic; attribute dont_touch of G34669: signal is true;
	signal G34670: std_logic; attribute dont_touch of G34670: signal is true;
	signal G34671: std_logic; attribute dont_touch of G34671: signal is true;
	signal G34672: std_logic; attribute dont_touch of G34672: signal is true;
	signal G34673: std_logic; attribute dont_touch of G34673: signal is true;
	signal G34674: std_logic; attribute dont_touch of G34674: signal is true;
	signal G34675: std_logic; attribute dont_touch of G34675: signal is true;
	signal G34676: std_logic; attribute dont_touch of G34676: signal is true;
	signal G34677: std_logic; attribute dont_touch of G34677: signal is true;
	signal G34678: std_logic; attribute dont_touch of G34678: signal is true;
	signal G34679: std_logic; attribute dont_touch of G34679: signal is true;
	signal G34680: std_logic; attribute dont_touch of G34680: signal is true;
	signal G34681: std_logic; attribute dont_touch of G34681: signal is true;
	signal G34682: std_logic; attribute dont_touch of G34682: signal is true;
	signal G34683: std_logic; attribute dont_touch of G34683: signal is true;
	signal G34684: std_logic; attribute dont_touch of G34684: signal is true;
	signal G34685: std_logic; attribute dont_touch of G34685: signal is true;
	signal G34686: std_logic; attribute dont_touch of G34686: signal is true;
	signal G34687: std_logic; attribute dont_touch of G34687: signal is true;
	signal G34688: std_logic; attribute dont_touch of G34688: signal is true;
	signal G34689: std_logic; attribute dont_touch of G34689: signal is true;
	signal G34690: std_logic; attribute dont_touch of G34690: signal is true;
	signal G34691: std_logic; attribute dont_touch of G34691: signal is true;
	signal G34692: std_logic; attribute dont_touch of G34692: signal is true;
	signal G34693: std_logic; attribute dont_touch of G34693: signal is true;
	signal G34694: std_logic; attribute dont_touch of G34694: signal is true;
	signal G34695: std_logic; attribute dont_touch of G34695: signal is true;
	signal G34696: std_logic; attribute dont_touch of G34696: signal is true;
	signal G34697: std_logic; attribute dont_touch of G34697: signal is true;
	signal G34698: std_logic; attribute dont_touch of G34698: signal is true;
	signal G34699: std_logic; attribute dont_touch of G34699: signal is true;
	signal G34700: std_logic; attribute dont_touch of G34700: signal is true;
	signal G34701: std_logic; attribute dont_touch of G34701: signal is true;
	signal G34702: std_logic; attribute dont_touch of G34702: signal is true;
	signal G34703: std_logic; attribute dont_touch of G34703: signal is true;
	signal G34706: std_logic; attribute dont_touch of G34706: signal is true;
	signal G34707: std_logic; attribute dont_touch of G34707: signal is true;
	signal G34708: std_logic; attribute dont_touch of G34708: signal is true;
	signal G34709: std_logic; attribute dont_touch of G34709: signal is true;
	signal G34710: std_logic; attribute dont_touch of G34710: signal is true;
	signal G34711: std_logic; attribute dont_touch of G34711: signal is true;
	signal G34712: std_logic; attribute dont_touch of G34712: signal is true;
	signal G34713: std_logic; attribute dont_touch of G34713: signal is true;
	signal G34714: std_logic; attribute dont_touch of G34714: signal is true;
	signal G34715: std_logic; attribute dont_touch of G34715: signal is true;
	signal G34716: std_logic; attribute dont_touch of G34716: signal is true;
	signal G34717: std_logic; attribute dont_touch of G34717: signal is true;
	signal G34718: std_logic; attribute dont_touch of G34718: signal is true;
	signal G34719: std_logic; attribute dont_touch of G34719: signal is true;
	signal G34720: std_logic; attribute dont_touch of G34720: signal is true;
	signal G34721: std_logic; attribute dont_touch of G34721: signal is true;
	signal G34722: std_logic; attribute dont_touch of G34722: signal is true;
	signal G34723: std_logic; attribute dont_touch of G34723: signal is true;
	signal G34724: std_logic; attribute dont_touch of G34724: signal is true;
	signal G34725: std_logic; attribute dont_touch of G34725: signal is true;
	signal G34726: std_logic; attribute dont_touch of G34726: signal is true;
	signal G34727: std_logic; attribute dont_touch of G34727: signal is true;
	signal G34728: std_logic; attribute dont_touch of G34728: signal is true;
	signal G34729: std_logic; attribute dont_touch of G34729: signal is true;
	signal G34730: std_logic; attribute dont_touch of G34730: signal is true;
	signal G34731: std_logic; attribute dont_touch of G34731: signal is true;
	signal G34732: std_logic; attribute dont_touch of G34732: signal is true;
	signal G34733: std_logic; attribute dont_touch of G34733: signal is true;
	signal G34734: std_logic; attribute dont_touch of G34734: signal is true;
	signal G34735: std_logic; attribute dont_touch of G34735: signal is true;
	signal G34736: std_logic; attribute dont_touch of G34736: signal is true;
	signal G34737: std_logic; attribute dont_touch of G34737: signal is true;
	signal G34738: std_logic; attribute dont_touch of G34738: signal is true;
	signal G34739: std_logic; attribute dont_touch of G34739: signal is true;
	signal G34740: std_logic; attribute dont_touch of G34740: signal is true;
	signal G34741: std_logic; attribute dont_touch of G34741: signal is true;
	signal G34742: std_logic; attribute dont_touch of G34742: signal is true;
	signal G34743: std_logic; attribute dont_touch of G34743: signal is true;
	signal G34744: std_logic; attribute dont_touch of G34744: signal is true;
	signal G34745: std_logic; attribute dont_touch of G34745: signal is true;
	signal G34746: std_logic; attribute dont_touch of G34746: signal is true;
	signal G34747: std_logic; attribute dont_touch of G34747: signal is true;
	signal G34748: std_logic; attribute dont_touch of G34748: signal is true;
	signal G34749: std_logic; attribute dont_touch of G34749: signal is true;
	signal G34750: std_logic; attribute dont_touch of G34750: signal is true;
	signal G34751: std_logic; attribute dont_touch of G34751: signal is true;
	signal G34752: std_logic; attribute dont_touch of G34752: signal is true;
	signal G34753: std_logic; attribute dont_touch of G34753: signal is true;
	signal G34754: std_logic; attribute dont_touch of G34754: signal is true;
	signal G34755: std_logic; attribute dont_touch of G34755: signal is true;
	signal G34756: std_logic; attribute dont_touch of G34756: signal is true;
	signal G34757: std_logic; attribute dont_touch of G34757: signal is true;
	signal G34758: std_logic; attribute dont_touch of G34758: signal is true;
	signal G34759: std_logic; attribute dont_touch of G34759: signal is true;
	signal G34760: std_logic; attribute dont_touch of G34760: signal is true;
	signal G34761: std_logic; attribute dont_touch of G34761: signal is true;
	signal G34762: std_logic; attribute dont_touch of G34762: signal is true;
	signal G34763: std_logic; attribute dont_touch of G34763: signal is true;
	signal G34764: std_logic; attribute dont_touch of G34764: signal is true;
	signal G34765: std_logic; attribute dont_touch of G34765: signal is true;
	signal G34766: std_logic; attribute dont_touch of G34766: signal is true;
	signal G34767: std_logic; attribute dont_touch of G34767: signal is true;
	signal G34768: std_logic; attribute dont_touch of G34768: signal is true;
	signal G34769: std_logic; attribute dont_touch of G34769: signal is true;
	signal G34770: std_logic; attribute dont_touch of G34770: signal is true;
	signal G34771: std_logic; attribute dont_touch of G34771: signal is true;
	signal G34772: std_logic; attribute dont_touch of G34772: signal is true;
	signal G34773: std_logic; attribute dont_touch of G34773: signal is true;
	signal G34774: std_logic; attribute dont_touch of G34774: signal is true;
	signal G34775: std_logic; attribute dont_touch of G34775: signal is true;
	signal G34776: std_logic; attribute dont_touch of G34776: signal is true;
	signal G34777: std_logic; attribute dont_touch of G34777: signal is true;
	signal G34778: std_logic; attribute dont_touch of G34778: signal is true;
	signal G34781: std_logic; attribute dont_touch of G34781: signal is true;
	signal G34782: std_logic; attribute dont_touch of G34782: signal is true;
	signal G34783: std_logic; attribute dont_touch of G34783: signal is true;
	signal G34784: std_logic; attribute dont_touch of G34784: signal is true;
	signal G34785: std_logic; attribute dont_touch of G34785: signal is true;
	signal G34786: std_logic; attribute dont_touch of G34786: signal is true;
	signal G34787: std_logic; attribute dont_touch of G34787: signal is true;
	signal G34789: std_logic; attribute dont_touch of G34789: signal is true;
	signal G34790: std_logic; attribute dont_touch of G34790: signal is true;
	signal G34791: std_logic; attribute dont_touch of G34791: signal is true;
	signal G34792: std_logic; attribute dont_touch of G34792: signal is true;
	signal G34793: std_logic; attribute dont_touch of G34793: signal is true;
	signal G34794: std_logic; attribute dont_touch of G34794: signal is true;
	signal G34795: std_logic; attribute dont_touch of G34795: signal is true;
	signal G34796: std_logic; attribute dont_touch of G34796: signal is true;
	signal G34797: std_logic; attribute dont_touch of G34797: signal is true;
	signal G34798: std_logic; attribute dont_touch of G34798: signal is true;
	signal G34799: std_logic; attribute dont_touch of G34799: signal is true;
	signal G34800: std_logic; attribute dont_touch of G34800: signal is true;
	signal G34801: std_logic; attribute dont_touch of G34801: signal is true;
	signal G34802: std_logic; attribute dont_touch of G34802: signal is true;
	signal G34803: std_logic; attribute dont_touch of G34803: signal is true;
	signal G34804: std_logic; attribute dont_touch of G34804: signal is true;
	signal G34805: std_logic; attribute dont_touch of G34805: signal is true;
	signal G34806: std_logic; attribute dont_touch of G34806: signal is true;
	signal G34807: std_logic; attribute dont_touch of G34807: signal is true;
	signal G34808: std_logic; attribute dont_touch of G34808: signal is true;
	signal G34809: std_logic; attribute dont_touch of G34809: signal is true;
	signal G34810: std_logic; attribute dont_touch of G34810: signal is true;
	signal G34811: std_logic; attribute dont_touch of G34811: signal is true;
	signal G34812: std_logic; attribute dont_touch of G34812: signal is true;
	signal G34813: std_logic; attribute dont_touch of G34813: signal is true;
	signal G34816: std_logic; attribute dont_touch of G34816: signal is true;
	signal G34819: std_logic; attribute dont_touch of G34819: signal is true;
	signal G34820: std_logic; attribute dont_touch of G34820: signal is true;
	signal G34823: std_logic; attribute dont_touch of G34823: signal is true;
	signal G34826: std_logic; attribute dont_touch of G34826: signal is true;
	signal G34827: std_logic; attribute dont_touch of G34827: signal is true;
	signal G34830: std_logic; attribute dont_touch of G34830: signal is true;
	signal G34833: std_logic; attribute dont_touch of G34833: signal is true;
	signal G34836: std_logic; attribute dont_touch of G34836: signal is true;
	signal G34840: std_logic; attribute dont_touch of G34840: signal is true;
	signal G34841: std_logic; attribute dont_touch of G34841: signal is true;
	signal G34842: std_logic; attribute dont_touch of G34842: signal is true;
	signal G34843: std_logic; attribute dont_touch of G34843: signal is true;
	signal G34844: std_logic; attribute dont_touch of G34844: signal is true;
	signal G34845: std_logic; attribute dont_touch of G34845: signal is true;
	signal G34846: std_logic; attribute dont_touch of G34846: signal is true;
	signal G34847: std_logic; attribute dont_touch of G34847: signal is true;
	signal G34848: std_logic; attribute dont_touch of G34848: signal is true;
	signal G34849: std_logic; attribute dont_touch of G34849: signal is true;
	signal G34850: std_logic; attribute dont_touch of G34850: signal is true;
	signal G34851: std_logic; attribute dont_touch of G34851: signal is true;
	signal G34852: std_logic; attribute dont_touch of G34852: signal is true;
	signal G34855: std_logic; attribute dont_touch of G34855: signal is true;
	signal G34856: std_logic; attribute dont_touch of G34856: signal is true;
	signal G34857: std_logic; attribute dont_touch of G34857: signal is true;
	signal G34858: std_logic; attribute dont_touch of G34858: signal is true;
	signal G34859: std_logic; attribute dont_touch of G34859: signal is true;
	signal G34860: std_logic; attribute dont_touch of G34860: signal is true;
	signal G34861: std_logic; attribute dont_touch of G34861: signal is true;
	signal G34862: std_logic; attribute dont_touch of G34862: signal is true;
	signal G34863: std_logic; attribute dont_touch of G34863: signal is true;
	signal G34864: std_logic; attribute dont_touch of G34864: signal is true;
	signal G34865: std_logic; attribute dont_touch of G34865: signal is true;
	signal G34866: std_logic; attribute dont_touch of G34866: signal is true;
	signal G34867: std_logic; attribute dont_touch of G34867: signal is true;
	signal G34868: std_logic; attribute dont_touch of G34868: signal is true;
	signal G34869: std_logic; attribute dont_touch of G34869: signal is true;
	signal G34870: std_logic; attribute dont_touch of G34870: signal is true;
	signal G34871: std_logic; attribute dont_touch of G34871: signal is true;
	signal G34872: std_logic; attribute dont_touch of G34872: signal is true;
	signal G34873: std_logic; attribute dont_touch of G34873: signal is true;
	signal G34874: std_logic; attribute dont_touch of G34874: signal is true;
	signal G34875: std_logic; attribute dont_touch of G34875: signal is true;
	signal G34876: std_logic; attribute dont_touch of G34876: signal is true;
	signal G34877: std_logic; attribute dont_touch of G34877: signal is true;
	signal G34878: std_logic; attribute dont_touch of G34878: signal is true;
	signal G34879: std_logic; attribute dont_touch of G34879: signal is true;
	signal G34880: std_logic; attribute dont_touch of G34880: signal is true;
	signal G34881: std_logic; attribute dont_touch of G34881: signal is true;
	signal G34882: std_logic; attribute dont_touch of G34882: signal is true;
	signal G34883: std_logic; attribute dont_touch of G34883: signal is true;
	signal G34884: std_logic; attribute dont_touch of G34884: signal is true;
	signal G34887: std_logic; attribute dont_touch of G34887: signal is true;
	signal G34890: std_logic; attribute dont_touch of G34890: signal is true;
	signal G34893: std_logic; attribute dont_touch of G34893: signal is true;
	signal G34894: std_logic; attribute dont_touch of G34894: signal is true;
	signal G34897: std_logic; attribute dont_touch of G34897: signal is true;
	signal G34900: std_logic; attribute dont_touch of G34900: signal is true;
	signal G34903: std_logic; attribute dont_touch of G34903: signal is true;
	signal G34906: std_logic; attribute dont_touch of G34906: signal is true;
	signal G34909: std_logic; attribute dont_touch of G34909: signal is true;
	signal G34910: std_logic; attribute dont_touch of G34910: signal is true;
	signal G34911: std_logic; attribute dont_touch of G34911: signal is true;
	signal G34912: std_logic; attribute dont_touch of G34912: signal is true;
	signal G34914: std_logic; attribute dont_touch of G34914: signal is true;
	signal G34916: std_logic; attribute dont_touch of G34916: signal is true;
	signal G34918: std_logic; attribute dont_touch of G34918: signal is true;
	signal G34920: std_logic; attribute dont_touch of G34920: signal is true;
	signal G34922: std_logic; attribute dont_touch of G34922: signal is true;
	signal G34924: std_logic; attribute dont_touch of G34924: signal is true;
	signal G34926: std_logic; attribute dont_touch of G34926: signal is true;
	signal G34928: std_logic; attribute dont_touch of G34928: signal is true;
	signal G34929: std_logic; attribute dont_touch of G34929: signal is true;
	signal G34930: std_logic; attribute dont_touch of G34930: signal is true;
	signal G34931: std_logic; attribute dont_touch of G34931: signal is true;
	signal G34932: std_logic; attribute dont_touch of G34932: signal is true;
	signal G34933: std_logic; attribute dont_touch of G34933: signal is true;
	signal G34934: std_logic; attribute dont_touch of G34934: signal is true;
	signal G34935: std_logic; attribute dont_touch of G34935: signal is true;
	signal G34938: std_logic; attribute dont_touch of G34938: signal is true;
	signal G34939: std_logic; attribute dont_touch of G34939: signal is true;
	signal G34940: std_logic; attribute dont_touch of G34940: signal is true;
	signal G34941: std_logic; attribute dont_touch of G34941: signal is true;
	signal G34942: std_logic; attribute dont_touch of G34942: signal is true;
	signal G34943: std_logic; attribute dont_touch of G34943: signal is true;
	signal G34944: std_logic; attribute dont_touch of G34944: signal is true;
	signal G34945: std_logic; attribute dont_touch of G34945: signal is true;
	signal G34946: std_logic; attribute dont_touch of G34946: signal is true;
	signal G34947: std_logic; attribute dont_touch of G34947: signal is true;
	signal G34948: std_logic; attribute dont_touch of G34948: signal is true;
	signal G34949: std_logic; attribute dont_touch of G34949: signal is true;
	signal G34950: std_logic; attribute dont_touch of G34950: signal is true;
	signal G34951: std_logic; attribute dont_touch of G34951: signal is true;
	signal G34952: std_logic; attribute dont_touch of G34952: signal is true;
	signal G34953: std_logic; attribute dont_touch of G34953: signal is true;
	signal G34954: std_logic; attribute dont_touch of G34954: signal is true;
	signal G34955: std_logic; attribute dont_touch of G34955: signal is true;
	signal G34957: std_logic; attribute dont_touch of G34957: signal is true;
	signal G34960: std_logic; attribute dont_touch of G34960: signal is true;
	signal G34961: std_logic; attribute dont_touch of G34961: signal is true;
	signal G34962: std_logic; attribute dont_touch of G34962: signal is true;
	signal G34963: std_logic; attribute dont_touch of G34963: signal is true;
	signal G34964: std_logic; attribute dont_touch of G34964: signal is true;
	signal G34965: std_logic; attribute dont_touch of G34965: signal is true;
	signal G34966: std_logic; attribute dont_touch of G34966: signal is true;
	signal G34967: std_logic; attribute dont_touch of G34967: signal is true;
	signal G34968: std_logic; attribute dont_touch of G34968: signal is true;
	signal G34969: std_logic; attribute dont_touch of G34969: signal is true;
	signal G34970: std_logic; attribute dont_touch of G34970: signal is true;
	signal G34971: std_logic; attribute dont_touch of G34971: signal is true;
	signal G34973: std_logic; attribute dont_touch of G34973: signal is true;
	signal G34974: std_logic; attribute dont_touch of G34974: signal is true;
	signal G34975: std_logic; attribute dont_touch of G34975: signal is true;
	signal G34976: std_logic; attribute dont_touch of G34976: signal is true;
	signal G34977: std_logic; attribute dont_touch of G34977: signal is true;
	signal G34978: std_logic; attribute dont_touch of G34978: signal is true;
	signal G34979: std_logic; attribute dont_touch of G34979: signal is true;
	signal G34980: std_logic; attribute dont_touch of G34980: signal is true;
	signal G34981: std_logic; attribute dont_touch of G34981: signal is true;
	signal G34982: std_logic; attribute dont_touch of G34982: signal is true;
	signal G34983: std_logic; attribute dont_touch of G34983: signal is true;
	signal G34984: std_logic; attribute dont_touch of G34984: signal is true;
	signal G34985: std_logic; attribute dont_touch of G34985: signal is true;
	signal G34986: std_logic; attribute dont_touch of G34986: signal is true;
	signal G34987: std_logic; attribute dont_touch of G34987: signal is true;
	signal G34988: std_logic; attribute dont_touch of G34988: signal is true;
	signal G34989: std_logic; attribute dont_touch of G34989: signal is true;
	signal G34990: std_logic; attribute dont_touch of G34990: signal is true;
	signal G34991: std_logic; attribute dont_touch of G34991: signal is true;
	signal G34992: std_logic; attribute dont_touch of G34992: signal is true;
	signal G34993: std_logic; attribute dont_touch of G34993: signal is true;
	signal G34994: std_logic; attribute dont_touch of G34994: signal is true;
	signal G34995: std_logic; attribute dont_touch of G34995: signal is true;
	signal G34996: std_logic; attribute dont_touch of G34996: signal is true;
	signal G34997: std_logic; attribute dont_touch of G34997: signal is true;
	signal G34998: std_logic; attribute dont_touch of G34998: signal is true;
	signal G34999: std_logic; attribute dont_touch of G34999: signal is true;
	signal G35000: std_logic; attribute dont_touch of G35000: signal is true;
	signal G35001: std_logic; attribute dont_touch of G35001: signal is true;
	signal G35002: std_logic; attribute dont_touch of G35002: signal is true;
	signal I11617: std_logic; attribute dont_touch of I11617: signal is true;
	signal I11620: std_logic; attribute dont_touch of I11620: signal is true;
	signal I11623: std_logic; attribute dont_touch of I11623: signal is true;
	signal I11626: std_logic; attribute dont_touch of I11626: signal is true;
	signal I11629: std_logic; attribute dont_touch of I11629: signal is true;
	signal I11632: std_logic; attribute dont_touch of I11632: signal is true;
	signal I11635: std_logic; attribute dont_touch of I11635: signal is true;
	signal I11655: std_logic; attribute dont_touch of I11655: signal is true;
	signal I11665: std_logic; attribute dont_touch of I11665: signal is true;
	signal I11682: std_logic; attribute dont_touch of I11682: signal is true;
	signal I11685: std_logic; attribute dont_touch of I11685: signal is true;
	signal I11688: std_logic; attribute dont_touch of I11688: signal is true;
	signal I11691: std_logic; attribute dont_touch of I11691: signal is true;
	signal I11697: std_logic; attribute dont_touch of I11697: signal is true;
	signal I11701: std_logic; attribute dont_touch of I11701: signal is true;
	signal I11708: std_logic; attribute dont_touch of I11708: signal is true;
	signal I11716: std_logic; attribute dont_touch of I11716: signal is true;
	signal I11721: std_logic; attribute dont_touch of I11721: signal is true;
	signal I11726: std_logic; attribute dont_touch of I11726: signal is true;
	signal I11734: std_logic; attribute dont_touch of I11734: signal is true;
	signal I11737: std_logic; attribute dont_touch of I11737: signal is true;
	signal I11740: std_logic; attribute dont_touch of I11740: signal is true;
	signal I11743: std_logic; attribute dont_touch of I11743: signal is true;
	signal I11746: std_logic; attribute dont_touch of I11746: signal is true;
	signal I11750: std_logic; attribute dont_touch of I11750: signal is true;
	signal I11753: std_logic; attribute dont_touch of I11753: signal is true;
	signal I11777: std_logic; attribute dont_touch of I11777: signal is true;
	signal I11785: std_logic; attribute dont_touch of I11785: signal is true;
	signal I11793: std_logic; attribute dont_touch of I11793: signal is true;
	signal I11801: std_logic; attribute dont_touch of I11801: signal is true;
	signal I11809: std_logic; attribute dont_touch of I11809: signal is true;
	signal I11816: std_logic; attribute dont_touch of I11816: signal is true;
	signal I11820: std_logic; attribute dont_touch of I11820: signal is true;
	signal I11824: std_logic; attribute dont_touch of I11824: signal is true;
	signal I11825: std_logic; attribute dont_touch of I11825: signal is true;
	signal I11826: std_logic; attribute dont_touch of I11826: signal is true;
	signal I11835: std_logic; attribute dont_touch of I11835: signal is true;
	signal I11843: std_logic; attribute dont_touch of I11843: signal is true;
	signal I11860: std_logic; attribute dont_touch of I11860: signal is true;
	signal I11864: std_logic; attribute dont_touch of I11864: signal is true;
	signal I11865: std_logic; attribute dont_touch of I11865: signal is true;
	signal I11866: std_logic; attribute dont_touch of I11866: signal is true;
	signal I11877: std_logic; attribute dont_touch of I11877: signal is true;
	signal I11878: std_logic; attribute dont_touch of I11878: signal is true;
	signal I11879: std_logic; attribute dont_touch of I11879: signal is true;
	signal I11892: std_logic; attribute dont_touch of I11892: signal is true;
	signal I11896: std_logic; attribute dont_touch of I11896: signal is true;
	signal I11903: std_logic; attribute dont_touch of I11903: signal is true;
	signal I11908: std_logic; attribute dont_touch of I11908: signal is true;
	signal I11980: std_logic; attribute dont_touch of I11980: signal is true;
	signal I11992: std_logic; attribute dont_touch of I11992: signal is true;
	signal I12000: std_logic; attribute dont_touch of I12000: signal is true;
	signal I12003: std_logic; attribute dont_touch of I12003: signal is true;
	signal I12013: std_logic; attribute dont_touch of I12013: signal is true;
	signal I12016: std_logic; attribute dont_touch of I12016: signal is true;
	signal I12026: std_logic; attribute dont_touch of I12026: signal is true;
	signal I12030: std_logic; attribute dont_touch of I12030: signal is true;
	signal I12033: std_logic; attribute dont_touch of I12033: signal is true;
	signal I12041: std_logic; attribute dont_touch of I12041: signal is true;
	signal I12046: std_logic; attribute dont_touch of I12046: signal is true;
	signal I12049: std_logic; attribute dont_touch of I12049: signal is true;
	signal I12056: std_logic; attribute dont_touch of I12056: signal is true;
	signal I12061: std_logic; attribute dont_touch of I12061: signal is true;
	signal I12064: std_logic; attribute dont_touch of I12064: signal is true;
	signal I12067: std_logic; attribute dont_touch of I12067: signal is true;
	signal I12070: std_logic; attribute dont_touch of I12070: signal is true;
	signal I12074: std_logic; attribute dont_touch of I12074: signal is true;
	signal I12075: std_logic; attribute dont_touch of I12075: signal is true;
	signal I12076: std_logic; attribute dont_touch of I12076: signal is true;
	signal I12083: std_logic; attribute dont_touch of I12083: signal is true;
	signal I12086: std_logic; attribute dont_touch of I12086: signal is true;
	signal I12089: std_logic; attribute dont_touch of I12089: signal is true;
	signal I12092: std_logic; attribute dont_touch of I12092: signal is true;
	signal I12096: std_logic; attribute dont_touch of I12096: signal is true;
	signal I12097: std_logic; attribute dont_touch of I12097: signal is true;
	signal I12098: std_logic; attribute dont_touch of I12098: signal is true;
	signal I12103: std_logic; attribute dont_touch of I12103: signal is true;
	signal I12106: std_logic; attribute dont_touch of I12106: signal is true;
	signal I12109: std_logic; attribute dont_touch of I12109: signal is true;
	signal I12112: std_logic; attribute dont_touch of I12112: signal is true;
	signal I12117: std_logic; attribute dont_touch of I12117: signal is true;
	signal I12120: std_logic; attribute dont_touch of I12120: signal is true;
	signal I12123: std_logic; attribute dont_touch of I12123: signal is true;
	signal I12128: std_logic; attribute dont_touch of I12128: signal is true;
	signal I12132: std_logic; attribute dont_touch of I12132: signal is true;
	signal I12135: std_logic; attribute dont_touch of I12135: signal is true;
	signal I12141: std_logic; attribute dont_touch of I12141: signal is true;
	signal I12144: std_logic; attribute dont_touch of I12144: signal is true;
	signal I12151: std_logic; attribute dont_touch of I12151: signal is true;
	signal I12159: std_logic; attribute dont_touch of I12159: signal is true;
	signal I12167: std_logic; attribute dont_touch of I12167: signal is true;
	signal I12172: std_logic; attribute dont_touch of I12172: signal is true;
	signal I12176: std_logic; attribute dont_touch of I12176: signal is true;
	signal I12183: std_logic; attribute dont_touch of I12183: signal is true;
	signal I12189: std_logic; attribute dont_touch of I12189: signal is true;
	signal I12199: std_logic; attribute dont_touch of I12199: signal is true;
	signal I12203: std_logic; attribute dont_touch of I12203: signal is true;
	signal I12204: std_logic; attribute dont_touch of I12204: signal is true;
	signal I12205: std_logic; attribute dont_touch of I12205: signal is true;
	signal I12214: std_logic; attribute dont_touch of I12214: signal is true;
	signal I12217: std_logic; attribute dont_touch of I12217: signal is true;
	signal I12218: std_logic; attribute dont_touch of I12218: signal is true;
	signal I12219: std_logic; attribute dont_touch of I12219: signal is true;
	signal I12227: std_logic; attribute dont_touch of I12227: signal is true;
	signal I12240: std_logic; attribute dont_touch of I12240: signal is true;
	signal I12241: std_logic; attribute dont_touch of I12241: signal is true;
	signal I12242: std_logic; attribute dont_touch of I12242: signal is true;
	signal I12251: std_logic; attribute dont_touch of I12251: signal is true;
	signal I12252: std_logic; attribute dont_touch of I12252: signal is true;
	signal I12253: std_logic; attribute dont_touch of I12253: signal is true;
	signal I12261: std_logic; attribute dont_touch of I12261: signal is true;
	signal I12262: std_logic; attribute dont_touch of I12262: signal is true;
	signal I12263: std_logic; attribute dont_touch of I12263: signal is true;
	signal I12269: std_logic; attribute dont_touch of I12269: signal is true;
	signal I12270: std_logic; attribute dont_touch of I12270: signal is true;
	signal I12271: std_logic; attribute dont_touch of I12271: signal is true;
	signal I12277: std_logic; attribute dont_touch of I12277: signal is true;
	signal I12278: std_logic; attribute dont_touch of I12278: signal is true;
	signal I12279: std_logic; attribute dont_touch of I12279: signal is true;
	signal I12287: std_logic; attribute dont_touch of I12287: signal is true;
	signal I12288: std_logic; attribute dont_touch of I12288: signal is true;
	signal I12289: std_logic; attribute dont_touch of I12289: signal is true;
	signal I12300: std_logic; attribute dont_touch of I12300: signal is true;
	signal I12314: std_logic; attribute dont_touch of I12314: signal is true;
	signal I12333: std_logic; attribute dont_touch of I12333: signal is true;
	signal I12336: std_logic; attribute dont_touch of I12336: signal is true;
	signal I12344: std_logic; attribute dont_touch of I12344: signal is true;
	signal I12345: std_logic; attribute dont_touch of I12345: signal is true;
	signal I12346: std_logic; attribute dont_touch of I12346: signal is true;
	signal I12355: std_logic; attribute dont_touch of I12355: signal is true;
	signal I12360: std_logic; attribute dont_touch of I12360: signal is true;
	signal I12372: std_logic; attribute dont_touch of I12372: signal is true;
	signal I12373: std_logic; attribute dont_touch of I12373: signal is true;
	signal I12374: std_logic; attribute dont_touch of I12374: signal is true;
	signal I12382: std_logic; attribute dont_touch of I12382: signal is true;
	signal I12401: std_logic; attribute dont_touch of I12401: signal is true;
	signal I12402: std_logic; attribute dont_touch of I12402: signal is true;
	signal I12403: std_logic; attribute dont_touch of I12403: signal is true;
	signal I12411: std_logic; attribute dont_touch of I12411: signal is true;
	signal I12415: std_logic; attribute dont_touch of I12415: signal is true;
	signal I12418: std_logic; attribute dont_touch of I12418: signal is true;
	signal I12437: std_logic; attribute dont_touch of I12437: signal is true;
	signal I12451: std_logic; attribute dont_touch of I12451: signal is true;
	signal I12463: std_logic; attribute dont_touch of I12463: signal is true;
	signal I12468: std_logic; attribute dont_touch of I12468: signal is true;
	signal I12469: std_logic; attribute dont_touch of I12469: signal is true;
	signal I12470: std_logic; attribute dont_touch of I12470: signal is true;
	signal I12483: std_logic; attribute dont_touch of I12483: signal is true;
	signal I12487: std_logic; attribute dont_touch of I12487: signal is true;
	signal I12493: std_logic; attribute dont_touch of I12493: signal is true;
	signal I12497: std_logic; attribute dont_touch of I12497: signal is true;
	signal I12503: std_logic; attribute dont_touch of I12503: signal is true;
	signal I12519: std_logic; attribute dont_touch of I12519: signal is true;
	signal I12523: std_logic; attribute dont_touch of I12523: signal is true;
	signal I12530: std_logic; attribute dont_touch of I12530: signal is true;
	signal I12534: std_logic; attribute dont_touch of I12534: signal is true;
	signal I12538: std_logic; attribute dont_touch of I12538: signal is true;
	signal I12541: std_logic; attribute dont_touch of I12541: signal is true;
	signal I12544: std_logic; attribute dont_touch of I12544: signal is true;
	signal I12545: std_logic; attribute dont_touch of I12545: signal is true;
	signal I12546: std_logic; attribute dont_touch of I12546: signal is true;
	signal I12563: std_logic; attribute dont_touch of I12563: signal is true;
	signal I12568: std_logic; attribute dont_touch of I12568: signal is true;
	signal I12572: std_logic; attribute dont_touch of I12572: signal is true;
	signal I12577: std_logic; attribute dont_touch of I12577: signal is true;
	signal I12580: std_logic; attribute dont_touch of I12580: signal is true;
	signal I12583: std_logic; attribute dont_touch of I12583: signal is true;
	signal I12605: std_logic; attribute dont_touch of I12605: signal is true;
	signal I12608: std_logic; attribute dont_touch of I12608: signal is true;
	signal I12611: std_logic; attribute dont_touch of I12611: signal is true;
	signal I12618: std_logic; attribute dont_touch of I12618: signal is true;
	signal I12631: std_logic; attribute dont_touch of I12631: signal is true;
	signal I12644: std_logic; attribute dont_touch of I12644: signal is true;
	signal I12654: std_logic; attribute dont_touch of I12654: signal is true;
	signal I12666: std_logic; attribute dont_touch of I12666: signal is true;
	signal I12709: std_logic; attribute dont_touch of I12709: signal is true;
	signal I12712: std_logic; attribute dont_touch of I12712: signal is true;
	signal I12719: std_logic; attribute dont_touch of I12719: signal is true;
	signal I12728: std_logic; attribute dont_touch of I12728: signal is true;
	signal I12729: std_logic; attribute dont_touch of I12729: signal is true;
	signal I12730: std_logic; attribute dont_touch of I12730: signal is true;
	signal I12735: std_logic; attribute dont_touch of I12735: signal is true;
	signal I12746: std_logic; attribute dont_touch of I12746: signal is true;
	signal I12749: std_logic; attribute dont_touch of I12749: signal is true;
	signal I12758: std_logic; attribute dont_touch of I12758: signal is true;
	signal I12761: std_logic; attribute dont_touch of I12761: signal is true;
	signal I12764: std_logic; attribute dont_touch of I12764: signal is true;
	signal I12767: std_logic; attribute dont_touch of I12767: signal is true;
	signal I12770: std_logic; attribute dont_touch of I12770: signal is true;
	signal I12773: std_logic; attribute dont_touch of I12773: signal is true;
	signal I12776: std_logic; attribute dont_touch of I12776: signal is true;
	signal I12779: std_logic; attribute dont_touch of I12779: signal is true;
	signal I12782: std_logic; attribute dont_touch of I12782: signal is true;
	signal I12783: std_logic; attribute dont_touch of I12783: signal is true;
	signal I12787: std_logic; attribute dont_touch of I12787: signal is true;
	signal I12790: std_logic; attribute dont_touch of I12790: signal is true;
	signal I12793: std_logic; attribute dont_touch of I12793: signal is true;
	signal I12799: std_logic; attribute dont_touch of I12799: signal is true;
	signal I12805: std_logic; attribute dont_touch of I12805: signal is true;
	signal I12808: std_logic; attribute dont_touch of I12808: signal is true;
	signal I12811: std_logic; attribute dont_touch of I12811: signal is true;
	signal I12819: std_logic; attribute dont_touch of I12819: signal is true;
	signal I12823: std_logic; attribute dont_touch of I12823: signal is true;
	signal I12826: std_logic; attribute dont_touch of I12826: signal is true;
	signal I12837: std_logic; attribute dont_touch of I12837: signal is true;
	signal I12840: std_logic; attribute dont_touch of I12840: signal is true;
	signal I12841: std_logic; attribute dont_touch of I12841: signal is true;
	signal I12842: std_logic; attribute dont_touch of I12842: signal is true;
	signal I12848: std_logic; attribute dont_touch of I12848: signal is true;
	signal I12849: std_logic; attribute dont_touch of I12849: signal is true;
	signal I12850: std_logic; attribute dont_touch of I12850: signal is true;
	signal I12855: std_logic; attribute dont_touch of I12855: signal is true;
	signal I12858: std_logic; attribute dont_touch of I12858: signal is true;
	signal I12861: std_logic; attribute dont_touch of I12861: signal is true;
	signal I12876: std_logic; attribute dont_touch of I12876: signal is true;
	signal I12877: std_logic; attribute dont_touch of I12877: signal is true;
	signal I12878: std_logic; attribute dont_touch of I12878: signal is true;
	signal I12884: std_logic; attribute dont_touch of I12884: signal is true;
	signal I12887: std_logic; attribute dont_touch of I12887: signal is true;
	signal I12890: std_logic; attribute dont_touch of I12890: signal is true;
	signal I12893: std_logic; attribute dont_touch of I12893: signal is true;
	signal I12896: std_logic; attribute dont_touch of I12896: signal is true;
	signal I12899: std_logic; attribute dont_touch of I12899: signal is true;
	signal I12902: std_logic; attribute dont_touch of I12902: signal is true;
	signal I12903: std_logic; attribute dont_touch of I12903: signal is true;
	signal I12907: std_logic; attribute dont_touch of I12907: signal is true;
	signal I12910: std_logic; attribute dont_touch of I12910: signal is true;
	signal I12927: std_logic; attribute dont_touch of I12927: signal is true;
	signal I12930: std_logic; attribute dont_touch of I12930: signal is true;
	signal I12935: std_logic; attribute dont_touch of I12935: signal is true;
	signal I12950: std_logic; attribute dont_touch of I12950: signal is true;
	signal I12954: std_logic; attribute dont_touch of I12954: signal is true;
	signal I12963: std_logic; attribute dont_touch of I12963: signal is true;
	signal I12987: std_logic; attribute dont_touch of I12987: signal is true;
	signal I12991: std_logic; attribute dont_touch of I12991: signal is true;
	signal I12994: std_logic; attribute dont_touch of I12994: signal is true;
	signal I12997: std_logic; attribute dont_touch of I12997: signal is true;
	signal I13007: std_logic; attribute dont_touch of I13007: signal is true;
	signal I13010: std_logic; attribute dont_touch of I13010: signal is true;
	signal I13020: std_logic; attribute dont_touch of I13020: signal is true;
	signal I13031: std_logic; attribute dont_touch of I13031: signal is true;
	signal I13037: std_logic; attribute dont_touch of I13037: signal is true;
	signal I13043: std_logic; attribute dont_touch of I13043: signal is true;
	signal I13044: std_logic; attribute dont_touch of I13044: signal is true;
	signal I13045: std_logic; attribute dont_touch of I13045: signal is true;
	signal I13054: std_logic; attribute dont_touch of I13054: signal is true;
	signal I13057: std_logic; attribute dont_touch of I13057: signal is true;
	signal I13065: std_logic; attribute dont_touch of I13065: signal is true;
	signal I13066: std_logic; attribute dont_touch of I13066: signal is true;
	signal I13067: std_logic; attribute dont_touch of I13067: signal is true;
	signal I13077: std_logic; attribute dont_touch of I13077: signal is true;
	signal I13078: std_logic; attribute dont_touch of I13078: signal is true;
	signal I13079: std_logic; attribute dont_touch of I13079: signal is true;
	signal I13094: std_logic; attribute dont_touch of I13094: signal is true;
	signal I13109: std_logic; attribute dont_touch of I13109: signal is true;
	signal I13110: std_logic; attribute dont_touch of I13110: signal is true;
	signal I13111: std_logic; attribute dont_touch of I13111: signal is true;
	signal I13124: std_logic; attribute dont_touch of I13124: signal is true;
	signal I13139: std_logic; attribute dont_touch of I13139: signal is true;
	signal I13140: std_logic; attribute dont_touch of I13140: signal is true;
	signal I13141: std_logic; attribute dont_touch of I13141: signal is true;
	signal I13149: std_logic; attribute dont_touch of I13149: signal is true;
	signal I13152: std_logic; attribute dont_touch of I13152: signal is true;
	signal I13166: std_logic; attribute dont_touch of I13166: signal is true;
	signal I13182: std_logic; attribute dont_touch of I13182: signal is true;
	signal I13183: std_logic; attribute dont_touch of I13183: signal is true;
	signal I13184: std_logic; attribute dont_touch of I13184: signal is true;
	signal I13202: std_logic; attribute dont_touch of I13202: signal is true;
	signal I13206: std_logic; attribute dont_touch of I13206: signal is true;
	signal I13236: std_logic; attribute dont_touch of I13236: signal is true;
	signal I13240: std_logic; attribute dont_touch of I13240: signal is true;
	signal I13252: std_logic; attribute dont_touch of I13252: signal is true;
	signal I13276: std_logic; attribute dont_touch of I13276: signal is true;
	signal I13280: std_logic; attribute dont_touch of I13280: signal is true;
	signal I13287: std_logic; attribute dont_touch of I13287: signal is true;
	signal I13317: std_logic; attribute dont_touch of I13317: signal is true;
	signal I13321: std_logic; attribute dont_touch of I13321: signal is true;
	signal I13326: std_logic; attribute dont_touch of I13326: signal is true;
	signal I13329: std_logic; attribute dont_touch of I13329: signal is true;
	signal I13334: std_logic; attribute dont_touch of I13334: signal is true;
	signal I13335: std_logic; attribute dont_touch of I13335: signal is true;
	signal I13336: std_logic; attribute dont_touch of I13336: signal is true;
	signal I13352: std_logic; attribute dont_touch of I13352: signal is true;
	signal I13360: std_logic; attribute dont_touch of I13360: signal is true;
	signal I13374: std_logic; attribute dont_touch of I13374: signal is true;
	signal I13382: std_logic; attribute dont_touch of I13382: signal is true;
	signal I13383: std_logic; attribute dont_touch of I13383: signal is true;
	signal I13384: std_logic; attribute dont_touch of I13384: signal is true;
	signal I13390: std_logic; attribute dont_touch of I13390: signal is true;
	signal I13391: std_logic; attribute dont_touch of I13391: signal is true;
	signal I13392: std_logic; attribute dont_touch of I13392: signal is true;
	signal I13401: std_logic; attribute dont_touch of I13401: signal is true;
	signal I13402: std_logic; attribute dont_touch of I13402: signal is true;
	signal I13403: std_logic; attribute dont_touch of I13403: signal is true;
	signal I13424: std_logic; attribute dont_touch of I13424: signal is true;
	signal I13442: std_logic; attribute dont_touch of I13442: signal is true;
	signal I13443: std_logic; attribute dont_touch of I13443: signal is true;
	signal I13444: std_logic; attribute dont_touch of I13444: signal is true;
	signal I13452: std_logic; attribute dont_touch of I13452: signal is true;
	signal I13453: std_logic; attribute dont_touch of I13453: signal is true;
	signal I13454: std_logic; attribute dont_touch of I13454: signal is true;
	signal I13462: std_logic; attribute dont_touch of I13462: signal is true;
	signal I13463: std_logic; attribute dont_touch of I13463: signal is true;
	signal I13464: std_logic; attribute dont_touch of I13464: signal is true;
	signal I13473: std_logic; attribute dont_touch of I13473: signal is true;
	signal I13483: std_logic; attribute dont_touch of I13483: signal is true;
	signal I13497: std_logic; attribute dont_touch of I13497: signal is true;
	signal I13498: std_logic; attribute dont_touch of I13498: signal is true;
	signal I13499: std_logic; attribute dont_touch of I13499: signal is true;
	signal I13509: std_logic; attribute dont_touch of I13509: signal is true;
	signal I13510: std_logic; attribute dont_touch of I13510: signal is true;
	signal I13511: std_logic; attribute dont_touch of I13511: signal is true;
	signal I13518: std_logic; attribute dont_touch of I13518: signal is true;
	signal I13519: std_logic; attribute dont_touch of I13519: signal is true;
	signal I13520: std_logic; attribute dont_touch of I13520: signal is true;
	signal I13539: std_logic; attribute dont_touch of I13539: signal is true;
	signal I13548: std_logic; attribute dont_touch of I13548: signal is true;
	signal I13552: std_logic; attribute dont_touch of I13552: signal is true;
	signal I13564: std_logic; attribute dont_touch of I13564: signal is true;
	signal I13565: std_logic; attribute dont_touch of I13565: signal is true;
	signal I13566: std_logic; attribute dont_touch of I13566: signal is true;
	signal I13581: std_logic; attribute dont_touch of I13581: signal is true;
	signal I13597: std_logic; attribute dont_touch of I13597: signal is true;
	signal I13606: std_logic; attribute dont_touch of I13606: signal is true;
	signal I13623: std_logic; attribute dont_touch of I13623: signal is true;
	signal I13634: std_logic; attribute dont_touch of I13634: signal is true;
	signal I13637: std_logic; attribute dont_touch of I13637: signal is true;
	signal I13672: std_logic; attribute dont_touch of I13672: signal is true;
	signal I13684: std_logic; attribute dont_touch of I13684: signal is true;
	signal I13694: std_logic; attribute dont_touch of I13694: signal is true;
	signal I13699: std_logic; attribute dont_touch of I13699: signal is true;
	signal I13705: std_logic; attribute dont_touch of I13705: signal is true;
	signal I13708: std_logic; attribute dont_touch of I13708: signal is true;
	signal I13715: std_logic; attribute dont_touch of I13715: signal is true;
	signal I13718: std_logic; attribute dont_touch of I13718: signal is true;
	signal I13723: std_logic; attribute dont_touch of I13723: signal is true;
	signal I13726: std_logic; attribute dont_touch of I13726: signal is true;
	signal I13729: std_logic; attribute dont_touch of I13729: signal is true;
	signal I13730: std_logic; attribute dont_touch of I13730: signal is true;
	signal I13731: std_logic; attribute dont_touch of I13731: signal is true;
	signal I13740: std_logic; attribute dont_touch of I13740: signal is true;
	signal I13744: std_logic; attribute dont_touch of I13744: signal is true;
	signal I13749: std_logic; attribute dont_touch of I13749: signal is true;
	signal I13750: std_logic; attribute dont_touch of I13750: signal is true;
	signal I13751: std_logic; attribute dont_touch of I13751: signal is true;
	signal I13759: std_logic; attribute dont_touch of I13759: signal is true;
	signal I13762: std_logic; attribute dont_touch of I13762: signal is true;
	signal I13779: std_logic; attribute dont_touch of I13779: signal is true;
	signal I13802: std_logic; attribute dont_touch of I13802: signal is true;
	signal I13805: std_logic; attribute dont_touch of I13805: signal is true;
	signal I13847: std_logic; attribute dont_touch of I13847: signal is true;
	signal I13850: std_logic; attribute dont_touch of I13850: signal is true;
	signal I13851: std_logic; attribute dont_touch of I13851: signal is true;
	signal I13852: std_logic; attribute dont_touch of I13852: signal is true;
	signal I13857: std_logic; attribute dont_touch of I13857: signal is true;
	signal I13862: std_logic; attribute dont_touch of I13862: signal is true;
	signal I13872: std_logic; attribute dont_touch of I13872: signal is true;
	signal I13875: std_logic; attribute dont_touch of I13875: signal is true;
	signal I13889: std_logic; attribute dont_touch of I13889: signal is true;
	signal I13892: std_logic; attribute dont_touch of I13892: signal is true;
	signal I13906: std_logic; attribute dont_touch of I13906: signal is true;
	signal I13937: std_logic; attribute dont_touch of I13937: signal is true;
	signal I13968: std_logic; attribute dont_touch of I13968: signal is true;
	signal I13979: std_logic; attribute dont_touch of I13979: signal is true;
	signal I13990: std_logic; attribute dont_touch of I13990: signal is true;
	signal I13995: std_logic; attribute dont_touch of I13995: signal is true;
	signal I14006: std_logic; attribute dont_touch of I14006: signal is true;
	signal I14016: std_logic; attribute dont_touch of I14016: signal is true;
	signal I14033: std_logic; attribute dont_touch of I14033: signal is true;
	signal I14046: std_logic; attribute dont_touch of I14046: signal is true;
	signal I14050: std_logic; attribute dont_touch of I14050: signal is true;
	signal I14054: std_logic; attribute dont_touch of I14054: signal is true;
	signal I14069: std_logic; attribute dont_touch of I14069: signal is true;
	signal I14079: std_logic; attribute dont_touch of I14079: signal is true;
	signal I14119: std_logic; attribute dont_touch of I14119: signal is true;
	signal I14158: std_logic; attribute dont_touch of I14158: signal is true;
	signal I14169: std_logic; attribute dont_touch of I14169: signal is true;
	signal I14170: std_logic; attribute dont_touch of I14170: signal is true;
	signal I14171: std_logic; attribute dont_touch of I14171: signal is true;
	signal I14185: std_logic; attribute dont_touch of I14185: signal is true;
	signal I14186: std_logic; attribute dont_touch of I14186: signal is true;
	signal I14187: std_logic; attribute dont_touch of I14187: signal is true;
	signal I14192: std_logic; attribute dont_touch of I14192: signal is true;
	signal I14198: std_logic; attribute dont_touch of I14198: signal is true;
	signal I14204: std_logic; attribute dont_touch of I14204: signal is true;
	signal I14205: std_logic; attribute dont_touch of I14205: signal is true;
	signal I14206: std_logic; attribute dont_touch of I14206: signal is true;
	signal I14211: std_logic; attribute dont_touch of I14211: signal is true;
	signal I14212: std_logic; attribute dont_touch of I14212: signal is true;
	signal I14213: std_logic; attribute dont_touch of I14213: signal is true;
	signal I14222: std_logic; attribute dont_touch of I14222: signal is true;
	signal I14225: std_logic; attribute dont_touch of I14225: signal is true;
	signal I14228: std_logic; attribute dont_touch of I14228: signal is true;
	signal I14229: std_logic; attribute dont_touch of I14229: signal is true;
	signal I14230: std_logic; attribute dont_touch of I14230: signal is true;
	signal I14241: std_logic; attribute dont_touch of I14241: signal is true;
	signal I14247: std_logic; attribute dont_touch of I14247: signal is true;
	signal I14248: std_logic; attribute dont_touch of I14248: signal is true;
	signal I14249: std_logic; attribute dont_touch of I14249: signal is true;
	signal I14257: std_logic; attribute dont_touch of I14257: signal is true;
	signal I14258: std_logic; attribute dont_touch of I14258: signal is true;
	signal I14259: std_logic; attribute dont_touch of I14259: signal is true;
	signal I14267: std_logic; attribute dont_touch of I14267: signal is true;
	signal I14271: std_logic; attribute dont_touch of I14271: signal is true;
	signal I14275: std_logic; attribute dont_touch of I14275: signal is true;
	signal I14276: std_logic; attribute dont_touch of I14276: signal is true;
	signal I14277: std_logic; attribute dont_touch of I14277: signal is true;
	signal I14289: std_logic; attribute dont_touch of I14289: signal is true;
	signal I14290: std_logic; attribute dont_touch of I14290: signal is true;
	signal I14291: std_logic; attribute dont_touch of I14291: signal is true;
	signal I14301: std_logic; attribute dont_touch of I14301: signal is true;
	signal I14305: std_logic; attribute dont_touch of I14305: signal is true;
	signal I14326: std_logic; attribute dont_touch of I14326: signal is true;
	signal I14330: std_logic; attribute dont_touch of I14330: signal is true;
	signal I14331: std_logic; attribute dont_touch of I14331: signal is true;
	signal I14332: std_logic; attribute dont_touch of I14332: signal is true;
	signal I14346: std_logic; attribute dont_touch of I14346: signal is true;
	signal I14350: std_logic; attribute dont_touch of I14350: signal is true;
	signal I14351: std_logic; attribute dont_touch of I14351: signal is true;
	signal I14352: std_logic; attribute dont_touch of I14352: signal is true;
	signal I14365: std_logic; attribute dont_touch of I14365: signal is true;
	signal I14368: std_logic; attribute dont_touch of I14368: signal is true;
	signal I14369: std_logic; attribute dont_touch of I14369: signal is true;
	signal I14370: std_logic; attribute dont_touch of I14370: signal is true;
	signal I14381: std_logic; attribute dont_touch of I14381: signal is true;
	signal I14395: std_logic; attribute dont_touch of I14395: signal is true;
	signal I14398: std_logic; attribute dont_touch of I14398: signal is true;
	signal I14399: std_logic; attribute dont_touch of I14399: signal is true;
	signal I14400: std_logic; attribute dont_touch of I14400: signal is true;
	signal I14409: std_logic; attribute dont_touch of I14409: signal is true;
	signal I14424: std_logic; attribute dont_touch of I14424: signal is true;
	signal I14427: std_logic; attribute dont_touch of I14427: signal is true;
	signal I14428: std_logic; attribute dont_touch of I14428: signal is true;
	signal I14429: std_logic; attribute dont_touch of I14429: signal is true;
	signal I14450: std_logic; attribute dont_touch of I14450: signal is true;
	signal I14455: std_logic; attribute dont_touch of I14455: signal is true;
	signal I14475: std_logic; attribute dont_touch of I14475: signal is true;
	signal I14480: std_logic; attribute dont_touch of I14480: signal is true;
	signal I14481: std_logic; attribute dont_touch of I14481: signal is true;
	signal I14482: std_logic; attribute dont_touch of I14482: signal is true;
	signal I14497: std_logic; attribute dont_touch of I14497: signal is true;
	signal I14498: std_logic; attribute dont_touch of I14498: signal is true;
	signal I14499: std_logic; attribute dont_touch of I14499: signal is true;
	signal I14505: std_logic; attribute dont_touch of I14505: signal is true;
	signal I14508: std_logic; attribute dont_touch of I14508: signal is true;
	signal I14509: std_logic; attribute dont_touch of I14509: signal is true;
	signal I14510: std_logic; attribute dont_touch of I14510: signal is true;
	signal I14516: std_logic; attribute dont_touch of I14516: signal is true;
	signal I14517: std_logic; attribute dont_touch of I14517: signal is true;
	signal I14518: std_logic; attribute dont_touch of I14518: signal is true;
	signal I14530: std_logic; attribute dont_touch of I14530: signal is true;
	signal I14531: std_logic; attribute dont_touch of I14531: signal is true;
	signal I14532: std_logic; attribute dont_touch of I14532: signal is true;
	signal I14537: std_logic; attribute dont_touch of I14537: signal is true;
	signal I14550: std_logic; attribute dont_touch of I14550: signal is true;
	signal I14563: std_logic; attribute dont_touch of I14563: signal is true;
	signal I14567: std_logic; attribute dont_touch of I14567: signal is true;
	signal I14570: std_logic; attribute dont_touch of I14570: signal is true;
	signal I14576: std_logic; attribute dont_touch of I14576: signal is true;
	signal I14579: std_logic; attribute dont_touch of I14579: signal is true;
	signal I14584: std_logic; attribute dont_touch of I14584: signal is true;
	signal I14589: std_logic; attribute dont_touch of I14589: signal is true;
	signal I14593: std_logic; attribute dont_touch of I14593: signal is true;
	signal I14602: std_logic; attribute dont_touch of I14602: signal is true;
	signal I14609: std_logic; attribute dont_touch of I14609: signal is true;
	signal I14610: std_logic; attribute dont_touch of I14610: signal is true;
	signal I14611: std_logic; attribute dont_touch of I14611: signal is true;
	signal I14619: std_logic; attribute dont_touch of I14619: signal is true;
	signal I14623: std_logic; attribute dont_touch of I14623: signal is true;
	signal I14630: std_logic; attribute dont_touch of I14630: signal is true;
	signal I14633: std_logic; attribute dont_touch of I14633: signal is true;
	signal I14644: std_logic; attribute dont_touch of I14644: signal is true;
	signal I14647: std_logic; attribute dont_touch of I14647: signal is true;
	signal I14650: std_logic; attribute dont_touch of I14650: signal is true;
	signal I14653: std_logic; attribute dont_touch of I14653: signal is true;
	signal I14660: std_logic; attribute dont_touch of I14660: signal is true;
	signal I14663: std_logic; attribute dont_touch of I14663: signal is true;
	signal I14668: std_logic; attribute dont_touch of I14668: signal is true;
	signal I14671: std_logic; attribute dont_touch of I14671: signal is true;
	signal I14679: std_logic; attribute dont_touch of I14679: signal is true;
	signal I14684: std_logic; attribute dont_touch of I14684: signal is true;
	signal I14687: std_logic; attribute dont_touch of I14687: signal is true;
	signal I14690: std_logic; attribute dont_touch of I14690: signal is true;
	signal I14702: std_logic; attribute dont_touch of I14702: signal is true;
	signal I14705: std_logic; attribute dont_touch of I14705: signal is true;
	signal I14708: std_logic; attribute dont_touch of I14708: signal is true;
	signal I14712: std_logic; attribute dont_touch of I14712: signal is true;
	signal I14713: std_logic; attribute dont_touch of I14713: signal is true;
	signal I14714: std_logic; attribute dont_touch of I14714: signal is true;
	signal I14727: std_logic; attribute dont_touch of I14727: signal is true;
	signal I14730: std_logic; attribute dont_touch of I14730: signal is true;
	signal I14733: std_logic; attribute dont_touch of I14733: signal is true;
	signal I14734: std_logic; attribute dont_touch of I14734: signal is true;
	signal I14735: std_logic; attribute dont_touch of I14735: signal is true;
	signal I14742: std_logic; attribute dont_touch of I14742: signal is true;
	signal I14745: std_logic; attribute dont_touch of I14745: signal is true;
	signal I14749: std_logic; attribute dont_touch of I14749: signal is true;
	signal I14761: std_logic; attribute dont_touch of I14761: signal is true;
	signal I14764: std_logic; attribute dont_touch of I14764: signal is true;
	signal I14765: std_logic; attribute dont_touch of I14765: signal is true;
	signal I14766: std_logic; attribute dont_touch of I14766: signal is true;
	signal I14773: std_logic; attribute dont_touch of I14773: signal is true;
	signal I14788: std_logic; attribute dont_touch of I14788: signal is true;
	signal I14789: std_logic; attribute dont_touch of I14789: signal is true;
	signal I14790: std_logic; attribute dont_touch of I14790: signal is true;
	signal I14797: std_logic; attribute dont_touch of I14797: signal is true;
	signal I14800: std_logic; attribute dont_touch of I14800: signal is true;
	signal I14816: std_logic; attribute dont_touch of I14816: signal is true;
	signal I14817: std_logic; attribute dont_touch of I14817: signal is true;
	signal I14818: std_logic; attribute dont_touch of I14818: signal is true;
	signal I14823: std_logic; attribute dont_touch of I14823: signal is true;
	signal I14827: std_logic; attribute dont_touch of I14827: signal is true;
	signal I14830: std_logic; attribute dont_touch of I14830: signal is true;
	signal I14833: std_logic; attribute dont_touch of I14833: signal is true;
	signal I14836: std_logic; attribute dont_touch of I14836: signal is true;
	signal I14839: std_logic; attribute dont_touch of I14839: signal is true;
	signal I14853: std_logic; attribute dont_touch of I14853: signal is true;
	signal I14854: std_logic; attribute dont_touch of I14854: signal is true;
	signal I14855: std_logic; attribute dont_touch of I14855: signal is true;
	signal I14862: std_logic; attribute dont_touch of I14862: signal is true;
	signal I14866: std_logic; attribute dont_touch of I14866: signal is true;
	signal I14883: std_logic; attribute dont_touch of I14883: signal is true;
	signal I14884: std_logic; attribute dont_touch of I14884: signal is true;
	signal I14885: std_logic; attribute dont_touch of I14885: signal is true;
	signal I14893: std_logic; attribute dont_touch of I14893: signal is true;
	signal I14896: std_logic; attribute dont_touch of I14896: signal is true;
	signal I14899: std_logic; attribute dont_touch of I14899: signal is true;
	signal I14902: std_logic; attribute dont_touch of I14902: signal is true;
	signal I14905: std_logic; attribute dont_touch of I14905: signal is true;
	signal I14923: std_logic; attribute dont_touch of I14923: signal is true;
	signal I14924: std_logic; attribute dont_touch of I14924: signal is true;
	signal I14925: std_logic; attribute dont_touch of I14925: signal is true;
	signal I14932: std_logic; attribute dont_touch of I14932: signal is true;
	signal I14935: std_logic; attribute dont_touch of I14935: signal is true;
	signal I14939: std_logic; attribute dont_touch of I14939: signal is true;
	signal I14955: std_logic; attribute dont_touch of I14955: signal is true;
	signal I14956: std_logic; attribute dont_touch of I14956: signal is true;
	signal I14957: std_logic; attribute dont_touch of I14957: signal is true;
	signal I14964: std_logic; attribute dont_touch of I14964: signal is true;
	signal I14967: std_logic; attribute dont_touch of I14967: signal is true;
	signal I14970: std_logic; attribute dont_touch of I14970: signal is true;
	signal I14991: std_logic; attribute dont_touch of I14991: signal is true;
	signal I14992: std_logic; attribute dont_touch of I14992: signal is true;
	signal I14993: std_logic; attribute dont_touch of I14993: signal is true;
	signal I14999: std_logic; attribute dont_touch of I14999: signal is true;
	signal I15002: std_logic; attribute dont_touch of I15002: signal is true;
	signal I15003: std_logic; attribute dont_touch of I15003: signal is true;
	signal I15004: std_logic; attribute dont_touch of I15004: signal is true;
	signal I15030: std_logic; attribute dont_touch of I15030: signal is true;
	signal I15033: std_logic; attribute dont_touch of I15033: signal is true;
	signal I15036: std_logic; attribute dont_touch of I15036: signal is true;
	signal I15041: std_logic; attribute dont_touch of I15041: signal is true;
	signal I15042: std_logic; attribute dont_touch of I15042: signal is true;
	signal I15043: std_logic; attribute dont_touch of I15043: signal is true;
	signal I15051: std_logic; attribute dont_touch of I15051: signal is true;
	signal I15052: std_logic; attribute dont_touch of I15052: signal is true;
	signal I15053: std_logic; attribute dont_touch of I15053: signal is true;
	signal I15070: std_logic; attribute dont_touch of I15070: signal is true;
	signal I15073: std_logic; attribute dont_touch of I15073: signal is true;
	signal I15078: std_logic; attribute dont_touch of I15078: signal is true;
	signal I15079: std_logic; attribute dont_touch of I15079: signal is true;
	signal I15080: std_logic; attribute dont_touch of I15080: signal is true;
	signal I15087: std_logic; attribute dont_touch of I15087: signal is true;
	signal I15088: std_logic; attribute dont_touch of I15088: signal is true;
	signal I15089: std_logic; attribute dont_touch of I15089: signal is true;
	signal I15102: std_logic; attribute dont_touch of I15102: signal is true;
	signal I15105: std_logic; attribute dont_touch of I15105: signal is true;
	signal I15106: std_logic; attribute dont_touch of I15106: signal is true;
	signal I15107: std_logic; attribute dont_touch of I15107: signal is true;
	signal I15121: std_logic; attribute dont_touch of I15121: signal is true;
	signal I15122: std_logic; attribute dont_touch of I15122: signal is true;
	signal I15123: std_logic; attribute dont_touch of I15123: signal is true;
	signal I15128: std_logic; attribute dont_touch of I15128: signal is true;
	signal I15129: std_logic; attribute dont_touch of I15129: signal is true;
	signal I15130: std_logic; attribute dont_touch of I15130: signal is true;
	signal I15144: std_logic; attribute dont_touch of I15144: signal is true;
	signal I15147: std_logic; attribute dont_touch of I15147: signal is true;
	signal I15148: std_logic; attribute dont_touch of I15148: signal is true;
	signal I15149: std_logic; attribute dont_touch of I15149: signal is true;
	signal I15162: std_logic; attribute dont_touch of I15162: signal is true;
	signal I15166: std_logic; attribute dont_touch of I15166: signal is true;
	signal I15167: std_logic; attribute dont_touch of I15167: signal is true;
	signal I15168: std_logic; attribute dont_touch of I15168: signal is true;
	signal I15174: std_logic; attribute dont_touch of I15174: signal is true;
	signal I15175: std_logic; attribute dont_touch of I15175: signal is true;
	signal I15176: std_logic; attribute dont_touch of I15176: signal is true;
	signal I15190: std_logic; attribute dont_touch of I15190: signal is true;
	signal I15193: std_logic; attribute dont_touch of I15193: signal is true;
	signal I15194: std_logic; attribute dont_touch of I15194: signal is true;
	signal I15195: std_logic; attribute dont_touch of I15195: signal is true;
	signal I15205: std_logic; attribute dont_touch of I15205: signal is true;
	signal I15208: std_logic; attribute dont_touch of I15208: signal is true;
	signal I15212: std_logic; attribute dont_touch of I15212: signal is true;
	signal I15213: std_logic; attribute dont_touch of I15213: signal is true;
	signal I15214: std_logic; attribute dont_touch of I15214: signal is true;
	signal I15223: std_logic; attribute dont_touch of I15223: signal is true;
	signal I15238: std_logic; attribute dont_touch of I15238: signal is true;
	signal I15241: std_logic; attribute dont_touch of I15241: signal is true;
	signal I15242: std_logic; attribute dont_touch of I15242: signal is true;
	signal I15243: std_logic; attribute dont_touch of I15243: signal is true;
	signal I15250: std_logic; attribute dont_touch of I15250: signal is true;
	signal I15253: std_logic; attribute dont_touch of I15253: signal is true;
	signal I15254: std_logic; attribute dont_touch of I15254: signal is true;
	signal I15255: std_logic; attribute dont_touch of I15255: signal is true;
	signal I15262: std_logic; attribute dont_touch of I15262: signal is true;
	signal I15263: std_logic; attribute dont_touch of I15263: signal is true;
	signal I15264: std_logic; attribute dont_touch of I15264: signal is true;
	signal I15284: std_logic; attribute dont_touch of I15284: signal is true;
	signal I15287: std_logic; attribute dont_touch of I15287: signal is true;
	signal I15288: std_logic; attribute dont_touch of I15288: signal is true;
	signal I15289: std_logic; attribute dont_touch of I15289: signal is true;
	signal I15295: std_logic; attribute dont_touch of I15295: signal is true;
	signal I15298: std_logic; attribute dont_touch of I15298: signal is true;
	signal I15299: std_logic; attribute dont_touch of I15299: signal is true;
	signal I15300: std_logic; attribute dont_touch of I15300: signal is true;
	signal I15306: std_logic; attribute dont_touch of I15306: signal is true;
	signal I15307: std_logic; attribute dont_touch of I15307: signal is true;
	signal I15308: std_logic; attribute dont_touch of I15308: signal is true;
	signal I15316: std_logic; attribute dont_touch of I15316: signal is true;
	signal I15333: std_logic; attribute dont_touch of I15333: signal is true;
	signal I15334: std_logic; attribute dont_touch of I15334: signal is true;
	signal I15335: std_logic; attribute dont_touch of I15335: signal is true;
	signal I15340: std_logic; attribute dont_touch of I15340: signal is true;
	signal I15341: std_logic; attribute dont_touch of I15341: signal is true;
	signal I15342: std_logic; attribute dont_touch of I15342: signal is true;
	signal I15363: std_logic; attribute dont_touch of I15363: signal is true;
	signal I15364: std_logic; attribute dont_touch of I15364: signal is true;
	signal I15365: std_logic; attribute dont_touch of I15365: signal is true;
	signal I15382: std_logic; attribute dont_touch of I15382: signal is true;
	signal I15448: std_logic; attribute dont_touch of I15448: signal is true;
	signal I15474: std_logic; attribute dont_touch of I15474: signal is true;
	signal I15494: std_logic; attribute dont_touch of I15494: signal is true;
	signal I15533: std_logic; attribute dont_touch of I15533: signal is true;
	signal I15536: std_logic; attribute dont_touch of I15536: signal is true;
	signal I15542: std_logic; attribute dont_touch of I15542: signal is true;
	signal I15550: std_logic; attribute dont_touch of I15550: signal is true;
	signal I15556: std_logic; attribute dont_touch of I15556: signal is true;
	signal I15564: std_logic; attribute dont_touch of I15564: signal is true;
	signal I15569: std_logic; attribute dont_touch of I15569: signal is true;
	signal I15572: std_logic; attribute dont_touch of I15572: signal is true;
	signal I15577: std_logic; attribute dont_touch of I15577: signal is true;
	signal I15587: std_logic; attribute dont_touch of I15587: signal is true;
	signal I15590: std_logic; attribute dont_touch of I15590: signal is true;
	signal I15593: std_logic; attribute dont_touch of I15593: signal is true;
	signal I15600: std_logic; attribute dont_touch of I15600: signal is true;
	signal I15609: std_logic; attribute dont_touch of I15609: signal is true;
	signal I15617: std_logic; attribute dont_touch of I15617: signal is true;
	signal I15620: std_logic; attribute dont_touch of I15620: signal is true;
	signal I15623: std_logic; attribute dont_touch of I15623: signal is true;
	signal I15626: std_logic; attribute dont_touch of I15626: signal is true;
	signal I15633: std_logic; attribute dont_touch of I15633: signal is true;
	signal I15636: std_logic; attribute dont_touch of I15636: signal is true;
	signal I15647: std_logic; attribute dont_touch of I15647: signal is true;
	signal I15650: std_logic; attribute dont_touch of I15650: signal is true;
	signal I15663: std_logic; attribute dont_touch of I15663: signal is true;
	signal I15667: std_logic; attribute dont_touch of I15667: signal is true;
	signal I15677: std_logic; attribute dont_touch of I15677: signal is true;
	signal I15682: std_logic; attribute dont_touch of I15682: signal is true;
	signal I15697: std_logic; attribute dont_touch of I15697: signal is true;
	signal I15702: std_logic; attribute dont_touch of I15702: signal is true;
	signal I15705: std_logic; attribute dont_touch of I15705: signal is true;
	signal I15717: std_logic; attribute dont_touch of I15717: signal is true;
	signal I15727: std_logic; attribute dont_touch of I15727: signal is true;
	signal I15732: std_logic; attribute dont_touch of I15732: signal is true;
	signal I15736: std_logic; attribute dont_touch of I15736: signal is true;
	signal I15765: std_logic; attribute dont_touch of I15765: signal is true;
	signal I15773: std_logic; attribute dont_touch of I15773: signal is true;
	signal I15782: std_logic; attribute dont_touch of I15782: signal is true;
	signal I15788: std_logic; attribute dont_touch of I15788: signal is true;
	signal I15800: std_logic; attribute dont_touch of I15800: signal is true;
	signal I15811: std_logic; attribute dont_touch of I15811: signal is true;
	signal I15814: std_logic; attribute dont_touch of I15814: signal is true;
	signal I15821: std_logic; attribute dont_touch of I15821: signal is true;
	signal I15824: std_logic; attribute dont_touch of I15824: signal is true;
	signal I15831: std_logic; attribute dont_touch of I15831: signal is true;
	signal I15834: std_logic; attribute dont_touch of I15834: signal is true;
	signal I15837: std_logic; attribute dont_touch of I15837: signal is true;
	signal I15843: std_logic; attribute dont_touch of I15843: signal is true;
	signal I15846: std_logic; attribute dont_touch of I15846: signal is true;
	signal I15862: std_logic; attribute dont_touch of I15862: signal is true;
	signal I15869: std_logic; attribute dont_touch of I15869: signal is true;
	signal I15872: std_logic; attribute dont_touch of I15872: signal is true;
	signal I15878: std_logic; attribute dont_touch of I15878: signal is true;
	signal I15893: std_logic; attribute dont_touch of I15893: signal is true;
	signal I15906: std_logic; attribute dont_touch of I15906: signal is true;
	signal I15915: std_logic; attribute dont_touch of I15915: signal is true;
	signal I15918: std_logic; attribute dont_touch of I15918: signal is true;
	signal I15921: std_logic; attribute dont_touch of I15921: signal is true;
	signal I15929: std_logic; attribute dont_touch of I15929: signal is true;
	signal I15932: std_logic; attribute dont_touch of I15932: signal is true;
	signal I15937: std_logic; attribute dont_touch of I15937: signal is true;
	signal I15942: std_logic; attribute dont_touch of I15942: signal is true;
	signal I15954: std_logic; attribute dont_touch of I15954: signal is true;
	signal I15981: std_logic; attribute dont_touch of I15981: signal is true;
	signal I15987: std_logic; attribute dont_touch of I15987: signal is true;
	signal I16010: std_logic; attribute dont_touch of I16010: signal is true;
	signal I16024: std_logic; attribute dont_touch of I16024: signal is true;
	signal I16028: std_logic; attribute dont_touch of I16028: signal is true;
	signal I16040: std_logic; attribute dont_touch of I16040: signal is true;
	signal I16057: std_logic; attribute dont_touch of I16057: signal is true;
	signal I16077: std_logic; attribute dont_touch of I16077: signal is true;
	signal I16090: std_logic; attribute dont_touch of I16090: signal is true;
	signal I16102: std_logic; attribute dont_touch of I16102: signal is true;
	signal I16111: std_logic; attribute dont_touch of I16111: signal is true;
	signal I16117: std_logic; attribute dont_touch of I16117: signal is true;
	signal I16120: std_logic; attribute dont_touch of I16120: signal is true;
	signal I16129: std_logic; attribute dont_touch of I16129: signal is true;
	signal I16135: std_logic; attribute dont_touch of I16135: signal is true;
	signal I16143: std_logic; attribute dont_touch of I16143: signal is true;
	signal I16150: std_logic; attribute dont_touch of I16150: signal is true;
	signal I16160: std_logic; attribute dont_touch of I16160: signal is true;
	signal I16163: std_logic; attribute dont_touch of I16163: signal is true;
	signal I16168: std_logic; attribute dont_touch of I16168: signal is true;
	signal I16181: std_logic; attribute dont_touch of I16181: signal is true;
	signal I16193: std_logic; attribute dont_touch of I16193: signal is true;
	signal I16201: std_logic; attribute dont_touch of I16201: signal is true;
	signal I16217: std_logic; attribute dont_touch of I16217: signal is true;
	signal I16231: std_logic; attribute dont_touch of I16231: signal is true;
	signal I16246: std_logic; attribute dont_touch of I16246: signal is true;
	signal I16289: std_logic; attribute dont_touch of I16289: signal is true;
	signal I16328: std_logic; attribute dont_touch of I16328: signal is true;
	signal I16345: std_logic; attribute dont_touch of I16345: signal is true;
	signal I16357: std_logic; attribute dont_touch of I16357: signal is true;
	signal I16371: std_logic; attribute dont_touch of I16371: signal is true;
	signal I16391: std_logic; attribute dont_touch of I16391: signal is true;
	signal I16401: std_logic; attribute dont_touch of I16401: signal is true;
	signal I16417: std_logic; attribute dont_touch of I16417: signal is true;
	signal I16438: std_logic; attribute dont_touch of I16438: signal is true;
	signal I16452: std_logic; attribute dont_touch of I16452: signal is true;
	signal I16455: std_logic; attribute dont_touch of I16455: signal is true;
	signal I16460: std_logic; attribute dont_touch of I16460: signal is true;
	signal I16468: std_logic; attribute dont_touch of I16468: signal is true;
	signal I16471: std_logic; attribute dont_touch of I16471: signal is true;
	signal I16476: std_logic; attribute dont_touch of I16476: signal is true;
	signal I16479: std_logic; attribute dont_touch of I16479: signal is true;
	signal I16486: std_logic; attribute dont_touch of I16486: signal is true;
	signal I16489: std_logic; attribute dont_touch of I16489: signal is true;
	signal I16492: std_logic; attribute dont_touch of I16492: signal is true;
	signal I16498: std_logic; attribute dont_touch of I16498: signal is true;
	signal I16502: std_logic; attribute dont_touch of I16502: signal is true;
	signal I16512: std_logic; attribute dont_touch of I16512: signal is true;
	signal I16515: std_logic; attribute dont_touch of I16515: signal is true;
	signal I16521: std_logic; attribute dont_touch of I16521: signal is true;
	signal I16526: std_logic; attribute dont_touch of I16526: signal is true;
	signal I16535: std_logic; attribute dont_touch of I16535: signal is true;
	signal I16538: std_logic; attribute dont_touch of I16538: signal is true;
	signal I16541: std_logic; attribute dont_touch of I16541: signal is true;
	signal I16544: std_logic; attribute dont_touch of I16544: signal is true;
	signal I16555: std_logic; attribute dont_touch of I16555: signal is true;
	signal I16564: std_logic; attribute dont_touch of I16564: signal is true;
	signal I16575: std_logic; attribute dont_touch of I16575: signal is true;
	signal I16579: std_logic; attribute dont_touch of I16579: signal is true;
	signal I16590: std_logic; attribute dont_touch of I16590: signal is true;
	signal I16593: std_logic; attribute dont_touch of I16593: signal is true;
	signal I16596: std_logic; attribute dont_touch of I16596: signal is true;
	signal I16606: std_logic; attribute dont_touch of I16606: signal is true;
	signal I16610: std_logic; attribute dont_touch of I16610: signal is true;
	signal I16613: std_logic; attribute dont_touch of I16613: signal is true;
	signal I16618: std_logic; attribute dont_touch of I16618: signal is true;
	signal I16626: std_logic; attribute dont_touch of I16626: signal is true;
	signal I16629: std_logic; attribute dont_touch of I16629: signal is true;
	signal I16639: std_logic; attribute dont_touch of I16639: signal is true;
	signal I16646: std_logic; attribute dont_touch of I16646: signal is true;
	signal I16651: std_logic; attribute dont_touch of I16651: signal is true;
	signal I16660: std_logic; attribute dont_touch of I16660: signal is true;
	signal I16663: std_logic; attribute dont_touch of I16663: signal is true;
	signal I16671: std_logic; attribute dont_touch of I16671: signal is true;
	signal I16676: std_logic; attribute dont_touch of I16676: signal is true;
	signal I16679: std_logic; attribute dont_touch of I16679: signal is true;
	signal I16688: std_logic; attribute dont_touch of I16688: signal is true;
	signal I16695: std_logic; attribute dont_touch of I16695: signal is true;
	signal I16698: std_logic; attribute dont_touch of I16698: signal is true;
	signal I16709: std_logic; attribute dont_touch of I16709: signal is true;
	signal I16713: std_logic; attribute dont_touch of I16713: signal is true;
	signal I16721: std_logic; attribute dont_touch of I16721: signal is true;
	signal I16724: std_logic; attribute dont_touch of I16724: signal is true;
	signal I16733: std_logic; attribute dont_touch of I16733: signal is true;
	signal I16741: std_logic; attribute dont_touch of I16741: signal is true;
	signal I16747: std_logic; attribute dont_touch of I16747: signal is true;
	signal I16755: std_logic; attribute dont_touch of I16755: signal is true;
	signal I16762: std_logic; attribute dont_touch of I16762: signal is true;
	signal I16770: std_logic; attribute dont_touch of I16770: signal is true;
	signal I16775: std_logic; attribute dont_touch of I16775: signal is true;
	signal I16778: std_logic; attribute dont_touch of I16778: signal is true;
	signal I16779: std_logic; attribute dont_touch of I16779: signal is true;
	signal I16780: std_logic; attribute dont_touch of I16780: signal is true;
	signal I16795: std_logic; attribute dont_touch of I16795: signal is true;
	signal I16803: std_logic; attribute dont_touch of I16803: signal is true;
	signal I16821: std_logic; attribute dont_touch of I16821: signal is true;
	signal I16829: std_logic; attribute dont_touch of I16829: signal is true;
	signal I16847: std_logic; attribute dont_touch of I16847: signal is true;
	signal I16855: std_logic; attribute dont_touch of I16855: signal is true;
	signal I16875: std_logic; attribute dont_touch of I16875: signal is true;
	signal I16898: std_logic; attribute dont_touch of I16898: signal is true;
	signal I16917: std_logic; attribute dont_touch of I16917: signal is true;
	signal I16969: std_logic; attribute dont_touch of I16969: signal is true;
	signal I17008: std_logic; attribute dont_touch of I17008: signal is true;
	signal I17094: std_logic; attribute dont_touch of I17094: signal is true;
	signal I17098: std_logic; attribute dont_touch of I17098: signal is true;
	signal I17101: std_logic; attribute dont_touch of I17101: signal is true;
	signal I17104: std_logic; attribute dont_touch of I17104: signal is true;
	signal I17108: std_logic; attribute dont_touch of I17108: signal is true;
	signal I17111: std_logic; attribute dont_touch of I17111: signal is true;
	signal I17114: std_logic; attribute dont_touch of I17114: signal is true;
	signal I17118: std_logic; attribute dont_touch of I17118: signal is true;
	signal I17121: std_logic; attribute dont_touch of I17121: signal is true;
	signal I17125: std_logic; attribute dont_touch of I17125: signal is true;
	signal I17128: std_logic; attribute dont_touch of I17128: signal is true;
	signal I17131: std_logic; attribute dont_touch of I17131: signal is true;
	signal I17136: std_logic; attribute dont_touch of I17136: signal is true;
	signal I17140: std_logic; attribute dont_touch of I17140: signal is true;
	signal I17143: std_logic; attribute dont_touch of I17143: signal is true;
	signal I17148: std_logic; attribute dont_touch of I17148: signal is true;
	signal I17154: std_logic; attribute dont_touch of I17154: signal is true;
	signal I17159: std_logic; attribute dont_touch of I17159: signal is true;
	signal I17166: std_logic; attribute dont_touch of I17166: signal is true;
	signal I17173: std_logic; attribute dont_touch of I17173: signal is true;
	signal I17181: std_logic; attribute dont_touch of I17181: signal is true;
	signal I17188: std_logic; attribute dont_touch of I17188: signal is true;
	signal I17198: std_logic; attribute dont_touch of I17198: signal is true;
	signal I17207: std_logic; attribute dont_touch of I17207: signal is true;
	signal I17228: std_logic; attribute dont_touch of I17228: signal is true;
	signal I17249: std_logic; attribute dont_touch of I17249: signal is true;
	signal I17276: std_logic; attribute dont_touch of I17276: signal is true;
	signal I17302: std_logic; attribute dont_touch of I17302: signal is true;
	signal I17314: std_logic; attribute dont_touch of I17314: signal is true;
	signal I17324: std_logic; attribute dont_touch of I17324: signal is true;
	signal I17355: std_logic; attribute dont_touch of I17355: signal is true;
	signal I17374: std_logic; attribute dont_touch of I17374: signal is true;
	signal I17379: std_logic; attribute dont_touch of I17379: signal is true;
	signal I17380: std_logic; attribute dont_touch of I17380: signal is true;
	signal I17381: std_logic; attribute dont_touch of I17381: signal is true;
	signal I17392: std_logic; attribute dont_touch of I17392: signal is true;
	signal I17395: std_logic; attribute dont_touch of I17395: signal is true;
	signal I17401: std_logic; attribute dont_touch of I17401: signal is true;
	signal I17404: std_logic; attribute dont_touch of I17404: signal is true;
	signal I17405: std_logic; attribute dont_touch of I17405: signal is true;
	signal I17406: std_logic; attribute dont_touch of I17406: signal is true;
	signal I17416: std_logic; attribute dont_touch of I17416: signal is true;
	signal I17420: std_logic; attribute dont_touch of I17420: signal is true;
	signal I17425: std_logic; attribute dont_touch of I17425: signal is true;
	signal I17436: std_logic; attribute dont_touch of I17436: signal is true;
	signal I17442: std_logic; attribute dont_touch of I17442: signal is true;
	signal I17446: std_logic; attribute dont_touch of I17446: signal is true;
	signal I17447: std_logic; attribute dont_touch of I17447: signal is true;
	signal I17448: std_logic; attribute dont_touch of I17448: signal is true;
	signal I17456: std_logic; attribute dont_touch of I17456: signal is true;
	signal I17460: std_logic; attribute dont_touch of I17460: signal is true;
	signal I17461: std_logic; attribute dont_touch of I17461: signal is true;
	signal I17462: std_logic; attribute dont_touch of I17462: signal is true;
	signal I17471: std_logic; attribute dont_touch of I17471: signal is true;
	signal I17474: std_logic; attribute dont_touch of I17474: signal is true;
	signal I17475: std_logic; attribute dont_touch of I17475: signal is true;
	signal I17476: std_logic; attribute dont_touch of I17476: signal is true;
	signal I17488: std_logic; attribute dont_touch of I17488: signal is true;
	signal I17491: std_logic; attribute dont_touch of I17491: signal is true;
	signal I17494: std_logic; attribute dont_touch of I17494: signal is true;
	signal I17495: std_logic; attribute dont_touch of I17495: signal is true;
	signal I17496: std_logic; attribute dont_touch of I17496: signal is true;
	signal I17507: std_logic; attribute dont_touch of I17507: signal is true;
	signal I17529: std_logic; attribute dont_touch of I17529: signal is true;
	signal I17542: std_logic; attribute dont_touch of I17542: signal is true;
	signal I17552: std_logic; attribute dont_touch of I17552: signal is true;
	signal I17557: std_logic; attribute dont_touch of I17557: signal is true;
	signal I17569: std_logic; attribute dont_touch of I17569: signal is true;
	signal I17575: std_logic; attribute dont_touch of I17575: signal is true;
	signal I17585: std_logic; attribute dont_touch of I17585: signal is true;
	signal I17590: std_logic; attribute dont_touch of I17590: signal is true;
	signal I17606: std_logic; attribute dont_touch of I17606: signal is true;
	signal I17609: std_logic; attribute dont_touch of I17609: signal is true;
	signal I17612: std_logic; attribute dont_touch of I17612: signal is true;
	signal I17615: std_logic; attribute dont_touch of I17615: signal is true;
	signal I17626: std_logic; attribute dont_touch of I17626: signal is true;
	signal I17633: std_logic; attribute dont_touch of I17633: signal is true;
	signal I17636: std_logic; attribute dont_touch of I17636: signal is true;
	signal I17639: std_logic; attribute dont_touch of I17639: signal is true;
	signal I17650: std_logic; attribute dont_touch of I17650: signal is true;
	signal I17653: std_logic; attribute dont_touch of I17653: signal is true;
	signal I17658: std_logic; attribute dont_touch of I17658: signal is true;
	signal I17661: std_logic; attribute dont_touch of I17661: signal is true;
	signal I17668: std_logic; attribute dont_touch of I17668: signal is true;
	signal I17671: std_logic; attribute dont_touch of I17671: signal is true;
	signal I17675: std_logic; attribute dont_touch of I17675: signal is true;
	signal I17679: std_logic; attribute dont_touch of I17679: signal is true;
	signal I17692: std_logic; attribute dont_touch of I17692: signal is true;
	signal I17695: std_logic; attribute dont_touch of I17695: signal is true;
	signal I17699: std_logic; attribute dont_touch of I17699: signal is true;
	signal I17704: std_logic; attribute dont_touch of I17704: signal is true;
	signal I17723: std_logic; attribute dont_touch of I17723: signal is true;
	signal I17733: std_logic; attribute dont_touch of I17733: signal is true;
	signal I17741: std_logic; attribute dont_touch of I17741: signal is true;
	signal I17744: std_logic; attribute dont_touch of I17744: signal is true;
	signal I17747: std_logic; attribute dont_touch of I17747: signal is true;
	signal I17750: std_logic; attribute dont_touch of I17750: signal is true;
	signal I17754: std_logic; attribute dont_touch of I17754: signal is true;
	signal I17763: std_logic; attribute dont_touch of I17763: signal is true;
	signal I17772: std_logic; attribute dont_touch of I17772: signal is true;
	signal I17780: std_logic; attribute dont_touch of I17780: signal is true;
	signal I17783: std_logic; attribute dont_touch of I17783: signal is true;
	signal I17787: std_logic; attribute dont_touch of I17787: signal is true;
	signal I17801: std_logic; attribute dont_touch of I17801: signal is true;
	signal I17808: std_logic; attribute dont_touch of I17808: signal is true;
	signal I17814: std_logic; attribute dont_touch of I17814: signal is true;
	signal I17819: std_logic; attribute dont_touch of I17819: signal is true;
	signal I17834: std_logic; attribute dont_touch of I17834: signal is true;
	signal I17839: std_logic; attribute dont_touch of I17839: signal is true;
	signal I17842: std_logic; attribute dont_touch of I17842: signal is true;
	signal I17852: std_logic; attribute dont_touch of I17852: signal is true;
	signal I17857: std_logic; attribute dont_touch of I17857: signal is true;
	signal I17873: std_logic; attribute dont_touch of I17873: signal is true;
	signal I17876: std_logic; attribute dont_touch of I17876: signal is true;
	signal I17879: std_logic; attribute dont_touch of I17879: signal is true;
	signal I17883: std_logic; attribute dont_touch of I17883: signal is true;
	signal I17884: std_logic; attribute dont_touch of I17884: signal is true;
	signal I17885: std_logic; attribute dont_touch of I17885: signal is true;
	signal I17892: std_logic; attribute dont_touch of I17892: signal is true;
	signal I17901: std_logic; attribute dont_touch of I17901: signal is true;
	signal I17916: std_logic; attribute dont_touch of I17916: signal is true;
	signal I17919: std_logic; attribute dont_touch of I17919: signal is true;
	signal I17923: std_logic; attribute dont_touch of I17923: signal is true;
	signal I17924: std_logic; attribute dont_touch of I17924: signal is true;
	signal I17925: std_logic; attribute dont_touch of I17925: signal is true;
	signal I17932: std_logic; attribute dont_touch of I17932: signal is true;
	signal I17938: std_logic; attribute dont_touch of I17938: signal is true;
	signal I17956: std_logic; attribute dont_touch of I17956: signal is true;
	signal I17964: std_logic; attribute dont_touch of I17964: signal is true;
	signal I17970: std_logic; attribute dont_touch of I17970: signal is true;
	signal I17976: std_logic; attribute dont_touch of I17976: signal is true;
	signal I17989: std_logic; attribute dont_touch of I17989: signal is true;
	signal I17999: std_logic; attribute dont_touch of I17999: signal is true;
	signal I18003: std_logic; attribute dont_touch of I18003: signal is true;
	signal I18006: std_logic; attribute dont_touch of I18006: signal is true;
	signal I18009: std_logic; attribute dont_touch of I18009: signal is true;
	signal I18028: std_logic; attribute dont_touch of I18028: signal is true;
	signal I18031: std_logic; attribute dont_touch of I18031: signal is true;
	signal I18034: std_logic; attribute dont_touch of I18034: signal is true;
	signal I18048: std_logic; attribute dont_touch of I18048: signal is true;
	signal I18051: std_logic; attribute dont_touch of I18051: signal is true;
	signal I18060: std_logic; attribute dont_touch of I18060: signal is true;
	signal I18063: std_logic; attribute dont_touch of I18063: signal is true;
	signal I18066: std_logic; attribute dont_touch of I18066: signal is true;
	signal I18071: std_logic; attribute dont_touch of I18071: signal is true;
	signal I18078: std_logic; attribute dont_touch of I18078: signal is true;
	signal I18083: std_logic; attribute dont_touch of I18083: signal is true;
	signal I18086: std_logic; attribute dont_touch of I18086: signal is true;
	signal I18089: std_logic; attribute dont_touch of I18089: signal is true;
	signal I18092: std_logic; attribute dont_touch of I18092: signal is true;
	signal I18101: std_logic; attribute dont_touch of I18101: signal is true;
	signal I18104: std_logic; attribute dont_touch of I18104: signal is true;
	signal I18107: std_logic; attribute dont_touch of I18107: signal is true;
	signal I18114: std_logic; attribute dont_touch of I18114: signal is true;
	signal I18117: std_logic; attribute dont_touch of I18117: signal is true;
	signal I18120: std_logic; attribute dont_touch of I18120: signal is true;
	signal I18125: std_logic; attribute dont_touch of I18125: signal is true;
	signal I18131: std_logic; attribute dont_touch of I18131: signal is true;
	signal I18135: std_logic; attribute dont_touch of I18135: signal is true;
	signal I18138: std_logic; attribute dont_touch of I18138: signal is true;
	signal I18143: std_logic; attribute dont_touch of I18143: signal is true;
	signal I18148: std_logic; attribute dont_touch of I18148: signal is true;
	signal I18151: std_logic; attribute dont_touch of I18151: signal is true;
	signal I18154: std_logic; attribute dont_touch of I18154: signal is true;
	signal I18160: std_logic; attribute dont_touch of I18160: signal is true;
	signal I18165: std_logic; attribute dont_touch of I18165: signal is true;
	signal I18168: std_logic; attribute dont_touch of I18168: signal is true;
	signal I18177: std_logic; attribute dont_touch of I18177: signal is true;
	signal I18180: std_logic; attribute dont_touch of I18180: signal is true;
	signal I18191: std_logic; attribute dont_touch of I18191: signal is true;
	signal I18205: std_logic; attribute dont_touch of I18205: signal is true;
	signal I18214: std_logic; attribute dont_touch of I18214: signal is true;
	signal I18221: std_logic; attribute dont_touch of I18221: signal is true;
	signal I18224: std_logic; attribute dont_touch of I18224: signal is true;
	signal I18233: std_logic; attribute dont_touch of I18233: signal is true;
	signal I18238: std_logic; attribute dont_touch of I18238: signal is true;
	signal I18245: std_logic; attribute dont_touch of I18245: signal is true;
	signal I18248: std_logic; attribute dont_touch of I18248: signal is true;
	signal I18252: std_logic; attribute dont_touch of I18252: signal is true;
	signal I18259: std_logic; attribute dont_touch of I18259: signal is true;
	signal I18262: std_logic; attribute dont_touch of I18262: signal is true;
	signal I18265: std_logic; attribute dont_touch of I18265: signal is true;
	signal I18270: std_logic; attribute dont_touch of I18270: signal is true;
	signal I18276: std_logic; attribute dont_touch of I18276: signal is true;
	signal I18280: std_logic; attribute dont_touch of I18280: signal is true;
	signal I18285: std_logic; attribute dont_touch of I18285: signal is true;
	signal I18293: std_logic; attribute dont_touch of I18293: signal is true;
	signal I18297: std_logic; attribute dont_touch of I18297: signal is true;
	signal I18301: std_logic; attribute dont_touch of I18301: signal is true;
	signal I18304: std_logic; attribute dont_touch of I18304: signal is true;
	signal I18307: std_logic; attribute dont_touch of I18307: signal is true;
	signal I18310: std_logic; attribute dont_touch of I18310: signal is true;
	signal I18313: std_logic; attribute dont_touch of I18313: signal is true;
	signal I18320: std_logic; attribute dont_touch of I18320: signal is true;
	signal I18323: std_logic; attribute dont_touch of I18323: signal is true;
	signal I18333: std_logic; attribute dont_touch of I18333: signal is true;
	signal I18337: std_logic; attribute dont_touch of I18337: signal is true;
	signal I18341: std_logic; attribute dont_touch of I18341: signal is true;
	signal I18344: std_logic; attribute dont_touch of I18344: signal is true;
	signal I18350: std_logic; attribute dont_touch of I18350: signal is true;
	signal I18360: std_logic; attribute dont_touch of I18360: signal is true;
	signal I18364: std_logic; attribute dont_touch of I18364: signal is true;
	signal I18367: std_logic; attribute dont_touch of I18367: signal is true;
	signal I18370: std_logic; attribute dont_touch of I18370: signal is true;
	signal I18373: std_logic; attribute dont_touch of I18373: signal is true;
	signal I18376: std_logic; attribute dont_touch of I18376: signal is true;
	signal I18379: std_logic; attribute dont_touch of I18379: signal is true;
	signal I18382: std_logic; attribute dont_touch of I18382: signal is true;
	signal I18385: std_logic; attribute dont_touch of I18385: signal is true;
	signal I18398: std_logic; attribute dont_touch of I18398: signal is true;
	signal I18408: std_logic; attribute dont_touch of I18408: signal is true;
	signal I18411: std_logic; attribute dont_touch of I18411: signal is true;
	signal I18414: std_logic; attribute dont_touch of I18414: signal is true;
	signal I18417: std_logic; attribute dont_touch of I18417: signal is true;
	signal I18421: std_logic; attribute dont_touch of I18421: signal is true;
	signal I18434: std_logic; attribute dont_touch of I18434: signal is true;
	signal I18443: std_logic; attribute dont_touch of I18443: signal is true;
	signal I18446: std_logic; attribute dont_touch of I18446: signal is true;
	signal I18449: std_logic; attribute dont_touch of I18449: signal is true;
	signal I18452: std_logic; attribute dont_touch of I18452: signal is true;
	signal I18460: std_logic; attribute dont_touch of I18460: signal is true;
	signal I18469: std_logic; attribute dont_touch of I18469: signal is true;
	signal I18476: std_logic; attribute dont_touch of I18476: signal is true;
	signal I18479: std_logic; attribute dont_touch of I18479: signal is true;
	signal I18482: std_logic; attribute dont_touch of I18482: signal is true;
	signal I18485: std_logic; attribute dont_touch of I18485: signal is true;
	signal I18486: std_logic; attribute dont_touch of I18486: signal is true;
	signal I18487: std_logic; attribute dont_touch of I18487: signal is true;
	signal I18492: std_logic; attribute dont_touch of I18492: signal is true;
	signal I18495: std_logic; attribute dont_touch of I18495: signal is true;
	signal I18504: std_logic; attribute dont_touch of I18504: signal is true;
	signal I18509: std_logic; attribute dont_touch of I18509: signal is true;
	signal I18518: std_logic; attribute dont_touch of I18518: signal is true;
	signal I18523: std_logic; attribute dont_touch of I18523: signal is true;
	signal I18526: std_logic; attribute dont_touch of I18526: signal is true;
	signal I18529: std_logic; attribute dont_touch of I18529: signal is true;
	signal I18530: std_logic; attribute dont_touch of I18530: signal is true;
	signal I18531: std_logic; attribute dont_touch of I18531: signal is true;
	signal I18536: std_logic; attribute dont_touch of I18536: signal is true;
	signal I18537: std_logic; attribute dont_touch of I18537: signal is true;
	signal I18538: std_logic; attribute dont_touch of I18538: signal is true;
	signal I18543: std_logic; attribute dont_touch of I18543: signal is true;
	signal I18555: std_logic; attribute dont_touch of I18555: signal is true;
	signal I18560: std_logic; attribute dont_touch of I18560: signal is true;
	signal I18568: std_logic; attribute dont_touch of I18568: signal is true;
	signal I18571: std_logic; attribute dont_touch of I18571: signal is true;
	signal I18574: std_logic; attribute dont_touch of I18574: signal is true;
	signal I18579: std_logic; attribute dont_touch of I18579: signal is true;
	signal I18580: std_logic; attribute dont_touch of I18580: signal is true;
	signal I18581: std_logic; attribute dont_touch of I18581: signal is true;
	signal I18587: std_logic; attribute dont_touch of I18587: signal is true;
	signal I18588: std_logic; attribute dont_touch of I18588: signal is true;
	signal I18589: std_logic; attribute dont_touch of I18589: signal is true;
	signal I18600: std_logic; attribute dont_touch of I18600: signal is true;
	signal I18609: std_logic; attribute dont_touch of I18609: signal is true;
	signal I18614: std_logic; attribute dont_touch of I18614: signal is true;
	signal I18620: std_logic; attribute dont_touch of I18620: signal is true;
	signal I18625: std_logic; attribute dont_touch of I18625: signal is true;
	signal I18626: std_logic; attribute dont_touch of I18626: signal is true;
	signal I18627: std_logic; attribute dont_touch of I18627: signal is true;
	signal I18633: std_logic; attribute dont_touch of I18633: signal is true;
	signal I18634: std_logic; attribute dont_touch of I18634: signal is true;
	signal I18635: std_logic; attribute dont_touch of I18635: signal is true;
	signal I18647: std_logic; attribute dont_touch of I18647: signal is true;
	signal I18653: std_logic; attribute dont_touch of I18653: signal is true;
	signal I18662: std_logic; attribute dont_touch of I18662: signal is true;
	signal I18667: std_logic; attribute dont_touch of I18667: signal is true;
	signal I18671: std_logic; attribute dont_touch of I18671: signal is true;
	signal I18674: std_logic; attribute dont_touch of I18674: signal is true;
	signal I18680: std_logic; attribute dont_touch of I18680: signal is true;
	signal I18681: std_logic; attribute dont_touch of I18681: signal is true;
	signal I18682: std_logic; attribute dont_touch of I18682: signal is true;
	signal I18694: std_logic; attribute dont_touch of I18694: signal is true;
	signal I18700: std_logic; attribute dont_touch of I18700: signal is true;
	signal I18709: std_logic; attribute dont_touch of I18709: signal is true;
	signal I18713: std_logic; attribute dont_touch of I18713: signal is true;
	signal I18716: std_logic; attribute dont_touch of I18716: signal is true;
	signal I18728: std_logic; attribute dont_touch of I18728: signal is true;
	signal I18734: std_logic; attribute dont_touch of I18734: signal is true;
	signal I18740: std_logic; attribute dont_touch of I18740: signal is true;
	signal I18752: std_logic; attribute dont_touch of I18752: signal is true;
	signal I18758: std_logic; attribute dont_touch of I18758: signal is true;
	signal I18762: std_logic; attribute dont_touch of I18762: signal is true;
	signal I18765: std_logic; attribute dont_touch of I18765: signal is true;
	signal I18778: std_logic; attribute dont_touch of I18778: signal is true;
	signal I18782: std_logic; attribute dont_touch of I18782: signal is true;
	signal I18785: std_logic; attribute dont_touch of I18785: signal is true;
	signal I18788: std_logic; attribute dont_touch of I18788: signal is true;
	signal I18795: std_logic; attribute dont_touch of I18795: signal is true;
	signal I18803: std_logic; attribute dont_touch of I18803: signal is true;
	signal I18810: std_logic; attribute dont_touch of I18810: signal is true;
	signal I18813: std_logic; attribute dont_touch of I18813: signal is true;
	signal I18819: std_logic; attribute dont_touch of I18819: signal is true;
	signal I18822: std_logic; attribute dont_touch of I18822: signal is true;
	signal I18825: std_logic; attribute dont_touch of I18825: signal is true;
	signal I18829: std_logic; attribute dont_touch of I18829: signal is true;
	signal I18832: std_logic; attribute dont_touch of I18832: signal is true;
	signal I18835: std_logic; attribute dont_touch of I18835: signal is true;
	signal I18839: std_logic; attribute dont_touch of I18839: signal is true;
	signal I18842: std_logic; attribute dont_touch of I18842: signal is true;
	signal I18845: std_logic; attribute dont_touch of I18845: signal is true;
	signal I18849: std_logic; attribute dont_touch of I18849: signal is true;
	signal I18852: std_logic; attribute dont_touch of I18852: signal is true;
	signal I18855: std_logic; attribute dont_touch of I18855: signal is true;
	signal I18858: std_logic; attribute dont_touch of I18858: signal is true;
	signal I18861: std_logic; attribute dont_touch of I18861: signal is true;
	signal I18865: std_logic; attribute dont_touch of I18865: signal is true;
	signal I18868: std_logic; attribute dont_touch of I18868: signal is true;
	signal I18872: std_logic; attribute dont_touch of I18872: signal is true;
	signal I18875: std_logic; attribute dont_touch of I18875: signal is true;
	signal I18879: std_logic; attribute dont_touch of I18879: signal is true;
	signal I18882: std_logic; attribute dont_touch of I18882: signal is true;
	signal I18885: std_logic; attribute dont_touch of I18885: signal is true;
	signal I18888: std_logic; attribute dont_touch of I18888: signal is true;
	signal I18891: std_logic; attribute dont_touch of I18891: signal is true;
	signal I18894: std_logic; attribute dont_touch of I18894: signal is true;
	signal I18897: std_logic; attribute dont_touch of I18897: signal is true;
	signal I18900: std_logic; attribute dont_touch of I18900: signal is true;
	signal I18903: std_logic; attribute dont_touch of I18903: signal is true;
	signal I18906: std_logic; attribute dont_touch of I18906: signal is true;
	signal I18909: std_logic; attribute dont_touch of I18909: signal is true;
	signal I18912: std_logic; attribute dont_touch of I18912: signal is true;
	signal I19012: std_logic; attribute dont_touch of I19012: signal is true;
	signal I19235: std_logic; attribute dont_touch of I19235: signal is true;
	signal I19238: std_logic; attribute dont_touch of I19238: signal is true;
	signal I19345: std_logic; attribute dont_touch of I19345: signal is true;
	signal I19348: std_logic; attribute dont_touch of I19348: signal is true;
	signal I19384: std_logic; attribute dont_touch of I19384: signal is true;
	signal I19484: std_logic; attribute dont_touch of I19484: signal is true;
	signal I19487: std_logic; attribute dont_touch of I19487: signal is true;
	signal I19661: std_logic; attribute dont_touch of I19661: signal is true;
	signal I19671: std_logic; attribute dont_touch of I19671: signal is true;
	signal I19674: std_logic; attribute dont_touch of I19674: signal is true;
	signal I19704: std_logic; attribute dont_touch of I19704: signal is true;
	signal I19707: std_logic; attribute dont_touch of I19707: signal is true;
	signal I19719: std_logic; attribute dont_touch of I19719: signal is true;
	signal I19734: std_logic; attribute dont_touch of I19734: signal is true;
	signal I19756: std_logic; attribute dont_touch of I19756: signal is true;
	signal I19759: std_logic; attribute dont_touch of I19759: signal is true;
	signal I19762: std_logic; attribute dont_touch of I19762: signal is true;
	signal I19772: std_logic; attribute dont_touch of I19772: signal is true;
	signal I19775: std_logic; attribute dont_touch of I19775: signal is true;
	signal I19778: std_logic; attribute dont_touch of I19778: signal is true;
	signal I19786: std_logic; attribute dont_touch of I19786: signal is true;
	signal I19789: std_logic; attribute dont_touch of I19789: signal is true;
	signal I19796: std_logic; attribute dont_touch of I19796: signal is true;
	signal I19799: std_logic; attribute dont_touch of I19799: signal is true;
	signal I19802: std_logic; attribute dont_touch of I19802: signal is true;
	signal I19813: std_logic; attribute dont_touch of I19813: signal is true;
	signal I19818: std_logic; attribute dont_touch of I19818: signal is true;
	signal I19831: std_logic; attribute dont_touch of I19831: signal is true;
	signal I19837: std_logic; attribute dont_touch of I19837: signal is true;
	signal I19843: std_logic; attribute dont_touch of I19843: signal is true;
	signal I19851: std_logic; attribute dont_touch of I19851: signal is true;
	signal I19857: std_logic; attribute dont_touch of I19857: signal is true;
	signal I19863: std_logic; attribute dont_touch of I19863: signal is true;
	signal I19917: std_logic; attribute dont_touch of I19917: signal is true;
	signal I19927: std_logic; attribute dont_touch of I19927: signal is true;
	signal I20035: std_logic; attribute dont_touch of I20035: signal is true;
	signal I20116: std_logic; attribute dont_touch of I20116: signal is true;
	signal I20130: std_logic; attribute dont_touch of I20130: signal is true;
	signal I20165: std_logic; attribute dont_touch of I20165: signal is true;
	signal I20166: std_logic; attribute dont_touch of I20166: signal is true;
	signal I20167: std_logic; attribute dont_touch of I20167: signal is true;
	signal I20187: std_logic; attribute dont_touch of I20187: signal is true;
	signal I20188: std_logic; attribute dont_touch of I20188: signal is true;
	signal I20189: std_logic; attribute dont_touch of I20189: signal is true;
	signal I20203: std_logic; attribute dont_touch of I20203: signal is true;
	signal I20204: std_logic; attribute dont_touch of I20204: signal is true;
	signal I20205: std_logic; attribute dont_touch of I20205: signal is true;
	signal I20216: std_logic; attribute dont_touch of I20216: signal is true;
	signal I20221: std_logic; attribute dont_touch of I20221: signal is true;
	signal I20222: std_logic; attribute dont_touch of I20222: signal is true;
	signal I20223: std_logic; attribute dont_touch of I20223: signal is true;
	signal I20233: std_logic; attribute dont_touch of I20233: signal is true;
	signal I20318: std_logic; attribute dont_touch of I20318: signal is true;
	signal I20321: std_logic; attribute dont_touch of I20321: signal is true;
	signal I20355: std_logic; attribute dont_touch of I20355: signal is true;
	signal I20369: std_logic; attribute dont_touch of I20369: signal is true;
	signal I20385: std_logic; attribute dont_touch of I20385: signal is true;
	signal I20388: std_logic; attribute dont_touch of I20388: signal is true;
	signal I20399: std_logic; attribute dont_touch of I20399: signal is true;
	signal I20412: std_logic; attribute dont_touch of I20412: signal is true;
	signal I20433: std_logic; attribute dont_touch of I20433: signal is true;
	signal I20447: std_logic; attribute dont_touch of I20447: signal is true;
	signal I20460: std_logic; attribute dont_touch of I20460: signal is true;
	signal I20461: std_logic; attribute dont_touch of I20461: signal is true;
	signal I20462: std_logic; attribute dont_touch of I20462: signal is true;
	signal I20467: std_logic; attribute dont_touch of I20467: signal is true;
	signal I20468: std_logic; attribute dont_touch of I20468: signal is true;
	signal I20469: std_logic; attribute dont_touch of I20469: signal is true;
	signal I20486: std_logic; attribute dont_touch of I20486: signal is true;
	signal I20487: std_logic; attribute dont_touch of I20487: signal is true;
	signal I20488: std_logic; attribute dont_touch of I20488: signal is true;
	signal I20495: std_logic; attribute dont_touch of I20495: signal is true;
	signal I20499: std_logic; attribute dont_touch of I20499: signal is true;
	signal I20529: std_logic; attribute dont_touch of I20529: signal is true;
	signal I20542: std_logic; attribute dont_touch of I20542: signal is true;
	signal I20562: std_logic; attribute dont_touch of I20562: signal is true;
	signal I20569: std_logic; attribute dont_touch of I20569: signal is true;
	signal I20584: std_logic; attribute dont_touch of I20584: signal is true;
	signal I20609: std_logic; attribute dont_touch of I20609: signal is true;
	signal I20647: std_logic; attribute dont_touch of I20647: signal is true;
	signal I20650: std_logic; attribute dont_touch of I20650: signal is true;
	signal I20690: std_logic; attribute dont_touch of I20690: signal is true;
	signal I20744: std_logic; attribute dont_touch of I20744: signal is true;
	signal I20747: std_logic; attribute dont_touch of I20747: signal is true;
	signal I20750: std_logic; attribute dont_touch of I20750: signal is true;
	signal I20753: std_logic; attribute dont_touch of I20753: signal is true;
	signal I20781: std_logic; attribute dont_touch of I20781: signal is true;
	signal I20793: std_logic; attribute dont_touch of I20793: signal is true;
	signal I20816: std_logic; attribute dont_touch of I20816: signal is true;
	signal I20819: std_logic; attribute dont_touch of I20819: signal is true;
	signal I20830: std_logic; attribute dont_touch of I20830: signal is true;
	signal I20840: std_logic; attribute dont_touch of I20840: signal is true;
	signal I20846: std_logic; attribute dont_touch of I20846: signal is true;
	signal I20861: std_logic; attribute dont_touch of I20861: signal is true;
	signal I20864: std_logic; attribute dont_touch of I20864: signal is true;
	signal I20867: std_logic; attribute dont_touch of I20867: signal is true;
	signal I20870: std_logic; attribute dont_touch of I20870: signal is true;
	signal I20882: std_logic; attribute dont_touch of I20882: signal is true;
	signal I20891: std_logic; attribute dont_touch of I20891: signal is true;
	signal I20895: std_logic; attribute dont_touch of I20895: signal is true;
	signal I20910: std_logic; attribute dont_touch of I20910: signal is true;
	signal I20913: std_logic; attribute dont_touch of I20913: signal is true;
	signal I20929: std_logic; attribute dont_touch of I20929: signal is true;
	signal I20937: std_logic; attribute dont_touch of I20937: signal is true;
	signal I20951: std_logic; attribute dont_touch of I20951: signal is true;
	signal I20954: std_logic; attribute dont_touch of I20954: signal is true;
	signal I20957: std_logic; attribute dont_touch of I20957: signal is true;
	signal I20982: std_logic; attribute dont_touch of I20982: signal is true;
	signal I20985: std_logic; attribute dont_touch of I20985: signal is true;
	signal I20999: std_logic; attribute dont_touch of I20999: signal is true;
	signal I21002: std_logic; attribute dont_touch of I21002: signal is true;
	signal I21006: std_logic; attribute dont_touch of I21006: signal is true;
	signal I21013: std_logic; attribute dont_touch of I21013: signal is true;
	signal I21019: std_logic; attribute dont_touch of I21019: signal is true;
	signal I21029: std_logic; attribute dont_touch of I21029: signal is true;
	signal I21033: std_logic; attribute dont_touch of I21033: signal is true;
	signal I21036: std_logic; attribute dont_touch of I21036: signal is true;
	signal I21042: std_logic; attribute dont_touch of I21042: signal is true;
	signal I21047: std_logic; attribute dont_touch of I21047: signal is true;
	signal I21058: std_logic; attribute dont_touch of I21058: signal is true;
	signal I21067: std_logic; attribute dont_touch of I21067: signal is true;
	signal I21074: std_logic; attribute dont_touch of I21074: signal is true;
	signal I21100: std_logic; attribute dont_touch of I21100: signal is true;
	signal I21115: std_logic; attribute dont_touch of I21115: signal is true;
	signal I21162: std_logic; attribute dont_touch of I21162: signal is true;
	signal I21181: std_logic; attribute dont_touch of I21181: signal is true;
	signal I21189: std_logic; attribute dont_touch of I21189: signal is true;
	signal I21199: std_logic; attribute dont_touch of I21199: signal is true;
	signal I21210: std_logic; attribute dont_touch of I21210: signal is true;
	signal I21222: std_logic; attribute dont_touch of I21222: signal is true;
	signal I21226: std_logic; attribute dont_touch of I21226: signal is true;
	signal I21230: std_logic; attribute dont_touch of I21230: signal is true;
	signal I21234: std_logic; attribute dont_touch of I21234: signal is true;
	signal I21238: std_logic; attribute dont_touch of I21238: signal is true;
	signal I21242: std_logic; attribute dont_touch of I21242: signal is true;
	signal I21246: std_logic; attribute dont_touch of I21246: signal is true;
	signal I21250: std_logic; attribute dont_touch of I21250: signal is true;
	signal I21254: std_logic; attribute dont_touch of I21254: signal is true;
	signal I21258: std_logic; attribute dont_touch of I21258: signal is true;
	signal I21285: std_logic; attribute dont_touch of I21285: signal is true;
	signal I21288: std_logic; attribute dont_touch of I21288: signal is true;
	signal I21291: std_logic; attribute dont_touch of I21291: signal is true;
	signal I21294: std_logic; attribute dont_touch of I21294: signal is true;
	signal I21297: std_logic; attribute dont_touch of I21297: signal is true;
	signal I21300: std_logic; attribute dont_touch of I21300: signal is true;
	signal I21477: std_logic; attribute dont_touch of I21477: signal is true;
	signal I21480: std_logic; attribute dont_touch of I21480: signal is true;
	signal I21483: std_logic; attribute dont_touch of I21483: signal is true;
	signal I21486: std_logic; attribute dont_touch of I21486: signal is true;
	signal I21722: std_logic; attribute dont_touch of I21722: signal is true;
	signal I21734: std_logic; attribute dont_touch of I21734: signal is true;
	signal I21744: std_logic; attribute dont_touch of I21744: signal is true;
	signal I21757: std_logic; attribute dont_touch of I21757: signal is true;
	signal I21766: std_logic; attribute dont_touch of I21766: signal is true;
	signal I21769: std_logic; attribute dont_touch of I21769: signal is true;
	signal I21776: std_logic; attribute dont_touch of I21776: signal is true;
	signal I21784: std_logic; attribute dont_touch of I21784: signal is true;
	signal I21787: std_logic; attribute dont_touch of I21787: signal is true;
	signal I21792: std_logic; attribute dont_touch of I21792: signal is true;
	signal I21802: std_logic; attribute dont_touch of I21802: signal is true;
	signal I21810: std_logic; attribute dont_touch of I21810: signal is true;
	signal I21815: std_logic; attribute dont_touch of I21815: signal is true;
	signal I21831: std_logic; attribute dont_touch of I21831: signal is true;
	signal I21838: std_logic; attribute dont_touch of I21838: signal is true;
	signal I21849: std_logic; attribute dont_touch of I21849: signal is true;
	signal I21860: std_logic; attribute dont_touch of I21860: signal is true;
	signal I21911: std_logic; attribute dont_touch of I21911: signal is true;
	signal I21918: std_logic; attribute dont_touch of I21918: signal is true;
	signal I21922: std_logic; attribute dont_touch of I21922: signal is true;
	signal I21930: std_logic; attribute dont_touch of I21930: signal is true;
	signal I21934: std_logic; attribute dont_touch of I21934: signal is true;
	signal I21941: std_logic; attribute dont_touch of I21941: signal is true;
	signal I21959: std_logic; attribute dont_touch of I21959: signal is true;
	signal I21969: std_logic; attribute dont_touch of I21969: signal is true;
	signal I21976: std_logic; attribute dont_touch of I21976: signal is true;
	signal I21977: std_logic; attribute dont_touch of I21977: signal is true;
	signal I21978: std_logic; attribute dont_touch of I21978: signal is true;
	signal I21992: std_logic; attribute dont_touch of I21992: signal is true;
	signal I21993: std_logic; attribute dont_touch of I21993: signal is true;
	signal I21994: std_logic; attribute dont_touch of I21994: signal is true;
	signal I22000: std_logic; attribute dont_touch of I22000: signal is true;
	signal I22009: std_logic; attribute dont_touch of I22009: signal is true;
	signal I22024: std_logic; attribute dont_touch of I22024: signal is true;
	signal I22028: std_logic; attribute dont_touch of I22028: signal is true;
	signal I22031: std_logic; attribute dont_touch of I22031: signal is true;
	signal I22046: std_logic; attribute dont_touch of I22046: signal is true;
	signal I22096: std_logic; attribute dont_touch of I22096: signal is true;
	signal I22111: std_logic; attribute dont_touch of I22111: signal is true;
	signal I22114: std_logic; attribute dont_touch of I22114: signal is true;
	signal I22124: std_logic; attribute dont_touch of I22124: signal is true;
	signal I22128: std_logic; attribute dont_touch of I22128: signal is true;
	signal I22131: std_logic; attribute dont_touch of I22131: signal is true;
	signal I22143: std_logic; attribute dont_touch of I22143: signal is true;
	signal I22149: std_logic; attribute dont_touch of I22149: signal is true;
	signal I22153: std_logic; attribute dont_touch of I22153: signal is true;
	signal I22177: std_logic; attribute dont_touch of I22177: signal is true;
	signal I22180: std_logic; attribute dont_touch of I22180: signal is true;
	signal I22211: std_logic; attribute dont_touch of I22211: signal is true;
	signal I22240: std_logic; attribute dont_touch of I22240: signal is true;
	signal I22264: std_logic; attribute dont_touch of I22264: signal is true;
	signal I22267: std_logic; attribute dont_touch of I22267: signal is true;
	signal I22275: std_logic; attribute dont_touch of I22275: signal is true;
	signal I22280: std_logic; attribute dont_touch of I22280: signal is true;
	signal I22286: std_logic; attribute dont_touch of I22286: signal is true;
	signal I22289: std_logic; attribute dont_touch of I22289: signal is true;
	signal I22298: std_logic; attribute dont_touch of I22298: signal is true;
	signal I22302: std_logic; attribute dont_touch of I22302: signal is true;
	signal I22316: std_logic; attribute dont_touch of I22316: signal is true;
	signal I22327: std_logic; attribute dont_touch of I22327: signal is true;
	signal I22331: std_logic; attribute dont_touch of I22331: signal is true;
	signal I22343: std_logic; attribute dont_touch of I22343: signal is true;
	signal I22353: std_logic; attribute dont_touch of I22353: signal is true;
	signal I22366: std_logic; attribute dont_touch of I22366: signal is true;
	signal I22380: std_logic; attribute dont_touch of I22380: signal is true;
	signal I22400: std_logic; attribute dont_touch of I22400: signal is true;
	signal I22419: std_logic; attribute dont_touch of I22419: signal is true;
	signal I22422: std_logic; attribute dont_touch of I22422: signal is true;
	signal I22425: std_logic; attribute dont_touch of I22425: signal is true;
	signal I22444: std_logic; attribute dont_touch of I22444: signal is true;
	signal I22458: std_logic; attribute dont_touch of I22458: signal is true;
	signal I22461: std_logic; attribute dont_touch of I22461: signal is true;
	signal I22464: std_logic; attribute dont_touch of I22464: signal is true;
	signal I22467: std_logic; attribute dont_touch of I22467: signal is true;
	signal I22470: std_logic; attribute dont_touch of I22470: signal is true;
	signal I22485: std_logic; attribute dont_touch of I22485: signal is true;
	signal I22488: std_logic; attribute dont_touch of I22488: signal is true;
	signal I22499: std_logic; attribute dont_touch of I22499: signal is true;
	signal I22502: std_logic; attribute dont_touch of I22502: signal is true;
	signal I22512: std_logic; attribute dont_touch of I22512: signal is true;
	signal I22525: std_logic; attribute dont_touch of I22525: signal is true;
	signal I22539: std_logic; attribute dont_touch of I22539: signal is true;
	signal I22542: std_logic; attribute dont_touch of I22542: signal is true;
	signal I22547: std_logic; attribute dont_touch of I22547: signal is true;
	signal I22557: std_logic; attribute dont_touch of I22557: signal is true;
	signal I22561: std_logic; attribute dont_touch of I22561: signal is true;
	signal I22564: std_logic; attribute dont_touch of I22564: signal is true;
	signal I22571: std_logic; attribute dont_touch of I22571: signal is true;
	signal I22576: std_logic; attribute dont_touch of I22576: signal is true;
	signal I22580: std_logic; attribute dont_touch of I22580: signal is true;
	signal I22583: std_logic; attribute dont_touch of I22583: signal is true;
	signal I22589: std_logic; attribute dont_touch of I22589: signal is true;
	signal I22601: std_logic; attribute dont_touch of I22601: signal is true;
	signal I22604: std_logic; attribute dont_touch of I22604: signal is true;
	signal I22619: std_logic; attribute dont_touch of I22619: signal is true;
	signal I22622: std_logic; attribute dont_touch of I22622: signal is true;
	signal I22640: std_logic; attribute dont_touch of I22640: signal is true;
	signal I22665: std_logic; attribute dont_touch of I22665: signal is true;
	signal I22683: std_logic; attribute dont_touch of I22683: signal is true;
	signal I22684: std_logic; attribute dont_touch of I22684: signal is true;
	signal I22685: std_logic; attribute dont_touch of I22685: signal is true;
	signal I22692: std_logic; attribute dont_touch of I22692: signal is true;
	signal I22710: std_logic; attribute dont_touch of I22710: signal is true;
	signal I22711: std_logic; attribute dont_touch of I22711: signal is true;
	signal I22712: std_logic; attribute dont_touch of I22712: signal is true;
	signal I22717: std_logic; attribute dont_touch of I22717: signal is true;
	signal I22718: std_logic; attribute dont_touch of I22718: signal is true;
	signal I22719: std_logic; attribute dont_touch of I22719: signal is true;
	signal I22725: std_logic; attribute dont_touch of I22725: signal is true;
	signal I22729: std_logic; attribute dont_touch of I22729: signal is true;
	signal I22745: std_logic; attribute dont_touch of I22745: signal is true;
	signal I22748: std_logic; attribute dont_touch of I22748: signal is true;
	signal I22753: std_logic; attribute dont_touch of I22753: signal is true;
	signal I22754: std_logic; attribute dont_touch of I22754: signal is true;
	signal I22755: std_logic; attribute dont_touch of I22755: signal is true;
	signal I22760: std_logic; attribute dont_touch of I22760: signal is true;
	signal I22761: std_logic; attribute dont_touch of I22761: signal is true;
	signal I22762: std_logic; attribute dont_touch of I22762: signal is true;
	signal I22769: std_logic; attribute dont_touch of I22769: signal is true;
	signal I22785: std_logic; attribute dont_touch of I22785: signal is true;
	signal I22788: std_logic; attribute dont_touch of I22788: signal is true;
	signal I22792: std_logic; attribute dont_touch of I22792: signal is true;
	signal I22793: std_logic; attribute dont_touch of I22793: signal is true;
	signal I22794: std_logic; attribute dont_touch of I22794: signal is true;
	signal I22799: std_logic; attribute dont_touch of I22799: signal is true;
	signal I22800: std_logic; attribute dont_touch of I22800: signal is true;
	signal I22801: std_logic; attribute dont_touch of I22801: signal is true;
	signal I22816: std_logic; attribute dont_touch of I22816: signal is true;
	signal I22819: std_logic; attribute dont_touch of I22819: signal is true;
	signal I22822: std_logic; attribute dont_touch of I22822: signal is true;
	signal I22823: std_logic; attribute dont_touch of I22823: signal is true;
	signal I22824: std_logic; attribute dont_touch of I22824: signal is true;
	signal I22830: std_logic; attribute dont_touch of I22830: signal is true;
	signal I22844: std_logic; attribute dont_touch of I22844: signal is true;
	signal I22845: std_logic; attribute dont_touch of I22845: signal is true;
	signal I22846: std_logic; attribute dont_touch of I22846: signal is true;
	signal I22852: std_logic; attribute dont_touch of I22852: signal is true;
	signal I22864: std_logic; attribute dont_touch of I22864: signal is true;
	signal I22865: std_logic; attribute dont_touch of I22865: signal is true;
	signal I22866: std_logic; attribute dont_touch of I22866: signal is true;
	signal I22871: std_logic; attribute dont_touch of I22871: signal is true;
	signal I22872: std_logic; attribute dont_touch of I22872: signal is true;
	signal I22873: std_logic; attribute dont_touch of I22873: signal is true;
	signal I22880: std_logic; attribute dont_touch of I22880: signal is true;
	signal I22886: std_logic; attribute dont_touch of I22886: signal is true;
	signal I22889: std_logic; attribute dont_touch of I22889: signal is true;
	signal I22892: std_logic; attribute dont_touch of I22892: signal is true;
	signal I22893: std_logic; attribute dont_touch of I22893: signal is true;
	signal I22894: std_logic; attribute dont_touch of I22894: signal is true;
	signal I22899: std_logic; attribute dont_touch of I22899: signal is true;
	signal I22900: std_logic; attribute dont_touch of I22900: signal is true;
	signal I22901: std_logic; attribute dont_touch of I22901: signal is true;
	signal I22912: std_logic; attribute dont_touch of I22912: signal is true;
	signal I22918: std_logic; attribute dont_touch of I22918: signal is true;
	signal I22921: std_logic; attribute dont_touch of I22921: signal is true;
	signal I22922: std_logic; attribute dont_touch of I22922: signal is true;
	signal I22923: std_logic; attribute dont_touch of I22923: signal is true;
	signal I22929: std_logic; attribute dont_touch of I22929: signal is true;
	signal I22930: std_logic; attribute dont_touch of I22930: signal is true;
	signal I22931: std_logic; attribute dont_touch of I22931: signal is true;
	signal I22936: std_logic; attribute dont_touch of I22936: signal is true;
	signal I22937: std_logic; attribute dont_touch of I22937: signal is true;
	signal I22938: std_logic; attribute dont_touch of I22938: signal is true;
	signal I22944: std_logic; attribute dont_touch of I22944: signal is true;
	signal I22945: std_logic; attribute dont_touch of I22945: signal is true;
	signal I22946: std_logic; attribute dont_touch of I22946: signal is true;
	signal I22958: std_logic; attribute dont_touch of I22958: signal is true;
	signal I22965: std_logic; attribute dont_touch of I22965: signal is true;
	signal I22966: std_logic; attribute dont_touch of I22966: signal is true;
	signal I22967: std_logic; attribute dont_touch of I22967: signal is true;
	signal I22972: std_logic; attribute dont_touch of I22972: signal is true;
	signal I22973: std_logic; attribute dont_touch of I22973: signal is true;
	signal I22974: std_logic; attribute dont_touch of I22974: signal is true;
	signal I22989: std_logic; attribute dont_touch of I22989: signal is true;
	signal I23099: std_logic; attribute dont_touch of I23099: signal is true;
	signal I23118: std_logic; attribute dont_touch of I23118: signal is true;
	signal I23119: std_logic; attribute dont_touch of I23119: signal is true;
	signal I23120: std_logic; attribute dont_touch of I23120: signal is true;
	signal I23149: std_logic; attribute dont_touch of I23149: signal is true;
	signal I23162: std_logic; attribute dont_touch of I23162: signal is true;
	signal I23163: std_logic; attribute dont_touch of I23163: signal is true;
	signal I23300: std_logic; attribute dont_touch of I23300: signal is true;
	signal I23303: std_logic; attribute dont_touch of I23303: signal is true;
	signal I23306: std_logic; attribute dont_touch of I23306: signal is true;
	signal I23309: std_logic; attribute dont_touch of I23309: signal is true;
	signal I23312: std_logic; attribute dont_touch of I23312: signal is true;
	signal I23315: std_logic; attribute dont_touch of I23315: signal is true;
	signal I23318: std_logic; attribute dont_touch of I23318: signal is true;
	signal I23321: std_logic; attribute dont_touch of I23321: signal is true;
	signal I23324: std_logic; attribute dont_touch of I23324: signal is true;
	signal I23327: std_logic; attribute dont_touch of I23327: signal is true;
	signal I23330: std_logic; attribute dont_touch of I23330: signal is true;
	signal I23333: std_logic; attribute dont_touch of I23333: signal is true;
	signal I23336: std_logic; attribute dont_touch of I23336: signal is true;
	signal I23339: std_logic; attribute dont_touch of I23339: signal is true;
	signal I23342: std_logic; attribute dont_touch of I23342: signal is true;
	signal I23345: std_logic; attribute dont_touch of I23345: signal is true;
	signal I23348: std_logic; attribute dont_touch of I23348: signal is true;
	signal I23351: std_logic; attribute dont_touch of I23351: signal is true;
	signal I23354: std_logic; attribute dont_touch of I23354: signal is true;
	signal I23357: std_logic; attribute dont_touch of I23357: signal is true;
	signal I23360: std_logic; attribute dont_touch of I23360: signal is true;
	signal I23363: std_logic; attribute dont_touch of I23363: signal is true;
	signal I23366: std_logic; attribute dont_touch of I23366: signal is true;
	signal I23369: std_logic; attribute dont_touch of I23369: signal is true;
	signal I23372: std_logic; attribute dont_touch of I23372: signal is true;
	signal I23375: std_logic; attribute dont_touch of I23375: signal is true;
	signal I23378: std_logic; attribute dont_touch of I23378: signal is true;
	signal I23381: std_logic; attribute dont_touch of I23381: signal is true;
	signal I23384: std_logic; attribute dont_touch of I23384: signal is true;
	signal I23387: std_logic; attribute dont_touch of I23387: signal is true;
	signal I23390: std_logic; attribute dont_touch of I23390: signal is true;
	signal I23393: std_logic; attribute dont_touch of I23393: signal is true;
	signal I23396: std_logic; attribute dont_touch of I23396: signal is true;
	signal I23399: std_logic; attribute dont_touch of I23399: signal is true;
	signal I23585: std_logic; attribute dont_touch of I23585: signal is true;
	signal I23586: std_logic; attribute dont_touch of I23586: signal is true;
	signal I23587: std_logic; attribute dont_touch of I23587: signal is true;
	signal I23600: std_logic; attribute dont_touch of I23600: signal is true;
	signal I23601: std_logic; attribute dont_touch of I23601: signal is true;
	signal I23602: std_logic; attribute dont_touch of I23602: signal is true;
	signal I23671: std_logic; attribute dont_touch of I23671: signal is true;
	signal I23680: std_logic; attribute dont_touch of I23680: signal is true;
	signal I23684: std_logic; attribute dont_touch of I23684: signal is true;
	signal I23688: std_logic; attribute dont_touch of I23688: signal is true;
	signal I23694: std_logic; attribute dont_touch of I23694: signal is true;
	signal I23711: std_logic; attribute dont_touch of I23711: signal is true;
	signal I23755: std_logic; attribute dont_touch of I23755: signal is true;
	signal I23756: std_logic; attribute dont_touch of I23756: signal is true;
	signal I23917: std_logic; attribute dont_touch of I23917: signal is true;
	signal I23918: std_logic; attribute dont_touch of I23918: signal is true;
	signal I23919: std_logic; attribute dont_touch of I23919: signal is true;
	signal I23949: std_logic; attribute dont_touch of I23949: signal is true;
	signal I23950: std_logic; attribute dont_touch of I23950: signal is true;
	signal I23951: std_logic; attribute dont_touch of I23951: signal is true;
	signal I23961: std_logic; attribute dont_touch of I23961: signal is true;
	signal I23962: std_logic; attribute dont_touch of I23962: signal is true;
	signal I23963: std_logic; attribute dont_touch of I23963: signal is true;
	signal I23969: std_logic; attribute dont_touch of I23969: signal is true;
	signal I23970: std_logic; attribute dont_touch of I23970: signal is true;
	signal I23971: std_logic; attribute dont_touch of I23971: signal is true;
	signal I23978: std_logic; attribute dont_touch of I23978: signal is true;
	signal I23979: std_logic; attribute dont_touch of I23979: signal is true;
	signal I23980: std_logic; attribute dont_touch of I23980: signal is true;
	signal I23985: std_logic; attribute dont_touch of I23985: signal is true;
	signal I23986: std_logic; attribute dont_touch of I23986: signal is true;
	signal I23987: std_logic; attribute dont_touch of I23987: signal is true;
	signal I23998: std_logic; attribute dont_touch of I23998: signal is true;
	signal I24003: std_logic; attribute dont_touch of I24003: signal is true;
	signal I24008: std_logic; attribute dont_touch of I24008: signal is true;
	signal I24015: std_logic; attribute dont_touch of I24015: signal is true;
	signal I24018: std_logic; attribute dont_touch of I24018: signal is true;
	signal I24022: std_logic; attribute dont_touch of I24022: signal is true;
	signal I24027: std_logic; attribute dont_touch of I24027: signal is true;
	signal I24030: std_logic; attribute dont_touch of I24030: signal is true;
	signal I24033: std_logic; attribute dont_touch of I24033: signal is true;
	signal I24038: std_logic; attribute dont_touch of I24038: signal is true;
	signal I24041: std_logic; attribute dont_touch of I24041: signal is true;
	signal I24048: std_logic; attribute dont_touch of I24048: signal is true;
	signal I24051: std_logic; attribute dont_touch of I24051: signal is true;
	signal I24054: std_logic; attribute dont_touch of I24054: signal is true;
	signal I24060: std_logic; attribute dont_touch of I24060: signal is true;
	signal I24064: std_logic; attribute dont_touch of I24064: signal is true;
	signal I24067: std_logic; attribute dont_touch of I24067: signal is true;
	signal I24075: std_logic; attribute dont_touch of I24075: signal is true;
	signal I24078: std_logic; attribute dont_touch of I24078: signal is true;
	signal I24089: std_logic; attribute dont_touch of I24089: signal is true;
	signal I24117: std_logic; attribute dont_touch of I24117: signal is true;
	signal I24128: std_logic; attribute dont_touch of I24128: signal is true;
	signal I24191: std_logic; attribute dont_touch of I24191: signal is true;
	signal I24215: std_logic; attribute dont_touch of I24215: signal is true;
	signal I24228: std_logic; attribute dont_touch of I24228: signal is true;
	signal I24237: std_logic; attribute dont_touch of I24237: signal is true;
	signal I24278: std_logic; attribute dont_touch of I24278: signal is true;
	signal I24281: std_logic; attribute dont_touch of I24281: signal is true;
	signal I24331: std_logic; attribute dont_touch of I24331: signal is true;
	signal I24334: std_logic; attribute dont_touch of I24334: signal is true;
	signal I24363: std_logic; attribute dont_touch of I24363: signal is true;
	signal I24364: std_logic; attribute dont_touch of I24364: signal is true;
	signal I24365: std_logic; attribute dont_touch of I24365: signal is true;
	signal I24383: std_logic; attribute dont_touch of I24383: signal is true;
	signal I24384: std_logic; attribute dont_touch of I24384: signal is true;
	signal I24385: std_logic; attribute dont_touch of I24385: signal is true;
	signal I24393: std_logic; attribute dont_touch of I24393: signal is true;
	signal I24396: std_logic; attribute dont_touch of I24396: signal is true;
	signal I24400: std_logic; attribute dont_touch of I24400: signal is true;
	signal I24414: std_logic; attribute dont_touch of I24414: signal is true;
	signal I24415: std_logic; attribute dont_touch of I24415: signal is true;
	signal I24416: std_logic; attribute dont_touch of I24416: signal is true;
	signal I24434: std_logic; attribute dont_touch of I24434: signal is true;
	signal I24438: std_logic; attribute dont_touch of I24438: signal is true;
	signal I24439: std_logic; attribute dont_touch of I24439: signal is true;
	signal I24440: std_logic; attribute dont_touch of I24440: signal is true;
	signal I24445: std_logic; attribute dont_touch of I24445: signal is true;
	signal I24448: std_logic; attribute dont_touch of I24448: signal is true;
	signal I24455: std_logic; attribute dont_touch of I24455: signal is true;
	signal I24461: std_logic; attribute dont_touch of I24461: signal is true;
	signal I24462: std_logic; attribute dont_touch of I24462: signal is true;
	signal I24463: std_logic; attribute dont_touch of I24463: signal is true;
	signal I24474: std_logic; attribute dont_touch of I24474: signal is true;
	signal I24482: std_logic; attribute dont_touch of I24482: signal is true;
	signal I24497: std_logic; attribute dont_touch of I24497: signal is true;
	signal I24505: std_logic; attribute dont_touch of I24505: signal is true;
	signal I24508: std_logic; attribute dont_touch of I24508: signal is true;
	signal I24524: std_logic; attribute dont_touch of I24524: signal is true;
	signal I24527: std_logic; attribute dont_touch of I24527: signal is true;
	signal I24530: std_logic; attribute dont_touch of I24530: signal is true;
	signal I24546: std_logic; attribute dont_touch of I24546: signal is true;
	signal I24549: std_logic; attribute dont_touch of I24549: signal is true;
	signal I24552: std_logic; attribute dont_touch of I24552: signal is true;
	signal I24555: std_logic; attribute dont_touch of I24555: signal is true;
	signal I24558: std_logic; attribute dont_touch of I24558: signal is true;
	signal I24576: std_logic; attribute dont_touch of I24576: signal is true;
	signal I24579: std_logic; attribute dont_touch of I24579: signal is true;
	signal I24582: std_logic; attribute dont_touch of I24582: signal is true;
	signal I24585: std_logic; attribute dont_touch of I24585: signal is true;
	signal I24597: std_logic; attribute dont_touch of I24597: signal is true;
	signal I24600: std_logic; attribute dont_touch of I24600: signal is true;
	signal I24603: std_logic; attribute dont_touch of I24603: signal is true;
	signal I24616: std_logic; attribute dont_touch of I24616: signal is true;
	signal I24619: std_logic; attribute dont_touch of I24619: signal is true;
	signal I24625: std_logic; attribute dont_touch of I24625: signal is true;
	signal I24674: std_logic; attribute dont_touch of I24674: signal is true;
	signal I24675: std_logic; attribute dont_touch of I24675: signal is true;
	signal I24679: std_logic; attribute dont_touch of I24679: signal is true;
	signal I24680: std_logic; attribute dont_touch of I24680: signal is true;
	signal I24684: std_logic; attribute dont_touch of I24684: signal is true;
	signal I24685: std_logic; attribute dont_touch of I24685: signal is true;
	signal I24689: std_logic; attribute dont_touch of I24689: signal is true;
	signal I24690: std_logic; attribute dont_touch of I24690: signal is true;
	signal I24694: std_logic; attribute dont_touch of I24694: signal is true;
	signal I24695: std_logic; attribute dont_touch of I24695: signal is true;
	signal I24699: std_logic; attribute dont_touch of I24699: signal is true;
	signal I24700: std_logic; attribute dont_touch of I24700: signal is true;
	signal I24704: std_logic; attribute dont_touch of I24704: signal is true;
	signal I24705: std_logic; attribute dont_touch of I24705: signal is true;
	signal I24709: std_logic; attribute dont_touch of I24709: signal is true;
	signal I24710: std_logic; attribute dont_touch of I24710: signal is true;
	signal I24759: std_logic; attribute dont_touch of I24759: signal is true;
	signal I24781: std_logic; attribute dont_touch of I24781: signal is true;
	signal I24784: std_logic; attribute dont_touch of I24784: signal is true;
	signal I24787: std_logic; attribute dont_touch of I24787: signal is true;
	signal I24839: std_logic; attribute dont_touch of I24839: signal is true;
	signal I24920: std_logic; attribute dont_touch of I24920: signal is true;
	signal I25005: std_logic; attribute dont_touch of I25005: signal is true;
	signal I25028: std_logic; attribute dont_touch of I25028: signal is true;
	signal I25095: std_logic; attribute dont_touch of I25095: signal is true;
	signal I25105: std_logic; attribute dont_touch of I25105: signal is true;
	signal I25115: std_logic; attribute dont_touch of I25115: signal is true;
	signal I25146: std_logic; attribute dont_touch of I25146: signal is true;
	signal I25161: std_logic; attribute dont_touch of I25161: signal is true;
	signal I25190: std_logic; attribute dont_touch of I25190: signal is true;
	signal I25219: std_logic; attribute dont_touch of I25219: signal is true;
	signal I25220: std_logic; attribute dont_touch of I25220: signal is true;
	signal I25221: std_logic; attribute dont_touch of I25221: signal is true;
	signal I25242: std_logic; attribute dont_touch of I25242: signal is true;
	signal I25243: std_logic; attribute dont_touch of I25243: signal is true;
	signal I25244: std_logic; attribute dont_touch of I25244: signal is true;
	signal I25327: std_logic; attribute dont_touch of I25327: signal is true;
	signal I25351: std_logic; attribute dont_touch of I25351: signal is true;
	signal I25356: std_logic; attribute dont_touch of I25356: signal is true;
	signal I25359: std_logic; attribute dont_touch of I25359: signal is true;
	signal I25366: std_logic; attribute dont_touch of I25366: signal is true;
	signal I25369: std_logic; attribute dont_touch of I25369: signal is true;
	signal I25380: std_logic; attribute dont_touch of I25380: signal is true;
	signal I25391: std_logic; attribute dont_touch of I25391: signal is true;
	signal I25399: std_logic; attribute dont_touch of I25399: signal is true;
	signal I25511: std_logic; attribute dont_touch of I25511: signal is true;
	signal I25514: std_logic; attribute dont_touch of I25514: signal is true;
	signal I25530: std_logic; attribute dont_touch of I25530: signal is true;
	signal I25534: std_logic; attribute dont_touch of I25534: signal is true;
	signal I25541: std_logic; attribute dont_touch of I25541: signal is true;
	signal I25552: std_logic; attribute dont_touch of I25552: signal is true;
	signal I25555: std_logic; attribute dont_touch of I25555: signal is true;
	signal I25562: std_logic; attribute dont_touch of I25562: signal is true;
	signal I25567: std_logic; attribute dont_touch of I25567: signal is true;
	signal I25576: std_logic; attribute dont_touch of I25576: signal is true;
	signal I25579: std_logic; attribute dont_touch of I25579: signal is true;
	signal I25586: std_logic; attribute dont_touch of I25586: signal is true;
	signal I25591: std_logic; attribute dont_touch of I25591: signal is true;
	signal I25594: std_logic; attribute dont_touch of I25594: signal is true;
	signal I25598: std_logic; attribute dont_touch of I25598: signal is true;
	signal I25606: std_logic; attribute dont_touch of I25606: signal is true;
	signal I25612: std_logic; attribute dont_touch of I25612: signal is true;
	signal I25613: std_logic; attribute dont_touch of I25613: signal is true;
	signal I25677: std_logic; attribute dont_touch of I25677: signal is true;
	signal I25680: std_logic; attribute dont_touch of I25680: signal is true;
	signal I25683: std_logic; attribute dont_touch of I25683: signal is true;
	signal I25689: std_logic; attribute dont_touch of I25689: signal is true;
	signal I25692: std_logic; attribute dont_touch of I25692: signal is true;
	signal I25695: std_logic; attribute dont_touch of I25695: signal is true;
	signal I25736: std_logic; attribute dont_touch of I25736: signal is true;
	signal I25743: std_logic; attribute dont_touch of I25743: signal is true;
	signal I25750: std_logic; attribute dont_touch of I25750: signal is true;
	signal I25779: std_logic; attribute dont_touch of I25779: signal is true;
	signal I25786: std_logic; attribute dont_touch of I25786: signal is true;
	signal I25790: std_logic; attribute dont_touch of I25790: signal is true;
	signal I25845: std_logic; attribute dont_touch of I25845: signal is true;
	signal I25846: std_logic; attribute dont_touch of I25846: signal is true;
	signal I25847: std_logic; attribute dont_touch of I25847: signal is true;
	signal I25869: std_logic; attribute dont_touch of I25869: signal is true;
	signal I25882: std_logic; attribute dont_touch of I25882: signal is true;
	signal I25907: std_logic; attribute dont_touch of I25907: signal is true;
	signal I25908: std_logic; attribute dont_touch of I25908: signal is true;
	signal I25909: std_logic; attribute dont_touch of I25909: signal is true;
	signal I26004: std_logic; attribute dont_touch of I26004: signal is true;
	signal I26049: std_logic; attribute dont_touch of I26049: signal is true;
	signal I26050: std_logic; attribute dont_touch of I26050: signal is true;
	signal I26051: std_logic; attribute dont_touch of I26051: signal is true;
	signal I26070: std_logic; attribute dont_touch of I26070: signal is true;
	signal I26071: std_logic; attribute dont_touch of I26071: signal is true;
	signal I26072: std_logic; attribute dont_touch of I26072: signal is true;
	signal I26093: std_logic; attribute dont_touch of I26093: signal is true;
	signal I26094: std_logic; attribute dont_touch of I26094: signal is true;
	signal I26095: std_logic; attribute dont_touch of I26095: signal is true;
	signal I26100: std_logic; attribute dont_touch of I26100: signal is true;
	signal I26130: std_logic; attribute dont_touch of I26130: signal is true;
	signal I26195: std_logic; attribute dont_touch of I26195: signal is true;
	signal I26296: std_logic; attribute dont_touch of I26296: signal is true;
	signal I26309: std_logic; attribute dont_touch of I26309: signal is true;
	signal I26334: std_logic; attribute dont_touch of I26334: signal is true;
	signal I26337: std_logic; attribute dont_touch of I26337: signal is true;
	signal I26356: std_logic; attribute dont_touch of I26356: signal is true;
	signal I26366: std_logic; attribute dont_touch of I26366: signal is true;
	signal I26367: std_logic; attribute dont_touch of I26367: signal is true;
	signal I26368: std_logic; attribute dont_touch of I26368: signal is true;
	signal I26378: std_logic; attribute dont_touch of I26378: signal is true;
	signal I26381: std_logic; attribute dont_touch of I26381: signal is true;
	signal I26393: std_logic; attribute dont_touch of I26393: signal is true;
	signal I26394: std_logic; attribute dont_touch of I26394: signal is true;
	signal I26395: std_logic; attribute dont_touch of I26395: signal is true;
	signal I26406: std_logic; attribute dont_touch of I26406: signal is true;
	signal I26409: std_logic; attribute dont_touch of I26409: signal is true;
	signal I26417: std_logic; attribute dont_touch of I26417: signal is true;
	signal I26418: std_logic; attribute dont_touch of I26418: signal is true;
	signal I26419: std_logic; attribute dont_touch of I26419: signal is true;
	signal I26427: std_logic; attribute dont_touch of I26427: signal is true;
	signal I26430: std_logic; attribute dont_touch of I26430: signal is true;
	signal I26438: std_logic; attribute dont_touch of I26438: signal is true;
	signal I26439: std_logic; attribute dont_touch of I26439: signal is true;
	signal I26440: std_logic; attribute dont_touch of I26440: signal is true;
	signal I26448: std_logic; attribute dont_touch of I26448: signal is true;
	signal I26451: std_logic; attribute dont_touch of I26451: signal is true;
	signal I26459: std_logic; attribute dont_touch of I26459: signal is true;
	signal I26460: std_logic; attribute dont_touch of I26460: signal is true;
	signal I26461: std_logic; attribute dont_touch of I26461: signal is true;
	signal I26466: std_logic; attribute dont_touch of I26466: signal is true;
	signal I26479: std_logic; attribute dont_touch of I26479: signal is true;
	signal I26503: std_logic; attribute dont_touch of I26503: signal is true;
	signal I26508: std_logic; attribute dont_touch of I26508: signal is true;
	signal I26512: std_logic; attribute dont_touch of I26512: signal is true;
	signal I26516: std_logic; attribute dont_touch of I26516: signal is true;
	signal I26522: std_logic; attribute dont_touch of I26522: signal is true;
	signal I26523: std_logic; attribute dont_touch of I26523: signal is true;
	signal I26530: std_logic; attribute dont_touch of I26530: signal is true;
	signal I26531: std_logic; attribute dont_touch of I26531: signal is true;
	signal I26578: std_logic; attribute dont_touch of I26578: signal is true;
	signal I26581: std_logic; attribute dont_touch of I26581: signal is true;
	signal I26584: std_logic; attribute dont_touch of I26584: signal is true;
	signal I26638: std_logic; attribute dont_touch of I26638: signal is true;
	signal I26643: std_logic; attribute dont_touch of I26643: signal is true;
	signal I26644: std_logic; attribute dont_touch of I26644: signal is true;
	signal I26649: std_logic; attribute dont_touch of I26649: signal is true;
	signal I26654: std_logic; attribute dont_touch of I26654: signal is true;
	signal I26664: std_logic; attribute dont_touch of I26664: signal is true;
	signal I26667: std_logic; attribute dont_touch of I26667: signal is true;
	signal I26670: std_logic; attribute dont_touch of I26670: signal is true;
	signal I26676: std_logic; attribute dont_touch of I26676: signal is true;
	signal I26679: std_logic; attribute dont_touch of I26679: signal is true;
	signal I26682: std_logic; attribute dont_touch of I26682: signal is true;
	signal I26687: std_logic; attribute dont_touch of I26687: signal is true;
	signal I26693: std_logic; attribute dont_touch of I26693: signal is true;
	signal I26700: std_logic; attribute dont_touch of I26700: signal is true;
	signal I26705: std_logic; attribute dont_touch of I26705: signal is true;
	signal I26710: std_logic; attribute dont_touch of I26710: signal is true;
	signal I26741: std_logic; attribute dont_touch of I26741: signal is true;
	signal I26742: std_logic; attribute dont_touch of I26742: signal is true;
	signal I26785: std_logic; attribute dont_touch of I26785: signal is true;
	signal I26799: std_logic; attribute dont_touch of I26799: signal is true;
	signal I26880: std_logic; attribute dont_touch of I26880: signal is true;
	signal I26925: std_logic; attribute dont_touch of I26925: signal is true;
	signal I26929: std_logic; attribute dont_touch of I26929: signal is true;
	signal I26936: std_logic; attribute dont_touch of I26936: signal is true;
	signal I26948: std_logic; attribute dont_touch of I26948: signal is true;
	signal I26952: std_logic; attribute dont_touch of I26952: signal is true;
	signal I26960: std_logic; attribute dont_touch of I26960: signal is true;
	signal I26972: std_logic; attribute dont_touch of I26972: signal is true;
	signal I26989: std_logic; attribute dont_touch of I26989: signal is true;
	signal I27192: std_logic; attribute dont_touch of I27192: signal is true;
	signal I27232: std_logic; attribute dont_touch of I27232: signal is true;
	signal I27235: std_logic; attribute dont_touch of I27235: signal is true;
	signal I27238: std_logic; attribute dont_touch of I27238: signal is true;
	signal I27253: std_logic; attribute dont_touch of I27253: signal is true;
	signal I27271: std_logic; attribute dont_touch of I27271: signal is true;
	signal I27314: std_logic; attribute dont_touch of I27314: signal is true;
	signal I27349: std_logic; attribute dont_touch of I27349: signal is true;
	signal I27364: std_logic; attribute dont_touch of I27364: signal is true;
	signal I27368: std_logic; attribute dont_touch of I27368: signal is true;
	signal I27381: std_logic; attribute dont_touch of I27381: signal is true;
	signal I27385: std_logic; attribute dont_touch of I27385: signal is true;
	signal I27388: std_logic; attribute dont_touch of I27388: signal is true;
	signal I27391: std_logic; attribute dont_touch of I27391: signal is true;
	signal I27401: std_logic; attribute dont_touch of I27401: signal is true;
	signal I27409: std_logic; attribute dont_touch of I27409: signal is true;
	signal I27429: std_logic; attribute dont_touch of I27429: signal is true;
	signal I27449: std_logic; attribute dont_touch of I27449: signal is true;
	signal I27481: std_logic; attribute dont_touch of I27481: signal is true;
	signal I27492: std_logic; attribute dont_touch of I27492: signal is true;
	signal I27495: std_logic; attribute dont_touch of I27495: signal is true;
	signal I27503: std_logic; attribute dont_touch of I27503: signal is true;
	signal I27504: std_logic; attribute dont_touch of I27504: signal is true;
	signal I27508: std_logic; attribute dont_touch of I27508: signal is true;
	signal I27509: std_logic; attribute dont_touch of I27509: signal is true;
	signal I27513: std_logic; attribute dont_touch of I27513: signal is true;
	signal I27514: std_logic; attribute dont_touch of I27514: signal is true;
	signal I27518: std_logic; attribute dont_touch of I27518: signal is true;
	signal I27519: std_logic; attribute dont_touch of I27519: signal is true;
	signal I27523: std_logic; attribute dont_touch of I27523: signal is true;
	signal I27524: std_logic; attribute dont_touch of I27524: signal is true;
	signal I27528: std_logic; attribute dont_touch of I27528: signal is true;
	signal I27529: std_logic; attribute dont_touch of I27529: signal is true;
	signal I27533: std_logic; attribute dont_touch of I27533: signal is true;
	signal I27534: std_logic; attribute dont_touch of I27534: signal is true;
	signal I27538: std_logic; attribute dont_touch of I27538: signal is true;
	signal I27539: std_logic; attribute dont_touch of I27539: signal is true;
	signal I27543: std_logic; attribute dont_touch of I27543: signal is true;
	signal I27546: std_logic; attribute dont_touch of I27546: signal is true;
	signal I27549: std_logic; attribute dont_touch of I27549: signal is true;
	signal I27552: std_logic; attribute dont_touch of I27552: signal is true;
	signal I27555: std_logic; attribute dont_touch of I27555: signal is true;
	signal I27558: std_logic; attribute dont_touch of I27558: signal is true;
	signal I27561: std_logic; attribute dont_touch of I27561: signal is true;
	signal I27564: std_logic; attribute dont_touch of I27564: signal is true;
	signal I27567: std_logic; attribute dont_touch of I27567: signal is true;
	signal I27570: std_logic; attribute dont_touch of I27570: signal is true;
	signal I27573: std_logic; attribute dont_touch of I27573: signal is true;
	signal I27576: std_logic; attribute dont_touch of I27576: signal is true;
	signal I27579: std_logic; attribute dont_touch of I27579: signal is true;
	signal I27677: std_logic; attribute dont_touch of I27677: signal is true;
	signal I27713: std_logic; attribute dont_touch of I27713: signal is true;
	signal I27718: std_logic; attribute dont_touch of I27718: signal is true;
	signal I27730: std_logic; attribute dont_touch of I27730: signal is true;
	signal I27735: std_logic; attribute dont_touch of I27735: signal is true;
	signal I27738: std_logic; attribute dont_touch of I27738: signal is true;
	signal I27742: std_logic; attribute dont_touch of I27742: signal is true;
	signal I27749: std_logic; attribute dont_touch of I27749: signal is true;
	signal I27758: std_logic; attribute dont_touch of I27758: signal is true;
	signal I27777: std_logic; attribute dont_touch of I27777: signal is true;
	signal I27784: std_logic; attribute dont_touch of I27784: signal is true;
	signal I27927: std_logic; attribute dont_touch of I27927: signal is true;
	signal I27941: std_logic; attribute dont_touch of I27941: signal is true;
	signal I27954: std_logic; attribute dont_touch of I27954: signal is true;
	signal I27970: std_logic; attribute dont_touch of I27970: signal is true;
	signal I28002: std_logic; attribute dont_touch of I28002: signal is true;
	signal I28014: std_logic; attribute dont_touch of I28014: signal is true;
	signal I28062: std_logic; attribute dont_touch of I28062: signal is true;
	signal I28128: std_logic; attribute dont_touch of I28128: signal is true;
	signal I28147: std_logic; attribute dont_touch of I28147: signal is true;
	signal I28162: std_logic; attribute dont_touch of I28162: signal is true;
	signal I28174: std_logic; attribute dont_touch of I28174: signal is true;
	signal I28185: std_logic; attribute dont_touch of I28185: signal is true;
	signal I28199: std_logic; attribute dont_touch of I28199: signal is true;
	signal I28241: std_logic; attribute dont_touch of I28241: signal is true;
	signal I28301: std_logic; attribute dont_touch of I28301: signal is true;
	signal I28336: std_logic; attribute dont_touch of I28336: signal is true;
	signal I28349: std_logic; attribute dont_touch of I28349: signal is true;
	signal I28390: std_logic; attribute dont_touch of I28390: signal is true;
	signal I28419: std_logic; attribute dont_touch of I28419: signal is true;
	signal I28434: std_logic; attribute dont_touch of I28434: signal is true;
	signal I28458: std_logic; attribute dont_touch of I28458: signal is true;
	signal I28480: std_logic; attribute dont_touch of I28480: signal is true;
	signal I28540: std_logic; attribute dont_touch of I28540: signal is true;
	signal I28548: std_logic; attribute dont_touch of I28548: signal is true;
	signal I28566: std_logic; attribute dont_touch of I28566: signal is true;
	signal I28567: std_logic; attribute dont_touch of I28567: signal is true;
	signal I28572: std_logic; attribute dont_touch of I28572: signal is true;
	signal I28576: std_logic; attribute dont_touch of I28576: signal is true;
	signal I28579: std_logic; attribute dont_touch of I28579: signal is true;
	signal I28582: std_logic; attribute dont_touch of I28582: signal is true;
	signal I28585: std_logic; attribute dont_touch of I28585: signal is true;
	signal I28588: std_logic; attribute dont_touch of I28588: signal is true;
	signal I28591: std_logic; attribute dont_touch of I28591: signal is true;
	signal I28594: std_logic; attribute dont_touch of I28594: signal is true;
	signal I28597: std_logic; attribute dont_touch of I28597: signal is true;
	signal I28832: std_logic; attribute dont_touch of I28832: signal is true;
	signal I28838: std_logic; attribute dont_touch of I28838: signal is true;
	signal I28851: std_logic; attribute dont_touch of I28851: signal is true;
	signal I28866: std_logic; attribute dont_touch of I28866: signal is true;
	signal I28872: std_logic; attribute dont_touch of I28872: signal is true;
	signal I28883: std_logic; attribute dont_touch of I28883: signal is true;
	signal I28897: std_logic; attribute dont_touch of I28897: signal is true;
	signal I28908: std_logic; attribute dont_touch of I28908: signal is true;
	signal I28913: std_logic; attribute dont_touch of I28913: signal is true;
	signal I28925: std_logic; attribute dont_touch of I28925: signal is true;
	signal I29002: std_logic; attribute dont_touch of I29002: signal is true;
	signal I29013: std_logic; attribute dont_touch of I29013: signal is true;
	signal I29139: std_logic; attribute dont_touch of I29139: signal is true;
	signal I29149: std_logic; attribute dont_touch of I29149: signal is true;
	signal I29182: std_logic; attribute dont_touch of I29182: signal is true;
	signal I29185: std_logic; attribute dont_touch of I29185: signal is true;
	signal I29199: std_logic; attribute dont_touch of I29199: signal is true;
	signal I29204: std_logic; attribute dont_touch of I29204: signal is true;
	signal I29207: std_logic; attribute dont_touch of I29207: signal is true;
	signal I29211: std_logic; attribute dont_touch of I29211: signal is true;
	signal I29214: std_logic; attribute dont_touch of I29214: signal is true;
	signal I29218: std_logic; attribute dont_touch of I29218: signal is true;
	signal I29221: std_logic; attribute dont_touch of I29221: signal is true;
	signal I29225: std_logic; attribute dont_touch of I29225: signal is true;
	signal I29228: std_logic; attribute dont_touch of I29228: signal is true;
	signal I29233: std_logic; attribute dont_touch of I29233: signal is true;
	signal I29236: std_logic; attribute dont_touch of I29236: signal is true;
	signal I29239: std_logic; attribute dont_touch of I29239: signal is true;
	signal I29242: std_logic; attribute dont_touch of I29242: signal is true;
	signal I29245: std_logic; attribute dont_touch of I29245: signal is true;
	signal I29248: std_logic; attribute dont_touch of I29248: signal is true;
	signal I29253: std_logic; attribute dont_touch of I29253: signal is true;
	signal I29254: std_logic; attribute dont_touch of I29254: signal is true;
	signal I29255: std_logic; attribute dont_touch of I29255: signal is true;
	signal I29261: std_logic; attribute dont_touch of I29261: signal is true;
	signal I29262: std_logic; attribute dont_touch of I29262: signal is true;
	signal I29263: std_logic; attribute dont_touch of I29263: signal is true;
	signal I29269: std_logic; attribute dont_touch of I29269: signal is true;
	signal I29270: std_logic; attribute dont_touch of I29270: signal is true;
	signal I29271: std_logic; attribute dont_touch of I29271: signal is true;
	signal I29277: std_logic; attribute dont_touch of I29277: signal is true;
	signal I29278: std_logic; attribute dont_touch of I29278: signal is true;
	signal I29279: std_logic; attribute dont_touch of I29279: signal is true;
	signal I29284: std_logic; attribute dont_touch of I29284: signal is true;
	signal I29285: std_logic; attribute dont_touch of I29285: signal is true;
	signal I29286: std_logic; attribute dont_touch of I29286: signal is true;
	signal I29295: std_logic; attribute dont_touch of I29295: signal is true;
	signal I29296: std_logic; attribute dont_touch of I29296: signal is true;
	signal I29297: std_logic; attribute dont_touch of I29297: signal is true;
	signal I29302: std_logic; attribute dont_touch of I29302: signal is true;
	signal I29303: std_logic; attribute dont_touch of I29303: signal is true;
	signal I29304: std_logic; attribute dont_touch of I29304: signal is true;
	signal I29313: std_logic; attribute dont_touch of I29313: signal is true;
	signal I29314: std_logic; attribute dont_touch of I29314: signal is true;
	signal I29315: std_logic; attribute dont_touch of I29315: signal is true;
	signal I29337: std_logic; attribute dont_touch of I29337: signal is true;
	signal I29351: std_logic; attribute dont_touch of I29351: signal is true;
	signal I29352: std_logic; attribute dont_touch of I29352: signal is true;
	signal I29363: std_logic; attribute dont_touch of I29363: signal is true;
	signal I29368: std_logic; attribute dont_touch of I29368: signal is true;
	signal I29371: std_logic; attribute dont_touch of I29371: signal is true;
	signal I29438: std_logic; attribute dont_touch of I29438: signal is true;
	signal I29441: std_logic; attribute dont_touch of I29441: signal is true;
	signal I29444: std_logic; attribute dont_touch of I29444: signal is true;
	signal I29447: std_logic; attribute dont_touch of I29447: signal is true;
	signal I29571: std_logic; attribute dont_touch of I29571: signal is true;
	signal I29579: std_logic; attribute dont_touch of I29579: signal is true;
	signal I29582: std_logic; attribute dont_touch of I29582: signal is true;
	signal I29585: std_logic; attribute dont_touch of I29585: signal is true;
	signal I29717: std_logic; attribute dont_touch of I29717: signal is true;
	signal I29720: std_logic; attribute dont_touch of I29720: signal is true;
	signal I29891: std_logic; attribute dont_touch of I29891: signal is true;
	signal I29894: std_logic; attribute dont_touch of I29894: signal is true;
	signal I29909: std_logic; attribute dont_touch of I29909: signal is true;
	signal I29913: std_logic; attribute dont_touch of I29913: signal is true;
	signal I29936: std_logic; attribute dont_touch of I29936: signal is true;
	signal I29939: std_logic; attribute dont_touch of I29939: signal is true;
	signal I29961: std_logic; attribute dont_touch of I29961: signal is true;
	signal I29965: std_logic; attribute dont_touch of I29965: signal is true;
	signal I29969: std_logic; attribute dont_touch of I29969: signal is true;
	signal I29973: std_logic; attribute dont_touch of I29973: signal is true;
	signal I29977: std_logic; attribute dont_touch of I29977: signal is true;
	signal I29981: std_logic; attribute dont_touch of I29981: signal is true;
	signal I29985: std_logic; attribute dont_touch of I29985: signal is true;
	signal I29986: std_logic; attribute dont_touch of I29986: signal is true;
	signal I30054: std_logic; attribute dont_touch of I30054: signal is true;
	signal I30055: std_logic; attribute dont_touch of I30055: signal is true;
	signal I30123: std_logic; attribute dont_touch of I30123: signal is true;
	signal I30124: std_logic; attribute dont_touch of I30124: signal is true;
	signal I30192: std_logic; attribute dont_touch of I30192: signal is true;
	signal I30193: std_logic; attribute dont_touch of I30193: signal is true;
	signal I30261: std_logic; attribute dont_touch of I30261: signal is true;
	signal I30262: std_logic; attribute dont_touch of I30262: signal is true;
	signal I30330: std_logic; attribute dont_touch of I30330: signal is true;
	signal I30331: std_logic; attribute dont_touch of I30331: signal is true;
	signal I30399: std_logic; attribute dont_touch of I30399: signal is true;
	signal I30400: std_logic; attribute dont_touch of I30400: signal is true;
	signal I30468: std_logic; attribute dont_touch of I30468: signal is true;
	signal I30469: std_logic; attribute dont_touch of I30469: signal is true;
	signal I30537: std_logic; attribute dont_touch of I30537: signal is true;
	signal I30641: std_logic; attribute dont_touch of I30641: signal is true;
	signal I30644: std_logic; attribute dont_touch of I30644: signal is true;
	signal I30686: std_logic; attribute dont_touch of I30686: signal is true;
	signal I30717: std_logic; attribute dont_touch of I30717: signal is true;
	signal I30718: std_logic; attribute dont_touch of I30718: signal is true;
	signal I30727: std_logic; attribute dont_touch of I30727: signal is true;
	signal I30728: std_logic; attribute dont_touch of I30728: signal is true;
	signal I30734: std_logic; attribute dont_touch of I30734: signal is true;
	signal I30735: std_logic; attribute dont_touch of I30735: signal is true;
	signal I30740: std_logic; attribute dont_touch of I30740: signal is true;
	signal I30741: std_logic; attribute dont_touch of I30741: signal is true;
	signal I30745: std_logic; attribute dont_touch of I30745: signal is true;
	signal I30746: std_logic; attribute dont_touch of I30746: signal is true;
	signal I30750: std_logic; attribute dont_touch of I30750: signal is true;
	signal I30751: std_logic; attribute dont_touch of I30751: signal is true;
	signal I30755: std_logic; attribute dont_touch of I30755: signal is true;
	signal I30756: std_logic; attribute dont_touch of I30756: signal is true;
	signal I30760: std_logic; attribute dont_touch of I30760: signal is true;
	signal I30761: std_logic; attribute dont_touch of I30761: signal is true;
	signal I30766: std_logic; attribute dont_touch of I30766: signal is true;
	signal I30861: std_logic; attribute dont_touch of I30861: signal is true;
	signal I30901: std_logic; attribute dont_touch of I30901: signal is true;
	signal I30904: std_logic; attribute dont_touch of I30904: signal is true;
	signal I30959: std_logic; attribute dont_touch of I30959: signal is true;
	signal I30962: std_logic; attribute dont_touch of I30962: signal is true;
	signal I30971: std_logic; attribute dont_touch of I30971: signal is true;
	signal I30980: std_logic; attribute dont_touch of I30980: signal is true;
	signal I30983: std_logic; attribute dont_touch of I30983: signal is true;
	signal I30986: std_logic; attribute dont_touch of I30986: signal is true;
	signal I30989: std_logic; attribute dont_touch of I30989: signal is true;
	signal I30992: std_logic; attribute dont_touch of I30992: signal is true;
	signal I30995: std_logic; attribute dont_touch of I30995: signal is true;
	signal I30998: std_logic; attribute dont_touch of I30998: signal is true;
	signal I31001: std_logic; attribute dont_touch of I31001: signal is true;
	signal I31002: std_logic; attribute dont_touch of I31002: signal is true;
	signal I31006: std_logic; attribute dont_touch of I31006: signal is true;
	signal I31007: std_logic; attribute dont_touch of I31007: signal is true;
	signal I31011: std_logic; attribute dont_touch of I31011: signal is true;
	signal I31012: std_logic; attribute dont_touch of I31012: signal is true;
	signal I31016: std_logic; attribute dont_touch of I31016: signal is true;
	signal I31017: std_logic; attribute dont_touch of I31017: signal is true;
	signal I31021: std_logic; attribute dont_touch of I31021: signal is true;
	signal I31022: std_logic; attribute dont_touch of I31022: signal is true;
	signal I31026: std_logic; attribute dont_touch of I31026: signal is true;
	signal I31027: std_logic; attribute dont_touch of I31027: signal is true;
	signal I31031: std_logic; attribute dont_touch of I31031: signal is true;
	signal I31032: std_logic; attribute dont_touch of I31032: signal is true;
	signal I31036: std_logic; attribute dont_touch of I31036: signal is true;
	signal I31037: std_logic; attribute dont_touch of I31037: signal is true;
	signal I31041: std_logic; attribute dont_touch of I31041: signal is true;
	signal I31042: std_logic; attribute dont_touch of I31042: signal is true;
	signal I31046: std_logic; attribute dont_touch of I31046: signal is true;
	signal I31047: std_logic; attribute dont_touch of I31047: signal is true;
	signal I31051: std_logic; attribute dont_touch of I31051: signal is true;
	signal I31052: std_logic; attribute dont_touch of I31052: signal is true;
	signal I31056: std_logic; attribute dont_touch of I31056: signal is true;
	signal I31057: std_logic; attribute dont_touch of I31057: signal is true;
	signal I31061: std_logic; attribute dont_touch of I31061: signal is true;
	signal I31062: std_logic; attribute dont_touch of I31062: signal is true;
	signal I31066: std_logic; attribute dont_touch of I31066: signal is true;
	signal I31067: std_logic; attribute dont_touch of I31067: signal is true;
	signal I31071: std_logic; attribute dont_touch of I31071: signal is true;
	signal I31072: std_logic; attribute dont_touch of I31072: signal is true;
	signal I31076: std_logic; attribute dont_touch of I31076: signal is true;
	signal I31077: std_logic; attribute dont_touch of I31077: signal is true;
	signal I31081: std_logic; attribute dont_touch of I31081: signal is true;
	signal I31082: std_logic; attribute dont_touch of I31082: signal is true;
	signal I31086: std_logic; attribute dont_touch of I31086: signal is true;
	signal I31087: std_logic; attribute dont_touch of I31087: signal is true;
	signal I31091: std_logic; attribute dont_touch of I31091: signal is true;
	signal I31092: std_logic; attribute dont_touch of I31092: signal is true;
	signal I31096: std_logic; attribute dont_touch of I31096: signal is true;
	signal I31097: std_logic; attribute dont_touch of I31097: signal is true;
	signal I31101: std_logic; attribute dont_touch of I31101: signal is true;
	signal I31102: std_logic; attribute dont_touch of I31102: signal is true;
	signal I31106: std_logic; attribute dont_touch of I31106: signal is true;
	signal I31107: std_logic; attribute dont_touch of I31107: signal is true;
	signal I31111: std_logic; attribute dont_touch of I31111: signal is true;
	signal I31112: std_logic; attribute dont_touch of I31112: signal is true;
	signal I31116: std_logic; attribute dont_touch of I31116: signal is true;
	signal I31117: std_logic; attribute dont_touch of I31117: signal is true;
	signal I31121: std_logic; attribute dont_touch of I31121: signal is true;
	signal I31122: std_logic; attribute dont_touch of I31122: signal is true;
	signal I31126: std_logic; attribute dont_touch of I31126: signal is true;
	signal I31127: std_logic; attribute dont_touch of I31127: signal is true;
	signal I31131: std_logic; attribute dont_touch of I31131: signal is true;
	signal I31132: std_logic; attribute dont_touch of I31132: signal is true;
	signal I31136: std_logic; attribute dont_touch of I31136: signal is true;
	signal I31137: std_logic; attribute dont_touch of I31137: signal is true;
	signal I31141: std_logic; attribute dont_touch of I31141: signal is true;
	signal I31142: std_logic; attribute dont_touch of I31142: signal is true;
	signal I31146: std_logic; attribute dont_touch of I31146: signal is true;
	signal I31147: std_logic; attribute dont_touch of I31147: signal is true;
	signal I31151: std_logic; attribute dont_touch of I31151: signal is true;
	signal I31152: std_logic; attribute dont_touch of I31152: signal is true;
	signal I31156: std_logic; attribute dont_touch of I31156: signal is true;
	signal I31157: std_logic; attribute dont_touch of I31157: signal is true;
	signal I31161: std_logic; attribute dont_touch of I31161: signal is true;
	signal I31162: std_logic; attribute dont_touch of I31162: signal is true;
	signal I31166: std_logic; attribute dont_touch of I31166: signal is true;
	signal I31167: std_logic; attribute dont_touch of I31167: signal is true;
	signal I31171: std_logic; attribute dont_touch of I31171: signal is true;
	signal I31172: std_logic; attribute dont_touch of I31172: signal is true;
	signal I31176: std_logic; attribute dont_touch of I31176: signal is true;
	signal I31177: std_logic; attribute dont_touch of I31177: signal is true;
	signal I31181: std_logic; attribute dont_touch of I31181: signal is true;
	signal I31182: std_logic; attribute dont_touch of I31182: signal is true;
	signal I31186: std_logic; attribute dont_touch of I31186: signal is true;
	signal I31187: std_logic; attribute dont_touch of I31187: signal is true;
	signal I31191: std_logic; attribute dont_touch of I31191: signal is true;
	signal I31192: std_logic; attribute dont_touch of I31192: signal is true;
	signal I31196: std_logic; attribute dont_touch of I31196: signal is true;
	signal I31197: std_logic; attribute dont_touch of I31197: signal is true;
	signal I31201: std_logic; attribute dont_touch of I31201: signal is true;
	signal I31202: std_logic; attribute dont_touch of I31202: signal is true;
	signal I31206: std_logic; attribute dont_touch of I31206: signal is true;
	signal I31207: std_logic; attribute dont_touch of I31207: signal is true;
	signal I31211: std_logic; attribute dont_touch of I31211: signal is true;
	signal I31212: std_logic; attribute dont_touch of I31212: signal is true;
	signal I31216: std_logic; attribute dont_touch of I31216: signal is true;
	signal I31217: std_logic; attribute dont_touch of I31217: signal is true;
	signal I31221: std_logic; attribute dont_touch of I31221: signal is true;
	signal I31222: std_logic; attribute dont_touch of I31222: signal is true;
	signal I31226: std_logic; attribute dont_touch of I31226: signal is true;
	signal I31227: std_logic; attribute dont_touch of I31227: signal is true;
	signal I31231: std_logic; attribute dont_touch of I31231: signal is true;
	signal I31232: std_logic; attribute dont_touch of I31232: signal is true;
	signal I31236: std_logic; attribute dont_touch of I31236: signal is true;
	signal I31237: std_logic; attribute dont_touch of I31237: signal is true;
	signal I31241: std_logic; attribute dont_touch of I31241: signal is true;
	signal I31242: std_logic; attribute dont_touch of I31242: signal is true;
	signal I31246: std_logic; attribute dont_touch of I31246: signal is true;
	signal I31247: std_logic; attribute dont_touch of I31247: signal is true;
	signal I31251: std_logic; attribute dont_touch of I31251: signal is true;
	signal I31252: std_logic; attribute dont_touch of I31252: signal is true;
	signal I31256: std_logic; attribute dont_touch of I31256: signal is true;
	signal I31257: std_logic; attribute dont_touch of I31257: signal is true;
	signal I31261: std_logic; attribute dont_touch of I31261: signal is true;
	signal I31262: std_logic; attribute dont_touch of I31262: signal is true;
	signal I31266: std_logic; attribute dont_touch of I31266: signal is true;
	signal I31267: std_logic; attribute dont_touch of I31267: signal is true;
	signal I31271: std_logic; attribute dont_touch of I31271: signal is true;
	signal I31272: std_logic; attribute dont_touch of I31272: signal is true;
	signal I31276: std_logic; attribute dont_touch of I31276: signal is true;
	signal I31277: std_logic; attribute dont_touch of I31277: signal is true;
	signal I31281: std_logic; attribute dont_touch of I31281: signal is true;
	signal I31282: std_logic; attribute dont_touch of I31282: signal is true;
	signal I31286: std_logic; attribute dont_touch of I31286: signal is true;
	signal I31287: std_logic; attribute dont_touch of I31287: signal is true;
	signal I31291: std_logic; attribute dont_touch of I31291: signal is true;
	signal I31292: std_logic; attribute dont_touch of I31292: signal is true;
	signal I31296: std_logic; attribute dont_touch of I31296: signal is true;
	signal I31297: std_logic; attribute dont_touch of I31297: signal is true;
	signal I31301: std_logic; attribute dont_touch of I31301: signal is true;
	signal I31302: std_logic; attribute dont_touch of I31302: signal is true;
	signal I31306: std_logic; attribute dont_touch of I31306: signal is true;
	signal I31307: std_logic; attribute dont_touch of I31307: signal is true;
	signal I31311: std_logic; attribute dont_touch of I31311: signal is true;
	signal I31312: std_logic; attribute dont_touch of I31312: signal is true;
	signal I31316: std_logic; attribute dont_touch of I31316: signal is true;
	signal I31317: std_logic; attribute dont_touch of I31317: signal is true;
	signal I31321: std_logic; attribute dont_touch of I31321: signal is true;
	signal I31322: std_logic; attribute dont_touch of I31322: signal is true;
	signal I31326: std_logic; attribute dont_touch of I31326: signal is true;
	signal I31327: std_logic; attribute dont_touch of I31327: signal is true;
	signal I31331: std_logic; attribute dont_touch of I31331: signal is true;
	signal I31332: std_logic; attribute dont_touch of I31332: signal is true;
	signal I31336: std_logic; attribute dont_touch of I31336: signal is true;
	signal I31337: std_logic; attribute dont_touch of I31337: signal is true;
	signal I31341: std_logic; attribute dont_touch of I31341: signal is true;
	signal I31342: std_logic; attribute dont_touch of I31342: signal is true;
	signal I31346: std_logic; attribute dont_touch of I31346: signal is true;
	signal I31347: std_logic; attribute dont_touch of I31347: signal is true;
	signal I31351: std_logic; attribute dont_touch of I31351: signal is true;
	signal I31352: std_logic; attribute dont_touch of I31352: signal is true;
	signal I31356: std_logic; attribute dont_touch of I31356: signal is true;
	signal I31357: std_logic; attribute dont_touch of I31357: signal is true;
	signal I31361: std_logic; attribute dont_touch of I31361: signal is true;
	signal I31459: std_logic; attribute dont_touch of I31459: signal is true;
	signal I31463: std_logic; attribute dont_touch of I31463: signal is true;
	signal I31466: std_logic; attribute dont_touch of I31466: signal is true;
	signal I31469: std_logic; attribute dont_touch of I31469: signal is true;
	signal I31474: std_logic; attribute dont_touch of I31474: signal is true;
	signal I31477: std_logic; attribute dont_touch of I31477: signal is true;
	signal I31482: std_logic; attribute dont_touch of I31482: signal is true;
	signal I31486: std_logic; attribute dont_touch of I31486: signal is true;
	signal I31491: std_logic; attribute dont_touch of I31491: signal is true;
	signal I31494: std_logic; attribute dont_touch of I31494: signal is true;
	signal I31497: std_logic; attribute dont_touch of I31497: signal is true;
	signal I31500: std_logic; attribute dont_touch of I31500: signal is true;
	signal I31504: std_logic; attribute dont_touch of I31504: signal is true;
	signal I31515: std_logic; attribute dont_touch of I31515: signal is true;
	signal I31523: std_logic; attribute dont_touch of I31523: signal is true;
	signal I31528: std_logic; attribute dont_touch of I31528: signal is true;
	signal I31535: std_logic; attribute dont_touch of I31535: signal is true;
	signal I31539: std_logic; attribute dont_touch of I31539: signal is true;
	signal I31545: std_logic; attribute dont_touch of I31545: signal is true;
	signal I31550: std_logic; attribute dont_touch of I31550: signal is true;
	signal I31555: std_logic; attribute dont_touch of I31555: signal is true;
	signal I31561: std_logic; attribute dont_touch of I31561: signal is true;
	signal I31564: std_logic; attribute dont_touch of I31564: signal is true;
	signal I31569: std_logic; attribute dont_touch of I31569: signal is true;
	signal I31581: std_logic; attribute dont_touch of I31581: signal is true;
	signal I31586: std_logic; attribute dont_touch of I31586: signal is true;
	signal I31593: std_logic; attribute dont_touch of I31593: signal is true;
	signal I31597: std_logic; attribute dont_touch of I31597: signal is true;
	signal I31600: std_logic; attribute dont_touch of I31600: signal is true;
	signal I31604: std_logic; attribute dont_touch of I31604: signal is true;
	signal I31607: std_logic; attribute dont_touch of I31607: signal is true;
	signal I31610: std_logic; attribute dont_touch of I31610: signal is true;
	signal I31616: std_logic; attribute dont_touch of I31616: signal is true;
	signal I31619: std_logic; attribute dont_touch of I31619: signal is true;
	signal I31622: std_logic; attribute dont_touch of I31622: signal is true;
	signal I31625: std_logic; attribute dont_touch of I31625: signal is true;
	signal I31642: std_logic; attribute dont_touch of I31642: signal is true;
	signal I31650: std_logic; attribute dont_touch of I31650: signal is true;
	signal I31659: std_logic; attribute dont_touch of I31659: signal is true;
	signal I31672: std_logic; attribute dont_touch of I31672: signal is true;
	signal I31686: std_logic; attribute dont_touch of I31686: signal is true;
	signal I31694: std_logic; attribute dont_touch of I31694: signal is true;
	signal I31701: std_logic; attribute dont_touch of I31701: signal is true;
	signal I31724: std_logic; attribute dont_touch of I31724: signal is true;
	signal I31727: std_logic; attribute dont_touch of I31727: signal is true;
	signal I31748: std_logic; attribute dont_touch of I31748: signal is true;
	signal I31751: std_logic; attribute dont_touch of I31751: signal is true;
	signal I31770: std_logic; attribute dont_touch of I31770: signal is true;
	signal I31776: std_logic; attribute dont_touch of I31776: signal is true;
	signal I31779: std_logic; attribute dont_touch of I31779: signal is true;
	signal I31782: std_logic; attribute dont_touch of I31782: signal is true;
	signal I31786: std_logic; attribute dont_touch of I31786: signal is true;
	signal I31791: std_logic; attribute dont_touch of I31791: signal is true;
	signal I31796: std_logic; attribute dont_touch of I31796: signal is true;
	signal I31800: std_logic; attribute dont_touch of I31800: signal is true;
	signal I31803: std_logic; attribute dont_touch of I31803: signal is true;
	signal I31807: std_logic; attribute dont_touch of I31807: signal is true;
	signal I31810: std_logic; attribute dont_touch of I31810: signal is true;
	signal I31814: std_logic; attribute dont_touch of I31814: signal is true;
	signal I31817: std_logic; attribute dont_touch of I31817: signal is true;
	signal I31820: std_logic; attribute dont_touch of I31820: signal is true;
	signal I31823: std_logic; attribute dont_touch of I31823: signal is true;
	signal I31829: std_logic; attribute dont_touch of I31829: signal is true;
	signal I31838: std_logic; attribute dont_touch of I31838: signal is true;
	signal I31839: std_logic; attribute dont_touch of I31839: signal is true;
	signal I31843: std_logic; attribute dont_touch of I31843: signal is true;
	signal I31844: std_logic; attribute dont_touch of I31844: signal is true;
	signal I31848: std_logic; attribute dont_touch of I31848: signal is true;
	signal I31849: std_logic; attribute dont_touch of I31849: signal is true;
	signal I31853: std_logic; attribute dont_touch of I31853: signal is true;
	signal I31854: std_logic; attribute dont_touch of I31854: signal is true;
	signal I31858: std_logic; attribute dont_touch of I31858: signal is true;
	signal I31859: std_logic; attribute dont_touch of I31859: signal is true;
	signal I31863: std_logic; attribute dont_touch of I31863: signal is true;
	signal I31864: std_logic; attribute dont_touch of I31864: signal is true;
	signal I31868: std_logic; attribute dont_touch of I31868: signal is true;
	signal I31869: std_logic; attribute dont_touch of I31869: signal is true;
	signal I31873: std_logic; attribute dont_touch of I31873: signal is true;
	signal I31874: std_logic; attribute dont_touch of I31874: signal is true;
	signal I31878: std_logic; attribute dont_touch of I31878: signal is true;
	signal I31972: std_logic; attribute dont_touch of I31972: signal is true;
	signal I31973: std_logic; attribute dont_touch of I31973: signal is true;
	signal I31974: std_logic; attribute dont_touch of I31974: signal is true;
	signal I31983: std_logic; attribute dont_touch of I31983: signal is true;
	signal I31984: std_logic; attribute dont_touch of I31984: signal is true;
	signal I31985: std_logic; attribute dont_touch of I31985: signal is true;
	signal I32051: std_logic; attribute dont_touch of I32051: signal is true;
	signal I32056: std_logic; attribute dont_touch of I32056: signal is true;
	signal I32059: std_logic; attribute dont_touch of I32059: signal is true;
	signal I32062: std_logic; attribute dont_touch of I32062: signal is true;
	signal I32067: std_logic; attribute dont_touch of I32067: signal is true;
	signal I32071: std_logic; attribute dont_touch of I32071: signal is true;
	signal I32074: std_logic; attribute dont_touch of I32074: signal is true;
	signal I32079: std_logic; attribute dont_touch of I32079: signal is true;
	signal I32089: std_logic; attribute dont_touch of I32089: signal is true;
	signal I32093: std_logic; attribute dont_touch of I32093: signal is true;
	signal I32096: std_logic; attribute dont_touch of I32096: signal is true;
	signal I32103: std_logic; attribute dont_touch of I32103: signal is true;
	signal I32106: std_logic; attribute dont_touch of I32106: signal is true;
	signal I32109: std_logic; attribute dont_touch of I32109: signal is true;
	signal I32116: std_logic; attribute dont_touch of I32116: signal is true;
	signal I32119: std_logic; attribute dont_touch of I32119: signal is true;
	signal I32150: std_logic; attribute dont_touch of I32150: signal is true;
	signal I32158: std_logic; attribute dont_touch of I32158: signal is true;
	signal I32161: std_logic; attribute dont_touch of I32161: signal is true;
	signal I32170: std_logic; attribute dont_touch of I32170: signal is true;
	signal I32173: std_logic; attribute dont_touch of I32173: signal is true;
	signal I32185: std_logic; attribute dont_touch of I32185: signal is true;
	signal I32186: std_logic; attribute dont_touch of I32186: signal is true;
	signal I32187: std_logic; attribute dont_touch of I32187: signal is true;
	signal I32192: std_logic; attribute dont_touch of I32192: signal is true;
	signal I32195: std_logic; attribute dont_touch of I32195: signal is true;
	signal I32202: std_logic; attribute dont_touch of I32202: signal is true;
	signal I32203: std_logic; attribute dont_touch of I32203: signal is true;
	signal I32204: std_logic; attribute dont_touch of I32204: signal is true;
	signal I32222: std_logic; attribute dont_touch of I32222: signal is true;
	signal I32225: std_logic; attribute dont_touch of I32225: signal is true;
	signal I32228: std_logic; attribute dont_touch of I32228: signal is true;
	signal I32231: std_logic; attribute dont_touch of I32231: signal is true;
	signal I32234: std_logic; attribute dont_touch of I32234: signal is true;
	signal I32237: std_logic; attribute dont_touch of I32237: signal is true;
	signal I32240: std_logic; attribute dont_touch of I32240: signal is true;
	signal I32243: std_logic; attribute dont_touch of I32243: signal is true;
	signal I32274: std_logic; attribute dont_touch of I32274: signal is true;
	signal I32284: std_logic; attribute dont_touch of I32284: signal is true;
	signal I32297: std_logic; attribute dont_touch of I32297: signal is true;
	signal I32305: std_logic; attribute dont_touch of I32305: signal is true;
	signal I32309: std_logic; attribute dont_touch of I32309: signal is true;
	signal I32352: std_logic; attribute dont_touch of I32352: signal is true;
	signal I32364: std_logic; attribute dont_touch of I32364: signal is true;
	signal I32388: std_logic; attribute dont_touch of I32388: signal is true;
	signal I32391: std_logic; attribute dont_touch of I32391: signal is true;
	signal I32431: std_logic; attribute dont_touch of I32431: signal is true;
	signal I32432: std_logic; attribute dont_touch of I32432: signal is true;
	signal I32433: std_logic; attribute dont_touch of I32433: signal is true;
	signal I32439: std_logic; attribute dont_touch of I32439: signal is true;
	signal I32440: std_logic; attribute dont_touch of I32440: signal is true;
	signal I32441: std_logic; attribute dont_touch of I32441: signal is true;
	signal I32446: std_logic; attribute dont_touch of I32446: signal is true;
	signal I32449: std_logic; attribute dont_touch of I32449: signal is true;
	signal I32452: std_logic; attribute dont_touch of I32452: signal is true;
	signal I32455: std_logic; attribute dont_touch of I32455: signal is true;
	signal I32458: std_logic; attribute dont_touch of I32458: signal is true;
	signal I32461: std_logic; attribute dont_touch of I32461: signal is true;
	signal I32464: std_logic; attribute dont_touch of I32464: signal is true;
	signal I32467: std_logic; attribute dont_touch of I32467: signal is true;
	signal I32470: std_logic; attribute dont_touch of I32470: signal is true;
	signal I32473: std_logic; attribute dont_touch of I32473: signal is true;
	signal I32476: std_logic; attribute dont_touch of I32476: signal is true;
	signal I32479: std_logic; attribute dont_touch of I32479: signal is true;
	signal I32482: std_logic; attribute dont_touch of I32482: signal is true;
	signal I32516: std_logic; attribute dont_touch of I32516: signal is true;
	signal I32517: std_logic; attribute dont_touch of I32517: signal is true;
	signal I32518: std_logic; attribute dont_touch of I32518: signal is true;
	signal I32525: std_logic; attribute dont_touch of I32525: signal is true;
	signal I32535: std_logic; attribute dont_touch of I32535: signal is true;
	signal I32547: std_logic; attribute dont_touch of I32547: signal is true;
	signal I32550: std_logic; attribute dont_touch of I32550: signal is true;
	signal I32591: std_logic; attribute dont_touch of I32591: signal is true;
	signal I32594: std_logic; attribute dont_touch of I32594: signal is true;
	signal I32601: std_logic; attribute dont_touch of I32601: signal is true;
	signal I32607: std_logic; attribute dont_touch of I32607: signal is true;
	signal I32613: std_logic; attribute dont_touch of I32613: signal is true;
	signal I32617: std_logic; attribute dont_touch of I32617: signal is true;
	signal I32621: std_logic; attribute dont_touch of I32621: signal is true;
	signal I32639: std_logic; attribute dont_touch of I32639: signal is true;
	signal I32645: std_logic; attribute dont_touch of I32645: signal is true;
	signal I32648: std_logic; attribute dont_touch of I32648: signal is true;
	signal I32651: std_logic; attribute dont_touch of I32651: signal is true;
	signal I32654: std_logic; attribute dont_touch of I32654: signal is true;
	signal I32659: std_logic; attribute dont_touch of I32659: signal is true;
	signal I32665: std_logic; attribute dont_touch of I32665: signal is true;
	signal I32671: std_logic; attribute dont_touch of I32671: signal is true;
	signal I32675: std_logic; attribute dont_touch of I32675: signal is true;
	signal I32678: std_logic; attribute dont_touch of I32678: signal is true;
	signal I32681: std_logic; attribute dont_touch of I32681: signal is true;
	signal I32684: std_logic; attribute dont_touch of I32684: signal is true;
	signal I32687: std_logic; attribute dont_touch of I32687: signal is true;
	signal I32690: std_logic; attribute dont_touch of I32690: signal is true;
	signal I32693: std_logic; attribute dont_touch of I32693: signal is true;
	signal I32696: std_logic; attribute dont_touch of I32696: signal is true;
	signal I32699: std_logic; attribute dont_touch of I32699: signal is true;
	signal I32752: std_logic; attribute dont_touch of I32752: signal is true;
	signal I32756: std_logic; attribute dont_touch of I32756: signal is true;
	signal I32757: std_logic; attribute dont_touch of I32757: signal is true;
	signal I32758: std_logic; attribute dont_touch of I32758: signal is true;
	signal I32763: std_logic; attribute dont_touch of I32763: signal is true;
	signal I32766: std_logic; attribute dont_touch of I32766: signal is true;
	signal I32770: std_logic; attribute dont_touch of I32770: signal is true;
	signal I32775: std_logic; attribute dont_touch of I32775: signal is true;
	signal I32782: std_logic; attribute dont_touch of I32782: signal is true;
	signal I32788: std_logic; attribute dont_touch of I32788: signal is true;
	signal I32791: std_logic; attribute dont_touch of I32791: signal is true;
	signal I32794: std_logic; attribute dont_touch of I32794: signal is true;
	signal I32797: std_logic; attribute dont_touch of I32797: signal is true;
	signal I32800: std_logic; attribute dont_touch of I32800: signal is true;
	signal I32803: std_logic; attribute dont_touch of I32803: signal is true;
	signal I32806: std_logic; attribute dont_touch of I32806: signal is true;
	signal I32809: std_logic; attribute dont_touch of I32809: signal is true;
	signal I32812: std_logic; attribute dont_touch of I32812: signal is true;
	signal I32815: std_logic; attribute dont_touch of I32815: signal is true;
	signal I32820: std_logic; attribute dont_touch of I32820: signal is true;
	signal I32824: std_logic; attribute dont_touch of I32824: signal is true;
	signal I32827: std_logic; attribute dont_touch of I32827: signal is true;
	signal I32834: std_logic; attribute dont_touch of I32834: signal is true;
	signal I32837: std_logic; attribute dont_touch of I32837: signal is true;
	signal I32840: std_logic; attribute dont_touch of I32840: signal is true;
	signal I32843: std_logic; attribute dont_touch of I32843: signal is true;
	signal I32846: std_logic; attribute dont_touch of I32846: signal is true;
	signal I32855: std_logic; attribute dont_touch of I32855: signal is true;
	signal I32868: std_logic; attribute dont_touch of I32868: signal is true;
	signal I32871: std_logic; attribute dont_touch of I32871: signal is true;
	signal I32874: std_logic; attribute dont_touch of I32874: signal is true;
	signal I32878: std_logic; attribute dont_touch of I32878: signal is true;
	signal I32881: std_logic; attribute dont_touch of I32881: signal is true;
	signal I32884: std_logic; attribute dont_touch of I32884: signal is true;
	signal I32904: std_logic; attribute dont_touch of I32904: signal is true;
	signal I32909: std_logic; attribute dont_touch of I32909: signal is true;
	signal I32921: std_logic; attribute dont_touch of I32921: signal is true;
	signal I32929: std_logic; attribute dont_touch of I32929: signal is true;
	signal I32935: std_logic; attribute dont_touch of I32935: signal is true;
	signal I32938: std_logic; attribute dont_touch of I32938: signal is true;
	signal I32947: std_logic; attribute dont_touch of I32947: signal is true;
	signal I32950: std_logic; attribute dont_touch of I32950: signal is true;
	signal I32953: std_logic; attribute dont_touch of I32953: signal is true;
	signal I32956: std_logic; attribute dont_touch of I32956: signal is true;
	signal I32960: std_logic; attribute dont_touch of I32960: signal is true;
	signal I32963: std_logic; attribute dont_touch of I32963: signal is true;
	signal I32967: std_logic; attribute dont_touch of I32967: signal is true;
	signal I32970: std_logic; attribute dont_touch of I32970: signal is true;
	signal I32973: std_logic; attribute dont_touch of I32973: signal is true;
	signal I32976: std_logic; attribute dont_touch of I32976: signal is true;
	signal I32982: std_logic; attribute dont_touch of I32982: signal is true;
	signal I32985: std_logic; attribute dont_touch of I32985: signal is true;
	signal I32988: std_logic; attribute dont_touch of I32988: signal is true;
	signal I32991: std_logic; attribute dont_touch of I32991: signal is true;
	signal I32994: std_logic; attribute dont_touch of I32994: signal is true;
	signal I32997: std_logic; attribute dont_touch of I32997: signal is true;
	signal I33020: std_logic; attribute dont_touch of I33020: signal is true;
	signal I33024: std_logic; attribute dont_touch of I33024: signal is true;
	signal I33027: std_logic; attribute dont_touch of I33027: signal is true;
	signal I33030: std_logic; attribute dont_touch of I33030: signal is true;
	signal I33034: std_logic; attribute dont_touch of I33034: signal is true;
	signal I33037: std_logic; attribute dont_touch of I33037: signal is true;
	signal I33041: std_logic; attribute dont_touch of I33041: signal is true;
	signal I33044: std_logic; attribute dont_touch of I33044: signal is true;
	signal I33047: std_logic; attribute dont_touch of I33047: signal is true;
	signal I33050: std_logic; attribute dont_touch of I33050: signal is true;
	signal I33053: std_logic; attribute dont_touch of I33053: signal is true;
	signal I33056: std_logic; attribute dont_touch of I33056: signal is true;
	signal I33064: std_logic; attribute dont_touch of I33064: signal is true;
	signal I33067: std_logic; attribute dont_touch of I33067: signal is true;
	signal I33070: std_logic; attribute dont_touch of I33070: signal is true;
	signal I33075: std_logic; attribute dont_touch of I33075: signal is true;
	signal I33079: std_logic; attribute dont_touch of I33079: signal is true;
	signal I33103: std_logic; attribute dont_touch of I33103: signal is true;
	signal I33106: std_logic; attribute dont_touch of I33106: signal is true;
	signal I33109: std_logic; attribute dont_touch of I33109: signal is true;
	signal I33119: std_logic; attribute dont_touch of I33119: signal is true;
	signal I33131: std_logic; attribute dont_touch of I33131: signal is true;
	signal I33134: std_logic; attribute dont_touch of I33134: signal is true;
	signal I33137: std_logic; attribute dont_touch of I33137: signal is true;
	signal I33140: std_logic; attribute dont_touch of I33140: signal is true;
	signal I33143: std_logic; attribute dont_touch of I33143: signal is true;
	signal I33146: std_logic; attribute dont_touch of I33146: signal is true;
	signal I33149: std_logic; attribute dont_touch of I33149: signal is true;
	signal I33152: std_logic; attribute dont_touch of I33152: signal is true;
	signal I33155: std_logic; attribute dont_touch of I33155: signal is true;
	signal I33158: std_logic; attribute dont_touch of I33158: signal is true;
	signal I33161: std_logic; attribute dont_touch of I33161: signal is true;
	signal I33164: std_logic; attribute dont_touch of I33164: signal is true;
	signal I33167: std_logic; attribute dont_touch of I33167: signal is true;
	signal I33170: std_logic; attribute dont_touch of I33170: signal is true;
	signal I33173: std_logic; attribute dont_touch of I33173: signal is true;
	signal I33176: std_logic; attribute dont_touch of I33176: signal is true;
	signal I33179: std_logic; attribute dont_touch of I33179: signal is true;
	signal I33182: std_logic; attribute dont_touch of I33182: signal is true;
	signal I33189: std_logic; attribute dont_touch of I33189: signal is true;
	signal I33197: std_logic; attribute dont_touch of I33197: signal is true;
	signal I33210: std_logic; attribute dont_touch of I33210: signal is true;
	signal I33214: std_logic; attribute dont_touch of I33214: signal is true;
	signal I33218: std_logic; attribute dont_touch of I33218: signal is true;
	signal I33232: std_logic; attribute dont_touch of I33232: signal is true;
	signal I33235: std_logic; attribute dont_touch of I33235: signal is true;
	signal I33246: std_logic; attribute dont_touch of I33246: signal is true;
	signal I33249: std_logic; attribute dont_touch of I33249: signal is true;
	signal I33252: std_logic; attribute dont_touch of I33252: signal is true;
	signal I33255: std_logic; attribute dont_touch of I33255: signal is true;
	signal I33258: std_logic; attribute dont_touch of I33258: signal is true;
	signal I33261: std_logic; attribute dont_touch of I33261: signal is true;
	signal I33264: std_logic; attribute dont_touch of I33264: signal is true;
	signal I33267: std_logic; attribute dont_touch of I33267: signal is true;
	signal I33270: std_logic; attribute dont_touch of I33270: signal is true;
	signal I33273: std_logic; attribute dont_touch of I33273: signal is true;
	signal I33276: std_logic; attribute dont_touch of I33276: signal is true;
	signal I33279: std_logic; attribute dont_touch of I33279: signal is true;
	signal I33282: std_logic; attribute dont_touch of I33282: signal is true;
	signal I33285: std_logic; attribute dont_touch of I33285: signal is true;
	signal I33288: std_logic; attribute dont_touch of I33288: signal is true;
	signal I33291: std_logic; attribute dont_touch of I33291: signal is true;
	signal I33297: std_logic; attribute dont_touch of I33297: signal is true;
	signal I33300: std_logic; attribute dont_touch of I33300: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			G1<=G26958;
			G6<=G34589;
			G7<=G34590;
			G8<=G34591;
			G9<=G34592;
			G12<=G30326;
			G16<=G34593;
			G19<=G34594;
			G22<=G29209;
			G25<=G15048;
			G28<=G34595;
			G31<=G34596;
			G34<=G34877;
			G37<=G34613;
			G43<=G34789;
			G45<=G34990;
			G46<=G34991;
			G47<=G34992;
			G48<=G34993;
			G49<=G34994;
			G50<=G34995;
			G51<=G34996;
			G52<=G34997;
			G55<=G35002;
			G58<=G30328;
			G59<=G29277;
			G63<=G34847;
			G65<=G34785;
			G66<=G24334;
			G70<=G18093;
			G71<=G34786;
			G74<=G26893;
			G79<=G26896;
			G85<=G34717;
			G86<=G25699;
			G93<=G34878;
			G94<=G34614;
			G101<=G34787;
			G102<=G33962;
			G106<=G26889;
			G110<=G34848;
			G111<=G34718;
			G112<=G34879;
			G117<=G30390;
			G121<=G30389;
			G128<=G28093;
			G136<=G34598;
			G142<=G34250;
			G146<=G30333;
			G150<=G32976;
			G153<=G33534;
			G157<=G33960;
			G160<=G34249;
			G164<=G31864;
			G168<=G25600;
			G174<=G25601;
			G182<=G25602;
			G191<=G194;
			G194<=G25592;
			G199<=G34721;
			G203<=G25599;
			G209<=G25593;
			G215<=G25591;
			G218<=G215;
			G222<=G33537;
			G225<=G26901;
			G232<=G26903;
			G239<=G26905;
			G246<=G26907;
			G255<=G26902;
			G262<=G26904;
			G269<=G26906;
			G278<=G25594;
			G283<=G28043;
			G287<=G31865;
			G291<=G32977;
			G294<=G33535;
			G298<=G33961;
			G301<=G33536;
			G305<=G26880;
			G311<=G26881;
			G316<=G26883;
			G319<=G26882;
			G324<=G26887;
			G329<=G26885;
			G333<=G26884;
			G336<=G26886;
			G341<=G26888;
			G344<=G26890;
			G347<=G344;
			G351<=G26891;
			G355<=G26892;
			G358<=G365;
			G365<=G25595;
			G370<=G25597;
			G376<=G25596;
			G385<=G25598;
			G391<=G26911;
			G392<=G24200;
			G401<=G24203;
			G405<=G24201;
			G411<=G29222;
			G417<=G24209;
			G424<=G24202;
			G429<=G24204;
			G433<=G24205;
			G437<=G24206;
			G441<=G24207;
			G446<=G26908;
			G452<=G25604;
			G457<=G25603;
			G460<=G25605;
			G464<=G25607;
			G468<=G25606;
			G471<=G25608;
			G475<=G24208;
			G479<=G24210;
			G482<=G28044;
			G490<=G29223;
			G496<=G33963;
			G499<=G25609;
			G504<=G25610;
			G513<=G25611;
			G518<=G25612;
			G528<=G26894;
			G534<=G34723;
			G538<=G34719;
			G542<=G24211;
			G546<=G34722;
			G550<=G34720;
			G554<=G34911;
			G559<=G640;
			G562<=G25613;
			G568<=G26895;
			G572<=G28045;
			G577<=G30334;
			G582<=G31866;
			G586<=G29224;
			G590<=G32978;
			G595<=G33538;
			G599<=G33964;
			G604<=G34251;
			G608<=G34438;
			G613<=G34599;
			G617<=G34724;
			G622<=G34790;
			G626<=G34849;
			G632<=G34880;
			G637<=G24212;
			G640<=G637;
			G645<=G28046;
			G650<=G28049;
			G655<=G28050;
			G661<=G28052;
			G667<=G25615;
			G671<=G29225;
			G676<=G29226;
			G681<=G28047;
			G686<=G25614;
			G691<=G28048;
			G699<=G28053;
			G703<=G24214;
			G714<=G29227;
			G718<=G28051;
			G723<=G29229;
			G728<=G28054;
			G732<=G25616;
			G736<=G802;
			G739<=G29228;
			G744<=G30335;
			G749<=G31867;
			G753<=G26897;
			G758<=G32979;
			G763<=G33539;
			G767<=G33965;
			G772<=G34252;
			G776<=G34439;
			G781<=G34600;
			G785<=G34725;
			G790<=G34791;
			G794<=G34850;
			G799<=G24213;
			G802<=G799;
			G807<=G34881;
			G812<=G26898;
			G817<=G25617;
			G822<=G26899;
			G827<=G28055;
			G832<=G25618;
			G837<=G24215;
			G843<=G25619;
			G847<=G24216;
			G854<=G32980;
			G859<=G26900;
			G862<=G26909;
			G869<=G859;
			G872<=G887;
			G875<=G869;
			G878<=G875;
			G881<=G878;
			G884<=G881;
			G887<=G884;
			G890<=G34440;
			G896<=G26910;
			G901<=G25620;
			G904<=G24231;
			G907<=G28056;
			G911<=G29230;
			G914<=G30336;
			G918<=G31868;
			G921<=G25621;
			G925<=G32981;
			G929<=G21725;
			G930<=G33540;
			G933<=G32982;
			G936<=G26912;
			G939<=G34727;
			G943<=G34728;
			G947<=G34601;
			G952<=G34726;
			G956<=G25626;
			G962<=G25627;
			G967<=G21722;
			G968<=G21723;
			G969<=G25622;
			G976<=G24232;
			G979<=G1116;
			G990<=G1239;
			G996<=G24243;
			G1002<=G28057;
			G1008<=G25623;
			G1018<=G30337;
			G1024<=G31869;
			G1030<=G32983;
			G1036<=G33541;
			G1041<=G25624;
			G1046<=G26913;
			G1052<=G25625;
			G1056<=G24241;
			G1061<=G26914;
			G1070<=G30341;
			G1075<=G24238;
			G1079<=G1075;
			G1083<=G1079;
			G1087<=G1083;
			G1094<=G29231;
			G1099<=G24235;
			G1105<=G26915;
			G1111<=G29234;
			G1116<=G1056;
			G1124<=G29232;
			G1129<=G26916;
			G1135<=G26917;
			G1141<=G29233;
			G1146<=G24233;
			G1152<=G24234;
			G1157<=G24240;
			G1171<=G30338;
			G1178<=G24236;
			G1183<=G30339;
			G1189<=G24237;
			G1193<=G26918;
			G1199<=G30340;
			G1205<=G24244;
			G1211<=G25628;
			G1216<=G25629;
			G1221<=G24246;
			G1227<=G24242;
			G1233<=G24239;
			G1236<=G1233;
			G1239<=G1157;
			G1242<=G1227;
			G1246<=G24245;
			G1249<=G24247;
			G1252<=G28058;
			G1256<=G29235;
			G1259<=G30342;
			G1263<=G31870;
			G1266<=G25630;
			G1270<=G32984;
			G1274<=G33542;
			G1277<=G32985;
			G1280<=G26919;
			G1283<=G34730;
			G1287<=G34731;
			G1291<=G34602;
			G1296<=G34729;
			G1300<=G25635;
			G1306<=G25636;
			G1311<=G21724;
			G1312<=G25631;
			G1319<=G24248;
			G1322<=G1459;
			G1333<=G1582;
			G1339<=G24259;
			G1345<=G28059;
			G1351<=G25632;
			G1361<=G30343;
			G1367<=G31871;
			G1373<=G32986;
			G1379<=G33543;
			G1384<=G25633;
			G1389<=G26920;
			G1395<=G25634;
			G1399<=G24257;
			G1404<=G26921;
			G1413<=G30347;
			G1418<=G24254;
			G1422<=G1418;
			G1426<=G1422;
			G1430<=G1426;
			G1437<=G29236;
			G1442<=G24251;
			G1448<=G26922;
			G1454<=G29239;
			G1459<=G1399;
			G1467<=G29237;
			G1472<=G26923;
			G1478<=G26924;
			G1484<=G29238;
			G1489<=G24249;
			G1495<=G24250;
			G1500<=G24256;
			G1514<=G30344;
			G1521<=G24252;
			G1526<=G30345;
			G1532<=G24253;
			G1536<=G26925;
			G1542<=G30346;
			G1548<=G24260;
			G1554<=G25637;
			G1559<=G25638;
			G1564<=G24262;
			G1570<=G24258;
			G1576<=G24255;
			G1579<=G1576;
			G1582<=G1500;
			G1585<=G1570;
			G1589<=G24261;
			G1592<=G33544;
			G1600<=G33966;
			G1604<=G33972;
			G1608<=G33967;
			G1612<=G33968;
			G1616<=G33969;
			G1620<=G33970;
			G1624<=G32987;
			G1632<=G30348;
			G1636<=G33545;
			G1644<=G33551;
			G1648<=G32988;
			G1657<=G32989;
			G1664<=G32990;
			G1668<=G33546;
			G1677<=G29240;
			G1682<=G33971;
			G1687<=G33547;
			G1691<=G29241;
			G1696<=G30349;
			G1700<=G30350;
			G1706<=G33548;
			G1710<=G33549;
			G1714<=G33550;
			G1720<=G30351;
			G1724<=G30352;
			G1728<=G33552;
			G1736<=G33973;
			G1740<=G33979;
			G1744<=G33974;
			G1748<=G33975;
			G1752<=G33976;
			G1756<=G33977;
			G1760<=G32991;
			G1768<=G30353;
			G1772<=G33553;
			G1779<=G33559;
			G1783<=G32992;
			G1792<=G32993;
			G1798<=G32994;
			G1802<=G33554;
			G1811<=G29242;
			G1816<=G33978;
			G1821<=G33555;
			G1825<=G29243;
			G1830<=G30354;
			G1834<=G30355;
			G1840<=G33556;
			G1844<=G33557;
			G1848<=G33558;
			G1854<=G30356;
			G1858<=G30357;
			G1862<=G33560;
			G1870<=G33980;
			G1874<=G33986;
			G1878<=G33981;
			G1882<=G33982;
			G1886<=G33983;
			G1890<=G33984;
			G1894<=G32995;
			G1902<=G30358;
			G1906<=G33561;
			G1913<=G33567;
			G1917<=G32996;
			G1926<=G32997;
			G1932<=G32998;
			G1936<=G33562;
			G1945<=G29244;
			G1950<=G33985;
			G1955<=G33563;
			G1959<=G29245;
			G1964<=G30359;
			G1968<=G30360;
			G1974<=G33564;
			G1978<=G33565;
			G1982<=G33566;
			G1988<=G30361;
			G1992<=G30362;
			G1996<=G33568;
			G2004<=G33987;
			G2008<=G33993;
			G2012<=G33988;
			G2016<=G33989;
			G2020<=G33990;
			G2024<=G33991;
			G2028<=G32999;
			G2036<=G30363;
			G2040<=G33569;
			G2047<=G33575;
			G2051<=G33000;
			G2060<=G33001;
			G2066<=G33002;
			G2070<=G33570;
			G2079<=G29246;
			G2084<=G33992;
			G2089<=G33571;
			G2093<=G29247;
			G2098<=G30364;
			G2102<=G30365;
			G2108<=G33572;
			G2112<=G33573;
			G2116<=G33574;
			G2122<=G30366;
			G2126<=G30367;
			G2130<=G34603;
			G2138<=G34604;
			G2145<=G34605;
			G2151<=G18421;
			G2152<=G18422;
			G2153<=G33576;
			G2161<=G33994;
			G2165<=G34000;
			G2169<=G33995;
			G2173<=G33996;
			G2177<=G33997;
			G2181<=G33998;
			G2185<=G33003;
			G2193<=G30368;
			G2197<=G33577;
			G2204<=G33583;
			G2208<=G33004;
			G2217<=G33005;
			G2223<=G33006;
			G2227<=G33578;
			G2236<=G29248;
			G2241<=G33999;
			G2246<=G33579;
			G2250<=G29249;
			G2255<=G30369;
			G2259<=G30370;
			G2265<=G33580;
			G2269<=G33581;
			G2273<=G33582;
			G2279<=G30371;
			G2283<=G30372;
			G2287<=G33584;
			G2295<=G34001;
			G2299<=G34007;
			G2303<=G34002;
			G2307<=G34003;
			G2311<=G34004;
			G2315<=G34005;
			G2319<=G33007;
			G2327<=G30373;
			G2331<=G33585;
			G2338<=G33591;
			G2342<=G33008;
			G2351<=G33009;
			G2357<=G33010;
			G2361<=G33586;
			G2370<=G29250;
			G2375<=G34006;
			G2380<=G33587;
			G2384<=G29251;
			G2389<=G30374;
			G2393<=G30375;
			G2399<=G33588;
			G2403<=G33589;
			G2407<=G33590;
			G2413<=G30376;
			G2417<=G30377;
			G2421<=G33592;
			G2429<=G34008;
			G2433<=G34014;
			G2437<=G34009;
			G2441<=G34010;
			G2445<=G34011;
			G2449<=G34012;
			G2453<=G33011;
			G2461<=G30378;
			G2465<=G33593;
			G2472<=G33599;
			G2476<=G33012;
			G2485<=G33013;
			G2491<=G33014;
			G2495<=G33594;
			G2504<=G29252;
			G2509<=G34013;
			G2514<=G33595;
			G2518<=G29253;
			G2523<=G30379;
			G2527<=G30380;
			G2533<=G33596;
			G2537<=G33597;
			G2541<=G33598;
			G2547<=G30381;
			G2551<=G30382;
			G2555<=G33600;
			G2563<=G34015;
			G2567<=G34021;
			G2571<=G34016;
			G2575<=G34017;
			G2579<=G34018;
			G2583<=G34019;
			G2587<=G33015;
			G2595<=G30383;
			G2599<=G33601;
			G2606<=G33607;
			G2610<=G33016;
			G2619<=G33017;
			G2625<=G33018;
			G2629<=G33602;
			G2638<=G29254;
			G2643<=G34020;
			G2648<=G33603;
			G2652<=G29255;
			G2657<=G30384;
			G2661<=G30385;
			G2667<=G33604;
			G2671<=G33605;
			G2675<=G33606;
			G2681<=G30386;
			G2685<=G30387;
			G2689<=G34606;
			G2697<=G34607;
			G2704<=G34608;
			G2710<=G18527;
			G2711<=G18528;
			G2712<=G26937;
			G2715<=G24263;
			G2719<=G25639;
			G2724<=G26926;
			G2729<=G28060;
			G2735<=G29256;
			G2741<=G30388;
			G2748<=G31872;
			G2756<=G33019;
			G2759<=G33608;
			G2763<=G34022;
			G2767<=G26927;
			G2771<=G34441;
			G2775<=G34443;
			G2779<=G26928;
			G2783<=G34442;
			G2787<=G34444;
			G2791<=G26929;
			G2795<=G26930;
			G2799<=G26931;
			G2803<=G34445;
			G2807<=G34447;
			G2811<=G26932;
			G2815<=G34446;
			G2819<=G34448;
			G2823<=G26933;
			G2827<=G26934;
			G2831<=G30391;
			G2834<=G30392;
			G2837<=G26935;
			G2841<=G26936;
			G2844<=G34609;
			G2848<=G34792;
			G2852<=G34610;
			G2856<=G34793;
			G2860<=G34611;
			G2864<=G34794;
			G2868<=G34616;
			G2873<=G34615;
			G2878<=G34797;
			G2882<=G34796;
			G2886<=G34798;
			G2890<=G34799;
			G2894<=G34612;
			G2898<=G34795;
			G2902<=G34801;
			G2907<=G34617;
			G2912<=G34618;
			G2917<=G34802;
			G2922<=G34619;
			G2927<=G34803;
			G2932<=G24282;
			G2936<=G34620;
			G2941<=G34806;
			G2946<=G21899;
			G2950<=G34621;
			G2955<=G34807;
			G2960<=G34622;
			G2965<=G34808;
			G2970<=G34623;
			G2975<=G34804;
			G2980<=G34800;
			G2984<=G34980;
			G2988<=G34624;
			G2994<=G34732;
			G2999<=G34805;
			G3003<=G21726;
			G3004<=G31873;
			G3010<=G25651;
			G3017<=G31877;
			G3021<=G31879;
			G3025<=G31874;
			G3029<=G31875;
			G3034<=G31876;
			G3040<=G31878;
			G3045<=G33020;
			G3050<=G25650;
			G3057<=G28062;
			G3061<=G28061;
			G3065<=G25652;
			G3068<=G25643;
			G3072<=G25644;
			G3080<=G25645;
			G3085<=G25646;
			G3089<=G25647;
			G3092<=G25648;
			G3096<=G25649;
			G3100<=G3092;
			G3103<=G3096;
			G3106<=G29257;
			G3111<=G25656;
			G3115<=G29258;
			G3119<=G25653;
			G3125<=G29259;
			G3129<=G29260;
			G3133<=G29261;
			G3139<=G25654;
			G3143<=G25655;
			G3147<=G29262;
			G3151<=G34625;
			G3155<=G30393;
			G3161<=G33021;
			G3167<=G33022;
			G3171<=G33023;
			G3179<=G33024;
			G3187<=G30394;
			G3191<=G30395;
			G3195<=G30410;
			G3199<=G30396;
			G3203<=G30411;
			G3207<=G30397;
			G3211<=G30412;
			G3215<=G30398;
			G3219<=G30399;
			G3223<=G30400;
			G3227<=G30401;
			G3231<=G30402;
			G3235<=G30403;
			G3239<=G30404;
			G3243<=G30405;
			G3247<=G30406;
			G3251<=G30407;
			G3255<=G30408;
			G3259<=G30409;
			G3263<=G30413;
			G3267<=G3310;
			G3274<=G3267;
			G3281<=G3303;
			G3288<=G33610;
			G3298<=G3274;
			G3303<=G24267;
			G3310<=G3281;
			G3317<=G3298;
			G3321<=G3317;
			G3325<=G3321;
			G3329<=G3325;
			G3333<=G28063;
			G3338<=G24268;
			G3343<=G24269;
			G3347<=G24270;
			G3352<=G33609;
			G3355<=G31880;
			G3361<=G25665;
			G3368<=G31884;
			G3372<=G31886;
			G3376<=G31881;
			G3380<=G31882;
			G3385<=G31883;
			G3391<=G31885;
			G3396<=G33025;
			G3401<=G25664;
			G3408<=G28065;
			G3412<=G28064;
			G3416<=G25666;
			G3419<=G25657;
			G3423<=G25658;
			G3431<=G25659;
			G3436<=G25660;
			G3440<=G25661;
			G3443<=G25662;
			G3447<=G25663;
			G3451<=G3443;
			G3454<=G3447;
			G3457<=G29263;
			G3462<=G25670;
			G3466<=G29264;
			G3470<=G25667;
			G3476<=G29265;
			G3480<=G29266;
			G3484<=G29267;
			G3490<=G25668;
			G3494<=G25669;
			G3498<=G29268;
			G3502<=G34626;
			G3506<=G30414;
			G3512<=G33026;
			G3518<=G33027;
			G3522<=G33028;
			G3530<=G33029;
			G3538<=G30415;
			G3542<=G30416;
			G3546<=G30431;
			G3550<=G30417;
			G3554<=G30432;
			G3558<=G30418;
			G3562<=G30433;
			G3566<=G30419;
			G3570<=G30420;
			G3574<=G30421;
			G3578<=G30422;
			G3582<=G30423;
			G3586<=G30424;
			G3590<=G30425;
			G3594<=G30426;
			G3598<=G30427;
			G3602<=G30428;
			G3606<=G30429;
			G3610<=G30430;
			G3614<=G30434;
			G3618<=G3661;
			G3625<=G3618;
			G3632<=G3654;
			G3639<=G33612;
			G3649<=G3625;
			G3654<=G24271;
			G3661<=G3632;
			G3668<=G3649;
			G3672<=G3668;
			G3676<=G3672;
			G3680<=G3676;
			G3684<=G28066;
			G3689<=G24272;
			G3694<=G24273;
			G3698<=G24274;
			G3703<=G33611;
			G3706<=G31887;
			G3712<=G25679;
			G3719<=G31891;
			G3723<=G31893;
			G3727<=G31888;
			G3731<=G31889;
			G3736<=G31890;
			G3742<=G31892;
			G3747<=G33030;
			G3752<=G25678;
			G3759<=G28068;
			G3763<=G28067;
			G3767<=G25680;
			G3770<=G25671;
			G3774<=G25672;
			G3782<=G25673;
			G3787<=G25674;
			G3791<=G25675;
			G3794<=G25676;
			G3798<=G25677;
			G3802<=G3794;
			G3805<=G3798;
			G3808<=G29269;
			G3813<=G25684;
			G3817<=G29270;
			G3821<=G25681;
			G3827<=G29271;
			G3831<=G29272;
			G3835<=G29273;
			G3841<=G25682;
			G3845<=G25683;
			G3849<=G29274;
			G3853<=G34627;
			G3857<=G30435;
			G3863<=G33031;
			G3869<=G33032;
			G3873<=G33033;
			G3881<=G33034;
			G3889<=G30436;
			G3893<=G30437;
			G3897<=G30452;
			G3901<=G30438;
			G3905<=G30453;
			G3909<=G30439;
			G3913<=G30454;
			G3917<=G30440;
			G3921<=G30441;
			G3925<=G30442;
			G3929<=G30443;
			G3933<=G30444;
			G3937<=G30445;
			G3941<=G30446;
			G3945<=G30447;
			G3949<=G30448;
			G3953<=G30449;
			G3957<=G30450;
			G3961<=G30451;
			G3965<=G30455;
			G3969<=G4012;
			G3976<=G3969;
			G3983<=G4005;
			G3990<=G33614;
			G4000<=G3976;
			G4005<=G24275;
			G4012<=G3983;
			G4019<=G4000;
			G4023<=G4019;
			G4027<=G4023;
			G4031<=G4027;
			G4035<=G28069;
			G4040<=G24276;
			G4045<=G24277;
			G4049<=G24278;
			G4054<=G33613;
			G4057<=G25686;
			G4064<=G25685;
			G4072<=G25691;
			G4076<=G28070;
			G4082<=G26938;
			G4087<=G29275;
			G4093<=G30456;
			G4098<=G31894;
			G4104<=G33615;
			G4108<=G33035;
			G4112<=G28071;
			G4116<=G28072;
			G4119<=G28073;
			G4122<=G28074;
			G4125<=G28081;
			G4129<=G28075;
			G4132<=G28076;
			G4135<=G28077;
			G4138<=G28078;
			G4141<=G25687;
			G4145<=G26939;
			G4146<=G34628;
			G4153<=G30457;
			G4157<=G34629;
			G4164<=G26940;
			G4165<=G28079;
			G4169<=G28080;
			G4172<=G34733;
			G4176<=G34734;
			G4180<=G4210;
			G4185<=G21891;
			G4188<=G4191;
			G4191<=G21901;
			G4194<=G4188;
			G4197<=G4194;
			G4200<=G4197;
			G4204<=G4200;
			G4207<=G4204;
			G4210<=G4207;
			G4213<=G4185;
			G4216<=G4213;
			G4219<=G4216;
			G4222<=G4219;
			G4226<=G4222;
			G4229<=G4226;
			G4232<=G4229;
			G4235<=G4232;
			G4239<=G21892;
			G4242<=G24279;
			G4245<=G34632;
			G4249<=G34631;
			G4253<=G34630;
			G4258<=G21893;
			G4264<=G21894;
			G4269<=G21895;
			G4273<=G24280;
			G4277<=G21896;
			G4281<=G4277;
			G4284<=G21897;
			G4287<=G21898;
			G4291<=G4287;
			G4294<=G21900;
			G4297<=G4294;
			G4300<=G34735;
			G4304<=G24281;
			G4308<=G4304;
			G4311<=G34449;
			G4322<=G34450;
			G4332<=G34455;
			G4340<=G34459;
			G4349<=G34257;
			G4358<=G34258;
			G4366<=G26944;
			G4369<=G26970;
			G4372<=G34882;
			G4375<=G26951;
			G4382<=G26947;
			G4388<=G26949;
			G4392<=G26950;
			G4401<=G26948;
			G4405<=G4408;
			G4408<=G26945;
			G4411<=G4414;
			G4414<=G26946;
			G4417<=G31895;
			G4420<=G26965;
			G4423<=G4537;
			G4427<=G26952;
			G4430<=G26957;
			G4434<=G26956;
			G4438<=G26953;
			G4443<=G4449;
			G4446<=G26954;
			G4449<=G26955;
			G4452<=G4446;
			G4455<=G26959;
			G4456<=G25692;
			G4459<=G34253;
			G4462<=G34254;
			G4467<=G34255;
			G4473<=G34256;
			G4474<=G10384;
			G4477<=G26960;
			G4480<=G31896;
			G4483<=G4520;
			G4486<=G26961;
			G4489<=G26962;
			G4492<=G26963;
			G4495<=G33036;
			G4498<=G33037;
			G4501<=G33038;
			G4504<=G33039;
			G4507<=G30458;
			G4512<=G33040;
			G4515<=G26964;
			G4519<=G33616;
			G4520<=G6972;
			G4521<=G26971;
			G4527<=G28082;
			G4531<=G24335;
			G4534<=G34023;
			G4537<=G34024;
			G4540<=G31897;
			G4543<=G33042;
			G4546<=G33045;
			G4549<=G33041;
			G4552<=G33044;
			G4555<=G4571;
			G4558<=G26966;
			G4561<=G26968;
			G4564<=G26967;
			G4567<=G33043;
			G4570<=G33617;
			G4571<=G6974;
			G4572<=G29279;
			G4575<=G29276;
			G4578<=G29278;
			G4581<=G26969;
			G4584<=G34451;
			G4593<=G34452;
			G4601<=G34453;
			G4608<=G34454;
			G4616<=G34456;
			G4621<=G34460;
			G4628<=G34457;
			G4633<=G34458;
			G4639<=G34025;
			G4643<=G34259;
			G4646<=G34260;
			G4653<=G34462;
			G4659<=G34461;
			G4664<=G34463;
			G4669<=G34464;
			G4674<=G34026;
			G4681<=G34027;
			G4688<=G34028;
			G4698<=G34261;
			G4704<=G28083;
			G4709<=G34032;
			G4717<=G34635;
			G4722<=G34636;
			G4727<=G34633;
			G4732<=G34634;
			G4737<=G34637;
			G4741<=G21902;
			G4742<=G21903;
			G4743<=G34262;
			G4749<=G28084;
			G4754<=G34263;
			G4760<=G28085;
			G4765<=G34264;
			G4771<=G28086;
			G4776<=G34031;
			G4785<=G34029;
			G4793<=G34033;
			G4801<=G34030;
			G4809<=G25693;
			G4812<=G4809;
			G4815<=G4812;
			G4818<=G4815;
			G4821<=G28096;
			G4826<=G28102;
			G4831<=G28099;
			G4836<=G34265;
			G4843<=G34466;
			G4849<=G34465;
			G4854<=G34467;
			G4859<=G34468;
			G4864<=G34034;
			G4871<=G34035;
			G4878<=G34036;
			G4888<=G34266;
			G4894<=G28087;
			G4899<=G34040;
			G4907<=G34640;
			G4912<=G34641;
			G4917<=G34638;
			G4922<=G34639;
			G4927<=G34642;
			G4931<=G21904;
			G4932<=G21905;
			G4933<=G34267;
			G4939<=G28088;
			G4944<=G34268;
			G4950<=G28089;
			G4955<=G34269;
			G4961<=G28090;
			G4966<=G34039;
			G4975<=G34037;
			G4983<=G34041;
			G4991<=G34038;
			G4999<=G25694;
			G5002<=G4999;
			G5005<=G5002;
			G5008<=G5005;
			G5011<=G28105;
			G5016<=G31898;
			G5022<=G25703;
			G5029<=G31902;
			G5033<=G31904;
			G5037<=G31899;
			G5041<=G31900;
			G5046<=G31901;
			G5052<=G31903;
			G5057<=G33046;
			G5062<=G25702;
			G5069<=G28092;
			G5073<=G28091;
			G5077<=G25704;
			G5080<=G25695;
			G5084<=G25696;
			G5092<=G25697;
			G5097<=G25698;
			G5101<=G25700;
			G5105<=G25701;
			G5109<=G5101;
			G5112<=G5105;
			G5115<=G29280;
			G5120<=G25708;
			G5124<=G29281;
			G5128<=G25705;
			G5134<=G29282;
			G5138<=G29283;
			G5142<=G29284;
			G5148<=G25706;
			G5152<=G25707;
			G5156<=G29285;
			G5160<=G34643;
			G5164<=G30459;
			G5170<=G33047;
			G5176<=G33048;
			G5180<=G33049;
			G5188<=G33050;
			G5196<=G30460;
			G5200<=G30461;
			G5204<=G30476;
			G5208<=G30462;
			G5212<=G30477;
			G5216<=G30463;
			G5220<=G30478;
			G5224<=G30464;
			G5228<=G30465;
			G5232<=G30466;
			G5236<=G30467;
			G5240<=G30468;
			G5244<=G30469;
			G5248<=G30470;
			G5252<=G30471;
			G5256<=G30472;
			G5260<=G30473;
			G5264<=G30474;
			G5268<=G30475;
			G5272<=G30479;
			G5276<=G5320;
			G5283<=G5276;
			G5290<=G5313;
			G5297<=G33619;
			G5308<=G5283;
			G5313<=G24336;
			G5320<=G5290;
			G5327<=G5308;
			G5331<=G5327;
			G5335<=G5331;
			G5339<=G5335;
			G5343<=G24337;
			G5348<=G24338;
			G5352<=G24339;
			G5357<=G33618;
			G5360<=G31905;
			G5366<=G25717;
			G5373<=G31909;
			G5377<=G31911;
			G5381<=G31906;
			G5385<=G31907;
			G5390<=G31908;
			G5396<=G31910;
			G5401<=G33051;
			G5406<=G25716;
			G5413<=G28095;
			G5417<=G28094;
			G5421<=G25718;
			G5424<=G25709;
			G5428<=G25710;
			G5436<=G25711;
			G5441<=G25712;
			G5445<=G25713;
			G5448<=G25714;
			G5452<=G25715;
			G5456<=G5448;
			G5459<=G5452;
			G5462<=G29286;
			G5467<=G25722;
			G5471<=G29287;
			G5475<=G25719;
			G5481<=G29288;
			G5485<=G29289;
			G5489<=G29290;
			G5495<=G25720;
			G5499<=G25721;
			G5503<=G29291;
			G5507<=G34644;
			G5511<=G30480;
			G5517<=G33052;
			G5523<=G33053;
			G5527<=G33054;
			G5535<=G33055;
			G5543<=G30481;
			G5547<=G30482;
			G5551<=G30497;
			G5555<=G30483;
			G5559<=G30498;
			G5563<=G30484;
			G5567<=G30499;
			G5571<=G30485;
			G5575<=G30486;
			G5579<=G30487;
			G5583<=G30488;
			G5587<=G30489;
			G5591<=G30490;
			G5595<=G30491;
			G5599<=G30492;
			G5603<=G30493;
			G5607<=G30494;
			G5611<=G30495;
			G5615<=G30496;
			G5619<=G30500;
			G5623<=G5666;
			G5630<=G5623;
			G5637<=G5659;
			G5644<=G33621;
			G5654<=G5630;
			G5659<=G24340;
			G5666<=G5637;
			G5673<=G5654;
			G5677<=G5673;
			G5681<=G5677;
			G5685<=G5681;
			G5689<=G24341;
			G5694<=G24342;
			G5698<=G24343;
			G5703<=G33620;
			G5706<=G31912;
			G5712<=G25731;
			G5719<=G31916;
			G5723<=G31918;
			G5727<=G31913;
			G5731<=G31914;
			G5736<=G31915;
			G5742<=G31917;
			G5747<=G33056;
			G5752<=G25730;
			G5759<=G28098;
			G5763<=G28097;
			G5767<=G25732;
			G5770<=G25723;
			G5774<=G25724;
			G5782<=G25725;
			G5787<=G25726;
			G5791<=G25727;
			G5794<=G25728;
			G5798<=G25729;
			G5802<=G5794;
			G5805<=G5798;
			G5808<=G29292;
			G5813<=G25736;
			G5817<=G29293;
			G5821<=G25733;
			G5827<=G29294;
			G5831<=G29295;
			G5835<=G29296;
			G5841<=G25734;
			G5845<=G25735;
			G5849<=G29297;
			G5853<=G34645;
			G5857<=G30501;
			G5863<=G33057;
			G5869<=G33058;
			G5873<=G33059;
			G5881<=G33060;
			G5889<=G30502;
			G5893<=G30503;
			G5897<=G30518;
			G5901<=G30504;
			G5905<=G30519;
			G5909<=G30505;
			G5913<=G30520;
			G5917<=G30506;
			G5921<=G30507;
			G5925<=G30508;
			G5929<=G30509;
			G5933<=G30510;
			G5937<=G30511;
			G5941<=G30512;
			G5945<=G30513;
			G5949<=G30514;
			G5953<=G30515;
			G5957<=G30516;
			G5961<=G30517;
			G5965<=G30521;
			G5969<=G6012;
			G5976<=G5969;
			G5983<=G6005;
			G5990<=G33623;
			G6000<=G5976;
			G6005<=G24344;
			G6012<=G5983;
			G6019<=G6000;
			G6023<=G6019;
			G6027<=G6023;
			G6031<=G6027;
			G6035<=G24345;
			G6040<=G24346;
			G6044<=G24347;
			G6049<=G33622;
			G6052<=G31919;
			G6058<=G25745;
			G6065<=G31923;
			G6069<=G31925;
			G6073<=G31920;
			G6077<=G31921;
			G6082<=G31922;
			G6088<=G31924;
			G6093<=G33061;
			G6098<=G25744;
			G6105<=G28101;
			G6109<=G28100;
			G6113<=G25746;
			G6116<=G25737;
			G6120<=G25738;
			G6128<=G25739;
			G6133<=G25740;
			G6137<=G25741;
			G6140<=G25742;
			G6144<=G25743;
			G6148<=G6140;
			G6151<=G6144;
			G6154<=G29298;
			G6159<=G25750;
			G6163<=G29299;
			G6167<=G25747;
			G6173<=G29300;
			G6177<=G29301;
			G6181<=G29302;
			G6187<=G25748;
			G6191<=G25749;
			G6195<=G29303;
			G6199<=G34646;
			G6203<=G30522;
			G6209<=G33062;
			G6215<=G33063;
			G6219<=G33064;
			G6227<=G33065;
			G6235<=G30523;
			G6239<=G30524;
			G6243<=G30539;
			G6247<=G30525;
			G6251<=G30540;
			G6255<=G30526;
			G6259<=G30541;
			G6263<=G30527;
			G6267<=G30528;
			G6271<=G30529;
			G6275<=G30530;
			G6279<=G30531;
			G6283<=G30532;
			G6287<=G30533;
			G6291<=G30534;
			G6295<=G30535;
			G6299<=G30536;
			G6303<=G30537;
			G6307<=G30538;
			G6311<=G30542;
			G6315<=G6358;
			G6322<=G6315;
			G6329<=G6351;
			G6336<=G33625;
			G6346<=G6322;
			G6351<=G24348;
			G6358<=G6329;
			G6365<=G6346;
			G6369<=G6365;
			G6373<=G6369;
			G6377<=G6373;
			G6381<=G24349;
			G6386<=G24350;
			G6390<=G24351;
			G6395<=G33624;
			G6398<=G31926;
			G6404<=G25759;
			G6411<=G31930;
			G6415<=G31932;
			G6419<=G31927;
			G6423<=G31928;
			G6428<=G31929;
			G6434<=G31931;
			G6439<=G33066;
			G6444<=G25758;
			G6451<=G28104;
			G6455<=G28103;
			G6459<=G25760;
			G6462<=G25751;
			G6466<=G25752;
			G6474<=G25753;
			G6479<=G25754;
			G6483<=G25755;
			G6486<=G25756;
			G6490<=G25757;
			G6494<=G6486;
			G6497<=G6490;
			G6500<=G29304;
			G6505<=G25764;
			G6509<=G29305;
			G6513<=G25761;
			G6519<=G29306;
			G6523<=G29307;
			G6527<=G29308;
			G6533<=G25762;
			G6537<=G25763;
			G6541<=G29309;
			G6545<=G34647;
			G6549<=G30543;
			G6555<=G33067;
			G6561<=G33068;
			G6565<=G33069;
			G6573<=G33070;
			G6581<=G30544;
			G6585<=G30545;
			G6589<=G30560;
			G6593<=G30546;
			G6597<=G30561;
			G6601<=G30547;
			G6605<=G30562;
			G6609<=G30548;
			G6613<=G30549;
			G6617<=G30550;
			G6621<=G30551;
			G6625<=G30552;
			G6629<=G30553;
			G6633<=G30554;
			G6637<=G30555;
			G6641<=G30556;
			G6645<=G30557;
			G6649<=G30558;
			G6653<=G30559;
			G6657<=G30563;
			G6661<=G6704;
			G6668<=G6661;
			G6675<=G6697;
			G6682<=G33627;
			G6692<=G6668;
			G6697<=G24352;
			G6704<=G6675;
			G6711<=G6692;
			G6715<=G6711;
			G6719<=G6715;
			G6723<=G6719;
			G6727<=G24353;
			G6732<=G24354;
			G6736<=G24355;
			G6741<=G33626;
		end if;
	end process;
	G6754<= not I11617;
	G6755<= not I11620;
	G6756<= not I11623;
	G6767<= not I11626;
	G6772<= not I11629;
	G6782<= not I11632;
	G6789<= not I11635;
	G6799<= not G199;
	G6800<= not G203;
	G6801<= not G391;
	G6802<= not G468;
	G6803<= not G496;
	G6804<= not G490;
	G6808<= not G554;
	G6809<= not G341;
	G6810<= not G723;
	G6811<= not G714;
	G6814<= not G632;
	G6815<= not G929;
	G6816<= not G933;
	G6817<= not G956;
	G6818<= not G976;
	G6819<= not G1046;
	G6820<= not G1070;
	G6821<= not I11655;
	G6825<= not G979;
	G6826<= not G218;
	G6827<= not G1277;
	G6828<= not G1300;
	G6829<= not G1319;
	G6830<= not G1389;
	G6831<= not G1413;
	G6832<= not I11665;
	G6836<= not G1322;
	G6837<= not G968;
	G6838<= not G1724;
	G6839<= not G1858;
	G6840<= not G1992;
	G6841<= not G2145;
	G6845<= not G2126;
	G6846<= not G2152;
	G6847<= not G2283;
	G6848<= not G2417;
	G6849<= not G2551;
	G6850<= not G2704;
	G6854<= not G2685;
	G6855<= not G2711;
	G6856<= not I11682;
	G6867<= not I11685;
	G6868<= not I11688;
	G6869<= not I11691;
	G6870<= not G3089;
	G6873<= not G3151;
	G6874<= not G3143;
	G6875<= not I11697;
	G6887<= not G3333;
	G6888<= not I11701;
	G6895<= not G3288;
	G6900<= not G3440;
	G6903<= not G3502;
	G6904<= not G3494;
	G6905<= not I11708;
	G6917<= not G3684;
	G6918<= not G3639;
	G6923<= not G3791;
	G6926<= not G3853;
	G6927<= not G3845;
	G6928<= not I11716;
	G6940<= not G4035;
	G6941<= not G3990;
	G6946<= not I11721;
	G6953<= not G4157;
	G6954<= not G4138;
	G6955<= not I11726;
	G6956<= not G4242;
	G6957<= not G2932;
	G6958<= not G4372;
	G6959<= not G4420;
	G6960<= not G1;
	G6961<= not I11734;
	G6971<= not I11737;
	G6972<= not I11740;
	G6973<= not I11743;
	G6974<= not I11746;
	G6975<= not G4507;
	G6976<= not I11750;
	G6977<= not I11753;
	G6978<= not G4616;
	G6982<= not G4531;
	G6983<= not G4698;
	G6984<= not G4709;
	G6985<= not G4669;
	G6986<= not G4743;
	G6987<= not G4754;
	G6988<= not G4765;
	G6989<= not G4575;
	G6990<= not G4742;
	G6991<= not G4888;
	G6992<= not G4899;
	G6993<= not G4859;
	G6994<= not G4933;
	G6995<= not G4944;
	G6996<= not G4955;
	G6997<= not G4578;
	G6998<= not G4932;
	G6999<= not G86;
	G7002<= not G5160;
	G7003<= not G5152;
	G7004<= not I11777;
	G7017<= not G128;
	G7018<= not G5297;
	G7023<= not G5445;
	G7026<= not G5507;
	G7027<= not G5499;
	G7028<= not I11785;
	G7040<= not G4821;
	G7041<= not G5644;
	G7046<= not G5791;
	G7049<= not G5853;
	G7050<= not G5845;
	G7051<= not I11793;
	G7063<= not G4831;
	G7064<= not G5990;
	G7069<= not G6137;
	G7072<= not G6199;
	G7073<= not G6191;
	G7074<= not I11801;
	G7086<= not G4826;
	G7087<= not G6336;
	G7092<= not G6483;
	G7095<= not G6545;
	G7096<= not G6537;
	G7097<= not I11809;
	G7109<= not G5011;
	G7110<= not G6682;
	G7115<= not G12;
	G7116<= not G22;
	G7117<= not I11816;
	G7118<= not G832;
	G7121<= not I11820;
	G7132<= not G4558;
	G7134<= not G5029;
	G7138<= not G5360;
	G7148<= not I11835;
	G7149<= not G4564;
	G7153<= not G5373;
	G7157<= not G5706;
	G7161<= not I11843;
	G7162<= not G4521;
	G7163<= not G4593;
	G7166<= not G4311;
	G7170<= not G5719;
	G7174<= not G6052;
	G7178<= not G4392;
	G7183<= not G4608;
	G7187<= not G6065;
	G7191<= not G6398;
	G7195<= not G25;
	G7196<= not I11860;
	G7197<= not G812;
	G7202<= not G4639;
	G7212<= not G6411;
	G7216<= not G822;
	G7219<= not G4405;
	G7222<= not G4427;
	G7224<= not G4601;
	G7231<= not G5;
	G7232<= not G4411;
	G7235<= not G4521;
	G7236<= not G4608;
	G7239<= not G5033;
	G7243<= not I11892;
	G7244<= not G4408;
	G7245<= not I11896;
	G7246<= not G4446;
	G7247<= not G5377;
	G7252<= not G1592;
	G7257<= not I11903;
	G7258<= not G4414;
	G7259<= not G4375;
	G7260<= not I11908;
	G7261<= not G4449;
	G7262<= not G5723;
	G7266<= not G35;
	G7267<= not G1604;
	G7268<= not G1636;
	G7275<= not G1728;
	G7280<= not G2153;
	G7285<= not G4643;
	G7289<= not G4382;
	G7293<= not G4452;
	G7296<= not G5313;
	G7297<= not G6069;
	G7301<= not G925;
	G7308<= not G1668;
	G7314<= not G1740;
	G7315<= not G1772;
	G7322<= not G1862;
	G7327<= not G2165;
	G7328<= not G2197;
	G7335<= not G2287;
	G7340<= not G4443;
	G7343<= not G5290;
	G7344<= not G5659;
	G7345<= not G6415;
	G7349<= not G1270;
	G7356<= not G1802;
	G7361<= not G1874;
	G7362<= not G1906;
	G7369<= not G1996;
	G7374<= not G2227;
	G7379<= not G2299;
	G7380<= not G2331;
	G7387<= not G2421;
	G7392<= not G4438;
	G7393<= not G5320;
	G7394<= not G5637;
	G7395<= not G6005;
	G7397<= not G890;
	G7400<= not G911;
	G7405<= not G1936;
	G7410<= not G2008;
	G7411<= not G2040;
	G7418<= not G2361;
	G7423<= not G2433;
	G7424<= not G2465;
	G7431<= not G2555;
	G7436<= not G5276;
	G7437<= not G5666;
	G7438<= not G5983;
	G7439<= not G6351;
	G7440<= not G329;
	G7441<= not G862;
	G7443<= not G914;
	G7446<= not G1256;
	G7451<= not G2070;
	G7456<= not G2495;
	G7461<= not G2567;
	G7462<= not G2599;
	G7470<= not G5623;
	G7471<= not G6012;
	G7472<= not G6329;
	G7473<= not G6697;
	G7474<= not I11980;
	G7475<= not G896;
	G7479<= not G1008;
	G7487<= not G1259;
	G7490<= not G2629;
	G7495<= not G4375;
	G7496<= not G5969;
	G7497<= not G6358;
	G7498<= not G6675;
	G7502<= not I11992;
	G7503<= not G1351;
	G7512<= not G5283;
	G7513<= not G6315;
	G7514<= not G6704;
	G7515<= not I12000;
	G7516<= not I12003;
	G7517<= not G962;
	G7518<= not G1024;
	G7519<= not G1157;
	G7521<= not G5630;
	G7522<= not G6661;
	G7523<= not G305;
	G7526<= not I12013;
	G7527<= not I12016;
	G7528<= not G930;
	G7532<= not G1157;
	G7533<= not G1306;
	G7534<= not G1367;
	G7535<= not G1500;
	G7536<= not G5976;
	G7537<= not G311;
	G7540<= not I12026;
	G7541<= not G344;
	G7542<= not I12030;
	G7543<= not I12033;
	G7544<= not G918;
	G7548<= not G1036;
	G7553<= not G1274;
	G7557<= not G1500;
	G7558<= not I12041;
	G7563<= not G6322;
	G7564<= not G336;
	G7565<= not I12046;
	G7566<= not I12049;
	G7577<= not G1263;
	G7581<= not G1379;
	G7586<= not I12056;
	G7591<= not G6668;
	G7592<= not G347;
	G7593<= not I12061;
	G7594<= not I12064;
	G7595<= not I12067;
	G7596<= not I12070;
	G7597<= not G952;
	G7615<= not I12083;
	G7616<= not I12086;
	G7617<= not I12089;
	G7618<= not I12092;
	G7619<= not G1296;
	G7623<= not I12103;
	G7624<= not I12106;
	G7625<= not I12109;
	G7626<= not I12112;
	G7627<= not G4311;
	G7631<= not G74;
	G7632<= not I12117;
	G7633<= not I12120;
	G7634<= not I12123;
	G7635<= not G1002;
	G7636<= not G4098;
	G7640<= not I12128;
	G7643<= not G4322;
	G7647<= not I12132;
	G7648<= not I12135;
	G7649<= not G1345;
	G7650<= not G4064;
	G7655<= not G4332;
	G7659<= not I12141;
	G7660<= not I12144;
	G7666<= not G4076;
	G7670<= not G4104;
	G7674<= not I12151;
	G7680<= not G4108;
	G7686<= not G4659;
	G7689<= not I12159;
	G7693<= not G4849;
	G7697<= not G4087;
	G7704<= not I12167;
	G7715<= not G1178;
	G7716<= not G1199;
	G7717<= not I12172;
	G7733<= not G4093;
	G7738<= not I12176;
	G7749<= not G996;
	G7750<= not G1070;
	G7751<= not G1521;
	G7752<= not G1542;
	G7753<= not I12183;
	G7765<= not G4165;
	G7766<= not I12189;
	G7778<= not G1339;
	G7779<= not G1413;
	G7780<= not G2878;
	G7785<= not G4621;
	G7788<= not G4674;
	G7791<= not I12199;
	G7802<= not G324;
	G7805<= not G4366;
	G7806<= not G4681;
	G7809<= not G4864;
	G7812<= not I12214;
	G7824<= not G4169;
	G7827<= not G4688;
	G7828<= not G4871;
	G7831<= not I12227;
	G7835<= not G4125;
	G7840<= not G4878;
	G7841<= not G904;
	G7845<= not G1146;
	G7851<= not G921;
	G7854<= not G1152;
	G7858<= not G947;
	G7863<= not G1249;
	G7867<= not G1489;
	G7868<= not G1099;
	G7870<= not G1193;
	G7873<= not G1266;
	G7876<= not G1495;
	G7880<= not G1291;
	G7886<= not G1442;
	G7888<= not G1536;
	G7891<= not G2994;
	G7892<= not G4801;
	G7898<= not G4991;
	G7903<= not G969;
	G7907<= not G3072;
	G7908<= not G4157;
	G7909<= not G936;
	G7913<= not G1052;
	G7916<= not I12300;
	G7917<= not G1157;
	G7922<= not G1312;
	G7926<= not G3423;
	G7927<= not G4064;
	G7928<= not G4776;
	G7933<= not G907;
	G7936<= not G1061;
	G7939<= not G1280;
	G7943<= not G1395;
	G7946<= not I12314;
	G7947<= not G1500;
	G7952<= not G3774;
	G7953<= not G4966;
	G7957<= not G1252;
	G7960<= not G1404;
	G7963<= not G4146;
	G7964<= not G3155;
	G7970<= not G4688;
	G7971<= not G4818;
	G7972<= not G1046;
	G7975<= not G3040;
	G7980<= not G3161;
	G7985<= not G3506;
	G7991<= not G4878;
	G7992<= not G5008;
	G7993<= not I12333;
	G7994<= not I12336;
	G7995<= not G153;
	G7998<= not G392;
	G8002<= not G1389;
	G8005<= not G3025;
	G8009<= not G3106;
	G8011<= not G3167;
	G8016<= not G3391;
	G8021<= not G3512;
	G8026<= not G3857;
	G8032<= not I12355;
	G8033<= not G157;
	G8037<= not G405;
	G8038<= not I12360;
	G8046<= not G528;
	G8052<= not G1211;
	G8055<= not G1236;
	G8056<= not G1246;
	G8057<= not G3068;
	G8058<= not G3115;
	G8059<= not G3171;
	G8064<= not G3376;
	G8068<= not G3457;
	G8070<= not G3518;
	G8075<= not G3742;
	G8080<= not G3863;
	G8085<= not I12382;
	G8087<= not G1157;
	G8088<= not G1554;
	G8091<= not G1579;
	G8092<= not G1589;
	G8093<= not G1624;
	G8097<= not G3029;
	G8102<= not G3072;
	G8106<= not G3133;
	G8107<= not G3179;
	G8112<= not G3419;
	G8113<= not G3466;
	G8114<= not G3522;
	G8119<= not G3727;
	G8123<= not G3808;
	G8125<= not G3869;
	G8130<= not G4515;
	G8132<= not I12411;
	G8133<= not G4809;
	G8134<= not I12415;
	G8135<= not I12418;
	G8136<= not G269;
	G8137<= not G411;
	G8138<= not G1500;
	G8139<= not G1648;
	G8146<= not G1760;
	G8150<= not G2185;
	G8154<= not G3139;
	G8155<= not G3380;
	G8160<= not G3423;
	G8164<= not G3484;
	G8165<= not G3530;
	G8170<= not G3770;
	G8171<= not G3817;
	G8172<= not G3873;
	G8178<= not I12437;
	G8179<= not G4999;
	G8180<= not G262;
	G8181<= not G424;
	G8183<= not G482;
	G8186<= not G990;
	G8187<= not G1657;
	G8195<= not G1783;
	G8201<= not G1894;
	G8205<= not G2208;
	G8211<= not G2319;
	G8215<= not I12451;
	G8216<= not G3092;
	G8217<= not G3143;
	G8218<= not G3490;
	G8219<= not G3731;
	G8224<= not G3774;
	G8228<= not G3835;
	G8229<= not G3881;
	G8235<= not I12463;
	G8236<= not G4812;
	G8237<= not G255;
	G8239<= not G1056;
	G8240<= not G1333;
	G8241<= not G1792;
	G8249<= not G1917;
	G8255<= not G2028;
	G8259<= not G2217;
	G8267<= not G2342;
	G8273<= not G2453;
	G8277<= not I12483;
	G8278<= not G3096;
	G8279<= not I12487;
	G8280<= not G3443;
	G8281<= not G3494;
	G8282<= not G3841;
	G8283<= not I12493;
	G8284<= not G5002;
	G8285<= not I12497;
	G8286<= not G53;
	G8287<= not G160;
	G8290<= not G218;
	G8291<= not I12503;
	G8296<= not G246;
	G8297<= not G142;
	G8300<= not G1242;
	G8301<= not G1399;
	G8302<= not G1926;
	G8310<= not G2051;
	G8316<= not G2351;
	G8324<= not G2476;
	G8330<= not G2587;
	G8334<= not G3034;
	G8340<= not G3050;
	G8341<= not G3119;
	G8342<= not I12519;
	G8343<= not G3447;
	G8344<= not I12523;
	G8345<= not G3794;
	G8346<= not G3845;
	G8350<= not G4646;
	G8353<= not I12530;
	G8354<= not G4815;
	G8355<= not I12534;
	G8356<= not G54;
	G8357<= not I12538;
	G8358<= not I12541;
	G8362<= not G194;
	G8363<= not G239;
	G8364<= not G1585;
	G8365<= not G2060;
	G8373<= not G2485;
	G8381<= not G2610;
	G8387<= not G3080;
	G8388<= not G3010;
	G8389<= not G3125;
	G8390<= not G3385;
	G8396<= not G3401;
	G8397<= not G3470;
	G8398<= not I12563;
	G8399<= not G3798;
	G8400<= not G4836;
	G8403<= not I12568;
	G8404<= not G5005;
	G8405<= not I12572;
	G8406<= not G232;
	G8407<= not G1171;
	G8411<= not I12577;
	G8416<= not I12580;
	G8418<= not G2619;
	G8426<= not G3045;
	G8431<= not G3085;
	G8438<= not G3100;
	G8439<= not G3129;
	G8440<= not G3431;
	G8441<= not G3361;
	G8442<= not G3476;
	G8443<= not G3736;
	G8449<= not G3752;
	G8450<= not G3821;
	G8451<= not G4057;
	G8456<= not G56;
	G8457<= not G225;
	G8458<= not G294;
	G8462<= not G1183;
	G8466<= not G1514;
	G8470<= not I12605;
	G8475<= not I12608;
	G8477<= not G3061;
	G8478<= not G3103;
	G8479<= not G3057;
	G8480<= not G3147;
	G8481<= not I12618;
	G8492<= not G3396;
	G8497<= not G3436;
	G8504<= not G3451;
	G8505<= not G3480;
	G8506<= not G3782;
	G8507<= not G3712;
	G8508<= not G3827;
	G8509<= not G4141;
	G8514<= not G4258;
	G8515<= not I12631;
	G8519<= not G287;
	G8522<= not G298;
	G8526<= not G1526;
	G8531<= not G3288;
	G8534<= not G3338;
	G8538<= not G3412;
	G8539<= not G3454;
	G8540<= not G3408;
	G8541<= not G3498;
	G8542<= not I12644;
	G8553<= not G3747;
	G8558<= not G3787;
	G8565<= not G3802;
	G8566<= not G3831;
	G8567<= not G4082;
	G8571<= not G57;
	G8572<= not I12654;
	G8575<= not G291;
	G8579<= not G2771;
	G8584<= not G3639;
	G8587<= not G3689;
	G8591<= not G3763;
	G8592<= not G3805;
	G8593<= not G3759;
	G8594<= not G3849;
	G8595<= not I12666;
	G8606<= not G4653;
	G8607<= not G37;
	G8608<= not G278;
	G8612<= not G2775;
	G8616<= not G2803;
	G8620<= not G3065;
	G8623<= not G3990;
	G8626<= not G4040;
	G8630<= not G4843;
	G8631<= not G283;
	G8635<= not G2783;
	G8639<= not G2807;
	G8644<= not G3352;
	G8647<= not G3416;
	G8650<= not G4664;
	G8651<= not G758;
	G8654<= not G1087;
	G8655<= not G2787;
	G8659<= not G2815;
	G8663<= not G3343;
	G8666<= not G3703;
	G8669<= not G3767;
	G8672<= not G4669;
	G8673<= not G4737;
	G8676<= not G4821;
	G8677<= not G4854;
	G8680<= not G686;
	G8681<= not G763;
	G8685<= not G1430;
	G8686<= not G2819;
	G8696<= not G3347;
	G8697<= not G3694;
	G8700<= not G4054;
	G8703<= not I12709;
	G8712<= not I12712;
	G8713<= not G4826;
	G8714<= not G4859;
	G8715<= not G4927;
	G8718<= not G3333;
	G8719<= not I12719;
	G8725<= not G739;
	G8733<= not G3698;
	G8734<= not G4045;
	G8740<= not I12735;
	G8741<= not G4821;
	G8742<= not G4035;
	G8743<= not G550;
	G8744<= not G691;
	G8745<= not G744;
	G8748<= not G776;
	G8756<= not G4049;
	G8757<= not I12746;
	G8763<= not I12749;
	G8764<= not G4826;
	G8765<= not G3333;
	G8766<= not G572;
	G8770<= not G749;
	G8774<= not G781;
	G8778<= not I12758;
	G8783<= not I12761;
	G8784<= not I12764;
	G8785<= not I12767;
	G8786<= not I12770;
	G8787<= not I12773;
	G8788<= not I12776;
	G8789<= not I12779;
	G8791<= not I12787;
	G8792<= not I12790;
	G8795<= not I12793;
	G8796<= not G4785;
	G8804<= not G4035;
	G8805<= not I12799;
	G8807<= not G79;
	G8808<= not G595;
	G8812<= not I12805;
	G8818<= not I12808;
	G8821<= not I12811;
	G8822<= not G4975;
	G8830<= not G767;
	G8833<= not G794;
	G8836<= not G736;
	G8839<= not I12819;
	G8840<= not G4277;
	G8841<= not I12823;
	G8844<= not I12826;
	G8848<= not G358;
	G8851<= not G590;
	G8854<= not G613;
	G8858<= not G671;
	G8859<= not G772;
	G8870<= not I12837;
	G8872<= not G4258;
	G8876<= not I12855;
	G8879<= not I12858;
	G8880<= not I12861;
	G8883<= not G4709;
	G8890<= not G376;
	G8891<= not G582;
	G8895<= not G599;
	G8898<= not G676;
	G8899<= not G807;
	G8903<= not G1075;
	G8912<= not G4180;
	G8914<= not G4264;
	G8915<= not I12884;
	G8916<= not I12887;
	G8917<= not I12890;
	G8918<= not I12893;
	G8919<= not I12896;
	G8920<= not I12899;
	G8922<= not I12907;
	G8925<= not I12910;
	G8928<= not G4340;
	G8938<= not G4899;
	G8944<= not G370;
	G8945<= not G608;
	G8948<= not G785;
	G8951<= not G554;
	G8954<= not G1079;
	G8955<= not G1418;
	G8964<= not G4269;
	G8971<= not I12927;
	G8974<= not I12930;
	G8977<= not G4349;
	G8989<= not I12935;
	G8990<= not G146;
	G8993<= not G385;
	G8997<= not G577;
	G9000<= not G632;
	G9003<= not G790;
	G9007<= not G1083;
	G9011<= not G1422;
	G9014<= not G3004;
	G9018<= not G4273;
	G9019<= not I12950;
	G9020<= not G4287;
	G9021<= not I12954;
	G9024<= not G4358;
	G9030<= not G4793;
	G9036<= not G5084;
	G9037<= not G164;
	G9040<= not G499;
	G9044<= not G604;
	G9048<= not I12963;
	G9049<= not G640;
	G9050<= not G1087;
	G9051<= not G1426;
	G9056<= not G3017;
	G9060<= not G3355;
	G9064<= not G4983;
	G9070<= not G5428;
	G9071<= not G2831;
	G9072<= not G2994;
	G9073<= not G150;
	G9077<= not G504;
	G9083<= not G626;
	G9086<= not G847;
	G9091<= not G1430;
	G9095<= not G3368;
	G9099<= not G3706;
	G9103<= not G5774;
	G9104<= not I12987;
	G9152<= not G2834;
	G9153<= not I12991;
	G9154<= not I12994;
	G9155<= not I12997;
	G9158<= not G513;
	G9162<= not G622;
	G9166<= not G837;
	G9174<= not G1205;
	G9180<= not G3719;
	G9184<= not G6120;
	G9185<= not I13007;
	G9186<= not I13010;
	G9187<= not G518;
	G9194<= not G827;
	G9197<= not G1221;
	G9200<= not G1548;
	G9206<= not G5164;
	G9212<= not G6466;
	G9213<= not I13020;
	G9214<= not G617;
	G9220<= not G843;
	G9223<= not G1216;
	G9226<= not G1564;
	G9229<= not G5052;
	G9234<= not G5170;
	G9239<= not G5511;
	G9245<= not I13031;
	G9247<= not G1559;
	G9250<= not G1600;
	G9251<= not I13037;
	G9252<= not G4304;
	G9253<= not G5037;
	G9257<= not G5115;
	G9259<= not G5176;
	G9264<= not G5396;
	G9269<= not G5517;
	G9274<= not G5857;
	G9280<= not I13054;
	G9281<= not I13057;
	G9282<= not G723;
	G9283<= not G1736;
	G9284<= not G2161;
	G9285<= not G2715;
	G9291<= not G3021;
	G9298<= not G5080;
	G9299<= not G5124;
	G9300<= not G5180;
	G9305<= not G5381;
	G9309<= not G5462;
	G9311<= not G5523;
	G9316<= not G5742;
	G9321<= not G5863;
	G9326<= not G6203;
	G9332<= not G64;
	G9333<= not G417;
	G9337<= not G1608;
	G9338<= not G1870;
	G9339<= not G2295;
	G9340<= not I13094;
	G9354<= not G2719;
	G9360<= not G3372;
	G9364<= not G5041;
	G9369<= not G5084;
	G9373<= not G5142;
	G9374<= not G5188;
	G9379<= not G5424;
	G9380<= not G5471;
	G9381<= not G5527;
	G9386<= not G5727;
	G9390<= not G5808;
	G9392<= not G5869;
	G9397<= not G6088;
	G9402<= not G6209;
	G9407<= not G6549;
	G9413<= not G1744;
	G9414<= not G2004;
	G9415<= not G2169;
	G9416<= not G2429;
	G9417<= not I13124;
	G9429<= not G3723;
	G9433<= not G5148;
	G9434<= not G5385;
	G9439<= not G5428;
	G9443<= not G5489;
	G9444<= not G5535;
	G9449<= not G5770;
	G9450<= not G5817;
	G9451<= not G5873;
	G9456<= not G6073;
	G9460<= not G6154;
	G9462<= not G6215;
	G9467<= not G6434;
	G9472<= not G6555;
	G9477<= not I13149;
	G9478<= not I13152;
	G9480<= not G559;
	G9484<= not G1612;
	G9488<= not G1878;
	G9489<= not G2303;
	G9490<= not G2563;
	G9491<= not G2729;
	G9492<= not G2759;
	G9496<= not G3303;
	G9497<= not I13166;
	G9498<= not G5101;
	G9499<= not G5152;
	G9500<= not G5495;
	G9501<= not G5731;
	G9506<= not G5774;
	G9510<= not G5835;
	G9511<= not G5881;
	G9516<= not G6116;
	G9517<= not G6163;
	G9518<= not G6219;
	G9523<= not G6419;
	G9527<= not G6500;
	G9529<= not G6561;
	G9534<= not G90;
	G9537<= not G1748;
	G9541<= not G2012;
	G9542<= not G2173;
	G9546<= not G2437;
	G9547<= not G2735;
	G9551<= not G3281;
	G9552<= not G3654;
	G9553<= not I13202;
	G9554<= not G5105;
	G9555<= not I13206;
	G9556<= not G5448;
	G9557<= not G5499;
	G9558<= not G5841;
	G9559<= not G6077;
	G9564<= not G6120;
	G9568<= not G6181;
	G9569<= not G6227;
	G9574<= not G6462;
	G9575<= not G6509;
	G9576<= not G6565;
	G9581<= not G91;
	G9582<= not G703;
	G9585<= not G1616;
	G9590<= not G1882;
	G9594<= not G2307;
	G9598<= not G2571;
	G9599<= not G3310;
	G9600<= not G3632;
	G9601<= not G4005;
	G9607<= not G5046;
	G9613<= not G5062;
	G9614<= not G5128;
	G9615<= not I13236;
	G9616<= not G5452;
	G9617<= not I13240;
	G9618<= not G5794;
	G9619<= not G5845;
	G9620<= not G6187;
	G9621<= not G6423;
	G9626<= not G6466;
	G9630<= not G6527;
	G9631<= not G6573;
	G9636<= not G72;
	G9637<= not I13252;
	G9638<= not G1620;
	G9639<= not G1752;
	G9644<= not G2016;
	G9648<= not G2177;
	G9653<= not G2441;
	G9657<= not G2763;
	G9660<= not G3267;
	G9661<= not G3661;
	G9662<= not G3983;
	G9669<= not G5092;
	G9670<= not G5022;
	G9671<= not G5134;
	G9672<= not G5390;
	G9678<= not G5406;
	G9679<= not G5475;
	G9680<= not I13276;
	G9681<= not G5798;
	G9682<= not I13280;
	G9683<= not G6140;
	G9684<= not G6191;
	G9685<= not G6533;
	G9686<= not G73;
	G9687<= not I13287;
	G9688<= not G113;
	G9689<= not G124;
	G9690<= not G732;
	G9691<= not G1706;
	G9692<= not G1756;
	G9693<= not G1886;
	G9698<= not G2181;
	G9699<= not G2311;
	G9704<= not G2575;
	G9708<= not G2741;
	G9713<= not G3618;
	G9714<= not G4012;
	G9716<= not G5057;
	G9721<= not G5097;
	G9728<= not G5109;
	G9729<= not G5138;
	G9730<= not G5436;
	G9731<= not G5366;
	G9732<= not G5481;
	G9733<= not G5736;
	G9739<= not G5752;
	G9740<= not G5821;
	G9741<= not I13317;
	G9742<= not G6144;
	G9743<= not I13321;
	G9744<= not G6486;
	G9745<= not G6537;
	G9746<= not I13326;
	G9747<= not I13329;
	G9748<= not G114;
	G9749<= not G1691;
	G9751<= not G1710;
	G9752<= not G1840;
	G9753<= not G1890;
	G9754<= not G2020;
	G9759<= not G2265;
	G9760<= not G2315;
	G9761<= not G2445;
	G9766<= not G2748;
	G9771<= not G3969;
	G9772<= not I13352;
	G9776<= not G5073;
	G9777<= not G5112;
	G9778<= not G5069;
	G9779<= not G5156;
	G9780<= not I13360;
	G9792<= not G5401;
	G9797<= not G5441;
	G9804<= not G5456;
	G9805<= not G5485;
	G9806<= not G5782;
	G9807<= not G5712;
	G9808<= not G5827;
	G9809<= not G6082;
	G9815<= not G6098;
	G9816<= not G6167;
	G9817<= not I13374;
	G9818<= not G6490;
	G9819<= not G92;
	G9820<= not G99;
	G9821<= not G115;
	G9822<= not G125;
	G9824<= not G1825;
	G9826<= not G1844;
	G9827<= not G1974;
	G9828<= not G2024;
	G9829<= not G2250;
	G9831<= not G2269;
	G9832<= not G2399;
	G9833<= not G2449;
	G9834<= not G2579;
	G9839<= not G2724;
	G9842<= not G3274;
	G9843<= not G4311;
	G9848<= not G4462;
	G9853<= not G5297;
	G9856<= not G5343;
	G9860<= not G5417;
	G9861<= not G5459;
	G9862<= not G5413;
	G9863<= not G5503;
	G9864<= not I13424;
	G9875<= not G5747;
	G9880<= not G5787;
	G9887<= not G5802;
	G9888<= not G5831;
	G9889<= not G6128;
	G9890<= not G6058;
	G9891<= not G6173;
	G9892<= not G6428;
	G9898<= not G6444;
	G9899<= not G6513;
	G9900<= not G6;
	G9901<= not G84;
	G9902<= not G100;
	G9903<= not G681;
	G9905<= not G802;
	G9907<= not G1959;
	G9909<= not G1978;
	G9910<= not G2108;
	G9911<= not G2384;
	G9913<= not G2403;
	G9914<= not G2533;
	G9915<= not G2583;
	G9916<= not G3625;
	G9917<= not I13473;
	G9920<= not G4322;
	G9924<= not G5644;
	G9927<= not G5689;
	G9931<= not G5763;
	G9932<= not G5805;
	G9933<= not G5759;
	G9934<= not G5849;
	G9935<= not I13483;
	G9946<= not G6093;
	G9951<= not G6133;
	G9958<= not G6148;
	G9959<= not G6177;
	G9960<= not G6474;
	G9961<= not G6404;
	G9962<= not G6519;
	G9963<= not G7;
	G9964<= not G126;
	G9965<= not G127;
	G9969<= not G1682;
	G9970<= not G1714;
	G9971<= not G2093;
	G9973<= not G2112;
	G9974<= not G2518;
	G9976<= not G2537;
	G9977<= not G2667;
	G9978<= not G2756;
	G9982<= not G3976;
	G9983<= not G4239;
	G9985<= not G4332;
	G9989<= not G5077;
	G9992<= not G5990;
	G9995<= not G6035;
	G9999<= not G6109;
	G10000<= not G6151;
	G10001<= not G6105;
	G10002<= not G6195;
	G10003<= not I13539;
	G10014<= not G6439;
	G10019<= not G6479;
	G10026<= not G6494;
	G10027<= not G6523;
	G10028<= not G8;
	G10029<= not I13548;
	G10030<= not G116;
	G10031<= not I13552;
	G10032<= not G562;
	G10033<= not G655;
	G10035<= not G1720;
	G10036<= not G1816;
	G10037<= not G1848;
	G10038<= not G2241;
	G10039<= not G2273;
	G10040<= not G2652;
	G10042<= not G2671;
	G10043<= not G1632;
	G10044<= not G5357;
	G10047<= not G5421;
	G10050<= not G6336;
	G10053<= not G6381;
	G10057<= not G6455;
	G10058<= not G6497;
	G10059<= not G6451;
	G10060<= not G6541;
	G10061<= not I13581;
	G10072<= not G9;
	G10073<= not G134;
	G10074<= not G718;
	G10077<= not G1724;
	G10078<= not G1854;
	G10079<= not G1950;
	G10080<= not G1982;
	G10081<= not G2279;
	G10082<= not G2375;
	G10083<= not G2407;
	G10084<= not G2837;
	G10085<= not G1768;
	G10086<= not G2193;
	G10087<= not I13597;
	G10090<= not G5348;
	G10093<= not G5703;
	G10096<= not G5767;
	G10099<= not G6682;
	G10102<= not G6727;
	G10106<= not G16;
	G10107<= not I13606;
	G10108<= not G120;
	G10109<= not G135;
	G10110<= not G661;
	G10111<= not G1858;
	G10112<= not G1988;
	G10113<= not G2084;
	G10114<= not G2116;
	G10115<= not G2283;
	G10116<= not G2413;
	G10117<= not G2509;
	G10118<= not G2541;
	G10119<= not G2841;
	G10120<= not G1902;
	G10121<= not G2327;
	G10122<= not I13623;
	G10129<= not G5352;
	G10130<= not G5694;
	G10133<= not G6049;
	G10136<= not G6113;
	G10139<= not G136;
	G10140<= not G19;
	G10141<= not I13634;
	G10142<= not I13637;
	G10143<= not G568;
	G10147<= not G728;
	G10150<= not G1700;
	G10151<= not G1992;
	G10152<= not G2122;
	G10153<= not G2417;
	G10154<= not G2547;
	G10155<= not G2643;
	G10156<= not G2675;
	G10157<= not G2036;
	G10158<= not G2461;
	G10159<= not G4477;
	G10165<= not G5698;
	G10166<= not G6040;
	G10169<= not G6395;
	G10172<= not G6459;
	G10175<= not G28;
	G10176<= not G44;
	G10177<= not G1834;
	G10178<= not G2126;
	G10180<= not G2259;
	G10181<= not G2551;
	G10182<= not G2681;
	G10183<= not G2595;
	G10184<= not G4486;
	G10190<= not G6044;
	G10191<= not G6386;
	G10194<= not G6741;
	G10197<= not G31;
	G10198<= not I13672;
	G10199<= not G1968;
	G10200<= not G2138;
	G10203<= not G2393;
	G10204<= not G2685;
	G10206<= not G4489;
	G10212<= not G6390;
	G10213<= not G6732;
	G10216<= not I13684;
	G10217<= not G2102;
	G10218<= not G2527;
	G10219<= not G2697;
	G10222<= not G4492;
	G10223<= not G4561;
	G10229<= not G6736;
	G10230<= not I13694;
	G10231<= not G2661;
	G10232<= not G4527;
	G10233<= not I13699;
	G10261<= not G4555;
	G10262<= not G586;
	G10272<= not I13705;
	G10273<= not I13708;
	G10274<= not G976;
	G10275<= not G4584;
	G10278<= not G4628;
	G10287<= not I13715;
	G10288<= not I13718;
	G10289<= not G1319;
	G10295<= not I13723;
	G10306<= not I13726;
	G10308<= not G4459;
	G10311<= not G4633;
	G10319<= not I13740;
	G10320<= not G817;
	G10323<= not I13744;
	G10334<= not G4420;
	G10335<= not G4483;
	G10337<= not G5016;
	G10347<= not I13759;
	G10348<= not I13762;
	G10349<= not G6956;
	G10350<= not G6800;
	G10351<= not G6802;
	G10352<= not G6804;
	G10353<= not G6803;
	G10354<= not G6811;
	G10355<= not G6816;
	G10356<= not G6819;
	G10357<= not G6825;
	G10358<= not G6827;
	G10359<= not G6830;
	G10360<= not G6836;
	G10361<= not G6841;
	G10362<= not G6850;
	G10363<= not I13779;
	G10364<= not G6869;
	G10365<= not G6867;
	G10366<= not G6895;
	G10367<= not G6870;
	G10368<= not G6887;
	G10369<= not G6873;
	G10370<= not G7095;
	G10371<= not G6918;
	G10372<= not G6900;
	G10373<= not G6917;
	G10374<= not G6903;
	G10375<= not G6941;
	G10376<= not G6923;
	G10377<= not G6940;
	G10378<= not G6926;
	G10379<= not G6953;
	G10380<= not G6960;
	G10381<= not G6957;
	G10382<= not G6958;
	G10383<= not G6978;
	G10384<= not I13802;
	G10385<= not I13805;
	G10386<= not G6982;
	G10387<= not G6996;
	G10388<= not G6983;
	G10389<= not G6986;
	G10390<= not G6987;
	G10391<= not G6988;
	G10392<= not G6989;
	G10393<= not G6991;
	G10394<= not G6994;
	G10395<= not G6995;
	G10396<= not G6997;
	G10397<= not G7018;
	G10398<= not G6999;
	G10399<= not G7017;
	G10400<= not G7002;
	G10401<= not G7041;
	G10402<= not G7023;
	G10403<= not G7040;
	G10404<= not G7026;
	G10405<= not G7064;
	G10406<= not G7046;
	G10407<= not G7063;
	G10408<= not G7049;
	G10409<= not G7087;
	G10410<= not G7069;
	G10411<= not G7086;
	G10412<= not G7072;
	G10413<= not G7110;
	G10414<= not G7092;
	G10415<= not G7109;
	G10416<= not G10318;
	G10417<= not G7117;
	G10418<= not G8818;
	G10419<= not G8821;
	G10420<= not G9239;
	G10427<= not G10053;
	G10428<= not G9631;
	G10429<= not G7148;
	G10430<= not I13847;
	G10473<= not I13857;
	G10474<= not G8841;
	G10475<= not G8844;
	G10487<= not G10233;
	G10489<= not G9259;
	G10490<= not G9274;
	G10497<= not G10102;
	G10498<= not G7161;
	G10499<= not I13872;
	G10500<= not I13875;
	G10502<= not G8876;
	G10503<= not G8879;
	G10504<= not G8763;
	G10509<= not G10233;
	G10518<= not G9311;
	G10519<= not G9326;
	G10521<= not I13889;
	G10527<= not I13892;
	G10530<= not G8922;
	G10531<= not G8925;
	G10532<= not G10233;
	G10533<= not G8795;
	G10540<= not G9392;
	G10541<= not G9407;
	G10542<= not G7196;
	G10544<= not I13906;
	G10553<= not G8971;
	G10554<= not G8974;
	G10564<= not G9462;
	G10570<= not G9021;
	G10571<= not G10233;
	G10572<= not G10233;
	G10581<= not G9529;
	G10582<= not G7116;
	G10597<= not G10233;
	G10606<= not G10233;
	G10607<= not G10233;
	G10608<= not G9155;
	G10612<= not G10233;
	G10613<= not G10233;
	G10620<= not G10233;
	G10621<= not G7567;
	G10627<= not I13968;
	G10652<= not G7601;
	G10658<= not I13979;
	G10664<= not G8928;
	G10678<= not I13990;
	G10685<= not I13995;
	G10708<= not G7836;
	G10710<= not I14006;
	G10725<= not G7846;
	G10727<= not I14016;
	G10741<= not G8411;
	G10761<= not G8411;
	G10762<= not G8470;
	G10776<= not I14033;
	G10794<= not G8470;
	G10795<= not G7202;
	G10804<= not G9772;
	G10805<= not I14046;
	G10812<= not I14050;
	G10815<= not G9917;
	G10816<= not I14054;
	G10830<= not G10087;
	G10851<= not I14069;
	G10857<= not G8712;
	G10872<= not G7567;
	G10877<= not I14079;
	G10881<= not G7567;
	G10882<= not G7601;
	G10897<= not G7601;
	G10960<= not G9007;
	G10980<= not G9051;
	G10981<= not I14119;
	G11011<= not G10274;
	G11017<= not G10289;
	G11026<= not G8434;
	G11030<= not G8292;
	G11031<= not G8609;
	G11033<= not G8500;
	G11034<= not G7611;
	G11038<= not G8632;
	G11042<= not G8691;
	G11043<= not G8561;
	G11048<= not I14158;
	G11110<= not G8728;
	G11122<= not G8751;
	G11128<= not G7993;
	G11129<= not G7994;
	G11136<= not I14192;
	G11143<= not G8032;
	G11147<= not G8417;
	G11164<= not G8085;
	G11165<= not I14222;
	G11170<= not G8476;
	G11181<= not G8134;
	G11182<= not I14241;
	G11183<= not G8135;
	G11192<= not G8038;
	G11202<= not I14267;
	G11204<= not I14271;
	G11214<= not G9602;
	G11215<= not G8285;
	G11233<= not G9664;
	G11234<= not G8355;
	G11235<= not I14301;
	G11236<= not G8357;
	G11237<= not I14305;
	G11249<= not G8405;
	G11250<= not G7502;
	G11268<= not G7515;
	G11269<= not G7516;
	G11290<= not I14326;
	G11291<= not G7526;
	G11293<= not G7527;
	G11294<= not G7598;
	G11316<= not G8967;
	G11317<= not I14346;
	G11324<= not G7542;
	G11325<= not G7543;
	G11336<= not G7620;
	G11344<= not G9015;
	G11349<= not I14365;
	G11367<= not I14381;
	G11371<= not G7565;
	G11373<= not G7566;
	G11383<= not G9061;
	G11388<= not I14395;
	G11398<= not I14409;
	G11401<= not G7593;
	G11402<= not G7594;
	G11403<= not G7595;
	G11404<= not G7596;
	G11413<= not G9100;
	G11418<= not I14424;
	G11425<= not G7640;
	G11428<= not G7615;
	G11429<= not G7616;
	G11430<= not G7617;
	G11431<= not G7618;
	G11447<= not I14450;
	G11450<= not I14455;
	G11467<= not G7623;
	G11468<= not G7624;
	G11470<= not G7625;
	G11471<= not G7626;
	G11472<= not G7918;
	G11498<= not I14475;
	G11509<= not G7632;
	G11510<= not G7633;
	G11512<= not G7634;
	G11513<= not G7948;
	G11519<= not G8481;
	G11547<= not I14505;
	G11560<= not G7647;
	G11562<= not G7648;
	G11576<= not G8542;
	G11592<= not I14537;
	G11608<= not G7659;
	G11609<= not G7660;
	G11615<= not G6875;
	G11631<= not G8595;
	G11640<= not I14550;
	G11652<= not G7674;
	G11663<= not G6905;
	G11677<= not G7689;
	G11678<= not I14563;
	G11686<= not I14567;
	G11691<= not I14570;
	G11702<= not G6928;
	G11705<= not I14576;
	G11706<= not I14579;
	G11709<= not I14584;
	G11714<= not G8107;
	G11720<= not I14589;
	G11721<= not G10074;
	G11724<= not I14593;
	G11735<= not G8534;
	G11736<= not G8165;
	G11741<= not G10033;
	G11744<= not I14602;
	G11753<= not G8587;
	G11754<= not G8229;
	G11762<= not G7964;
	G11769<= not G8626;
	G11770<= not I14619;
	G11772<= not I14623;
	G11779<= not G9602;
	G11786<= not G7549;
	G11790<= not I14630;
	G11793<= not I14633;
	G11796<= not G7985;
	G11810<= not G9664;
	G11811<= not G9724;
	G11812<= not G7567;
	G11815<= not G7582;
	G11819<= not G7717;
	G11820<= not I14644;
	G11823<= not I14647;
	G11826<= not I14650;
	G11829<= not I14653;
	G11832<= not G8011;
	G11833<= not G8026;
	G11841<= not G9800;
	G11842<= not I14660;
	G11845<= not I14663;
	G11849<= not G7601;
	G11852<= not I14668;
	G11855<= not I14671;
	G11861<= not G8070;
	G11865<= not G10124;
	G11866<= not G9883;
	G11867<= not I14679;
	G11868<= not G9185;
	G11872<= not I14684;
	G11875<= not I14687;
	G11878<= not I14690;
	G11884<= not G8125;
	G11888<= not G10160;
	G11889<= not G9954;
	G11894<= not I14702;
	G11897<= not I14705;
	G11900<= not I14708;
	G11910<= not G10185;
	G11911<= not G10022;
	G11912<= not G8989;
	G11917<= not I14727;
	G11920<= not I14730;
	G11927<= not G10207;
	G11928<= not I14742;
	G11929<= not I14745;
	G11930<= not G9281;
	G11931<= not I14749;
	G11941<= not I14761;
	G11948<= not G10224;
	G11949<= not I14773;
	G11963<= not G9153;
	G11964<= not G9154;
	G11965<= not I14797;
	G11966<= not I14800;
	G11981<= not I14823;
	G11984<= not G9186;
	G11985<= not I14827;
	G11986<= not I14830;
	G11987<= not I14833;
	G11988<= not I14836;
	G11989<= not I14839;
	G11991<= not G9485;
	G12009<= not I14862;
	G12012<= not G9213;
	G12013<= not I14866;
	G12018<= not G9538;
	G12021<= not G9543;
	G12036<= not G9245;
	G12037<= not I14893;
	G12038<= not I14896;
	G12039<= not I14899;
	G12040<= not I14902;
	G12041<= not I14905;
	G12047<= not G9591;
	G12051<= not G9595;
	G12054<= not G7690;
	G12074<= not I14932;
	G12075<= not I14935;
	G12076<= not G9280;
	G12077<= not I14939;
	G12082<= not G9645;
	G12086<= not G9654;
	G12088<= not G7701;
	G12107<= not G9687;
	G12108<= not I14964;
	G12109<= not I14967;
	G12110<= not I14970;
	G12122<= not G9705;
	G12143<= not I14999;
	G12180<= not G9477;
	G12181<= not G9478;
	G12182<= not I15030;
	G12183<= not I15033;
	G12184<= not I15036;
	G12217<= not I15070;
	G12218<= not I15073;
	G12233<= not G10338;
	G12238<= not I15102;
	G12295<= not G7139;
	G12300<= not I15144;
	G12321<= not G9637;
	G12322<= not I15162;
	G12337<= not G9340;
	G12345<= not G7158;
	G12350<= not I15190;
	G12367<= not I15205;
	G12368<= not I15208;
	G12378<= not G9417;
	G12381<= not I15223;
	G12399<= not G9920;
	G12417<= not G7175;
	G12422<= not I15238;
	G12430<= not I15250;
	G12440<= not G9985;
	G12465<= not G7192;
	G12470<= not I15284;
	G12477<= not I15295;
	G12487<= not G9340;
	G12490<= not I15316;
	G12497<= not G9780;
	G12543<= not G9417;
	G12546<= not G8740;
	G12563<= not G9864;
	G12598<= not G7004;
	G12614<= not G9935;
	G12640<= not I15382;
	G12656<= not G7028;
	G12672<= not G10003;
	G12705<= not G7051;
	G12721<= not G10061;
	G12738<= not G9374;
	G12749<= not G7074;
	G12760<= not G10272;
	G12778<= not G9856;
	G12779<= not G9444;
	G12790<= not G7097;
	G12793<= not G10287;
	G12804<= not G9927;
	G12805<= not G9511;
	G12811<= not G10319;
	G12818<= not G8792;
	G12820<= not G10233;
	G12823<= not G9206;
	G12830<= not G9995;
	G12831<= not G9569;
	G12833<= not I15448;
	G12834<= not G10349;
	G12835<= not G10352;
	G12836<= not G10351;
	G12837<= not G10354;
	G12838<= not G10353;
	G12839<= not G10350;
	G12840<= not G10356;
	G12841<= not G10357;
	G12842<= not G10355;
	G12843<= not G10359;
	G12844<= not G10360;
	G12845<= not G10358;
	G12857<= not I15474;
	G12859<= not G10366;
	G12860<= not G10368;
	G12861<= not G10367;
	G12862<= not G10370;
	G12863<= not G10371;
	G12864<= not G10373;
	G12865<= not G10372;
	G12866<= not G10369;
	G12867<= not G10375;
	G12868<= not G10377;
	G12869<= not G10376;
	G12870<= not G10374;
	G12871<= not G10378;
	G12872<= not G10379;
	G12873<= not G10380;
	G12874<= not G10383;
	G12875<= not I15494;
	G12878<= not G10386;
	G12879<= not G10381;
	G12880<= not G10387;
	G12881<= not G10388;
	G12882<= not G10389;
	G12883<= not G10390;
	G12884<= not G10392;
	G12885<= not G10382;
	G12886<= not G10393;
	G12887<= not G10394;
	G12888<= not G10395;
	G12889<= not G10396;
	G12890<= not G10397;
	G12891<= not G10399;
	G12892<= not G10398;
	G12893<= not G10391;
	G12894<= not G10401;
	G12895<= not G10403;
	G12896<= not G10402;
	G12897<= not G10400;
	G12898<= not G10405;
	G12899<= not G10407;
	G12900<= not G10406;
	G12901<= not G10404;
	G12902<= not G10409;
	G12903<= not G10411;
	G12904<= not G10410;
	G12905<= not G10408;
	G12906<= not G10413;
	G12907<= not G10415;
	G12908<= not G10414;
	G12909<= not G10412;
	G12914<= not G12235;
	G12918<= not I15533;
	G12919<= not I15536;
	G12921<= not G12228;
	G12922<= not G12297;
	G12923<= not I15542;
	G12929<= not G12550;
	G12930<= not G12347;
	G12932<= not I15550;
	G12936<= not G12601;
	G12937<= not G12419;
	G12938<= not I15556;
	G12940<= not G11744;
	G12944<= not G12659;
	G12945<= not G12467;
	G12946<= not I15564;
	G12950<= not G12708;
	G12951<= not I15569;
	G12952<= not I15572;
	G12955<= not I15577;
	G12967<= not G11790;
	G12968<= not G11793;
	G12975<= not G12752;
	G12976<= not I15587;
	G12977<= not I15590;
	G12978<= not I15593;
	G12983<= not I15600;
	G12995<= not G11820;
	G12996<= not G11823;
	G12997<= not G11826;
	G12998<= not G11829;
	G13003<= not I15609;
	G13007<= not G11852;
	G13008<= not G11855;
	G13009<= not I15617;
	G13010<= not I15620;
	G13011<= not I15623;
	G13012<= not I15626;
	G13014<= not G11872;
	G13015<= not G11875;
	G13016<= not G11878;
	G13017<= not I15633;
	G13018<= not I15636;
	G13022<= not G11894;
	G13023<= not G11897;
	G13024<= not G11900;
	G13026<= not G11018;
	G13027<= not I15647;
	G13028<= not I15650;
	G13033<= not G11917;
	G13034<= not G11920;
	G13036<= not G10981;
	G13037<= not G10981;
	G13039<= not I15663;
	G13041<= not I15667;
	G13045<= not G11941;
	G13049<= not I15677;
	G13051<= not G11964;
	G13055<= not I15682;
	G13061<= not G10981;
	G13062<= not G10981;
	G13064<= not G11705;
	G13065<= not G10476;
	G13068<= not I15697;
	G13070<= not G11984;
	G13074<= not I15702;
	G13075<= not I15705;
	G13082<= not G10981;
	G13085<= not I15717;
	G13087<= not G12012;
	G13096<= not I15727;
	G13099<= not I15732;
	G13101<= not I15736;
	G13103<= not G10905;
	G13106<= not G10981;
	G13107<= not G10476;
	G13116<= not G10935;
	G13117<= not G10981;
	G13120<= not G10632;
	G13132<= not G10632;
	G13133<= not G11330;
	G13138<= not I15765;
	G13140<= not G10632;
	G13141<= not G11374;
	G13142<= not G10632;
	G13144<= not I15773;
	G13173<= not G10632;
	G13174<= not G10741;
	G13175<= not G10909;
	G13177<= not I15782;
	G13188<= not G10909;
	G13189<= not G10762;
	G13190<= not G10939;
	G13191<= not I15788;
	G13209<= not G10632;
	G13215<= not G10909;
	G13216<= not G10939;
	G13222<= not G10590;
	G13223<= not I15800;
	G13239<= not G10632;
	G13246<= not G10939;
	G13249<= not G10590;
	G13250<= not I15811;
	G13251<= not I15814;
	G13255<= not G10632;
	G13258<= not I15821;
	G13259<= not I15824;
	G13267<= not I15831;
	G13271<= not I15834;
	G13272<= not I15837;
	G13278<= not G10738;
	G13279<= not I15843;
	G13280<= not I15846;
	G13297<= not G10831;
	G13298<= not I15862;
	G13301<= not G10862;
	G13302<= not G12321;
	G13303<= not I15869;
	G13304<= not I15872;
	G13305<= not G11048;
	G13311<= not I15878;
	G13312<= not G11048;
	G13314<= not G10893;
	G13322<= not G10918;
	G13323<= not G11048;
	G13329<= not I15893;
	G13334<= not G11048;
	G13350<= not I15906;
	G13394<= not I15915;
	G13409<= not I15918;
	G13410<= not I15921;
	G13412<= not G11963;
	G13413<= not G11737;
	G13414<= not G11048;
	G13416<= not I15929;
	G13431<= not I15932;
	G13437<= not I15937;
	G13458<= not G11048;
	G13460<= not I15942;
	G13463<= not G10476;
	G13474<= not G11048;
	G13477<= not I15954;
	G13483<= not G11270;
	G13484<= not G10981;
	G13485<= not G10476;
	G13494<= not G11912;
	G13504<= not G11303;
	G13505<= not G10981;
	G13506<= not G10808;
	G13510<= not I15981;
	G13514<= not I15987;
	G13521<= not G11357;
	G13522<= not G10981;
	G13530<= not G12641;
	G13545<= not I16010;
	G13555<= not G12692;
	G13565<= not G11006;
	G13569<= not G10951;
	G13574<= not I16024;
	G13583<= not I16028;
	G13584<= not G12735;
	G13593<= not G10556;
	G13594<= not G11012;
	G13595<= not G10951;
	G13596<= not G10971;
	G13605<= not I16040;
	G13620<= not G10556;
	G13621<= not G10573;
	G13624<= not G10951;
	G13625<= not G10971;
	G13626<= not G11273;
	G13637<= not G10556;
	G13638<= not I16057;
	G13655<= not G10573;
	G13663<= not G10971;
	G13664<= not G11252;
	G13665<= not G11306;
	G13675<= not G10556;
	G13679<= not G10573;
	G13680<= not I16077;
	G13706<= not G11280;
	G13707<= not G11360;
	G13715<= not G10573;
	G13716<= not I16090;
	G13729<= not G10951;
	G13736<= not G11313;
	G13745<= not I16102;
	G13763<= not G10971;
	G13782<= not I16117;
	G13793<= not I16120;
	G13809<= not I16135;
	G13835<= not I16150;
	G13856<= not I16160;
	G13857<= not I16163;
	G13865<= not I16168;
	G13868<= not G11493;
	G13869<= not G10831;
	G13876<= not G11432;
	G13877<= not G11350;
	G13881<= not I16181;
	G13885<= not G10862;
	G13895<= not I16193;
	G13901<= not G11480;
	G13902<= not G11389;
	G13906<= not I16201;
	G13926<= not I16217;
	G13932<= not G11534;
	G13933<= not G11419;
	G13943<= not I16231;
	G13966<= not I16246;
	G13975<= not G11048;
	G13976<= not G11130;
	G13995<= not G11261;
	G13999<= not G11048;
	G14004<= not G11149;
	G14029<= not G11283;
	G14031<= not I16289;
	G14032<= not G11048;
	G14034<= not G11048;
	G14063<= not G11048;
	G14065<= not G11048;
	G14095<= not G11326;
	G14096<= not I16328;
	G14125<= not I16345;
	G14147<= not I16357;
	G14149<= not G12381;
	G14150<= not G12381;
	G14166<= not G11048;
	G14167<= not I16371;
	G14169<= not G12381;
	G14173<= not G12076;
	G14179<= not G11048;
	G14183<= not G12381;
	G14184<= not G12381;
	G14186<= not G11346;
	G14189<= not I16391;
	G14191<= not G12381;
	G14192<= not G11385;
	G14197<= not G12160;
	G14198<= not G12180;
	G14201<= not I16401;
	G14203<= not G12381;
	G14204<= not G12155;
	G14205<= not G12381;
	G14208<= not G11563;
	G14209<= not G11415;
	G14215<= not G12198;
	G14217<= not I16417;
	G14219<= not G12381;
	G14226<= not G11618;
	G14231<= not G12246;
	G14232<= not G11083;
	G14237<= not G11666;
	G14238<= not G10823;
	G14251<= not G12308;
	G14252<= not I16438;
	G14255<= not G12381;
	G14262<= not G10838;
	G14275<= not G12358;
	G14276<= not I16452;
	G14277<= not I16455;
	G14290<= not I16460;
	G14297<= not G10869;
	G14307<= not I16468;
	G14308<= not I16471;
	G14314<= not I16476;
	G14315<= not I16479;
	G14321<= not G10874;
	G14330<= not I16486;
	G14331<= not I16489;
	G14332<= not I16492;
	G14336<= not I16498;
	G14338<= not I16502;
	G14342<= not G12163;
	G14348<= not G10887;
	G14357<= not G12181;
	G14358<= not I16512;
	G14359<= not I16515;
	G14363<= not I16521;
	G14366<= not I16526;
	G14376<= not G12126;
	G14377<= not G12201;
	G14383<= not I16535;
	G14384<= not I16538;
	G14385<= not I16541;
	G14386<= not I16544;
	G14398<= not I16555;
	G14405<= not G12170;
	G14406<= not G12249;
	G14412<= not I16564;
	G14421<= not I16575;
	G14423<= not I16579;
	G14424<= not G11136;
	G14431<= not G12208;
	G14432<= not G12311;
	G14441<= not I16590;
	G14442<= not I16593;
	G14443<= not I16596;
	G14451<= not I16606;
	G14453<= not I16610;
	G14454<= not I16613;
	G14503<= not G12256;
	G14504<= not G12361;
	G14509<= not I16626;
	G14510<= not I16629;
	G14518<= not I16639;
	G14535<= not G12318;
	G14536<= not I16651;
	G14541<= not G11405;
	G14543<= not I16660;
	G14544<= not I16663;
	G14545<= not G12768;
	G14562<= not G12036;
	G14563<= not I16676;
	G14564<= not I16679;
	G14571<= not I16688;
	G14582<= not I16698;
	G14584<= not G11048;
	G14591<= not I16709;
	G14597<= not I16713;
	G14609<= not I16724;
	G14616<= not I16733;
	G14630<= not G12402;
	G14631<= not G12239;
	G14635<= not I16741;
	G14639<= not I16747;
	G14645<= not I16755;
	G14662<= not I16762;
	G14668<= not G12450;
	G14669<= not G12301;
	G14673<= not I16770;
	G14676<= not I16775;
	G14694<= not I16795;
	G14700<= not G12512;
	G14701<= not G12351;
	G14705<= not I16803;
	G14714<= not G11405;
	G14738<= not I16821;
	G14744<= not G12578;
	G14745<= not G12423;
	G14749<= not I16829;
	G14753<= not G11317;
	G14779<= not I16847;
	G14785<= not G12629;
	G14786<= not G12471;
	G14790<= not I16855;
	G14828<= not I16875;
	G14833<= not G11405;
	G14873<= not I16898;
	G14912<= not I16917;
	G15048<= not I16969;
	G15085<= not I17008;
	G15169<= not I17094;
	G15171<= not I17098;
	G15224<= not I17101;
	G15277<= not I17104;
	G15344<= not G14851;
	G15345<= not I17108;
	G15348<= not I17111;
	G15371<= not I17114;
	G15373<= not I17118;
	G15426<= not I17121;
	G15479<= not G14895;
	G15480<= not I17125;
	G15483<= not I17128;
	G15506<= not I17131;
	G15509<= not I17136;
	G15562<= not G14943;
	G15563<= not I17140;
	G15566<= not I17143;
	G15568<= not G14984;
	G15569<= not I17148;
	G15571<= not G13211;
	G15573<= not I17154;
	G15579<= not I17159;
	G15580<= not G13242;
	G15588<= not I17166;
	G15595<= not I17173;
	G15614<= not G14914;
	G15615<= not I17181;
	G15634<= not I17188;
	G15655<= not G13202;
	G15656<= not I17198;
	G15680<= not I17207;
	G15705<= not G13217;
	G15714<= not I17228;
	G15731<= not G13326;
	G15733<= not I17249;
	G15739<= not G13284;
	G15740<= not G13342;
	G15746<= not G13121;
	G15747<= not G13307;
	G15750<= not G13291;
	G15755<= not G13134;
	G15756<= not G13315;
	G15758<= not I17276;
	G15799<= not G13110;
	G15806<= not I17302;
	G15811<= not G13125;
	G15816<= not I17314;
	G15824<= not I17324;
	G15830<= not G13432;
	G15831<= not G13385;
	G15842<= not G13469;
	G15862<= not I17355;
	G15885<= not I17374;
	G15915<= not I17392;
	G15932<= not I17395;
	G15938<= not I17401;
	G15969<= not I17416;
	G15979<= not I17420;
	G16000<= not I17425;
	G16030<= not G13570;
	G16031<= not I17436;
	G16053<= not I17442;
	G16075<= not G13597;
	G16077<= not I17456;
	G16096<= not G13530;
	G16099<= not G13437;
	G16100<= not I17471;
	G16123<= not G13530;
	G16124<= not G13555;
	G16127<= not G13437;
	G16129<= not I17488;
	G16136<= not I17491;
	G16158<= not G13555;
	G16159<= not G13584;
	G16162<= not G13437;
	G16164<= not I17507;
	G16171<= not G13530;
	G16172<= not G13584;
	G16180<= not G13437;
	G16182<= not G13846;
	G16186<= not G13555;
	G16195<= not G13437;
	G16197<= not G13861;
	G16200<= not G13584;
	G16206<= not G13437;
	G16214<= not G13437;
	G16216<= not I17557;
	G16223<= not G13437;
	G16228<= not I17569;
	G16235<= not G13437;
	G16249<= not I17590;
	G16280<= not G13330;
	G16284<= not I17609;
	G16285<= not I17612;
	G16286<= not I17615;
	G16289<= not G13223;
	G16290<= not G13260;
	G16300<= not I17626;
	G16305<= not G13346;
	G16307<= not I17633;
	G16308<= not I17636;
	G16309<= not I17639;
	G16310<= not G13223;
	G16311<= not G13273;
	G16320<= not G14454;
	G16322<= not I17650;
	G16323<= not I17653;
	G16325<= not G13223;
	G16326<= not I17658;
	G16349<= not I17661;
	G16423<= not G14066;
	G16428<= not I17668;
	G16429<= not I17671;
	G16431<= not I17675;
	G16449<= not I17679;
	G16472<= not G14098;
	G16473<= not G13977;
	G16475<= not G14107;
	G16482<= not G13464;
	G16487<= not I17695;
	G16489<= not I17699;
	G16508<= not I17704;
	G16509<= not G13873;
	G16510<= not G14008;
	G16511<= not G14130;
	G16512<= not G14015;
	G16514<= not G14139;
	G16515<= not G13486;
	G16521<= not G13543;
	G16522<= not G13889;
	G16523<= not G14041;
	G16525<= not I17723;
	G16526<= not G13898;
	G16527<= not G14048;
	G16528<= not G14154;
	G16529<= not G14055;
	G16530<= not G14454;
	G16533<= not I17733;
	G16540<= not I17744;
	G16577<= not I17747;
	G16578<= not I17750;
	G16579<= not G13267;
	G16580<= not I17754;
	G16582<= not G13915;
	G16583<= not G14069;
	G16584<= not G13920;
	G16585<= not G14075;
	G16587<= not I17763;
	G16588<= not G13929;
	G16589<= not G14082;
	G16594<= not I17772;
	G16600<= not I17780;
	G16601<= not I17783;
	G16602<= not G14101;
	G16603<= not I17787;
	G16605<= not G13955;
	G16606<= not G14110;
	G16607<= not G13960;
	G16608<= not G14116;
	G16609<= not G14454;
	G16615<= not I17801;
	G16620<= not I17808;
	G16622<= not G14104;
	G16623<= not G14127;
	G16624<= not I17814;
	G16626<= not G14133;
	G16627<= not I17819;
	G16629<= not G13990;
	G16630<= not G14142;
	G16631<= not G14454;
	G16632<= not G14454;
	G16640<= not I17834;
	G16643<= not I17839;
	G16644<= not I17842;
	G16645<= not G13756;
	G16651<= not G14005;
	G16652<= not G13892;
	G16654<= not G14136;
	G16655<= not G14151;
	G16656<= not I17852;
	G16658<= not G14157;
	G16659<= not I17857;
	G16661<= not G14454;
	G16675<= not I17873;
	G16676<= not I17876;
	G16677<= not I17879;
	G16680<= not G13223;
	G16684<= not G14223;
	G16685<= not G14038;
	G16686<= not I17892;
	G16688<= not G14045;
	G16689<= not G13923;
	G16691<= not G14160;
	G16692<= not G14170;
	G16693<= not I17901;
	G16695<= not G14454;
	G16708<= not I17916;
	G16709<= not I17919;
	G16712<= not G13223;
	G16716<= not G13948;
	G16717<= not G13951;
	G16718<= not I17932;
	G16720<= not G14234;
	G16721<= not G14072;
	G16722<= not I17938;
	G16724<= not G14079;
	G16725<= not G13963;
	G16726<= not G14454;
	G16727<= not G14454;
	G16738<= not I17956;
	G16739<= not G13223;
	G16740<= not G13980;
	G16742<= not G13983;
	G16743<= not G13986;
	G16744<= not I17964;
	G16746<= not G14258;
	G16747<= not G14113;
	G16748<= not I17970;
	G16750<= not G14454;
	G16752<= not I17976;
	G16767<= not I17989;
	G16768<= not G13223;
	G16769<= not G13530;
	G16771<= not G14018;
	G16773<= not G14021;
	G16774<= not G14024;
	G16775<= not I17999;
	G16777<= not I18003;
	G16782<= not I18006;
	G16795<= not I18009;
	G16809<= not G14387;
	G16812<= not G13555;
	G16814<= not G14058;
	G16816<= not I18028;
	G16821<= not I18031;
	G16826<= not I18034;
	G16853<= not G13584;
	G16856<= not I18048;
	G16861<= not I18051;
	G16872<= not I18060;
	G16873<= not I18063;
	G16874<= not I18066;
	G16877<= not I18071;
	G16886<= not I18078;
	G16897<= not I18083;
	G16920<= not I18086;
	G16923<= not I18089;
	G16924<= not I18092;
	G16931<= not I18101;
	G16954<= not I18104;
	G16955<= not I18107;
	G16958<= not G14238;
	G16960<= not I18114;
	G16963<= not I18117;
	G16964<= not I18120;
	G16966<= not G14291;
	G16967<= not I18125;
	G16968<= not G14238;
	G16969<= not G14262;
	G16971<= not I18131;
	G16987<= not I18135;
	G17010<= not I18138;
	G17013<= not G14262;
	G17014<= not G14297;
	G17015<= not I18143;
	G17056<= not G13437;
	G17058<= not I18148;
	G17059<= not I18151;
	G17062<= not I18154;
	G17085<= not G14238;
	G17086<= not G14297;
	G17087<= not G14321;
	G17088<= not I18160;
	G17092<= not G14011;
	G17093<= not I18165;
	G17096<= not I18168;
	G17120<= not G14262;
	G17121<= not G14321;
	G17122<= not G14348;
	G17124<= not G14051;
	G17125<= not I18177;
	G17128<= not I18180;
	G17135<= not G14297;
	G17136<= not G14348;
	G17141<= not I18191;
	G17144<= not G14085;
	G17147<= not G14321;
	G17154<= not G14348;
	G17155<= not I18205;
	G17157<= not G13350;
	G17178<= not I18214;
	G17183<= not I18221;
	G17188<= not I18224;
	G17189<= not G14708;
	G17197<= not I18233;
	G17200<= not I18238;
	G17216<= not G14454;
	G17221<= not I18245;
	G17224<= not I18248;
	G17226<= not I18252;
	G17242<= not G14454;
	G17247<= not I18259;
	G17248<= not I18262;
	G17249<= not I18265;
	G17271<= not I18270;
	G17291<= not I18276;
	G17296<= not I18280;
	G17301<= not G14454;
	G17302<= not I18285;
	G17308<= not G14876;
	G17316<= not I18293;
	G17320<= not I18297;
	G17324<= not I18301;
	G17325<= not I18304;
	G17326<= not I18307;
	G17327<= not I18310;
	G17328<= not I18313;
	G17366<= not G14454;
	G17367<= not I18320;
	G17384<= not I18323;
	G17389<= not G14915;
	G17390<= not G14755;
	G17392<= not G14924;
	G17400<= not I18333;
	G17404<= not I18337;
	G17408<= not I18341;
	G17409<= not I18344;
	G17410<= not G12955;
	G17411<= not G14454;
	G17413<= not I18350;
	G17414<= not G14627;
	G17415<= not G14797;
	G17416<= not G14956;
	G17417<= not G14804;
	G17419<= not G14965;
	G17423<= not I18360;
	G17427<= not I18364;
	G17428<= not I18367;
	G17429<= not I18370;
	G17430<= not I18373;
	G17431<= not I18376;
	G17432<= not I18379;
	G17433<= not I18382;
	G17465<= not G12955;
	G17466<= not G12983;
	G17467<= not G14339;
	G17470<= not G14454;
	G17471<= not G14454;
	G17472<= not G14656;
	G17473<= not G14841;
	G17475<= not I18398;
	G17476<= not G14665;
	G17477<= not G14848;
	G17478<= not G14996;
	G17479<= not G14855;
	G17481<= not G15005;
	G17485<= not I18408;
	G17486<= not I18411;
	G17487<= not I18414;
	G17489<= not G12955;
	G17491<= not G12983;
	G17494<= not G14339;
	G17496<= not G14683;
	G17497<= not G14879;
	G17498<= not G14688;
	G17499<= not G14885;
	G17501<= not I18434;
	G17502<= not G14697;
	G17503<= not G14892;
	G17504<= not G15021;
	G17505<= not G14899;
	G17507<= not G15030;
	G17508<= not I18443;
	G17509<= not I18446;
	G17512<= not G12983;
	G17518<= not G14918;
	G17519<= not I18460;
	G17521<= not G14727;
	G17522<= not G14927;
	G17523<= not G14732;
	G17524<= not G14933;
	G17526<= not I18469;
	G17527<= not G14741;
	G17528<= not G14940;
	G17529<= not G15039;
	G17530<= not G14947;
	G17531<= not I18476;
	G17532<= not I18479;
	G17533<= not I18482;
	G17573<= not G12911;
	G17575<= not G14921;
	G17576<= not G14953;
	G17577<= not I18504;
	G17579<= not G14959;
	G17580<= not I18509;
	G17582<= not G14768;
	G17583<= not G14968;
	G17584<= not G14773;
	G17585<= not G14974;
	G17587<= not I18518;
	G17588<= not G14782;
	G17589<= not G14981;
	G17590<= not I18523;
	G17591<= not I18526;
	G17599<= not G14794;
	G17600<= not G14659;
	G17602<= not G14962;
	G17603<= not G14993;
	G17604<= not I18555;
	G17606<= not G14999;
	G17607<= not I18560;
	G17609<= not G14817;
	G17610<= not G15008;
	G17611<= not G14822;
	G17612<= not G15014;
	G17614<= not I18571;
	G17615<= not I18574;
	G17616<= not G14309;
	G17637<= not G12933;
	G17638<= not G14838;
	G17639<= not I18600;
	G17641<= not G14845;
	G17642<= not G14691;
	G17644<= not G15002;
	G17645<= not G15018;
	G17646<= not I18609;
	G17648<= not G15024;
	G17649<= not I18614;
	G17651<= not G14868;
	G17652<= not G15033;
	G17672<= not G14720;
	G17673<= not G14723;
	G17674<= not I18647;
	G17676<= not G12941;
	G17677<= not G14882;
	G17678<= not I18653;
	G17680<= not G14889;
	G17681<= not G14735;
	G17683<= not G15027;
	G17684<= not G15036;
	G17685<= not I18662;
	G17687<= not G15042;
	G17688<= not I18667;
	G17691<= not I18674;
	G17707<= not G14758;
	G17709<= not G14761;
	G17710<= not G14764;
	G17711<= not I18694;
	G17713<= not G12947;
	G17714<= not G14930;
	G17715<= not I18700;
	G17717<= not G14937;
	G17718<= not G14776;
	G17720<= not G15045;
	G17721<= not G12915;
	G17722<= not I18709;
	G17733<= not G14238;
	G17735<= not G14807;
	G17737<= not G14810;
	G17738<= not G14813;
	G17739<= not I18728;
	G17741<= not G12972;
	G17742<= not G14971;
	G17743<= not I18734;
	G17745<= not G14978;
	G17746<= not G14825;
	G17754<= not G14262;
	G17756<= not G14858;
	G17758<= not G14861;
	G17759<= not G14864;
	G17760<= not I18752;
	G17762<= not G13000;
	G17763<= not G15011;
	G17764<= not I18758;
	G17772<= not G14297;
	G17774<= not G14902;
	G17776<= not G14905;
	G17777<= not G14908;
	G17778<= not I18778;
	G17782<= not I18788;
	G17787<= not I18795;
	G17789<= not G14321;
	G17791<= not G14950;
	G17794<= not G13350;
	G17811<= not G12925;
	G17812<= not I18810;
	G17813<= not I18813;
	G17815<= not G14348;
	G17818<= not I18822;
	G17819<= not I18825;
	G17821<= not I18829;
	G17844<= not I18832;
	G17845<= not I18835;
	G17847<= not I18839;
	G17870<= not I18842;
	G17871<= not I18845;
	G17873<= not I18849;
	G17926<= not I18852;
	G17929<= not I18855;
	G17952<= not I18858;
	G17953<= not I18861;
	G17955<= not I18865;
	G18008<= not I18868;
	G18061<= not G14800;
	G18062<= not I18872;
	G18065<= not I18875;
	G18088<= not G13267;
	G18091<= not I18879;
	G18092<= not I18882;
	G18093<= not I18885;
	G18094<= not I18888;
	G18095<= not I18891;
	G18096<= not I18894;
	G18097<= not I18897;
	G18098<= not I18900;
	G18099<= not I18903;
	G18100<= not I18906;
	G18101<= not I18909;
	G18102<= not I18912;
	G18200<= not I19012;
	G18421<= not I19235;
	G18422<= not I19238;
	G18527<= not I19345;
	G18528<= not I19348;
	G18562<= not I19384;
	G18660<= not I19484;
	G18661<= not I19487;
	G18827<= not G16000;
	G18828<= not G17955;
	G18829<= not G15171;
	G18830<= not G18008;
	G18831<= not G15224;
	G18832<= not G15634;
	G18833<= not I19661;
	G18874<= not G15938;
	G18875<= not G15171;
	G18876<= not G15373;
	G18877<= not G15224;
	G18878<= not G15426;
	G18880<= not G15656;
	G18881<= not I19671;
	G18882<= not I19674;
	G18883<= not G15938;
	G18884<= not G15938;
	G18885<= not G15979;
	G18886<= not G16000;
	G18887<= not G15373;
	G18888<= not G15426;
	G18889<= not G15509;
	G18891<= not G16053;
	G18892<= not G15680;
	G18894<= not G16000;
	G18895<= not G16000;
	G18896<= not G16031;
	G18897<= not G15509;
	G18898<= not G15566;
	G18903<= not G15758;
	G18904<= not G16053;
	G18905<= not G16077;
	G18907<= not G15979;
	G18908<= not G16100;
	G18911<= not G15169;
	G18916<= not G16053;
	G18917<= not G16077;
	G18918<= not I19704;
	G18926<= not I19707;
	G18929<= not G16100;
	G18930<= not G15789;
	G18931<= not G16031;
	G18932<= not G16136;
	G18938<= not G16053;
	G18939<= not G16077;
	G18940<= not I19719;
	G18944<= not G15938;
	G18945<= not G16100;
	G18946<= not G16100;
	G18947<= not G16136;
	G18948<= not G15800;
	G18952<= not G16053;
	G18953<= not G16077;
	G18954<= not G17427;
	G18957<= not I19734;
	G18975<= not G15938;
	G18976<= not G16100;
	G18977<= not G16100;
	G18978<= not G16000;
	G18979<= not G16136;
	G18980<= not G16136;
	G18983<= not G16077;
	G18984<= not G17486;
	G18988<= not G15979;
	G18989<= not G16000;
	G18990<= not G16136;
	G18991<= not G16136;
	G18997<= not I19756;
	G19050<= not I19759;
	G19061<= not I19762;
	G19067<= not G15979;
	G19068<= not G16031;
	G19071<= not G15591;
	G19074<= not I19772;
	G19127<= not I19775;
	G19128<= not I19778;
	G19144<= not G16031;
	G19146<= not G15574;
	G19147<= not I19786;
	G19200<= not I19789;
	G19208<= not G17367;
	G19210<= not I19796;
	G19263<= not I19799;
	G19264<= not I19802;
	G19273<= not G16100;
	G19276<= not G17367;
	G19277<= not I19813;
	G19330<= not G17326;
	G19334<= not I19818;
	G19343<= not G16136;
	G19345<= not G17591;
	G19351<= not G17367;
	G19352<= not G15758;
	G19353<= not I19831;
	G19355<= not G16027;
	G19357<= not I19837;
	G19360<= not G16249;
	G19361<= not I19843;
	G19362<= not G16072;
	G19364<= not G15825;
	G19365<= not G16249;
	G19366<= not G15885;
	G19367<= not I19851;
	G19368<= not G16326;
	G19369<= not G15995;
	G19370<= not G15915;
	G19371<= not I19857;
	G19373<= not G16449;
	G19374<= not G16047;
	G19375<= not I19863;
	G19376<= not G17509;
	G19379<= not G17327;
	G19385<= not G16326;
	G19386<= not G16431;
	G19387<= not G16431;
	G19389<= not G17532;
	G19394<= not G16326;
	G19395<= not G16431;
	G19396<= not G16431;
	G19397<= not G16449;
	G19398<= not G16489;
	G19399<= not G16489;
	G19407<= not G16268;
	G19408<= not G16066;
	G19409<= not G16431;
	G19410<= not G16449;
	G19411<= not G16489;
	G19412<= not G16489;
	G19414<= not G16349;
	G19415<= not G15758;
	G19416<= not G15885;
	G19417<= not G17178;
	G19421<= not G16326;
	G19427<= not G16292;
	G19428<= not G16090;
	G19429<= not G16489;
	G19431<= not G16249;
	G19432<= not G15885;
	G19433<= not G15915;
	G19434<= not G16326;
	G19435<= not G16449;
	G19437<= not G16349;
	G19438<= not G16249;
	G19439<= not G15885;
	G19440<= not G15915;
	G19443<= not G16449;
	G19445<= not G15915;
	G19446<= not I19917;
	G19451<= not G15938;
	G19452<= not G16326;
	G19454<= not G16349;
	G19458<= not I19927;
	G19468<= not G15938;
	G19469<= not G16326;
	G19470<= not G16000;
	G19471<= not G16449;
	G19472<= not G16349;
	G19473<= not G16349;
	G19476<= not G16326;
	G19477<= not G16431;
	G19478<= not G16000;
	G19479<= not G16449;
	G19480<= not G16349;
	G19481<= not G16349;
	G19482<= not G16349;
	G19489<= not G16449;
	G19490<= not G16489;
	G19491<= not G16349;
	G19492<= not G16349;
	G19493<= not G16349;
	G19494<= not G16349;
	G19498<= not G16752;
	G19499<= not G16782;
	G19502<= not G15674;
	G19503<= not G16349;
	G19504<= not G16349;
	G19505<= not G16349;
	G19517<= not G16777;
	G19518<= not G16239;
	G19519<= not G16795;
	G19520<= not G16826;
	G19523<= not G16100;
	G19524<= not G15695;
	G19526<= not G16349;
	G19527<= not G16349;
	G19528<= not G16349;
	G19529<= not G16349;
	G19531<= not G16816;
	G19532<= not G16821;
	G19533<= not G16261;
	G19537<= not G15938;
	G19538<= not G16100;
	G19539<= not G16129;
	G19541<= not G16136;
	G19542<= not G16349;
	G19543<= not G16349;
	G19544<= not G16349;
	G19552<= not G16856;
	G19553<= not G16782;
	G19554<= not G16861;
	G19558<= not G15938;
	G19559<= not G16129;
	G19565<= not G16000;
	G19566<= not G16136;
	G19567<= not G16164;
	G19569<= not G16349;
	G19570<= not G16349;
	G19573<= not G16877;
	G19574<= not G16826;
	G19577<= not G16129;
	G19579<= not G16000;
	G19580<= not G16164;
	G19586<= not G16349;
	G19592<= not I20035;
	G19600<= not G16164;
	G19602<= not G16349;
	G19603<= not G16349;
	G19606<= not G17614;
	G19609<= not G16264;
	G19612<= not G16897;
	G19617<= not G16349;
	G19618<= not G16349;
	G19620<= not G17296;
	G19626<= not G17409;
	G19629<= not G17015;
	G19630<= not G16897;
	G19633<= not G16931;
	G19634<= not G16349;
	G19635<= not G16349;
	G19636<= not G16987;
	G19638<= not G17324;
	G19644<= not G17953;
	G19649<= not G17015;
	G19650<= not G16971;
	G19652<= not G16897;
	G19653<= not G16897;
	G19654<= not G16931;
	G19657<= not G16349;
	G19658<= not G16987;
	G19659<= not G17062;
	G19662<= not G17432;
	G19666<= not G17188;
	G19670<= not G16897;
	G19672<= not G16931;
	G19673<= not G16931;
	G19675<= not G16987;
	G19676<= not G17062;
	G19677<= not G17096;
	G19678<= not G16752;
	G19679<= not G16782;
	G19682<= not G17015;
	G19683<= not G16931;
	G19685<= not G16987;
	G19686<= not G17062;
	G19687<= not G17096;
	G19688<= not G16777;
	G19689<= not G16795;
	G19690<= not G16826;
	G19694<= not G16429;
	G19695<= not G17015;
	G19696<= not G17015;
	G19697<= not G16886;
	G19698<= not G16971;
	G19699<= not I20116;
	G19709<= not G16987;
	G19710<= not G17059;
	G19711<= not G17062;
	G19712<= not G17096;
	G19713<= not G16816;
	G19714<= not G16821;
	G19718<= not G17015;
	G19719<= not G16897;
	G19720<= not I20130;
	G19730<= not G17062;
	G19731<= not G17093;
	G19732<= not G17096;
	G19733<= not G16856;
	G19734<= not G16861;
	G19737<= not G17015;
	G19738<= not G15992;
	G19739<= not G16931;
	G19741<= not G16987;
	G19742<= not G17096;
	G19743<= not G17125;
	G19744<= not G15885;
	G19745<= not G16877;
	G19747<= not G17015;
	G19748<= not G17015;
	G19750<= not G16326;
	G19751<= not G16044;
	G19753<= not G16987;
	G19754<= not G17062;
	G19755<= not G15915;
	G19757<= not G17224;
	G19760<= not G17015;
	G19761<= not G17015;
	G19762<= not G16326;
	G19763<= not G16431;
	G19765<= not G16897;
	G19766<= not G16449;
	G19769<= not G16987;
	G19770<= not G17062;
	G19771<= not G17096;
	G19772<= not G17183;
	G19773<= not G17615;
	G19776<= not G17015;
	G19777<= not G17015;
	G19779<= not G16431;
	G19780<= not G16449;
	G19781<= not G16489;
	G19783<= not G16931;
	G19785<= not G16987;
	G19786<= not G17062;
	G19787<= not G17096;
	G19789<= not G17015;
	G19790<= not G16971;
	G19794<= not G16489;
	G19798<= not G17200;
	G19799<= not G17062;
	G19800<= not G17096;
	G19801<= not I20216;
	G19852<= not G17015;
	G19860<= not G17226;
	G19861<= not G17096;
	G19862<= not I20233;
	G19865<= not G15885;
	G19866<= not G16540;
	G19869<= not G16540;
	G19872<= not G17015;
	G19878<= not G17271;
	G19881<= not G15915;
	G19882<= not G16540;
	G19885<= not G17249;
	G19902<= not G17200;
	G19905<= not G15885;
	G19908<= not G16540;
	G19912<= not G17328;
	G19915<= not G16349;
	G19930<= not G17200;
	G19931<= not G17200;
	G19947<= not G17226;
	G19950<= not G15885;
	G19952<= not G15915;
	G19954<= not G16540;
	G19957<= not G16540;
	G19960<= not G17433;
	G19961<= not G17328;
	G19963<= not G16326;
	G19964<= not G17200;
	G19979<= not G17226;
	G19980<= not G17226;
	G19996<= not G17271;
	G19998<= not G15915;
	G20004<= not G17249;
	G20005<= not G17433;
	G20006<= not G17328;
	G20008<= not G16449;
	G20009<= not G16349;
	G20010<= not G17226;
	G20025<= not G17271;
	G20026<= not G17271;
	G20028<= not G15371;
	G20033<= not G16579;
	G20035<= not G16430;
	G20036<= not G17433;
	G20037<= not G17328;
	G20038<= not G17328;
	G20040<= not G17271;
	G20041<= not G15569;
	G20046<= not G16540;
	G20049<= not I20318;
	G20050<= not I20321;
	G20052<= not G17533;
	G20053<= not G17328;
	G20054<= not G17328;
	G20057<= not G16349;
	G20058<= not G16782;
	G20059<= not G17302;
	G20060<= not G16540;
	G20064<= not G17533;
	G20065<= not G16846;
	G20066<= not G17433;
	G20067<= not G17328;
	G20070<= not G16173;
	G20071<= not G16826;
	G20072<= not G17384;
	G20073<= not G16540;
	G20078<= not G16846;
	G20079<= not G17328;
	G20080<= not G17328;
	G20085<= not G16187;
	G20086<= not I20355;
	G20087<= not G17249;
	G20088<= not G17533;
	G20089<= not G17533;
	G20090<= not G17433;
	G20091<= not G17328;
	G20096<= not G16782;
	G20097<= not G17691;
	G20100<= not I20369;
	G20101<= not G17533;
	G20102<= not G17533;
	G20103<= not G17433;
	G20104<= not G17433;
	G20105<= not G17433;
	G20106<= not G17328;
	G20110<= not G16897;
	G20113<= not G16826;
	G20114<= not I20385;
	G20127<= not I20388;
	G20128<= not G17533;
	G20129<= not G17328;
	G20130<= not G17328;
	G20132<= not G16931;
	G20136<= not I20399;
	G20144<= not G17533;
	G20145<= not G17533;
	G20146<= not G17533;
	G20147<= not G17328;
	G20153<= not G16782;
	G20154<= not I20412;
	G20157<= not G16886;
	G20158<= not G16971;
	G20159<= not G17533;
	G20164<= not G16826;
	G20166<= not G16886;
	G20167<= not G16971;
	G20168<= not G17533;
	G20175<= not I20433;
	G20178<= not G16971;
	G20179<= not G17249;
	G20180<= not G17533;
	G20182<= not G16897;
	G20189<= not I20447;
	G20190<= not G16971;
	G20191<= not G17821;
	G20192<= not G17268;
	G20194<= not G16897;
	G20195<= not G16931;
	G20197<= not G16987;
	G20204<= not G16578;
	G20207<= not G17015;
	G20208<= not G17533;
	G20209<= not G17821;
	G20210<= not G16897;
	G20211<= not G16931;
	G20212<= not G17194;
	G20213<= not G17062;
	G20219<= not I20495;
	G20229<= not G17015;
	G20230<= not I20499;
	G20231<= not G17821;
	G20232<= not G16931;
	G20233<= not G17873;
	G20235<= not G15277;
	G20237<= not G17213;
	G20238<= not G17096;
	G20239<= not G17128;
	G20240<= not G17847;
	G20242<= not G16308;
	G20247<= not G17015;
	G20265<= not G17821;
	G20266<= not G17873;
	G20267<= not G17955;
	G20268<= not G18008;
	G20269<= not G15844;
	G20270<= not G15277;
	G20272<= not G17239;
	G20273<= not G17128;
	G20274<= not G17847;
	G20275<= not G17929;
	G20277<= not G16487;
	G20283<= not I20529;
	G20320<= not G17015;
	G20321<= not G17821;
	G20322<= not G17873;
	G20323<= not G17873;
	G20324<= not G17955;
	G20325<= not G15171;
	G20326<= not G18008;
	G20327<= not G15224;
	G20328<= not G15867;
	G20329<= not G15277;
	G20330<= not I20542;
	G20372<= not G17847;
	G20373<= not G17929;
	G20374<= not G18065;
	G20379<= not G17821;
	G20380<= not G17955;
	G20381<= not G17955;
	G20382<= not G15171;
	G20383<= not G15373;
	G20384<= not G18008;
	G20385<= not G18008;
	G20386<= not G15224;
	G20387<= not G15426;
	G20388<= not G17297;
	G20389<= not G15277;
	G20391<= not I20562;
	G20432<= not G17847;
	G20433<= not G17929;
	G20434<= not G18065;
	G20435<= not G15348;
	G20436<= not I20569;
	G20441<= not G17873;
	G20442<= not G15171;
	G20443<= not G15171;
	G20444<= not G15373;
	G20445<= not G15224;
	G20446<= not G15224;
	G20447<= not G15426;
	G20448<= not G15509;
	G20449<= not G15277;
	G20450<= not G15277;
	G20451<= not G15277;
	G20452<= not G17200;
	G20453<= not I20584;
	G20494<= not G17847;
	G20495<= not G17926;
	G20496<= not G17929;
	G20497<= not G18065;
	G20498<= not G15348;
	G20499<= not G15483;
	G20500<= not G17873;
	G20501<= not G17955;
	G20502<= not G15373;
	G20503<= not G15373;
	G20504<= not G18008;
	G20505<= not G15426;
	G20506<= not G15426;
	G20507<= not G15509;
	G20508<= not G15277;
	G20509<= not G15277;
	G20510<= not G17226;
	G20511<= not G17929;
	G20512<= not G18062;
	G20513<= not G18065;
	G20514<= not G15348;
	G20515<= not G15483;
	G20516<= not I20609;
	G20523<= not G17821;
	G20524<= not G17873;
	G20525<= not G17955;
	G20526<= not G15171;
	G20527<= not G18008;
	G20528<= not G15224;
	G20529<= not G15509;
	G20530<= not G15509;
	G20531<= not G15907;
	G20532<= not G15277;
	G20533<= not G17271;
	G20534<= not G17183;
	G20535<= not G17847;
	G20536<= not G18065;
	G20537<= not G15345;
	G20538<= not G15348;
	G20539<= not G15483;
	G20540<= not G16646;
	G20541<= not G17821;
	G20542<= not G17873;
	G20543<= not G17955;
	G20544<= not G15171;
	G20545<= not G15373;
	G20546<= not G18008;
	G20547<= not G15224;
	G20548<= not G15426;
	G20549<= not G15277;
	G20550<= not G15864;
	G20551<= not G17302;
	G20552<= not G17847;
	G20553<= not G17929;
	G20554<= not G15348;
	G20555<= not G15480;
	G20556<= not G15483;
	G20557<= not I20647;
	G20558<= not I20650;
	G20560<= not G17328;
	G20561<= not G17873;
	G20562<= not G17955;
	G20563<= not G15171;
	G20564<= not G15373;
	G20565<= not G18008;
	G20566<= not G15224;
	G20567<= not G15426;
	G20568<= not G15509;
	G20569<= not G15277;
	G20570<= not G15277;
	G20571<= not G15277;
	G20572<= not G15833;
	G20573<= not G17384;
	G20574<= not G17847;
	G20575<= not G17929;
	G20576<= not G18065;
	G20577<= not G15483;
	G20578<= not G15563;
	G20579<= not G17249;
	G20580<= not G17328;
	G20582<= not G17873;
	G20583<= not G17873;
	G20584<= not G17873;
	G20585<= not G17955;
	G20586<= not G15171;
	G20587<= not G15373;
	G20588<= not G18008;
	G20589<= not G15224;
	G20590<= not G15426;
	G20591<= not G15509;
	G20592<= not G15277;
	G20593<= not G15277;
	G20594<= not G15277;
	G20595<= not G15877;
	G20596<= not I20690;
	G20597<= not G17847;
	G20598<= not G17929;
	G20599<= not G18065;
	G20600<= not G15348;
	G20601<= not G17433;
	G20603<= not G17873;
	G20604<= not G17873;
	G20605<= not G17955;
	G20606<= not G17955;
	G20607<= not G17955;
	G20608<= not G15171;
	G20609<= not G15373;
	G20610<= not G18008;
	G20611<= not G18008;
	G20612<= not G18008;
	G20613<= not G15224;
	G20614<= not G15426;
	G20615<= not G15509;
	G20616<= not G15277;
	G20617<= not G15277;
	G20618<= not G15277;
	G20622<= not G15595;
	G20623<= not G17929;
	G20624<= not G18065;
	G20625<= not G15348;
	G20626<= not G15483;
	G20627<= not G17433;
	G20629<= not G17955;
	G20630<= not G17955;
	G20631<= not G15171;
	G20632<= not G15171;
	G20633<= not G15171;
	G20634<= not G15373;
	G20635<= not G18008;
	G20636<= not G18008;
	G20637<= not G15224;
	G20638<= not G15224;
	G20639<= not G15224;
	G20640<= not G15426;
	G20641<= not G15509;
	G20642<= not G15277;
	G20643<= not G15962;
	G20648<= not G15615;
	G20649<= not G18065;
	G20650<= not G15348;
	G20651<= not G15483;
	G20652<= not I20744;
	G20653<= not I20747;
	G20654<= not I20750;
	G20655<= not I20753;
	G20656<= not G17249;
	G20657<= not G17433;
	G20659<= not G17873;
	G20660<= not G17873;
	G20661<= not G15171;
	G20662<= not G15171;
	G20663<= not G15373;
	G20664<= not G15373;
	G20665<= not G15373;
	G20666<= not G15224;
	G20667<= not G15224;
	G20668<= not G15426;
	G20669<= not G15426;
	G20670<= not G15426;
	G20671<= not G15509;
	G20672<= not G15277;
	G20673<= not G15277;
	G20674<= not G15277;
	G20679<= not G15634;
	G20680<= not G15348;
	G20681<= not G15483;
	G20695<= not I20781;
	G20696<= not G17533;
	G20697<= not G17433;
	G20698<= not G17873;
	G20699<= not G17873;
	G20700<= not G17873;
	G20701<= not G17955;
	G20702<= not G17955;
	G20703<= not G15373;
	G20704<= not G15373;
	G20705<= not I20793;
	G20706<= not G18008;
	G20707<= not G18008;
	G20708<= not G15426;
	G20709<= not G15426;
	G20710<= not G15509;
	G20711<= not G15509;
	G20712<= not G15509;
	G20713<= not G15277;
	G20714<= not G15277;
	G20715<= not G15277;
	G20716<= not G15277;
	G20732<= not G15595;
	G20737<= not G15656;
	G20738<= not G15483;
	G20763<= not I20816;
	G20764<= not I20819;
	G20765<= not G17748;
	G20766<= not G17433;
	G20767<= not G17873;
	G20768<= not G17955;
	G20769<= not G17955;
	G20770<= not G17955;
	G20771<= not G15171;
	G20772<= not G15171;
	G20773<= not I20830;
	G20774<= not G18008;
	G20775<= not G18008;
	G20776<= not G18008;
	G20777<= not G15224;
	G20778<= not G15224;
	G20779<= not G15509;
	G20780<= not G15509;
	G20781<= not I20840;
	G20782<= not G15853;
	G20785<= not I20846;
	G20852<= not G15595;
	G20853<= not G15595;
	G20869<= not G15615;
	G20874<= not G15680;
	G20899<= not I20861;
	G20900<= not I20864;
	G20901<= not I20867;
	G20902<= not I20870;
	G20903<= not G17249;
	G20904<= not G17433;
	G20909<= not G17955;
	G20910<= not G15171;
	G20911<= not G15171;
	G20912<= not G15171;
	G20913<= not G15373;
	G20914<= not G15373;
	G20915<= not I20882;
	G20916<= not G18008;
	G20917<= not G15224;
	G20918<= not G15224;
	G20919<= not G15224;
	G20920<= not G15426;
	G20921<= not G15426;
	G20922<= not I20891;
	G20923<= not G15277;
	G20924<= not I20895;
	G20978<= not G15595;
	G20993<= not G15615;
	G20994<= not G15615;
	G21010<= not G15634;
	G21036<= not I20910;
	G21037<= not I20913;
	G21048<= not G17533;
	G21049<= not G17433;
	G21050<= not G17873;
	G21051<= not G15171;
	G21052<= not G15373;
	G21053<= not G15373;
	G21054<= not G15373;
	G21055<= not G15224;
	G21056<= not G15426;
	G21057<= not G15426;
	G21058<= not G15426;
	G21059<= not G15509;
	G21060<= not G15509;
	G21061<= not I20929;
	G21068<= not G15277;
	G21069<= not G15277;
	G21070<= not I20937;
	G21123<= not G15615;
	G21138<= not G15634;
	G21139<= not G15634;
	G21155<= not G15656;
	G21156<= not G17247;
	G21160<= not G17508;
	G21175<= not I20951;
	G21176<= not I20954;
	G21177<= not I20957;
	G21178<= not G17955;
	G21179<= not G15373;
	G21180<= not G18008;
	G21181<= not G15426;
	G21182<= not G15509;
	G21183<= not G15509;
	G21184<= not G15509;
	G21185<= not G15277;
	G21189<= not G15634;
	G21204<= not G15656;
	G21205<= not G15656;
	G21221<= not G15680;
	G21222<= not G17430;
	G21225<= not G17428;
	G21228<= not G17531;
	G21245<= not I20982;
	G21246<= not I20985;
	G21247<= not G15171;
	G21248<= not G15224;
	G21249<= not G15509;
	G21252<= not G15656;
	G21267<= not G15680;
	G21268<= not G15680;
	G21269<= not G15506;
	G21270<= not I20999;
	G21271<= not I21002;
	G21273<= not I21006;
	G21274<= not G15373;
	G21275<= not G15426;
	G21278<= not I21013;
	G21279<= not G15680;
	G21280<= not G16601;
	G21281<= not G16286;
	G21282<= not I21019;
	G21286<= not G15509;
	G21290<= not I21029;
	G21291<= not G16620;
	G21292<= not I21033;
	G21293<= not I21036;
	G21295<= not G17533;
	G21297<= not I21042;
	G21299<= not G16600;
	G21300<= not I21047;
	G21304<= not G17367;
	G21305<= not G15758;
	G21306<= not G15582;
	G21308<= not G17485;
	G21326<= not I21058;
	G21329<= not G16577;
	G21335<= not I21067;
	G21336<= not G17367;
	G21337<= not G15758;
	G21340<= not I21074;
	G21343<= not G16428;
	G21346<= not G17821;
	G21349<= not G15758;
	G21352<= not G16322;
	G21355<= not G17821;
	G21358<= not G16307;
	G21362<= not G17873;
	G21366<= not I21100;
	G21369<= not G16285;
	G21370<= not G16323;
	G21379<= not G17873;
	G21380<= not G17955;
	G21381<= not G18008;
	G21383<= not G17367;
	G21387<= not I21115;
	G21393<= not G17264;
	G21395<= not G17873;
	G21396<= not G17955;
	G21397<= not G15171;
	G21398<= not G18008;
	G21399<= not G15224;
	G21400<= not G17847;
	G21406<= not G17955;
	G21407<= not G15171;
	G21408<= not G15373;
	G21409<= not G18008;
	G21410<= not G15224;
	G21411<= not G15426;
	G21412<= not G15758;
	G21413<= not G15585;
	G21414<= not G17929;
	G21418<= not G17821;
	G21421<= not G15171;
	G21422<= not G15373;
	G21423<= not G15224;
	G21424<= not G15426;
	G21425<= not G15509;
	G21426<= not G15277;
	G21427<= not G17367;
	G21428<= not G15758;
	G21430<= not G15608;
	G21431<= not G18065;
	G21434<= not G17248;
	G21451<= not I21162;
	G21454<= not G15373;
	G21455<= not G15426;
	G21456<= not G15509;
	G21457<= not G17367;
	G21458<= not G15758;
	G21460<= not G15628;
	G21461<= not G15348;
	G21463<= not G15588;
	G21466<= not G15509;
	G21467<= not G15758;
	G21468<= not I21181;
	G21510<= not G15647;
	G21511<= not G15483;
	G21514<= not I21189;
	G21556<= not G15669;
	G21560<= not G17873;
	G21561<= not G15595;
	G21562<= not I21199;
	G21604<= not G15938;
	G21607<= not G17873;
	G21608<= not G17955;
	G21609<= not G18008;
	G21610<= not G15615;
	G21611<= not I21210;
	G21653<= not G17663;
	G21654<= not G17619;
	G21656<= not G17700;
	G21657<= not G17657;
	G21659<= not G17727;
	G21660<= not G17694;
	G21661<= not I21222;
	G21662<= not G16540;
	G21665<= not I21226;
	G21666<= not G16540;
	G21669<= not I21230;
	G21670<= not G16540;
	G21673<= not I21234;
	G21674<= not G16540;
	G21677<= not I21238;
	G21678<= not G16540;
	G21681<= not I21242;
	G21682<= not G16540;
	G21685<= not I21246;
	G21686<= not G16540;
	G21689<= not I21250;
	G21690<= not G16540;
	G21693<= not I21254;
	G21694<= not G16540;
	G21697<= not I21258;
	G21698<= not G18562;
	G21722<= not I21285;
	G21723<= not I21288;
	G21724<= not I21291;
	G21725<= not I21294;
	G21726<= not I21297;
	G21727<= not I21300;
	G21902<= not I21477;
	G21903<= not I21480;
	G21904<= not I21483;
	G21905<= not I21486;
	G22136<= not G20277;
	G22137<= not G21370;
	G22138<= not G21370;
	G22139<= not I21722;
	G22144<= not G18997;
	G22146<= not G18997;
	G22147<= not G18997;
	G22148<= not G19074;
	G22150<= not G21280;
	G22151<= not I21734;
	G22153<= not G18997;
	G22154<= not G19074;
	G22155<= not G19074;
	G22156<= not G19147;
	G22159<= not I21744;
	G22166<= not G18997;
	G22167<= not G19074;
	G22168<= not G19147;
	G22169<= not G19147;
	G22170<= not G19210;
	G22171<= not G18882;
	G22173<= not I21757;
	G22176<= not G18997;
	G22177<= not G19074;
	G22178<= not G19147;
	G22179<= not G19210;
	G22180<= not G19210;
	G22181<= not G19277;
	G22182<= not I21766;
	G22189<= not I21769;
	G22192<= not G19801;
	G22194<= not I21776;
	G22197<= not G19074;
	G22198<= not G19147;
	G22199<= not G19210;
	G22200<= not G19277;
	G22201<= not G19277;
	G22202<= not I21784;
	G22207<= not I21787;
	G22210<= not I21792;
	G22213<= not G19147;
	G22214<= not G19210;
	G22215<= not G19277;
	G22220<= not I21802;
	G22223<= not G19210;
	G22224<= not G19277;
	G22227<= not G19801;
	G22228<= not I21810;
	G22300<= not I21815;
	G22303<= not G19277;
	G22305<= not G19801;
	G22311<= not G18935;
	G22317<= not G19801;
	G22319<= not I21831;
	G22330<= not G19801;
	G22332<= not I21838;
	G22338<= not G19801;
	G22339<= not G19801;
	G22341<= not G19801;
	G22358<= not G19801;
	G22359<= not G19495;
	G22360<= not I21849;
	G22406<= not G19506;
	G22407<= not G19455;
	G22408<= not G19483;
	G22409<= not I21860;
	G22449<= not G19597;
	G22455<= not G19801;
	G22456<= not G19801;
	G22492<= not G19614;
	G22493<= not G19801;
	G22494<= not G19801;
	G22495<= not G19801;
	G22496<= not G19510;
	G22497<= not G19513;
	G22519<= not G19801;
	G22520<= not G19801;
	G22526<= not G19801;
	G22527<= not G19546;
	G22528<= not G19801;
	G22529<= not G19549;
	G22541<= not I21911;
	G22542<= not G19801;
	G22543<= not G19801;
	G22544<= not G19589;
	G22546<= not I21918;
	G22550<= not I21922;
	G22592<= not I21930;
	G22593<= not G19801;
	G22594<= not I21934;
	G22626<= not I21941;
	G22635<= not G19801;
	G22646<= not G19389;
	G22647<= not I21959;
	G22649<= not G19063;
	G22658<= not I21969;
	G22660<= not G19140;
	G22667<= not G21156;
	G22682<= not G19379;
	G22683<= not I22000;
	G22698<= not I22009;
	G22714<= not G20436;
	G22716<= not G19795;
	G22718<= not G20887;
	G22719<= not I22024;
	G22721<= not I22028;
	G22722<= not I22031;
	G22756<= not G20436;
	G22758<= not G20330;
	G22759<= not G19857;
	G22761<= not G21024;
	G22763<= not I22046;
	G22830<= not G20283;
	G22840<= not G20330;
	G22841<= not G20391;
	G22842<= not G19875;
	G22844<= not G21163;
	G22845<= not G20682;
	G22847<= not G20283;
	G22854<= not G20330;
	G22855<= not G20391;
	G22856<= not G20453;
	G22857<= not G20739;
	G22858<= not G20751;
	G22860<= not G20000;
	G22865<= not G20330;
	G22866<= not G20330;
	G22867<= not G20391;
	G22868<= not G20453;
	G22869<= not G20875;
	G22870<= not G20887;
	G22881<= not I22096;
	G22882<= not G20391;
	G22883<= not G20391;
	G22884<= not G20453;
	G22896<= not G21012;
	G22897<= not G21024;
	G22898<= not G20283;
	G22903<= not G20330;
	G22904<= not I22111;
	G22905<= not I22114;
	G22906<= not G20453;
	G22907<= not G20453;
	G22919<= not G21163;
	G22922<= not G20330;
	G22923<= not I22124;
	G22926<= not G20391;
	G22927<= not I22128;
	G22928<= not I22131;
	G22935<= not G20283;
	G22936<= not G20283;
	G22957<= not I22143;
	G22973<= not G20330;
	G22974<= not G20330;
	G22975<= not G20391;
	G22976<= not I22149;
	G22979<= not G20453;
	G22980<= not I22153;
	G22981<= not G20283;
	G22985<= not G20330;
	G22986<= not G20330;
	G22987<= not G20391;
	G22988<= not G20391;
	G22989<= not G20453;
	G22994<= not G20436;
	G22995<= not G20330;
	G22996<= not G20330;
	G22997<= not G20391;
	G22998<= not G20391;
	G22999<= not G20453;
	G23000<= not G20453;
	G23001<= not G19801;
	G23002<= not I22177;
	G23003<= not I22180;
	G23004<= not G20283;
	G23005<= not G20283;
	G23011<= not G20330;
	G23012<= not G20330;
	G23013<= not G20330;
	G23014<= not G20391;
	G23015<= not G20391;
	G23016<= not G20453;
	G23017<= not G20453;
	G23018<= not G19801;
	G23019<= not G19866;
	G23020<= not G19869;
	G23021<= not G20283;
	G23022<= not G20283;
	G23026<= not G20391;
	G23027<= not G20391;
	G23028<= not G20391;
	G23029<= not G20453;
	G23030<= not G20453;
	G23031<= not G19801;
	G23032<= not I22211;
	G23041<= not G19882;
	G23046<= not G20283;
	G23055<= not G20887;
	G23057<= not G20453;
	G23058<= not G20453;
	G23059<= not G20453;
	G23060<= not G19908;
	G23061<= not G20283;
	G23066<= not G20330;
	G23082<= not G21024;
	G23084<= not G19954;
	G23085<= not G19957;
	G23086<= not G20283;
	G23088<= not I22240;
	G23111<= not G20391;
	G23127<= not G21163;
	G23128<= not G20283;
	G23138<= not G20453;
	G23152<= not G20283;
	G23154<= not I22264;
	G23170<= not G20046;
	G23172<= not I22275;
	G23182<= not G21389;
	G23189<= not G20060;
	G23190<= not I22286;
	G23191<= not I22289;
	G23192<= not G20248;
	G23196<= not G20785;
	G23202<= not I22302;
	G23203<= not G20073;
	G23211<= not G21308;
	G23214<= not G20785;
	G23215<= not G20785;
	G23216<= not G20924;
	G23219<= not I22316;
	G23221<= not G20785;
	G23222<= not G20785;
	G23223<= not G21308;
	G23226<= not G20924;
	G23227<= not G20924;
	G23228<= not G21070;
	G23230<= not I22327;
	G23231<= not G20050;
	G23232<= not I22331;
	G23233<= not G21037;
	G23234<= not G20375;
	G23235<= not G20785;
	G23236<= not G20785;
	G23237<= not G20924;
	G23238<= not G20924;
	G23239<= not G21308;
	G23242<= not G21070;
	G23243<= not G21070;
	G23244<= not I22343;
	G23245<= not G20785;
	G23246<= not G20785;
	G23247<= not G20924;
	G23248<= not G20924;
	G23249<= not G21070;
	G23250<= not G21070;
	G23252<= not I22353;
	G23253<= not G21037;
	G23256<= not G20785;
	G23257<= not G20924;
	G23258<= not G20924;
	G23259<= not G21070;
	G23260<= not G21070;
	G23263<= not I22366;
	G23264<= not G21037;
	G23267<= not G20097;
	G23270<= not G20785;
	G23271<= not G20785;
	G23272<= not G20924;
	G23273<= not G21070;
	G23274<= not G21070;
	G23277<= not I22380;
	G23278<= not G20283;
	G23279<= not G21037;
	G23282<= not G20330;
	G23283<= not G20785;
	G23284<= not G20785;
	G23285<= not G20887;
	G23289<= not G20924;
	G23290<= not G20924;
	G23291<= not G21070;
	G23299<= not I22400;
	G23300<= not G20283;
	G23301<= not G21037;
	G23302<= not G20330;
	G23303<= not G20785;
	G23304<= not G20785;
	G23305<= not G20391;
	G23306<= not G20924;
	G23307<= not G20924;
	G23308<= not G21024;
	G23312<= not G21070;
	G23313<= not G21070;
	G23320<= not I22419;
	G23321<= not I22422;
	G23322<= not I22425;
	G23323<= not G20283;
	G23331<= not G20905;
	G23332<= not G20785;
	G23333<= not G20785;
	G23334<= not G20785;
	G23335<= not G20391;
	G23336<= not G20924;
	G23337<= not G20924;
	G23338<= not G20453;
	G23339<= not G21070;
	G23340<= not G21070;
	G23341<= not G21163;
	G23347<= not I22444;
	G23350<= not G20785;
	G23351<= not G20924;
	G23352<= not G20924;
	G23353<= not G20924;
	G23354<= not G20453;
	G23355<= not G21070;
	G23356<= not G21070;
	G23359<= not I22458;
	G23360<= not I22461;
	G23361<= not I22464;
	G23362<= not I22467;
	G23363<= not I22470;
	G23375<= not G20924;
	G23376<= not G21070;
	G23377<= not G21070;
	G23378<= not G21070;
	G23380<= not G20619;
	G23382<= not G20682;
	G23384<= not I22485;
	G23385<= not I22488;
	G23388<= not G21070;
	G23390<= not G21468;
	G23391<= not G20645;
	G23393<= not G20739;
	G23394<= not I22499;
	G23395<= not I22502;
	G23398<= not G21468;
	G23399<= not G21514;
	G23400<= not G20676;
	G23402<= not G20875;
	G23403<= not I22512;
	G23406<= not G20330;
	G23408<= not G21468;
	G23409<= not G21514;
	G23410<= not G21562;
	G23411<= not G20734;
	G23413<= not G21012;
	G23414<= not I22525;
	G23417<= not G20391;
	G23418<= not G21468;
	G23419<= not G21468;
	G23420<= not G21514;
	G23421<= not G21562;
	G23422<= not G21611;
	G23423<= not G20871;
	G23425<= not G20751;
	G23426<= not I22539;
	G23427<= not I22542;
	G23429<= not G20453;
	G23430<= not I22547;
	G23431<= not G21514;
	G23432<= not G21514;
	G23433<= not G21562;
	G23434<= not G21611;
	G23435<= not G18833;
	G23440<= not I22557;
	G23443<= not G21468;
	G23444<= not I22561;
	G23445<= not I22564;
	G23446<= not G21562;
	G23447<= not G21562;
	G23448<= not G21611;
	G23449<= not G18833;
	G23450<= not I22571;
	G23452<= not G21468;
	G23453<= not I22576;
	G23456<= not G21514;
	G23457<= not I22580;
	G23458<= not I22583;
	G23459<= not G21611;
	G23460<= not G21611;
	G23461<= not G18833;
	G23462<= not I22589;
	G23472<= not G21062;
	G23473<= not G20785;
	G23476<= not G21468;
	G23477<= not G21468;
	G23478<= not G21514;
	G23479<= not G21562;
	G23480<= not I22601;
	G23481<= not I22604;
	G23482<= not G18833;
	G23483<= not G18833;
	G23485<= not G20785;
	G23486<= not G20785;
	G23487<= not G20924;
	G23488<= not G21468;
	G23489<= not G21468;
	G23490<= not G21514;
	G23491<= not G21514;
	G23492<= not G21562;
	G23493<= not G21611;
	G23494<= not I22619;
	G23495<= not I22622;
	G23496<= not G20248;
	G23499<= not G20785;
	G23500<= not G20924;
	G23501<= not G20924;
	G23502<= not G21070;
	G23503<= not G21468;
	G23504<= not G21468;
	G23505<= not G21514;
	G23506<= not G21514;
	G23507<= not G21562;
	G23508<= not G21562;
	G23509<= not G21611;
	G23510<= not G18833;
	G23511<= not I22640;
	G23512<= not G20248;
	G23515<= not G20785;
	G23516<= not G20924;
	G23517<= not G21070;
	G23518<= not G21070;
	G23519<= not G21468;
	G23520<= not G21468;
	G23521<= not G21468;
	G23522<= not G21514;
	G23523<= not G21514;
	G23524<= not G21562;
	G23525<= not G21562;
	G23526<= not G21611;
	G23527<= not G21611;
	G23528<= not G18833;
	G23529<= not G20558;
	G23530<= not G20248;
	G23534<= not I22665;
	G23537<= not G20785;
	G23538<= not G20924;
	G23539<= not G21070;
	G23541<= not G21514;
	G23542<= not G21514;
	G23543<= not G21514;
	G23544<= not G21562;
	G23545<= not G21562;
	G23546<= not G21611;
	G23547<= not G21611;
	G23548<= not G18833;
	G23549<= not G18833;
	G23550<= not G20248;
	G23555<= not I22692;
	G23558<= not G20924;
	G23559<= not G21070;
	G23563<= not G20682;
	G23565<= not G21562;
	G23566<= not G21562;
	G23567<= not G21562;
	G23568<= not G21611;
	G23569<= not G21611;
	G23570<= not G18833;
	G23571<= not G18833;
	G23573<= not G20248;
	G23578<= not I22725;
	G23582<= not I22729;
	G23585<= not G21070;
	G23589<= not G21468;
	G23605<= not G20739;
	G23607<= not G21611;
	G23608<= not G21611;
	G23609<= not G21611;
	G23610<= not G18833;
	G23611<= not G18833;
	G23612<= not I22745;
	G23613<= not I22748;
	G23614<= not G20248;
	G23620<= not I22769;
	G23629<= not G21514;
	G23645<= not G20875;
	G23647<= not G18833;
	G23648<= not G18833;
	G23649<= not G18833;
	G23650<= not G20653;
	G23651<= not G20655;
	G23652<= not I22785;
	G23653<= not I22788;
	G23654<= not G20248;
	G23665<= not G21562;
	G23681<= not G21012;
	G23683<= not I22816;
	G23684<= not I22819;
	G23698<= not G21611;
	G23714<= not G20751;
	G23715<= not G20764;
	G23732<= not G18833;
	G23745<= not G20900;
	G23746<= not G20902;
	G23749<= not G18997;
	G23759<= not I22886;
	G23760<= not I22889;
	G23764<= not G21308;
	G23767<= not G18997;
	G23768<= not G18997;
	G23769<= not G19074;
	G23776<= not G21177;
	G23777<= not I22918;
	G23787<= not G18997;
	G23788<= not G18997;
	G23789<= not G21308;
	G23792<= not G19074;
	G23793<= not G19074;
	G23794<= not G19147;
	G23800<= not G21246;
	G23812<= not G18997;
	G23813<= not G18997;
	G23814<= not G19074;
	G23815<= not G19074;
	G23816<= not G21308;
	G23819<= not G19147;
	G23820<= not G19147;
	G23821<= not G19210;
	G23823<= not I22989;
	G23824<= not G21271;
	G23838<= not G18997;
	G23839<= not G18997;
	G23840<= not G19074;
	G23841<= not G19074;
	G23842<= not G19147;
	G23843<= not G19147;
	G23844<= not G21308;
	G23847<= not G19210;
	G23848<= not G19210;
	G23849<= not G19277;
	G23858<= not G18997;
	G23859<= not G19074;
	G23860<= not G19074;
	G23861<= not G19147;
	G23862<= not G19147;
	G23863<= not G19210;
	G23864<= not G19210;
	G23865<= not G21308;
	G23868<= not G19277;
	G23869<= not G19277;
	G23870<= not G21293;
	G23874<= not G18997;
	G23875<= not G18997;
	G23876<= not G19074;
	G23877<= not G19147;
	G23878<= not G19147;
	G23879<= not G19210;
	G23880<= not G19210;
	G23881<= not G19277;
	G23882<= not G19277;
	G23886<= not G21468;
	G23887<= not G18997;
	G23888<= not G18997;
	G23889<= not G20682;
	G23893<= not G19074;
	G23894<= not G19074;
	G23895<= not G19147;
	G23896<= not G19210;
	G23897<= not G19210;
	G23898<= not G19277;
	G23899<= not G19277;
	G23902<= not G21468;
	G23903<= not G18997;
	G23904<= not G18997;
	G23905<= not G21514;
	G23906<= not G19074;
	G23907<= not G19074;
	G23908<= not G20739;
	G23912<= not G19147;
	G23913<= not G19147;
	G23914<= not G19210;
	G23915<= not G19277;
	G23916<= not G19277;
	G23922<= not G18997;
	G23923<= not G18997;
	G23924<= not G18997;
	G23925<= not G21514;
	G23926<= not G19074;
	G23927<= not G19074;
	G23928<= not G21562;
	G23929<= not G19147;
	G23930<= not G19147;
	G23931<= not G20875;
	G23935<= not G19210;
	G23936<= not G19210;
	G23937<= not G19277;
	G23938<= not G18997;
	G23939<= not G19074;
	G23940<= not G19074;
	G23941<= not G19074;
	G23942<= not G21562;
	G23943<= not G19147;
	G23944<= not G19147;
	G23945<= not G21611;
	G23946<= not G19210;
	G23947<= not G19210;
	G23948<= not G21012;
	G23952<= not G19277;
	G23953<= not G19277;
	G23954<= not I23099;
	G23961<= not G19074;
	G23962<= not G19147;
	G23963<= not G19147;
	G23964<= not G19147;
	G23965<= not G21611;
	G23966<= not G19210;
	G23967<= not G19210;
	G23968<= not G18833;
	G23969<= not G19277;
	G23970<= not G19277;
	G23971<= not G20751;
	G23982<= not G19147;
	G23983<= not G19210;
	G23984<= not G19210;
	G23985<= not G19210;
	G23986<= not G18833;
	G23987<= not G19277;
	G23988<= not G19277;
	G23992<= not G19210;
	G23993<= not G19277;
	G23994<= not G19277;
	G23995<= not G19277;
	G23999<= not G21468;
	G24000<= not G19277;
	G24003<= not G21514;
	G24005<= not I23149;
	G24010<= not G21562;
	G24013<= not G21611;
	G24017<= not G18833;
	G24019<= not G19968;
	G24020<= not G20014;
	G24021<= not G20841;
	G24022<= not G20982;
	G24023<= not G21127;
	G24024<= not G21193;
	G24025<= not G21256;
	G24026<= not G19919;
	G24027<= not G20014;
	G24028<= not G20841;
	G24029<= not G20982;
	G24030<= not G21127;
	G24031<= not G21193;
	G24032<= not G21256;
	G24033<= not G19919;
	G24034<= not G19968;
	G24035<= not G20841;
	G24036<= not G20982;
	G24037<= not G21127;
	G24038<= not G21193;
	G24039<= not G21256;
	G24040<= not G19919;
	G24041<= not G19968;
	G24042<= not G20014;
	G24043<= not G20982;
	G24044<= not G21127;
	G24045<= not G21193;
	G24046<= not G21256;
	G24047<= not G19919;
	G24048<= not G19968;
	G24049<= not G20014;
	G24050<= not G20841;
	G24051<= not G21127;
	G24052<= not G21193;
	G24053<= not G21256;
	G24054<= not G19919;
	G24055<= not G19968;
	G24056<= not G20014;
	G24057<= not G20841;
	G24058<= not G20982;
	G24059<= not G21193;
	G24060<= not G21256;
	G24061<= not G19919;
	G24062<= not G19968;
	G24063<= not G20014;
	G24064<= not G20841;
	G24065<= not G20982;
	G24066<= not G21127;
	G24067<= not G21256;
	G24068<= not G19919;
	G24069<= not G19968;
	G24070<= not G20014;
	G24071<= not G20841;
	G24072<= not G20982;
	G24073<= not G21127;
	G24074<= not G21193;
	G24075<= not G19935;
	G24076<= not G19984;
	G24077<= not G20720;
	G24078<= not G20857;
	G24079<= not G20998;
	G24080<= not G21143;
	G24081<= not G21209;
	G24082<= not G19890;
	G24083<= not G19984;
	G24084<= not G20720;
	G24085<= not G20857;
	G24086<= not G20998;
	G24087<= not G21143;
	G24088<= not G21209;
	G24089<= not G19890;
	G24090<= not G19935;
	G24091<= not G20720;
	G24092<= not G20857;
	G24093<= not G20998;
	G24094<= not G21143;
	G24095<= not G21209;
	G24096<= not G19890;
	G24097<= not G19935;
	G24098<= not G19984;
	G24099<= not G20720;
	G24100<= not G20857;
	G24101<= not G20998;
	G24102<= not G21143;
	G24103<= not G21209;
	G24104<= not G19890;
	G24105<= not G19935;
	G24106<= not G19984;
	G24107<= not G20857;
	G24108<= not G20998;
	G24109<= not G21143;
	G24110<= not G21209;
	G24111<= not G19890;
	G24112<= not G19935;
	G24113<= not G19984;
	G24114<= not G20720;
	G24115<= not G20998;
	G24116<= not G21143;
	G24117<= not G21209;
	G24118<= not G19890;
	G24119<= not G19935;
	G24120<= not G19984;
	G24121<= not G20720;
	G24122<= not G20857;
	G24123<= not G21143;
	G24124<= not G21209;
	G24125<= not G19890;
	G24126<= not G19935;
	G24127<= not G19984;
	G24128<= not G20720;
	G24129<= not G20857;
	G24130<= not G20998;
	G24131<= not G21209;
	G24132<= not G19890;
	G24133<= not G19935;
	G24134<= not G19984;
	G24135<= not G20720;
	G24136<= not G20857;
	G24137<= not G20998;
	G24138<= not G21143;
	G24146<= not G19422;
	G24147<= not G19402;
	G24149<= not G19338;
	G24150<= not G19268;
	G24152<= not I23300;
	G24153<= not I23303;
	G24154<= not I23306;
	G24155<= not I23309;
	G24156<= not I23312;
	G24157<= not I23315;
	G24158<= not I23318;
	G24159<= not I23321;
	G24160<= not I23324;
	G24161<= not I23327;
	G24162<= not I23330;
	G24163<= not I23333;
	G24164<= not I23336;
	G24165<= not I23339;
	G24166<= not I23342;
	G24167<= not I23345;
	G24168<= not I23348;
	G24169<= not I23351;
	G24170<= not I23354;
	G24171<= not I23357;
	G24172<= not I23360;
	G24173<= not I23363;
	G24174<= not I23366;
	G24175<= not I23369;
	G24176<= not I23372;
	G24177<= not I23375;
	G24178<= not I23378;
	G24179<= not I23381;
	G24180<= not I23384;
	G24181<= not I23387;
	G24182<= not I23390;
	G24183<= not I23393;
	G24184<= not I23396;
	G24185<= not I23399;
	G24356<= not G22594;
	G24357<= not G22325;
	G24358<= not G22550;
	G24359<= not G22550;
	G24360<= not G22228;
	G24361<= not G22885;
	G24364<= not G22722;
	G24365<= not G22594;
	G24366<= not G22594;
	G24367<= not G22550;
	G24368<= not G22228;
	G24372<= not G22885;
	G24373<= not G22908;
	G24375<= not G22722;
	G24376<= not G22722;
	G24377<= not G22594;
	G24379<= not G22550;
	G24384<= not G22885;
	G24385<= not G22908;
	G24386<= not G22594;
	G24388<= not G22885;
	G24389<= not G22908;
	G24394<= not G22228;
	G24396<= not G22885;
	G24397<= not G22908;
	G24404<= not G22908;
	G24405<= not G22722;
	G24407<= not G22594;
	G24417<= not G22171;
	G24418<= not G22722;
	G24419<= not G22722;
	G24424<= not G22722;
	G24425<= not G22722;
	G24426<= not G22722;
	G24428<= not G22722;
	G24429<= not G22722;
	G24431<= not G22722;
	G24437<= not G22654;
	G24438<= not G22722;
	G24452<= not G22722;
	G24463<= not G23578;
	G24466<= not I23671;
	G24474<= not G23620;
	G24477<= not I23680;
	G24481<= not I23684;
	G24483<= not I23688;
	G24489<= not I23694;
	G24490<= not G22594;
	G24505<= not G22689;
	G24506<= not I23711;
	G24509<= not G22689;
	G24515<= not G22689;
	G24516<= not G22670;
	G24522<= not G22689;
	G24524<= not G22876;
	G24525<= not G22670;
	G24526<= not G22942;
	G24527<= not G22670;
	G24533<= not G22876;
	G24534<= not G22670;
	G24535<= not G22942;
	G24540<= not G22942;
	G24548<= not G22942;
	G24560<= not G22942;
	G24568<= not G22942;
	G24571<= not G22942;
	G24579<= not G23067;
	G24585<= not G23063;
	G24586<= not G23067;
	G24587<= not G23112;
	G24603<= not G23108;
	G24604<= not G23112;
	G24605<= not G23139;
	G24623<= not G23076;
	G24625<= not G23135;
	G24626<= not G23139;
	G24636<= not G23121;
	G24648<= not G23148;
	G24655<= not G23067;
	G24665<= not G23067;
	G24667<= not G23112;
	G24683<= not G23112;
	G24685<= not G23139;
	G24699<= not G23047;
	G24711<= not G23139;
	G24718<= not G22182;
	G24732<= not G23042;
	G24744<= not G22202;
	G24756<= not G22763;
	G24759<= not G23003;
	G24770<= not G22763;
	G24778<= not G23286;
	G24789<= not G23309;
	G24791<= not G23850;
	G24795<= not G23342;
	G24818<= not G23191;
	G24819<= not I23998;
	G24825<= not G23204;
	G24836<= not I24008;
	G24839<= not G23436;
	G24850<= not I24022;
	G24866<= not I24038;
	G24869<= not I24041;
	G24891<= not G23231;
	G24893<= not I24060;
	G24911<= not I24078;
	G24920<= not I24089;
	G24960<= not G23716;
	G24963<= not G22342;
	G24964<= not I24128;
	G24966<= not G22763;
	G24971<= not G23590;
	G24978<= not G22342;
	G24979<= not G22369;
	G24980<= not G22384;
	G24981<= not G22763;
	G24982<= not G22763;
	G24985<= not G23586;
	G24986<= not G23590;
	G24987<= not G23630;
	G24991<= not G22369;
	G24992<= not G22417;
	G24993<= not G22384;
	G24994<= not G22432;
	G24995<= not G22763;
	G24996<= not G22763;
	G24999<= not G23626;
	G25000<= not G23630;
	G25001<= not G23666;
	G25006<= not G22417;
	G25007<= not G22457;
	G25008<= not G22432;
	G25009<= not G22472;
	G25011<= not G22763;
	G25013<= not G23599;
	G25015<= not G23662;
	G25016<= not G23666;
	G25017<= not G23699;
	G25023<= not G22457;
	G25024<= not G22472;
	G25025<= not G22498;
	G25027<= not I24191;
	G25032<= not G23639;
	G25034<= not G23695;
	G25035<= not G23699;
	G25036<= not G23733;
	G25039<= not G22498;
	G25044<= not G23675;
	G25046<= not G23729;
	G25047<= not G23733;
	G25051<= not I24215;
	G25055<= not G23590;
	G25060<= not G23708;
	G25064<= not I24228;
	G25070<= not G23590;
	G25072<= not G23630;
	G25073<= not I24237;
	G25080<= not G23742;
	G25081<= not G22342;
	G25082<= not G22342;
	G25083<= not G23782;
	G25090<= not G23630;
	G25092<= not G23666;
	G25097<= not G22342;
	G25098<= not G22369;
	G25099<= not G22369;
	G25100<= not G22384;
	G25101<= not G22384;
	G25109<= not G23666;
	G25111<= not G23699;
	G25114<= not I24278;
	G25115<= not I24281;
	G25116<= not G22369;
	G25117<= not G22417;
	G25118<= not G22417;
	G25119<= not G22384;
	G25120<= not G22432;
	G25121<= not G22432;
	G25131<= not G23699;
	G25133<= not G23733;
	G25134<= not G22417;
	G25135<= not G22457;
	G25136<= not G22457;
	G25137<= not G22432;
	G25138<= not G22472;
	G25139<= not G22472;
	G25140<= not G22228;
	G25153<= not G23733;
	G25154<= not G22457;
	G25155<= not G22472;
	G25156<= not G22498;
	G25157<= not G22498;
	G25158<= not G22228;
	G25167<= not I24331;
	G25168<= not I24334;
	G25169<= not G22763;
	G25170<= not G22498;
	G25171<= not G22228;
	G25174<= not G23890;
	G25180<= not G23529;
	G25182<= not G22763;
	G25183<= not G22763;
	G25184<= not G22763;
	G25185<= not G22228;
	G25188<= not G23909;
	G25193<= not G22763;
	G25194<= not G22763;
	G25195<= not G22763;
	G25196<= not G22763;
	G25197<= not G23958;
	G25198<= not G22228;
	G25202<= not G23932;
	G25206<= not G23613;
	G25208<= not G22763;
	G25209<= not G22763;
	G25210<= not G23802;
	G25211<= not G22763;
	G25212<= not G22763;
	G25213<= not G23293;
	G25214<= not G22228;
	G25218<= not G23949;
	G25219<= not I24393;
	G25220<= not I24396;
	G25221<= not G23653;
	G25222<= not I24400;
	G25224<= not G22763;
	G25225<= not G23802;
	G25226<= not G22763;
	G25227<= not G22763;
	G25228<= not G23828;
	G25230<= not G23314;
	G25231<= not G22228;
	G25232<= not G22228;
	G25239<= not G23972;
	G25240<= not G23650;
	G25241<= not G23651;
	G25242<= not G23684;
	G25243<= not G22763;
	G25244<= not G23802;
	G25245<= not G22763;
	G25246<= not G23828;
	G25248<= not G22228;
	G25249<= not G22228;
	G25250<= not I24434;
	G25259<= not I24445;
	G25260<= not I24448;
	G25262<= not G22763;
	G25263<= not G22763;
	G25264<= not G23828;
	G25265<= not I24455;
	G25266<= not G22228;
	G25267<= not G22228;
	G25272<= not G23715;
	G25273<= not G23978;
	G25274<= not G22763;
	G25282<= not G22763;
	G25283<= not G22763;
	G25284<= not I24474;
	G25286<= not G22228;
	G25287<= not G22228;
	G25288<= not G22228;
	G25289<= not G22228;
	G25296<= not G23745;
	G25297<= not G23746;
	G25298<= not G23760;
	G25299<= not G22763;
	G25307<= not G22763;
	G25308<= not G22763;
	G25316<= not G22763;
	G25322<= not I24497;
	G25324<= not G22228;
	G25325<= not G22228;
	G25326<= not G22228;
	G25327<= not G22161;
	G25340<= not G22763;
	G25348<= not G22763;
	G25356<= not G22763;
	G25369<= not G22228;
	G25370<= not G22228;
	G25380<= not G23776;
	G25388<= not G22763;
	G25399<= not G22763;
	G25409<= not G22228;
	G25410<= not G22228;
	G25423<= not I24558;
	G25424<= not G23800;
	G25438<= not G22763;
	G25451<= not G22228;
	G25452<= not G22228;
	G25465<= not G23824;
	G25480<= not G22228;
	G25481<= not G22228;
	G25505<= not G22228;
	G25506<= not G22228;
	G25513<= not G23870;
	G25517<= not G22228;
	G25523<= not G22550;
	G25524<= not G22228;
	G25525<= not G22550;
	G25528<= not G22594;
	G25529<= not G22763;
	G25533<= not G22550;
	G25534<= not G22763;
	G25535<= not G22763;
	G25538<= not G22594;
	G25541<= not G22763;
	G25542<= not G22763;
	G25544<= not G22594;
	G25546<= not G22550;
	G25547<= not G22550;
	G25548<= not G22550;
	G25549<= not G22763;
	G25550<= not G22763;
	G25552<= not G22594;
	G25553<= not G22550;
	G25554<= not G22550;
	G25555<= not G22550;
	G25556<= not G22763;
	G25557<= not G22763;
	G25558<= not G22594;
	G25560<= not G22550;
	G25561<= not G22550;
	G25562<= not G22763;
	G25563<= not G22594;
	G25564<= not G22312;
	G25566<= not G22550;
	G25620<= not I24759;
	G25640<= not I24781;
	G25641<= not I24784;
	G25642<= not I24787;
	G25692<= not I24839;
	G25766<= not G24439;
	G25771<= not I24920;
	G25773<= not G24453;
	G25781<= not G24510;
	G25783<= not G25250;
	G25786<= not G24518;
	G25790<= not G25027;
	G25820<= not G25051;
	G25830<= not G24485;
	G25837<= not G25064;
	G25838<= not G25250;
	G25849<= not G24491;
	G25869<= not G25250;
	G25882<= not G25026;
	G25886<= not G24537;
	G25892<= not G24528;
	G25893<= not G24541;
	G25899<= not G24997;
	G25903<= not I25005;
	G25930<= not I25028;
	G25994<= not G24575;
	G25997<= not I25095;
	G26026<= not I25105;
	G26054<= not G24804;
	G26055<= not I25115;
	G26081<= not G24619;
	G26083<= not G24809;
	G26093<= not G24814;
	G26105<= not I25146;
	G26131<= not I25161;
	G26187<= not I25190;
	G26260<= not G24759;
	G26284<= not G24875;
	G26326<= not G24872;
	G26337<= not G24818;
	G26340<= not G24953;
	G26364<= not I25327;
	G26400<= not I25351;
	G26424<= not I25356;
	G26483<= not I25359;
	G26488<= not I25366;
	G26510<= not I25369;
	G26518<= not G25233;
	G26519<= not I25380;
	G26548<= not G25255;
	G26549<= not I25391;
	G26575<= not G25268;
	G26576<= not I25399;
	G26605<= not G25293;
	G26607<= not G25382;
	G26608<= not G25334;
	G26614<= not G25426;
	G26615<= not G25432;
	G26631<= not G25467;
	G26632<= not G25473;
	G26634<= not G25317;
	G26648<= not G25115;
	G26653<= not G25337;
	G26654<= not G25275;
	G26655<= not G25492;
	G26656<= not G25495;
	G26672<= not G25275;
	G26679<= not G25385;
	G26680<= not G25300;
	G26681<= not G25396;
	G26682<= not G25309;
	G26683<= not G25514;
	G26693<= not G25300;
	G26700<= not G25429;
	G26701<= not G25341;
	G26702<= not G25309;
	G26709<= not G25435;
	G26710<= not G25349;
	G26718<= not G25168;
	G26720<= not G25275;
	G26724<= not G25341;
	G26731<= not G25470;
	G26732<= not G25389;
	G26736<= not G25349;
	G26743<= not G25476;
	G26744<= not G25400;
	G26754<= not G25300;
	G26758<= not G25389;
	G26765<= not G25309;
	G26769<= not G25400;
	G26776<= not G25498;
	G26777<= not G25439;
	G26784<= not G25341;
	G26788<= not G25349;
	G26792<= not G25439;
	G26801<= not I25511;
	G26802<= not I25514;
	G26803<= not G25389;
	G26804<= not G25400;
	G26810<= not G25220;
	G26811<= not G25206;
	G26812<= not G25439;
	G26814<= not G25221;
	G26816<= not G25260;
	G26817<= not G25242;
	G26818<= not I25530;
	G26820<= not I25534;
	G26824<= not G25298;
	G26825<= not I25541;
	G26827<= not G24819;
	G26830<= not G24411;
	G26831<= not G24836;
	G26832<= not G24850;
	G26834<= not I25552;
	G26835<= not I25555;
	G26836<= not G24866;
	G26837<= not G24869;
	G26840<= not I25562;
	G26841<= not G24893;
	G26843<= not I25567;
	G26850<= not I25576;
	G26851<= not I25579;
	G26856<= not I25586;
	G26859<= not I25591;
	G26860<= not I25594;
	G26862<= not I25598;
	G26869<= not G24842;
	G26870<= not I25606;
	G26935<= not I25677;
	G26936<= not I25680;
	G26937<= not I25683;
	G26941<= not I25689;
	G26942<= not I25692;
	G26943<= not I25695;
	G26973<= not G26105;
	G26987<= not G26131;
	G26990<= not G26105;
	G27004<= not G26131;
	G27009<= not G25911;
	G27011<= not G25917;
	G27013<= not I25743;
	G27014<= not G25888;
	G27015<= not G26869;
	G27017<= not G25895;
	G27018<= not I25750;
	G27038<= not G25932;
	G27051<= not I25779;
	G27064<= not I25786;
	G27074<= not I25790;
	G27084<= not G26673;
	G27088<= not G26694;
	G27089<= not G26703;
	G27091<= not G26725;
	G27092<= not G26737;
	G27100<= not G26759;
	G27101<= not G26770;
	G27112<= not G26793;
	G27142<= not G26105;
	G27155<= not G26131;
	G27163<= not I25869;
	G27187<= not I25882;
	G27237<= not G26162;
	G27242<= not G26183;
	G27245<= not G26209;
	G27279<= not G26330;
	G27320<= not I26004;
	G27349<= not G26352;
	G27402<= not I26100;
	G27415<= not G26382;
	G27438<= not I26130;
	G27492<= not G26598;
	G27527<= not I26195;
	G27554<= not G26625;
	G27565<= not G26645;
	G27573<= not G26667;
	G27576<= not G26081;
	G27583<= not G26686;
	G27585<= not G25994;
	G27592<= not G26715;
	G27597<= not G26745;
	G27662<= not I26296;
	G27675<= not I26309;
	G27698<= not G26648;
	G27708<= not I26334;
	G27709<= not I26337;
	G27730<= not G26424;
	G27736<= not I26356;
	G27737<= not G26718;
	G27773<= not I26378;
	G27774<= not I26381;
	G27830<= not G26802;
	G27831<= not I26406;
	G27832<= not I26409;
	G27880<= not I26427;
	G27881<= not I26430;
	G27928<= not G26810;
	G27929<= not I26448;
	G27930<= not I26451;
	G27956<= not I26466;
	G27961<= not G26816;
	G27967<= not I26479;
	G27971<= not G26673;
	G27975<= not G26694;
	G27976<= not G26703;
	G27977<= not G26105;
	G27983<= not G26725;
	G27984<= not G26737;
	G27985<= not G26131;
	G27989<= not G26759;
	G27990<= not G26770;
	G27991<= not G25852;
	G27993<= not I26503;
	G27994<= not G26793;
	G27996<= not I26508;
	G27998<= not I26512;
	G28009<= not I26516;
	G28032<= not G26365;
	G28033<= not G26365;
	G28034<= not G26365;
	G28036<= not G26365;
	G28037<= not G26365;
	G28038<= not G26365;
	G28039<= not G26365;
	G28040<= not G26365;
	G28079<= not I26578;
	G28080<= not I26581;
	G28081<= not I26584;
	G28119<= not G27008;
	G28120<= not G27108;
	G28121<= not G27093;
	G28126<= not G27122;
	G28127<= not G27102;
	G28137<= not I26638;
	G28142<= not I26649;
	G28147<= not I26654;
	G28155<= not I26664;
	G28156<= not I26667;
	G28157<= not I26670;
	G28161<= not I26676;
	G28162<= not I26679;
	G28163<= not I26682;
	G28166<= not I26687;
	G28173<= not I26693;
	G28181<= not I26700;
	G28184<= not I26705;
	G28187<= not I26710;
	G28241<= not G27064;
	G28250<= not G27074;
	G28262<= not I26785;
	G28274<= not I26799;
	G28294<= not G27295;
	G28307<= not G27306;
	G28321<= not G27317;
	G28325<= not G27463;
	G28326<= not G27414;
	G28367<= not I26880;
	G28370<= not G27528;
	G28380<= not G27064;
	G28399<= not G27074;
	G28431<= not I26925;
	G28436<= not I26929;
	G28441<= not G27629;
	G28443<= not I26936;
	G28463<= not I26952;
	G28479<= not G27654;
	G28508<= not I26989;
	G28559<= not G27700;
	G28575<= not G27711;
	G28579<= not G27714;
	G28590<= not G27724;
	G28593<= not G27727;
	G28598<= not G27717;
	G28604<= not G27759;
	G28606<= not G27762;
	G28608<= not G27670;
	G28615<= not G27817;
	G28620<= not G27679;
	G28633<= not G27687;
	G28648<= not G27693;
	G28656<= not G27742;
	G28669<= not G27705;
	G28675<= not G27779;
	G28678<= not G27800;
	G28693<= not G27837;
	G28696<= not G27858;
	G28709<= not I27192;
	G28711<= not G27886;
	G28713<= not G27907;
	G28726<= not G27937;
	G28752<= not I27232;
	G28753<= not I27235;
	G28754<= not I27238;
	G28779<= not I27253;
	G28819<= not I27271;
	G28917<= not I27314;
	G28918<= not G27832;
	G28954<= not G27830;
	G29013<= not I27368;
	G29014<= not G27742;
	G29041<= not I27385;
	G29042<= not I27388;
	G29043<= not I27391;
	G29044<= not G27742;
	G29045<= not G27779;
	G29056<= not G27800;
	G29067<= not I27401;
	G29079<= not G27742;
	G29080<= not G27779;
	G29081<= not G27837;
	G29092<= not G27800;
	G29093<= not G27858;
	G29115<= not G27779;
	G29116<= not G27837;
	G29117<= not G27886;
	G29128<= not G27800;
	G29129<= not G27858;
	G29130<= not G27907;
	G29147<= not I27449;
	G29149<= not G27837;
	G29150<= not G27886;
	G29151<= not G27858;
	G29152<= not G27907;
	G29153<= not G27937;
	G29169<= not G27886;
	G29170<= not G27907;
	G29171<= not G27937;
	G29172<= not G27020;
	G29177<= not G27937;
	G29185<= not I27481;
	G29190<= not G27046;
	G29194<= not I27492;
	G29195<= not I27495;
	G29196<= not G27059;
	G29209<= not I27543;
	G29210<= not I27546;
	G29211<= not I27549;
	G29212<= not I27552;
	G29213<= not I27555;
	G29214<= not I27558;
	G29215<= not I27561;
	G29216<= not I27564;
	G29217<= not I27567;
	G29218<= not I27570;
	G29219<= not I27573;
	G29220<= not I27576;
	G29221<= not I27579;
	G29310<= not G28991;
	G29311<= not G28998;
	G29312<= not G28877;
	G29317<= not I27677;
	G29318<= not G29029;
	G29333<= not G28167;
	G29339<= not G28274;
	G29342<= not G28188;
	G29343<= not G28174;
	G29348<= not G28194;
	G29353<= not I27713;
	G29358<= not I27718;
	G29365<= not G29067;
	G29368<= not I27730;
	G29371<= not I27735;
	G29372<= not I27738;
	G29374<= not I27742;
	G29379<= not I27749;
	G29385<= not G28180;
	G29474<= not I27758;
	G29491<= not I27777;
	G29498<= not I27784;
	G29505<= not G29186;
	G29507<= not G28353;
	G29597<= not G28444;
	G29653<= not I27927;
	G29669<= not I27941;
	G29689<= not I27954;
	G29697<= not G28336;
	G29707<= not G28504;
	G29713<= not I27970;
	G29725<= not G28349;
	G29744<= not G28431;
	G29745<= not G28500;
	G29755<= not I28002;
	G29765<= not I28014;
	G29800<= not G28363;
	G29811<= not G28376;
	G29812<= not G28381;
	G29814<= not I28062;
	G29846<= not G28391;
	G29847<= not G28395;
	G29862<= not G28406;
	G29863<= not G28410;
	G29878<= not G28421;
	G29893<= not G28755;
	G29897<= not I28128;
	G29905<= not G28783;
	G29906<= not G28793;
	G29911<= not G28780;
	G29912<= not G28827;
	G29913<= not G28840;
	G29920<= not G28824;
	G29921<= not G28864;
	G29922<= not G28837;
	G29923<= not G28874;
	G29925<= not G28820;
	G29927<= not G28861;
	G29928<= not G28871;
	G29929<= not G28914;
	G29930<= not I28162;
	G29939<= not G28857;
	G29941<= not G28900;
	G29942<= not G28867;
	G29944<= not G28911;
	G29945<= not I28174;
	G29948<= not G28853;
	G29950<= not G28896;
	G29953<= not G28907;
	G29955<= not G28950;
	G29956<= not I28185;
	G29960<= not G28885;
	G29961<= not G28892;
	G29963<= not G28931;
	G29965<= not G28903;
	G29967<= not G28946;
	G29970<= not I28199;
	G29976<= not G29018;
	G29977<= not G28920;
	G29978<= not G28927;
	G29980<= not G28935;
	G29981<= not G28942;
	G29983<= not G28977;
	G29993<= not G29018;
	G29994<= not G29049;
	G29995<= not G28955;
	G29996<= not G28962;
	G29997<= not G29060;
	G29998<= not G28966;
	G29999<= not G28973;
	G30012<= not I28241;
	G30016<= not G29049;
	G30017<= not G29085;
	G30018<= not G28987;
	G30019<= not G29060;
	G30020<= not G29097;
	G30021<= not G28994;
	G30022<= not G29001;
	G30036<= not G29085;
	G30037<= not G29121;
	G30038<= not G29097;
	G30039<= not G29134;
	G30040<= not G29025;
	G30052<= not G29018;
	G30053<= not G29121;
	G30054<= not G29134;
	G30055<= not G29157;
	G30063<= not G29015;
	G30065<= not G29049;
	G30067<= not G29060;
	G30068<= not G29157;
	G30072<= not I28301;
	G30074<= not G29046;
	G30076<= not G29085;
	G30077<= not G29057;
	G30079<= not G29097;
	G30085<= not G29082;
	G30087<= not G29121;
	G30088<= not G29094;
	G30090<= not G29134;
	G30097<= not G29118;
	G30100<= not G29131;
	G30102<= not G29157;
	G30105<= not I28336;
	G30113<= not G29154;
	G30116<= not I28349;
	G30142<= not G28754;
	G30155<= not I28390;
	G30182<= not I28419;
	G30184<= not G28144;
	G30195<= not I28434;
	G30206<= not G28436;
	G30217<= not I28458;
	G30218<= not G28918;
	G30237<= not I28480;
	G30259<= not G28463;
	G30292<= not G28736;
	G30295<= not I28540;
	G30296<= not G28889;
	G30297<= not G28758;
	G30299<= not G28765;
	G30301<= not I28548;
	G30302<= not G28924;
	G30303<= not G28786;
	G30305<= not G28939;
	G30306<= not G28796;
	G30309<= not G28959;
	G30310<= not G28830;
	G30312<= not G28970;
	G30313<= not G28843;
	G30318<= not G28274;
	G30321<= not I28572;
	G30322<= not G28431;
	G30325<= not I28576;
	G30326<= not I28579;
	G30327<= not I28582;
	G30328<= not I28585;
	G30329<= not I28588;
	G30330<= not I28591;
	G30331<= not I28594;
	G30332<= not I28597;
	G30565<= not I28832;
	G30567<= not G29930;
	G30568<= not G29339;
	G30569<= not I28838;
	G30572<= not G29945;
	G30578<= not G29956;
	G30591<= not I28851;
	G30593<= not G29970;
	G30606<= not I28866;
	G30610<= not I28872;
	G30729<= not I28883;
	G30917<= not I28897;
	G30928<= not I28908;
	G30931<= not I28913;
	G30983<= not G29657;
	G30989<= not G29672;
	G30990<= not G29676;
	G30991<= not I28925;
	G30996<= not G29694;
	G30997<= not G29702;
	G30998<= not G29719;
	G30999<= not G29722;
	G31000<= not G29737;
	G31013<= not G29679;
	G31138<= not G29778;
	G31189<= not I29002;
	G31213<= not I29013;
	G31227<= not G29744;
	G31239<= not G29916;
	G31243<= not G29933;
	G31479<= not I29139;
	G31487<= not I29149;
	G31521<= not I29182;
	G31522<= not I29185;
	G31578<= not I29199;
	G31596<= not I29204;
	G31601<= not I29207;
	G31608<= not G29653;
	G31609<= not I29211;
	G31616<= not I29214;
	G31623<= not G29669;
	G31624<= not I29218;
	G31631<= not I29221;
	G31638<= not G29689;
	G31639<= not I29225;
	G31646<= not I29228;
	G31653<= not G29713;
	G31655<= not I29233;
	G31656<= not I29236;
	G31657<= not I29239;
	G31658<= not I29242;
	G31665<= not I29245;
	G31666<= not I29248;
	G31667<= not G30142;
	G31771<= not I29337;
	G31791<= not I29363;
	G31794<= not I29368;
	G31795<= not I29371;
	G31796<= not G29385;
	G31797<= not G29385;
	G31798<= not G29385;
	G31799<= not G29385;
	G31800<= not G29385;
	G31801<= not G29385;
	G31802<= not G29385;
	G31803<= not G29385;
	G31804<= not G29385;
	G31805<= not G29385;
	G31806<= not G29385;
	G31807<= not G29385;
	G31808<= not G29385;
	G31809<= not G29385;
	G31810<= not G29385;
	G31811<= not G29385;
	G31812<= not G29385;
	G31813<= not G29385;
	G31814<= not G29385;
	G31815<= not G29385;
	G31816<= not G29385;
	G31817<= not G29385;
	G31818<= not G29385;
	G31819<= not G29385;
	G31820<= not G29385;
	G31821<= not G29385;
	G31822<= not G29385;
	G31823<= not G29385;
	G31824<= not G29385;
	G31825<= not G29385;
	G31826<= not G29385;
	G31827<= not G29385;
	G31828<= not G29385;
	G31829<= not G29385;
	G31830<= not G29385;
	G31831<= not G29385;
	G31832<= not G29385;
	G31833<= not G29385;
	G31834<= not G29385;
	G31835<= not G29385;
	G31836<= not G29385;
	G31837<= not G29385;
	G31838<= not G29385;
	G31839<= not G29385;
	G31840<= not G29385;
	G31841<= not G29385;
	G31842<= not G29385;
	G31843<= not G29385;
	G31844<= not G29385;
	G31845<= not G29385;
	G31846<= not G29385;
	G31847<= not G29385;
	G31848<= not G29385;
	G31849<= not G29385;
	G31850<= not G29385;
	G31851<= not G29385;
	G31852<= not G29385;
	G31853<= not G29385;
	G31854<= not G29385;
	G31855<= not G29385;
	G31856<= not G29385;
	G31857<= not G29385;
	G31858<= not G29385;
	G31859<= not G29385;
	G31860<= not I29438;
	G31861<= not I29441;
	G31862<= not I29444;
	G31863<= not I29447;
	G31937<= not G30991;
	G31945<= not G31189;
	G32015<= not I29571;
	G32021<= not I29579;
	G32024<= not I29582;
	G32027<= not I29585;
	G32033<= not G30929;
	G32038<= not G30934;
	G32090<= not G31003;
	G32099<= not G31009;
	G32118<= not G31008;
	G32137<= not G31134;
	G32138<= not G31233;
	G32185<= not I29717;
	G32186<= not I29720;
	G32192<= not G31262;
	G32201<= not G31509;
	G32318<= not G31596;
	G32329<= not G31522;
	G32363<= not I29891;
	G32364<= not I29894;
	G32377<= not G30984;
	G32381<= not I29909;
	G32382<= not G31657;
	G32383<= not I29913;
	G32384<= not G31666;
	G32393<= not G30922;
	G32394<= not G30601;
	G32404<= not I29936;
	G32407<= not I29939;
	G32415<= not G31591;
	G32421<= not G31213;
	G32430<= not G30984;
	G32433<= not I29961;
	G32434<= not G31189;
	G32437<= not I29965;
	G32438<= not G30991;
	G32441<= not I29969;
	G32442<= not G31213;
	G32445<= not I29973;
	G32446<= not G31596;
	G32449<= not I29977;
	G32450<= not G31591;
	G32453<= not I29981;
	G32456<= not G31376;
	G32457<= not G30735;
	G32458<= not G30825;
	G32459<= not G31070;
	G32460<= not G31194;
	G32461<= not G30614;
	G32462<= not G30673;
	G32463<= not G31566;
	G32464<= not G30735;
	G32465<= not G30825;
	G32466<= not G31070;
	G32467<= not G31194;
	G32468<= not G30614;
	G32469<= not G30673;
	G32470<= not G31566;
	G32471<= not G31376;
	G32472<= not G30825;
	G32473<= not G31070;
	G32474<= not G31194;
	G32475<= not G30614;
	G32476<= not G30673;
	G32477<= not G31566;
	G32478<= not G31376;
	G32479<= not G30735;
	G32480<= not G31070;
	G32481<= not G31194;
	G32482<= not G30614;
	G32483<= not G30673;
	G32484<= not G31566;
	G32485<= not G31376;
	G32486<= not G30735;
	G32487<= not G30825;
	G32488<= not G31194;
	G32489<= not G30614;
	G32490<= not G30673;
	G32491<= not G31566;
	G32492<= not G31376;
	G32493<= not G30735;
	G32494<= not G30825;
	G32495<= not G31070;
	G32496<= not G30614;
	G32497<= not G30673;
	G32498<= not G31566;
	G32499<= not G31376;
	G32500<= not G30735;
	G32501<= not G30825;
	G32502<= not G31070;
	G32503<= not G31194;
	G32504<= not G30673;
	G32505<= not G31566;
	G32506<= not G31376;
	G32507<= not G30735;
	G32508<= not G30825;
	G32509<= not G31070;
	G32510<= not G31194;
	G32511<= not G30614;
	G32512<= not G31566;
	G32513<= not G31376;
	G32514<= not G30735;
	G32515<= not G30825;
	G32516<= not G31070;
	G32517<= not G31194;
	G32518<= not G30614;
	G32519<= not G30673;
	G32521<= not G31376;
	G32522<= not G30735;
	G32523<= not G30825;
	G32524<= not G31070;
	G32525<= not G31170;
	G32526<= not G30614;
	G32527<= not G30673;
	G32528<= not G31554;
	G32529<= not G30735;
	G32530<= not G30825;
	G32531<= not G31070;
	G32532<= not G31170;
	G32533<= not G30614;
	G32534<= not G30673;
	G32535<= not G31554;
	G32536<= not G31376;
	G32537<= not G30825;
	G32538<= not G31070;
	G32539<= not G31170;
	G32540<= not G30614;
	G32541<= not G30673;
	G32542<= not G31554;
	G32543<= not G31376;
	G32544<= not G30735;
	G32545<= not G31070;
	G32546<= not G31170;
	G32547<= not G30614;
	G32548<= not G30673;
	G32549<= not G31554;
	G32550<= not G31376;
	G32551<= not G30735;
	G32552<= not G30825;
	G32553<= not G31170;
	G32554<= not G30614;
	G32555<= not G30673;
	G32556<= not G31554;
	G32557<= not G31376;
	G32558<= not G30735;
	G32559<= not G30825;
	G32560<= not G31070;
	G32561<= not G30614;
	G32562<= not G30673;
	G32563<= not G31554;
	G32564<= not G31376;
	G32565<= not G30735;
	G32566<= not G30825;
	G32567<= not G31070;
	G32568<= not G31170;
	G32569<= not G30673;
	G32570<= not G31554;
	G32571<= not G31376;
	G32572<= not G30735;
	G32573<= not G30825;
	G32574<= not G31070;
	G32575<= not G31170;
	G32576<= not G30614;
	G32577<= not G31554;
	G32578<= not G31376;
	G32579<= not G30735;
	G32580<= not G30825;
	G32581<= not G31070;
	G32582<= not G31170;
	G32583<= not G30614;
	G32584<= not G30673;
	G32586<= not G31376;
	G32587<= not G30735;
	G32588<= not G30825;
	G32589<= not G31070;
	G32590<= not G31154;
	G32591<= not G30614;
	G32592<= not G30673;
	G32593<= not G31542;
	G32594<= not G30735;
	G32595<= not G30825;
	G32596<= not G31070;
	G32597<= not G31154;
	G32598<= not G30614;
	G32599<= not G30673;
	G32600<= not G31542;
	G32601<= not G31376;
	G32602<= not G30825;
	G32603<= not G31070;
	G32604<= not G31154;
	G32605<= not G30614;
	G32606<= not G30673;
	G32607<= not G31542;
	G32608<= not G31376;
	G32609<= not G30735;
	G32610<= not G31070;
	G32611<= not G31154;
	G32612<= not G30614;
	G32613<= not G30673;
	G32614<= not G31542;
	G32615<= not G31376;
	G32616<= not G30735;
	G32617<= not G30825;
	G32618<= not G31154;
	G32619<= not G30614;
	G32620<= not G30673;
	G32621<= not G31542;
	G32622<= not G31376;
	G32623<= not G30735;
	G32624<= not G30825;
	G32625<= not G31070;
	G32626<= not G30614;
	G32627<= not G30673;
	G32628<= not G31542;
	G32629<= not G31376;
	G32630<= not G30735;
	G32631<= not G30825;
	G32632<= not G31070;
	G32633<= not G31154;
	G32634<= not G30673;
	G32635<= not G31542;
	G32636<= not G31376;
	G32637<= not G30735;
	G32638<= not G30825;
	G32639<= not G31070;
	G32640<= not G31154;
	G32641<= not G30614;
	G32642<= not G31542;
	G32643<= not G31376;
	G32644<= not G30735;
	G32645<= not G30825;
	G32646<= not G31070;
	G32647<= not G31154;
	G32648<= not G30614;
	G32649<= not G30673;
	G32651<= not G31376;
	G32652<= not G30735;
	G32653<= not G30825;
	G32654<= not G31070;
	G32655<= not G30614;
	G32656<= not G30673;
	G32657<= not G31528;
	G32658<= not G31579;
	G32659<= not G30735;
	G32660<= not G30825;
	G32661<= not G31070;
	G32662<= not G30614;
	G32663<= not G30673;
	G32664<= not G31528;
	G32665<= not G31579;
	G32666<= not G31376;
	G32667<= not G30825;
	G32668<= not G31070;
	G32669<= not G30614;
	G32670<= not G30673;
	G32671<= not G31528;
	G32672<= not G31579;
	G32673<= not G31376;
	G32674<= not G30735;
	G32675<= not G31070;
	G32676<= not G30614;
	G32677<= not G30673;
	G32678<= not G31528;
	G32679<= not G31579;
	G32680<= not G31376;
	G32681<= not G30735;
	G32682<= not G30825;
	G32683<= not G30614;
	G32684<= not G30673;
	G32685<= not G31528;
	G32686<= not G31579;
	G32687<= not G31376;
	G32688<= not G30735;
	G32689<= not G30825;
	G32690<= not G31070;
	G32691<= not G30673;
	G32692<= not G31528;
	G32693<= not G31579;
	G32694<= not G31376;
	G32695<= not G30735;
	G32696<= not G30825;
	G32697<= not G31070;
	G32698<= not G30614;
	G32699<= not G31528;
	G32700<= not G31579;
	G32701<= not G31376;
	G32702<= not G30735;
	G32703<= not G30825;
	G32704<= not G31070;
	G32705<= not G30614;
	G32706<= not G30673;
	G32707<= not G31579;
	G32708<= not G31376;
	G32709<= not G30735;
	G32710<= not G30825;
	G32711<= not G31070;
	G32712<= not G30614;
	G32713<= not G30673;
	G32714<= not G31528;
	G32716<= not G31376;
	G32717<= not G30735;
	G32718<= not G30825;
	G32719<= not G31672;
	G32720<= not G31710;
	G32721<= not G31021;
	G32722<= not G30937;
	G32723<= not G31327;
	G32724<= not G30735;
	G32725<= not G30825;
	G32726<= not G31672;
	G32727<= not G31710;
	G32728<= not G31021;
	G32729<= not G30937;
	G32730<= not G31327;
	G32731<= not G31376;
	G32732<= not G30825;
	G32733<= not G31672;
	G32734<= not G31710;
	G32735<= not G31021;
	G32736<= not G30937;
	G32737<= not G31327;
	G32738<= not G31376;
	G32739<= not G30735;
	G32740<= not G31672;
	G32741<= not G31710;
	G32742<= not G31021;
	G32743<= not G30937;
	G32744<= not G31327;
	G32745<= not G31376;
	G32746<= not G30735;
	G32747<= not G30825;
	G32748<= not G31710;
	G32749<= not G31021;
	G32750<= not G30937;
	G32751<= not G31327;
	G32752<= not G31376;
	G32753<= not G30735;
	G32754<= not G30825;
	G32755<= not G31672;
	G32756<= not G31021;
	G32757<= not G30937;
	G32758<= not G31327;
	G32759<= not G31376;
	G32760<= not G30735;
	G32761<= not G30825;
	G32762<= not G31672;
	G32763<= not G31710;
	G32764<= not G30937;
	G32765<= not G31327;
	G32766<= not G31376;
	G32767<= not G30735;
	G32768<= not G30825;
	G32769<= not G31672;
	G32770<= not G31710;
	G32771<= not G31021;
	G32772<= not G31327;
	G32773<= not G31376;
	G32774<= not G30735;
	G32775<= not G30825;
	G32776<= not G31672;
	G32777<= not G31710;
	G32778<= not G31021;
	G32779<= not G30937;
	G32781<= not G31376;
	G32782<= not G30735;
	G32783<= not G30825;
	G32784<= not G31672;
	G32785<= not G31710;
	G32786<= not G31021;
	G32787<= not G30937;
	G32788<= not G31327;
	G32789<= not G30735;
	G32790<= not G30825;
	G32791<= not G31672;
	G32792<= not G31710;
	G32793<= not G31021;
	G32794<= not G30937;
	G32795<= not G31327;
	G32796<= not G31376;
	G32797<= not G30825;
	G32798<= not G31672;
	G32799<= not G31710;
	G32800<= not G31021;
	G32801<= not G30937;
	G32802<= not G31327;
	G32803<= not G31376;
	G32804<= not G30735;
	G32805<= not G31672;
	G32806<= not G31710;
	G32807<= not G31021;
	G32808<= not G30937;
	G32809<= not G31327;
	G32810<= not G31376;
	G32811<= not G30735;
	G32812<= not G30825;
	G32813<= not G31710;
	G32814<= not G31021;
	G32815<= not G30937;
	G32816<= not G31327;
	G32817<= not G31376;
	G32818<= not G30735;
	G32819<= not G30825;
	G32820<= not G31672;
	G32821<= not G31021;
	G32822<= not G30937;
	G32823<= not G31327;
	G32824<= not G31376;
	G32825<= not G30735;
	G32826<= not G30825;
	G32827<= not G31672;
	G32828<= not G31710;
	G32829<= not G30937;
	G32830<= not G31327;
	G32831<= not G31376;
	G32832<= not G30735;
	G32833<= not G30825;
	G32834<= not G31672;
	G32835<= not G31710;
	G32836<= not G31021;
	G32837<= not G31327;
	G32838<= not G31376;
	G32839<= not G30735;
	G32840<= not G30825;
	G32841<= not G31672;
	G32842<= not G31710;
	G32843<= not G31021;
	G32844<= not G30937;
	G32846<= not G31376;
	G32847<= not G30735;
	G32848<= not G30825;
	G32849<= not G31021;
	G32850<= not G30937;
	G32851<= not G31327;
	G32852<= not G30614;
	G32853<= not G30673;
	G32854<= not G30735;
	G32855<= not G30825;
	G32856<= not G31021;
	G32857<= not G30937;
	G32858<= not G31327;
	G32859<= not G30614;
	G32860<= not G30673;
	G32861<= not G31376;
	G32862<= not G30825;
	G32863<= not G31021;
	G32864<= not G30937;
	G32865<= not G31327;
	G32866<= not G30614;
	G32867<= not G30673;
	G32868<= not G31376;
	G32869<= not G30735;
	G32870<= not G31021;
	G32871<= not G30937;
	G32872<= not G31327;
	G32873<= not G30614;
	G32874<= not G30673;
	G32875<= not G31376;
	G32876<= not G30735;
	G32877<= not G30825;
	G32878<= not G30937;
	G32879<= not G31327;
	G32880<= not G30614;
	G32881<= not G30673;
	G32882<= not G31376;
	G32883<= not G30735;
	G32884<= not G30825;
	G32885<= not G31021;
	G32886<= not G31327;
	G32887<= not G30614;
	G32888<= not G30673;
	G32889<= not G31376;
	G32890<= not G30735;
	G32891<= not G30825;
	G32892<= not G31021;
	G32893<= not G30937;
	G32894<= not G30614;
	G32895<= not G30673;
	G32896<= not G31376;
	G32897<= not G30735;
	G32898<= not G30825;
	G32899<= not G31021;
	G32900<= not G30937;
	G32901<= not G31327;
	G32902<= not G30673;
	G32903<= not G31376;
	G32904<= not G30735;
	G32905<= not G30825;
	G32906<= not G31021;
	G32907<= not G30937;
	G32908<= not G31327;
	G32909<= not G30614;
	G32911<= not G31376;
	G32912<= not G30735;
	G32913<= not G30825;
	G32914<= not G31672;
	G32915<= not G31710;
	G32916<= not G31021;
	G32917<= not G30937;
	G32918<= not G31327;
	G32919<= not G30735;
	G32920<= not G30825;
	G32921<= not G31672;
	G32922<= not G31710;
	G32923<= not G31021;
	G32924<= not G30937;
	G32925<= not G31327;
	G32926<= not G31376;
	G32927<= not G30825;
	G32928<= not G31672;
	G32929<= not G31710;
	G32930<= not G31021;
	G32931<= not G30937;
	G32932<= not G31327;
	G32933<= not G31376;
	G32934<= not G30735;
	G32935<= not G31672;
	G32936<= not G31710;
	G32937<= not G31021;
	G32938<= not G30937;
	G32939<= not G31327;
	G32940<= not G31376;
	G32941<= not G30735;
	G32942<= not G30825;
	G32943<= not G31710;
	G32944<= not G31021;
	G32945<= not G30937;
	G32946<= not G31327;
	G32947<= not G31376;
	G32948<= not G30735;
	G32949<= not G30825;
	G32950<= not G31672;
	G32951<= not G31021;
	G32952<= not G30937;
	G32953<= not G31327;
	G32954<= not G31376;
	G32955<= not G30735;
	G32956<= not G30825;
	G32957<= not G31672;
	G32958<= not G31710;
	G32959<= not G30937;
	G32960<= not G31327;
	G32961<= not G31376;
	G32962<= not G30735;
	G32963<= not G30825;
	G32964<= not G31672;
	G32965<= not G31710;
	G32966<= not G31021;
	G32967<= not G31327;
	G32968<= not G31376;
	G32969<= not G30735;
	G32970<= not G30825;
	G32971<= not G31672;
	G32972<= not G31710;
	G32973<= not G31021;
	G32974<= not G30937;
	G32975<= not I30537;
	G33072<= not G31945;
	G33079<= not I30641;
	G33080<= not I30644;
	G33120<= not I30686;
	G33127<= not G31950;
	G33136<= not G32057;
	G33142<= not G32072;
	G33228<= not I30766;
	G33246<= not G32212;
	G33250<= not G32186;
	G33258<= not G32296;
	G33326<= not G32318;
	G33335<= not I30861;
	G33346<= not G32132;
	G33354<= not G32329;
	G33375<= not G32377;
	G33377<= not I30901;
	G33378<= not I30904;
	G33382<= not G32033;
	G33385<= not G32038;
	G33388<= not G32382;
	G33391<= not G32384;
	G33413<= not G31971;
	G33424<= not G32415;
	G33426<= not G32017;
	G33430<= not G32421;
	G33435<= not I30959;
	G33436<= not I30962;
	G33442<= not G31937;
	G33443<= not I30971;
	G33451<= not G32132;
	G33454<= not I30980;
	G33455<= not I30983;
	G33456<= not I30986;
	G33457<= not I30989;
	G33458<= not I30992;
	G33459<= not I30995;
	G33460<= not I30998;
	G33533<= not I31361;
	G33631<= not I31459;
	G33635<= not G33436;
	G33636<= not I31463;
	G33637<= not I31466;
	G33638<= not I31469;
	G33641<= not I31474;
	G33645<= not I31477;
	G33648<= not I31482;
	G33653<= not I31486;
	G33658<= not G33080;
	G33659<= not I31491;
	G33660<= not I31494;
	G33661<= not I31497;
	G33665<= not I31500;
	G33670<= not I31504;
	G33682<= not I31515;
	G33686<= not G33187;
	G33688<= not I31523;
	G33691<= not I31528;
	G33695<= not G33187;
	G33696<= not I31535;
	G33698<= not I31539;
	G33702<= not I31545;
	G33705<= not I31550;
	G33708<= not I31555;
	G33712<= not I31561;
	G33713<= not I31564;
	G33716<= not I31569;
	G33726<= not I31581;
	G33729<= not I31586;
	G33736<= not I31597;
	G33744<= not I31604;
	G33750<= not I31607;
	G33755<= not I31610;
	G33761<= not I31616;
	G33766<= not I31619;
	G33772<= not I31622;
	G33778<= not I31625;
	G33797<= not G33306;
	G33799<= not G33299;
	G33800<= not I31642;
	G33804<= not G33250;
	G33806<= not I31650;
	G33813<= not I31659;
	G33827<= not I31672;
	G33839<= not I31686;
	G33845<= not I31694;
	G33850<= not I31701;
	G33874<= not I31724;
	G33875<= not I31727;
	G33888<= not G33346;
	G33894<= not I31748;
	G33895<= not I31751;
	G33912<= not I31770;
	G33916<= not I31776;
	G33917<= not I31779;
	G33918<= not I31782;
	G33920<= not I31786;
	G33923<= not I31791;
	G33926<= not I31796;
	G33928<= not I31800;
	G33929<= not I31803;
	G33931<= not I31807;
	G33932<= not I31810;
	G33934<= not I31814;
	G33935<= not I31817;
	G33936<= not I31820;
	G33937<= not I31823;
	G33944<= not I31829;
	G33959<= not I31878;
	G34042<= not G33674;
	G34044<= not G33675;
	G34047<= not G33637;
	G34049<= not G33678;
	G34052<= not G33635;
	G34053<= not G33683;
	G34058<= not G33660;
	G34059<= not G33658;
	G34060<= not G33704;
	G34062<= not G33711;
	G34068<= not G33728;
	G34070<= not G33725;
	G34094<= not G33772;
	G34118<= not I32051;
	G34121<= not I32056;
	G34122<= not I32059;
	G34123<= not I32062;
	G34124<= not G33819;
	G34126<= not I32067;
	G34130<= not I32071;
	G34131<= not I32074;
	G34132<= not G33831;
	G34134<= not I32079;
	G34142<= not I32089;
	G34144<= not I32093;
	G34145<= not I32096;
	G34147<= not G33823;
	G34150<= not I32103;
	G34151<= not I32106;
	G34152<= not I32109;
	G34156<= not G33907;
	G34159<= not I32116;
	G34160<= not I32119;
	G34161<= not G33851;
	G34181<= not G33913;
	G34188<= not G33875;
	G34192<= not G33921;
	G34195<= not I32150;
	G34197<= not G33812;
	G34200<= not G33895;
	G34201<= not I32158;
	G34202<= not I32161;
	G34208<= not G33838;
	G34209<= not I32170;
	G34210<= not I32173;
	G34221<= not I32192;
	G34222<= not I32195;
	G34229<= not G33936;
	G34241<= not I32222;
	G34242<= not I32225;
	G34243<= not I32228;
	G34244<= not I32231;
	G34245<= not I32234;
	G34246<= not I32237;
	G34247<= not I32240;
	G34248<= not I32243;
	G34270<= not G34159;
	G34271<= not G34160;
	G34272<= not G34229;
	G34275<= not G34047;
	G34276<= not G34058;
	G34277<= not I32274;
	G34285<= not I32284;
	G34296<= not I32297;
	G34299<= not G34080;
	G34302<= not I32305;
	G34304<= not I32309;
	G34307<= not G34087;
	G34308<= not G34088;
	G34311<= not G34097;
	G34312<= not G34098;
	G34313<= not G34086;
	G34315<= not G34085;
	G34316<= not G34093;
	G34317<= not G34115;
	G34320<= not G34119;
	G34323<= not G34105;
	G34325<= not G34092;
	G34326<= not G34091;
	G34327<= not G34108;
	G34328<= not G34096;
	G34336<= not G34112;
	G34339<= not G34077;
	G34343<= not G34089;
	G34345<= not I32352;
	G34346<= not G34162;
	G34351<= not G34174;
	G34358<= not I32364;
	G34383<= not I32388;
	G34384<= not I32391;
	G34387<= not G34188;
	G34391<= not G34200;
	G34392<= not G34202;
	G34400<= not G34142;
	G34408<= not G34144;
	G34409<= not G34145;
	G34418<= not G34150;
	G34419<= not G34151;
	G34420<= not G34152;
	G34423<= not G34222;
	G34425<= not I32446;
	G34426<= not I32449;
	G34427<= not I32452;
	G34428<= not I32455;
	G34429<= not I32458;
	G34430<= not I32461;
	G34431<= not I32464;
	G34432<= not I32467;
	G34433<= not I32470;
	G34434<= not I32473;
	G34435<= not I32476;
	G34436<= not I32479;
	G34437<= not I32482;
	G34471<= not G34423;
	G34472<= not I32525;
	G34473<= not G34426;
	G34480<= not I32535;
	G34490<= not I32547;
	G34491<= not I32550;
	G34501<= not G34400;
	G34504<= not G34408;
	G34505<= not G34409;
	G34510<= not G34418;
	G34511<= not G34419;
	G34512<= not G34420;
	G34521<= not G34270;
	G34522<= not G34271;
	G34530<= not I32591;
	G34531<= not I32594;
	G34536<= not I32601;
	G34539<= not G34354;
	G34540<= not I32607;
	G34543<= not G34359;
	G34544<= not I32613;
	G34549<= not I32617;
	G34553<= not I32621;
	G34559<= not G34384;
	G34569<= not I32639;
	G34570<= not G34392;
	G34573<= not I32645;
	G34574<= not I32648;
	G34575<= not I32651;
	G34576<= not I32654;
	G34579<= not I32659;
	G34583<= not I32665;
	G34587<= not I32671;
	G34589<= not I32675;
	G34590<= not I32678;
	G34591<= not I32681;
	G34592<= not I32684;
	G34593<= not I32687;
	G34594<= not I32690;
	G34595<= not I32693;
	G34596<= not I32696;
	G34597<= not I32699;
	G34648<= not I32752;
	G34653<= not I32763;
	G34654<= not I32766;
	G34656<= not I32770;
	G34659<= not I32775;
	G34660<= not G34473;
	G34664<= not I32782;
	G34668<= not I32788;
	G34669<= not I32791;
	G34670<= not I32794;
	G34671<= not I32797;
	G34672<= not I32800;
	G34673<= not I32803;
	G34674<= not I32806;
	G34675<= not I32809;
	G34676<= not I32812;
	G34677<= not I32815;
	G34680<= not I32820;
	G34682<= not I32824;
	G34683<= not I32827;
	G34688<= not I32834;
	G34689<= not I32837;
	G34690<= not I32840;
	G34691<= not I32843;
	G34692<= not I32846;
	G34697<= not G34545;
	G34698<= not G34550;
	G34699<= not I32855;
	G34711<= not G34559;
	G34712<= not I32868;
	G34713<= not I32871;
	G34714<= not I32874;
	G34716<= not I32878;
	G34717<= not I32881;
	G34718<= not I32884;
	G34736<= not I32904;
	G34739<= not I32909;
	G34749<= not I32921;
	G34755<= not I32929;
	G34759<= not I32935;
	G34760<= not I32938;
	G34766<= not G34703;
	G34767<= not I32947;
	G34768<= not I32950;
	G34769<= not I32953;
	G34770<= not I32956;
	G34772<= not I32960;
	G34773<= not I32963;
	G34775<= not I32967;
	G34776<= not I32970;
	G34777<= not I32973;
	G34778<= not I32976;
	G34784<= not I32982;
	G34785<= not I32985;
	G34786<= not I32988;
	G34787<= not I32991;
	G34788<= not I32994;
	G34789<= not I32997;
	G34810<= not I33020;
	G34812<= not I33024;
	G34813<= not I33027;
	G34816<= not I33030;
	G34820<= not I33034;
	G34823<= not I33037;
	G34827<= not I33041;
	G34830<= not I33044;
	G34833<= not I33047;
	G34836<= not I33050;
	G34839<= not I33053;
	G34840<= not I33056;
	G34844<= not G34737;
	G34845<= not G34773;
	G34846<= not I33064;
	G34847<= not I33067;
	G34848<= not I33070;
	G34851<= not I33075;
	G34852<= not G34845;
	G34855<= not I33079;
	G34864<= not G34840;
	G34877<= not I33103;
	G34878<= not I33106;
	G34879<= not I33109;
	G34883<= not G34852;
	G34893<= not I33119;
	G34910<= not G34864;
	G34913<= not I33131;
	G34914<= not I33134;
	G34915<= not I33137;
	G34916<= not I33140;
	G34917<= not I33143;
	G34918<= not I33146;
	G34919<= not I33149;
	G34920<= not I33152;
	G34921<= not I33155;
	G34922<= not I33158;
	G34923<= not I33161;
	G34924<= not I33164;
	G34925<= not I33167;
	G34926<= not I33170;
	G34927<= not I33173;
	G34928<= not I33176;
	G34929<= not I33179;
	G34930<= not I33182;
	G34932<= not G34914;
	G34933<= not G34916;
	G34934<= not G34918;
	G34935<= not I33189;
	G34938<= not G34920;
	G34939<= not G34922;
	G34940<= not G34924;
	G34941<= not G34926;
	G34942<= not G34928;
	G34943<= not I33197;
	G34944<= not G34932;
	G34945<= not G34933;
	G34946<= not G34934;
	G34947<= not G34938;
	G34949<= not G34939;
	G34950<= not G34940;
	G34951<= not G34941;
	G34952<= not G34942;
	G34954<= not I33210;
	G34956<= not I33214;
	G34960<= not I33218;
	G34972<= not I33232;
	G34973<= not I33235;
	G34981<= not G34973;
	G34982<= not I33246;
	G34983<= not I33249;
	G34984<= not I33252;
	G34985<= not I33255;
	G34986<= not I33258;
	G34987<= not I33261;
	G34988<= not I33264;
	G34989<= not I33267;
	G34990<= not I33270;
	G34991<= not I33273;
	G34992<= not I33276;
	G34993<= not I33279;
	G34994<= not I33282;
	G34995<= not I33285;
	G34996<= not I33288;
	G34997<= not I33291;
	G34998<= not G34981;
	G35001<= not I33297;
	G35002<= not I33300;
	I11617<= not G1;
	I11620<= not G1;
	I11623<= not G28;
	I11626<= not G31;
	I11629<= not G19;
	I11632<= not G16;
	I11635<= not G9;
	I11655<= not G1246;
	I11665<= not G1589;
	I11682<= not G2756;
	I11685<= not G117;
	I11688<= not G70;
	I11691<= not G36;
	I11697<= not G3352;
	I11701<= not G4164;
	I11708<= not G3703;
	I11716<= not G4054;
	I11721<= not G4145;
	I11726<= not G4273;
	I11734<= not G4473;
	I11737<= not G4467;
	I11740<= not G4519;
	I11743<= not G4564;
	I11746<= not G4570;
	I11750<= not G4474;
	I11753<= not G4492;
	I11777<= not G5357;
	I11785<= not G5703;
	I11793<= not G6049;
	I11801<= not G6395;
	I11809<= not G6741;
	I11816<= not G93;
	I11820<= not G3869;
	I11835<= not G101;
	I11843<= not G111;
	I11860<= not G43;
	I11892<= not G4408;
	I11896<= not G4446;
	I11903<= not G4414;
	I11908<= not G4449;
	I11980<= not G66;
	I11992<= not G763;
	I12000<= not G582;
	I12003<= not G767;
	I12013<= not G590;
	I12016<= not G772;
	I12026<= not G344;
	I12030<= not G595;
	I12033<= not G776;
	I12041<= not G2741;
	I12046<= not G613;
	I12049<= not G781;
	I12056<= not G2748;
	I12061<= not G562;
	I12064<= not G617;
	I12067<= not G739;
	I12070<= not G785;
	I12083<= not G568;
	I12086<= not G622;
	I12089<= not G744;
	I12092<= not G790;
	I12103<= not G572;
	I12106<= not G626;
	I12109<= not G749;
	I12112<= not G794;
	I12117<= not G586;
	I12120<= not G632;
	I12123<= not G758;
	I12128<= not G4253;
	I12132<= not G577;
	I12135<= not G807;
	I12141<= not G599;
	I12144<= not G554;
	I12151<= not G604;
	I12159<= not G608;
	I12167<= not G5176;
	I12172<= not G2715;
	I12176<= not G5523;
	I12183<= not G2719;
	I12189<= not G5869;
	I12199<= not G6215;
	I12214<= not G6561;
	I12227<= not G34;
	I12300<= not G1157;
	I12314<= not G1500;
	I12333<= not G45;
	I12336<= not G52;
	I12355<= not G46;
	I12360<= not G528;
	I12382<= not G47;
	I12411<= not G4809;
	I12415<= not G48;
	I12418<= not G55;
	I12437<= not G4999;
	I12451<= not G3092;
	I12463<= not G4812;
	I12483<= not G3096;
	I12487<= not G3443;
	I12493<= not G5002;
	I12497<= not G49;
	I12503<= not G215;
	I12519<= not G3447;
	I12523<= not G3794;
	I12530<= not G4815;
	I12534<= not G50;
	I12538<= not G58;
	I12541<= not G194;
	I12563<= not G3798;
	I12568<= not G5005;
	I12572<= not G51;
	I12577<= not G1227;
	I12580<= not G1239;
	I12605<= not G1570;
	I12608<= not G1582;
	I12618<= not G3338;
	I12631<= not G1242;
	I12644<= not G3689;
	I12654<= not G1585;
	I12666<= not G4040;
	I12709<= not G4284;
	I12712<= not G59;
	I12719<= not G365;
	I12735<= not G4572;
	I12746<= not G4087;
	I12749<= not G4575;
	I12758<= not G4093;
	I12761<= not G4188;
	I12764<= not G4194;
	I12767<= not G4197;
	I12770<= not G4200;
	I12773<= not G4204;
	I12776<= not G4207;
	I12779<= not G4210;
	I12787<= not G4311;
	I12790<= not G4340;
	I12793<= not G4578;
	I12799<= not G59;
	I12805<= not G4098;
	I12808<= not G4322;
	I12811<= not G4340;
	I12819<= not G4277;
	I12823<= not G4311;
	I12826<= not G4349;
	I12837<= not G4222;
	I12855<= not G4311;
	I12858<= not G4340;
	I12861<= not G4372;
	I12884<= not G4213;
	I12887<= not G4216;
	I12890<= not G4219;
	I12893<= not G4226;
	I12896<= not G4229;
	I12899<= not G4232;
	I12907<= not G4322;
	I12910<= not G4340;
	I12927<= not G4332;
	I12930<= not G4349;
	I12935<= not G6753;
	I12950<= not G4287;
	I12954<= not G4358;
	I12963<= not G640;
	I12987<= not G12;
	I12991<= not G6752;
	I12994<= not G6748;
	I12997<= not G351;
	I13007<= not G65;
	I13010<= not G6749;
	I13020<= not G6750;
	I13031<= not G6747;
	I13037<= not G4304;
	I13054<= not G6744;
	I13057<= not G112;
	I13094<= not G2724;
	I13124<= not G2729;
	I13149<= not G6745;
	I13152<= not G6746;
	I13166<= not G5101;
	I13202<= not G5105;
	I13206<= not G5448;
	I13236<= not G5452;
	I13240<= not G5794;
	I13252<= not G6751;
	I13276<= not G5798;
	I13280<= not G6140;
	I13287<= not G110;
	I13317<= not G6144;
	I13321<= not G6486;
	I13326<= not G66;
	I13329<= not G86;
	I13352<= not G4146;
	I13360<= not G5343;
	I13374<= not G6490;
	I13424<= not G5689;
	I13473<= not G4157;
	I13483<= not G6035;
	I13539<= not G6381;
	I13548<= not G94;
	I13552<= not G121;
	I13581<= not G6727;
	I13597<= not G4417;
	I13606<= not G74;
	I13623<= not G4294;
	I13634<= not G79;
	I13637<= not G102;
	I13672<= not G106;
	I13684<= not G128;
	I13694<= not G117;
	I13699<= not G4581;
	I13705<= not G63;
	I13708<= not G136;
	I13715<= not G71;
	I13718<= not G890;
	I13723<= not G3167;
	I13726<= not G4537;
	I13740<= not G85;
	I13744<= not G3518;
	I13759<= not G6754;
	I13762<= not G6755;
	I13779<= not G6868;
	I13802<= not G6971;
	I13805<= not G6976;
	I13847<= not G7266;
	I13857<= not G9780;
	I13872<= not G7474;
	I13875<= not G1233;
	I13889<= not G7598;
	I13892<= not G1576;
	I13906<= not G7620;
	I13968<= not G7697;
	I13979<= not G7733;
	I13990<= not G7636;
	I13995<= not G8744;
	I14006<= not G9104;
	I14016<= not G9104;
	I14033<= not G8912;
	I14046<= not G9900;
	I14050<= not G9963;
	I14054<= not G10028;
	I14069<= not G9104;
	I14079<= not G7231;
	I14119<= not G7824;
	I14158<= not G8806;
	I14192<= not G10233;
	I14222<= not G8286;
	I14241<= not G8356;
	I14267<= not G7835;
	I14271<= not G8456;
	I14301<= not G8571;
	I14305<= not G8805;
	I14326<= not G8607;
	I14346<= not G10233;
	I14365<= not G3303;
	I14381<= not G8300;
	I14395<= not G3654;
	I14409<= not G8364;
	I14424<= not G4005;
	I14450<= not G4191;
	I14455<= not G10197;
	I14475<= not G10175;
	I14505<= not G10140;
	I14537<= not G10106;
	I14550<= not G10072;
	I14563<= not G802;
	I14567<= not G9708;
	I14570<= not G7932;
	I14576<= not G8791;
	I14579<= not G8792;
	I14584<= not G9766;
	I14589<= not G8818;
	I14593<= not G9978;
	I14602<= not G9340;
	I14619<= not G4185;
	I14623<= not G8925;
	I14630<= not G7717;
	I14633<= not G9340;
	I14644<= not G7717;
	I14647<= not G7717;
	I14650<= not G9340;
	I14653<= not G9417;
	I14660<= not G9746;
	I14663<= not G9747;
	I14668<= not G7753;
	I14671<= not G7717;
	I14679<= not G9332;
	I14684<= not G7717;
	I14687<= not G7753;
	I14690<= not G9340;
	I14702<= not G7717;
	I14705<= not G7717;
	I14708<= not G9417;
	I14727<= not G7753;
	I14730<= not G7717;
	I14742<= not G9534;
	I14745<= not G10029;
	I14749<= not G10031;
	I14761<= not G7753;
	I14773<= not G9581;
	I14797<= not G9636;
	I14800<= not G10107;
	I14823<= not G8056;
	I14827<= not G9686;
	I14830<= not G10141;
	I14833<= not G10142;
	I14836<= not G9688;
	I14839<= not G9689;
	I14862<= not G8092;
	I14866<= not G9748;
	I14893<= not G9819;
	I14896<= not G9820;
	I14899<= not G10198;
	I14902<= not G9821;
	I14905<= not G9822;
	I14932<= not G9901;
	I14935<= not G9902;
	I14939<= not G10216;
	I14964<= not G10230;
	I14967<= not G9964;
	I14970<= not G9965;
	I14999<= not G10030;
	I15030<= not G10073;
	I15033<= not G10273;
	I15036<= not G799;
	I15070<= not G10108;
	I15073<= not G10109;
	I15102<= not G5313;
	I15144<= not G5659;
	I15162<= not G10176;
	I15190<= not G6005;
	I15205<= not G10139;
	I15208<= not G637;
	I15223<= not G10119;
	I15238<= not G6351;
	I15250<= not G9152;
	I15284<= not G6697;
	I15295<= not G8515;
	I15316<= not G10087;
	I15382<= not G9071;
	I15448<= not G10877;
	I15474<= not G10364;
	I15494<= not G10385;
	I15533<= not G11867;
	I15536<= not G1227;
	I15542<= not G1570;
	I15550<= not G10430;
	I15556<= not G11928;
	I15564<= not G11949;
	I15569<= not G11965;
	I15572<= not G10499;
	I15577<= not G10430;
	I15587<= not G11985;
	I15590<= not G11988;
	I15593<= not G11989;
	I15600<= not G10430;
	I15609<= not G12013;
	I15617<= not G12037;
	I15620<= not G12038;
	I15623<= not G12040;
	I15626<= not G12041;
	I15633<= not G12074;
	I15636<= not G12075;
	I15647<= not G12109;
	I15650<= not G12110;
	I15663<= not G5308;
	I15667<= not G12143;
	I15677<= not G5654;
	I15682<= not G12182;
	I15697<= not G6000;
	I15702<= not G12217;
	I15705<= not G12218;
	I15717<= not G6346;
	I15727<= not G10981;
	I15732<= not G6692;
	I15736<= not G12322;
	I15765<= not G10823;
	I15773<= not G10430;
	I15782<= not G10430;
	I15788<= not G10430;
	I15800<= not G11607;
	I15811<= not G11128;
	I15814<= not G11129;
	I15821<= not G11143;
	I15824<= not G1116;
	I15831<= not G10416;
	I15834<= not G11164;
	I15837<= not G1459;
	I15843<= not G11181;
	I15846<= not G11183;
	I15862<= not G11215;
	I15869<= not G11234;
	I15872<= not G11236;
	I15878<= not G11249;
	I15893<= not G10430;
	I15906<= not G10430;
	I15915<= not G10430;
	I15918<= not G12381;
	I15921<= not G12381;
	I15929<= not G10430;
	I15932<= not G12381;
	I15937<= not G11676;
	I15942<= not G12381;
	I15954<= not G12381;
	I15981<= not G11290;
	I15987<= not G12381;
	I16010<= not G11148;
	I16024<= not G11171;
	I16028<= not G12381;
	I16040<= not G10430;
	I16057<= not G10430;
	I16077<= not G10430;
	I16090<= not G10430;
	I16102<= not G10430;
	I16117<= not G10430;
	I16120<= not G11868;
	I16135<= not G10430;
	I16150<= not G10430;
	I16160<= not G11237;
	I16163<= not G11930;
	I16168<= not G3321;
	I16181<= not G3672;
	I16193<= not G3281;
	I16201<= not G4023;
	I16217<= not G3632;
	I16231<= not G10520;
	I16246<= not G3983;
	I16289<= not G12107;
	I16328<= not G878;
	I16345<= not G881;
	I16357<= not G884;
	I16371<= not G887;
	I16391<= not G859;
	I16401<= not G869;
	I16417<= not G875;
	I16438<= not G11165;
	I16452<= not G11182;
	I16455<= not G11845;
	I16460<= not G10430;
	I16468<= not G12760;
	I16471<= not G12367;
	I16476<= not G10430;
	I16479<= not G10430;
	I16486<= not G11204;
	I16489<= not G12793;
	I16492<= not G12430;
	I16498<= not G10430;
	I16502<= not G10430;
	I16512<= not G12811;
	I16515<= not G12477;
	I16521<= not G10430;
	I16526<= not G10430;
	I16535<= not G11235;
	I16538<= not G10417;
	I16541<= not G11929;
	I16544<= not G11931;
	I16555<= not G10430;
	I16564<= not G10429;
	I16575<= not G3298;
	I16579<= not G10981;
	I16590<= not G11966;
	I16593<= not G10498;
	I16596<= not G12640;
	I16606<= not G3649;
	I16610<= not G10981;
	I16613<= not G10430;
	I16626<= not G11986;
	I16629<= not G11987;
	I16639<= not G4000;
	I16651<= not G10542;
	I16660<= not G10981;
	I16663<= not G10981;
	I16676<= not G10588;
	I16679<= not G12039;
	I16688<= not G10981;
	I16698<= not G12077;
	I16709<= not G10430;
	I16713<= not G5331;
	I16724<= not G12108;
	I16733<= not G12026;
	I16741<= not G5677;
	I16747<= not G12729;
	I16755<= not G12377;
	I16762<= not G5290;
	I16770<= not G6023;
	I16775<= not G12183;
	I16795<= not G5637;
	I16803<= not G6369;
	I16821<= not G5983;
	I16829<= not G6715;
	I16847<= not G6329;
	I16855<= not G10473;
	I16875<= not G6675;
	I16898<= not G10615;
	I16917<= not G10582;
	I16969<= not G13943;
	I17008<= not G12857;
	I17094<= not G14331;
	I17098<= not G14336;
	I17101<= not G14338;
	I17104<= not G12932;
	I17108<= not G13782;
	I17111<= not G13809;
	I17114<= not G14358;
	I17118<= not G14363;
	I17121<= not G14366;
	I17125<= not G13809;
	I17128<= not G13835;
	I17131<= not G14384;
	I17136<= not G14398;
	I17140<= not G13835;
	I17143<= not G14412;
	I17148<= not G14442;
	I17154<= not G13605;
	I17159<= not G13350;
	I17166<= not G14536;
	I17173<= not G13716;
	I17181<= not G13745;
	I17188<= not G13782;
	I17198<= not G13809;
	I17207<= not G13835;
	I17228<= not G13350;
	I17249<= not G13605;
	I17276<= not G13605;
	I17302<= not G14044;
	I17314<= not G14078;
	I17324<= not G14119;
	I17355<= not G14591;
	I17374<= not G13638;
	I17392<= not G13680;
	I17395<= not G12952;
	I17401<= not G13394;
	I17416<= not G13806;
	I17420<= not G13394;
	I17425<= not G13416;
	I17436<= not G13416;
	I17442<= not G13638;
	I17456<= not G13680;
	I17471<= not G13394;
	I17488<= not G13394;
	I17491<= not G13416;
	I17507<= not G13416;
	I17557<= not G14510;
	I17569<= not G14564;
	I17590<= not G14591;
	I17609<= not G13510;
	I17612<= not G13250;
	I17615<= not G13251;
	I17626<= not G14582;
	I17633<= not G13258;
	I17636<= not G14252;
	I17639<= not G13350;
	I17650<= not G13271;
	I17653<= not G14276;
	I17658<= not G13394;
	I17661<= not G13329;
	I17668<= not G13279;
	I17671<= not G13280;
	I17675<= not G13394;
	I17679<= not G13416;
	I17695<= not G14330;
	I17699<= not G13416;
	I17704<= not G13144;
	I17723<= not G13177;
	I17733<= not G14844;
	I17744<= not G14912;
	I17747<= not G13298;
	I17750<= not G14383;
	I17754<= not G13494;
	I17763<= not G13191;
	I17772<= not G14888;
	I17780<= not G13303;
	I17783<= not G13304;
	I17787<= not G3267;
	I17801<= not G14936;
	I17808<= not G13311;
	I17814<= not G3274;
	I17819<= not G3618;
	I17834<= not G14977;
	I17839<= not G13412;
	I17842<= not G13051;
	I17852<= not G3625;
	I17857<= not G3969;
	I17873<= not G15017;
	I17876<= not G13070;
	I17879<= not G14386;
	I17892<= not G3325;
	I17901<= not G3976;
	I17916<= not G13087;
	I17919<= not G14609;
	I17932<= not G3310;
	I17938<= not G3676;
	I17956<= not G14562;
	I17964<= not G3661;
	I17970<= not G4027;
	I17976<= not G13638;
	I17989<= not G14173;
	I17999<= not G4012;
	I18003<= not G13638;
	I18006<= not G13638;
	I18009<= not G13680;
	I18028<= not G13638;
	I18031<= not G13680;
	I18034<= not G13680;
	I18048<= not G13638;
	I18051<= not G13680;
	I18060<= not G14198;
	I18063<= not G14357;
	I18066<= not G3317;
	I18071<= not G13680;
	I18078<= not G13350;
	I18083<= not G13394;
	I18086<= not G13856;
	I18089<= not G13144;
	I18092<= not G3668;
	I18101<= not G13416;
	I18104<= not G13177;
	I18107<= not G4019;
	I18114<= not G14509;
	I18117<= not G13302;
	I18120<= not G13350;
	I18125<= not G13191;
	I18131<= not G13350;
	I18135<= not G13144;
	I18138<= not G14277;
	I18143<= not G13350;
	I18148<= not G13526;
	I18151<= not G13144;
	I18154<= not G13177;
	I18160<= not G14441;
	I18165<= not G13177;
	I18168<= not G13191;
	I18177<= not G13191;
	I18180<= not G13605;
	I18191<= not G14385;
	I18205<= not G14563;
	I18214<= not G12918;
	I18221<= not G13605;
	I18224<= not G13793;
	I18233<= not G14639;
	I18238<= not G13144;
	I18245<= not G14676;
	I18248<= not G12938;
	I18252<= not G13177;
	I18259<= not G12946;
	I18262<= not G13857;
	I18265<= not G13350;
	I18270<= not G13191;
	I18276<= not G1075;
	I18280<= not G12951;
	I18285<= not G13638;
	I18293<= not G1079;
	I18297<= not G1418;
	I18301<= not G12976;
	I18304<= not G14790;
	I18307<= not G12977;
	I18310<= not G12978;
	I18313<= not G13350;
	I18320<= not G13605;
	I18323<= not G13680;
	I18333<= not G1083;
	I18337<= not G1422;
	I18341<= not G14308;
	I18344<= not G13003;
	I18350<= not G13716;
	I18360<= not G1426;
	I18364<= not G13009;
	I18367<= not G13010;
	I18370<= not G14873;
	I18373<= not G13011;
	I18376<= not G14332;
	I18379<= not G13012;
	I18382<= not G13350;
	I18398<= not G13745;
	I18408<= not G13017;
	I18411<= not G13018;
	I18414<= not G14359;
	I18434<= not G13782;
	I18443<= not G13027;
	I18446<= not G13028;
	I18460<= not G5276;
	I18469<= not G13809;
	I18476<= not G14031;
	I18479<= not G13041;
	I18482<= not G13350;
	I18504<= not G5283;
	I18509<= not G5623;
	I18518<= not G13835;
	I18523<= not G14443;
	I18526<= not G13055;
	I18555<= not G5630;
	I18560<= not G5969;
	I18571<= not G13074;
	I18574<= not G13075;
	I18600<= not G5335;
	I18609<= not G5976;
	I18614<= not G6315;
	I18647<= not G5320;
	I18653<= not G5681;
	I18662<= not G6322;
	I18667<= not G6661;
	I18674<= not G13101;
	I18694<= not G5666;
	I18700<= not G6027;
	I18709<= not G6668;
	I18728<= not G6012;
	I18734<= not G6373;
	I18752<= not G6358;
	I18758<= not G6719;
	I18778<= not G6704;
	I18788<= not G13138;
	I18795<= not G5327;
	I18810<= not G13716;
	I18813<= not G5673;
	I18822<= not G13745;
	I18825<= not G6019;
	I18829<= not G13350;
	I18832<= not G13782;
	I18835<= not G6365;
	I18839<= not G13716;
	I18842<= not G13809;
	I18845<= not G6711;
	I18849<= not G14290;
	I18852<= not G13716;
	I18855<= not G13745;
	I18858<= not G13835;
	I18861<= not G14307;
	I18865<= not G14314;
	I18868<= not G14315;
	I18872<= not G13745;
	I18875<= not G13782;
	I18879<= not G13267;
	I18882<= not G16580;
	I18885<= not G16643;
	I18888<= not G16644;
	I18891<= not G16676;
	I18894<= not G16708;
	I18897<= not G16738;
	I18900<= not G16767;
	I18903<= not G16872;
	I18906<= not G16963;
	I18909<= not G16873;
	I18912<= not G15050;
	I19012<= not G15060;
	I19235<= not G15078;
	I19238<= not G15079;
	I19345<= not G15083;
	I19348<= not G15084;
	I19384<= not G15085;
	I19484<= not G15122;
	I19487<= not G15125;
	I19661<= not G17587;
	I19671<= not G15932;
	I19674<= not G15932;
	I19704<= not G17653;
	I19707<= not G17590;
	I19719<= not G17431;
	I19734<= not G17725;
	I19756<= not G17812;
	I19759<= not G17767;
	I19762<= not G15732;
	I19772<= not G17818;
	I19775<= not G17780;
	I19778<= not G17781;
	I19786<= not G17844;
	I19789<= not G17793;
	I19796<= not G17870;
	I19799<= not G17817;
	I19802<= not G15727;
	I19813<= not G17952;
	I19818<= not G1056;
	I19831<= not G16533;
	I19837<= not G1399;
	I19843<= not G16594;
	I19851<= not G16615;
	I19857<= not G16640;
	I19863<= not G16675;
	I19917<= not G18088;
	I19927<= not G17408;
	I20035<= not G15706;
	I20116<= not G15737;
	I20130<= not G15748;
	I20216<= not G15862;
	I20233<= not G17487;
	I20318<= not G16920;
	I20321<= not G16920;
	I20355<= not G17613;
	I20369<= not G17690;
	I20385<= not G16194;
	I20388<= not G17724;
	I20399<= not G16205;
	I20412<= not G16213;
	I20433<= not G16234;
	I20447<= not G16244;
	I20495<= not G16283;
	I20499<= not G16224;
	I20529<= not G16309;
	I20542<= not G16508;
	I20562<= not G16525;
	I20569<= not G16486;
	I20584<= not G16587;
	I20609<= not G16539;
	I20647<= not G17010;
	I20650<= not G17010;
	I20690<= not G15733;
	I20744<= not G17141;
	I20747<= not G17141;
	I20750<= not G16677;
	I20753<= not G16677;
	I20781<= not G17155;
	I20793<= not G17694;
	I20816<= not G17088;
	I20819<= not G17088;
	I20830<= not G17657;
	I20840<= not G17727;
	I20846<= not G16923;
	I20861<= not G16960;
	I20864<= not G16960;
	I20867<= not G16216;
	I20870<= not G16216;
	I20882<= not G17619;
	I20891<= not G17700;
	I20895<= not G16954;
	I20910<= not G17197;
	I20913<= not G16964;
	I20929<= not G17663;
	I20937<= not G16967;
	I20951<= not G17782;
	I20954<= not G16228;
	I20957<= not G16228;
	I20982<= not G16300;
	I20985<= not G16300;
	I20999<= not G16709;
	I21002<= not G16709;
	I21006<= not G15579;
	I21013<= not G15806;
	I21019<= not G17325;
	I21029<= not G15816;
	I21033<= not G17221;
	I21036<= not G17221;
	I21042<= not G15824;
	I21047<= not G17429;
	I21058<= not G17747;
	I21067<= not G15573;
	I21074<= not G17766;
	I21100<= not G16284;
	I21115<= not G15714;
	I21162<= not G17292;
	I21181<= not G17413;
	I21189<= not G17475;
	I21199<= not G17501;
	I21210<= not G17526;
	I21222<= not G18091;
	I21226<= not G16540;
	I21230<= not G16540;
	I21234<= not G16540;
	I21238<= not G16540;
	I21242<= not G16540;
	I21246<= not G16540;
	I21250<= not G16540;
	I21254<= not G16540;
	I21258<= not G16540;
	I21285<= not G18215;
	I21288<= not G18216;
	I21291<= not G18273;
	I21294<= not G18274;
	I21297<= not G18597;
	I21300<= not G18598;
	I21477<= not G18695;
	I21480<= not G18696;
	I21483<= not G18726;
	I21486<= not G18727;
	I21722<= not G19264;
	I21734<= not G19268;
	I21744<= not G19338;
	I21757<= not G21308;
	I21766<= not G19620;
	I21769<= not G19402;
	I21776<= not G21308;
	I21784<= not G19638;
	I21787<= not G19422;
	I21792<= not G21308;
	I21802<= not G21308;
	I21810<= not G20596;
	I21815<= not G21308;
	I21831<= not G19127;
	I21838<= not G19263;
	I21849<= not G19620;
	I21860<= not G19638;
	I21911<= not G21278;
	I21918<= not G21290;
	I21922<= not G21335;
	I21930<= not G21297;
	I21934<= not G21273;
	I21941<= not G18918;
	I21959<= not G20242;
	I21969<= not G21370;
	I22000<= not G20277;
	I22009<= not G21269;
	I22024<= not G19350;
	I22028<= not G20204;
	I22031<= not G21387;
	I22046<= not G19330;
	I22096<= not G19890;
	I22111<= not G19919;
	I22114<= not G19935;
	I22124<= not G21300;
	I22128<= not G19968;
	I22131<= not G19984;
	I22143<= not G20189;
	I22149<= not G21036;
	I22153<= not G20014;
	I22177<= not G21366;
	I22180<= not G21366;
	I22211<= not G21463;
	I22240<= not G20086;
	I22264<= not G20100;
	I22275<= not G20127;
	I22286<= not G19446;
	I22289<= not G19446;
	I22302<= not G19353;
	I22316<= not G19361;
	I22327<= not G19367;
	I22331<= not G19417;
	I22343<= not G19371;
	I22353<= not G19375;
	I22366<= not G19757;
	I22380<= not G21156;
	I22400<= not G19620;
	I22419<= not G19638;
	I22422<= not G19330;
	I22425<= not G19379;
	I22444<= not G19626;
	I22458<= not G18954;
	I22461<= not G21225;
	I22464<= not G21222;
	I22467<= not G19662;
	I22470<= not G21326;
	I22485<= not G21308;
	I22488<= not G18984;
	I22499<= not G21160;
	I22502<= not G19376;
	I22512<= not G19389;
	I22525<= not G19345;
	I22539<= not G19606;
	I22542<= not G19773;
	I22547<= not G20720;
	I22557<= not G20695;
	I22561<= not G20841;
	I22564<= not G20857;
	I22571<= not G20097;
	I22576<= not G21282;
	I22580<= not G20982;
	I22583<= not G20998;
	I22589<= not G21340;
	I22601<= not G21127;
	I22604<= not G21143;
	I22619<= not G21193;
	I22622<= not G21209;
	I22640<= not G21256;
	I22665<= not G21308;
	I22692<= not G21308;
	I22725<= not G21250;
	I22729<= not G21308;
	I22745<= not G19458;
	I22748<= not G19458;
	I22769<= not G21277;
	I22785<= not G18940;
	I22788<= not G18940;
	I22816<= not G19862;
	I22819<= not G19862;
	I22886<= not G18926;
	I22889<= not G18926;
	I22918<= not G21451;
	I22989<= not G21175;
	I23099<= not G20682;
	I23149<= not G19061;
	I23300<= not G21665;
	I23303<= not G21669;
	I23306<= not G21673;
	I23309<= not G21677;
	I23312<= not G21681;
	I23315<= not G21685;
	I23318<= not G21689;
	I23321<= not G21693;
	I23324<= not G21697;
	I23327<= not G22647;
	I23330<= not G22658;
	I23333<= not G22683;
	I23336<= not G22721;
	I23339<= not G23232;
	I23342<= not G23299;
	I23345<= not G23320;
	I23348<= not G23384;
	I23351<= not G23263;
	I23354<= not G23277;
	I23357<= not G23359;
	I23360<= not G23360;
	I23363<= not G23385;
	I23366<= not G23321;
	I23369<= not G23347;
	I23372<= not G23361;
	I23375<= not G23403;
	I23378<= not G23426;
	I23381<= not G23322;
	I23384<= not G23362;
	I23387<= not G23394;
	I23390<= not G23395;
	I23393<= not G23414;
	I23396<= not G23427;
	I23399<= not G23450;
	I23671<= not G23202;
	I23680<= not G23219;
	I23684<= not G23230;
	I23688<= not G23244;
	I23694<= not G23252;
	I23711<= not G23192;
	I23998<= not G22182;
	I24008<= not G22182;
	I24022<= not G22182;
	I24038<= not G22202;
	I24041<= not G22182;
	I24060<= not G22202;
	I24078<= not G22360;
	I24089<= not G22409;
	I24128<= not G23009;
	I24191<= not G22360;
	I24215<= not G22360;
	I24228<= not G22409;
	I24237<= not G23823;
	I24278<= not G23440;
	I24281<= not G23440;
	I24331<= not G22976;
	I24334<= not G22976;
	I24393<= not G23453;
	I24396<= not G23453;
	I24400<= not G23954;
	I24434<= not G22763;
	I24445<= not G22923;
	I24448<= not G22923;
	I24455<= not G22541;
	I24474<= not G22546;
	I24497<= not G22592;
	I24558<= not G23777;
	I24759<= not G24229;
	I24781<= not G24264;
	I24784<= not G24265;
	I24787<= not G24266;
	I24839<= not G24298;
	I24920<= not G25513;
	I25005<= not G24417;
	I25028<= not G24484;
	I25095<= not G25265;
	I25105<= not G25284;
	I25115<= not G25322;
	I25146<= not G24911;
	I25161<= not G24920;
	I25190<= not G25423;
	I25327<= not G24641;
	I25351<= not G24466;
	I25356<= not G24374;
	I25359<= not G24715;
	I25366<= not G24477;
	I25369<= not G24891;
	I25380<= not G24481;
	I25391<= not G24483;
	I25399<= not G24489;
	I25511<= not G25073;
	I25514<= not G25073;
	I25530<= not G25222;
	I25534<= not G25448;
	I25541<= not G25180;
	I25552<= not G25240;
	I25555<= not G25241;
	I25562<= not G25250;
	I25567<= not G25272;
	I25576<= not G25296;
	I25579<= not G25297;
	I25586<= not G25537;
	I25591<= not G25380;
	I25594<= not G25531;
	I25598<= not G25424;
	I25606<= not G25465;
	I25677<= not G25640;
	I25680<= not G25641;
	I25683<= not G25642;
	I25689<= not G25688;
	I25692<= not G25689;
	I25695<= not G25690;
	I25743<= not G25903;
	I25750<= not G26823;
	I25779<= not G26424;
	I25786<= not G26424;
	I25790<= not G26424;
	I25869<= not G25851;
	I25882<= not G25776;
	I26004<= not G26818;
	I26100<= not G26365;
	I26130<= not G26510;
	I26195<= not G26260;
	I26296<= not G26820;
	I26309<= not G26825;
	I26334<= not G26834;
	I26337<= not G26835;
	I26356<= not G26843;
	I26378<= not G26850;
	I26381<= not G26851;
	I26406<= not G26187;
	I26409<= not G26187;
	I26427<= not G26859;
	I26430<= not G26856;
	I26448<= not G26860;
	I26451<= not G26862;
	I26466<= not G26870;
	I26479<= not G25771;
	I26503<= not G26811;
	I26508<= not G26814;
	I26512<= not G26817;
	I26516<= not G26824;
	I26578<= not G26941;
	I26581<= not G26942;
	I26584<= not G26943;
	I26638<= not G27965;
	I26649<= not G27675;
	I26654<= not G27576;
	I26664<= not G27708;
	I26667<= not G27585;
	I26670<= not G27709;
	I26676<= not G27736;
	I26679<= not G27773;
	I26682<= not G27774;
	I26687<= not G27880;
	I26693<= not G27930;
	I26700<= not G27956;
	I26705<= not G27967;
	I26710<= not G27511;
	I26785<= not G27013;
	I26799<= not G27660;
	I26880<= not G27527;
	I26925<= not G27015;
	I26929<= not G27980;
	I26936<= not G27599;
	I26952<= not G27972;
	I26989<= not G27277;
	I27192<= not G27662;
	I27232<= not G27993;
	I27235<= not G27320;
	I27238<= not G27320;
	I27253<= not G27996;
	I27271<= not G27998;
	I27314<= not G28009;
	I27368<= not G27881;
	I27385<= not G27438;
	I27388<= not G27698;
	I27391<= not G27929;
	I27401<= not G27051;
	I27449<= not G27737;
	I27481<= not G27928;
	I27492<= not G27511;
	I27495<= not G27961;
	I27543<= not G28187;
	I27546<= not G29041;
	I27549<= not G28161;
	I27552<= not G28162;
	I27555<= not G28142;
	I27558<= not G28155;
	I27561<= not G28163;
	I27564<= not G28166;
	I27567<= not G28181;
	I27570<= not G28262;
	I27573<= not G28157;
	I27576<= not G28173;
	I27579<= not G28184;
	I27677<= not G28156;
	I27713<= not G28224;
	I27718<= not G28231;
	I27730<= not G28752;
	I27735<= not G28779;
	I27738<= not G28140;
	I27742<= not G28819;
	I27749<= not G28917;
	I27758<= not G28119;
	I27777<= not G29043;
	I27784<= not G29013;
	I27927<= not G28803;
	I27941<= not G28803;
	I27954<= not G28803;
	I27970<= not G28803;
	I28002<= not G28153;
	I28014<= not G28158;
	I28062<= not G29194;
	I28128<= not G28314;
	I28162<= not G28803;
	I28174<= not G28803;
	I28185<= not G28803;
	I28199<= not G28803;
	I28241<= not G28709;
	I28301<= not G29042;
	I28336<= not G29147;
	I28349<= not G28367;
	I28390<= not G29185;
	I28419<= not G29195;
	I28434<= not G28114;
	I28458<= not G28443;
	I28480<= not G28652;
	I28540<= not G28954;
	I28548<= not G28147;
	I28572<= not G28274;
	I28576<= not G28431;
	I28579<= not G29474;
	I28582<= not G30116;
	I28585<= not G30217;
	I28588<= not G29368;
	I28591<= not G29371;
	I28594<= not G29379;
	I28597<= not G29374;
	I28832<= not G30301;
	I28838<= not G29372;
	I28851<= not G29317;
	I28866<= not G29730;
	I28872<= not G30072;
	I28883<= not G30105;
	I28897<= not G30155;
	I28908<= not G30182;
	I28913<= not G30322;
	I28925<= not G29987;
	I29002<= not G29675;
	I29013<= not G29705;
	I29139<= not G29382;
	I29149<= not G29384;
	I29182<= not G30012;
	I29185<= not G30012;
	I29199<= not G30237;
	I29204<= not G29505;
	I29207<= not G30293;
	I29211<= not G30298;
	I29214<= not G30300;
	I29218<= not G30304;
	I29221<= not G30307;
	I29225<= not G30311;
	I29228<= not G30314;
	I29233<= not G30295;
	I29236<= not G29498;
	I29239<= not G29498;
	I29242<= not G29313;
	I29245<= not G29491;
	I29248<= not G29491;
	I29337<= not G30286;
	I29363<= not G30218;
	I29368<= not G30321;
	I29371<= not G30325;
	I29438<= not G30610;
	I29441<= not G30917;
	I29444<= not G30928;
	I29447<= not G30729;
	I29571<= not G31783;
	I29579<= not G30565;
	I29582<= not G30591;
	I29585<= not G31655;
	I29717<= not G30931;
	I29720<= not G30931;
	I29891<= not G31578;
	I29894<= not G31771;
	I29909<= not G31791;
	I29913<= not G30605;
	I29936<= not G30606;
	I29939<= not G31667;
	I29961<= not G30984;
	I29965<= not G31189;
	I29969<= not G30991;
	I29973<= not G31213;
	I29977<= not G31596;
	I29981<= not G31591;
	I30537<= not G32027;
	I30641<= not G32024;
	I30644<= not G32024;
	I30686<= not G32381;
	I30766<= not G32363;
	I30861<= not G32383;
	I30901<= not G32407;
	I30904<= not G32424;
	I30959<= not G32021;
	I30962<= not G32021;
	I30971<= not G32015;
	I30980<= not G32132;
	I30983<= not G32433;
	I30986<= not G32437;
	I30989<= not G32441;
	I30992<= not G32445;
	I30995<= not G32449;
	I30998<= not G32453;
	I31361<= not G33120;
	I31459<= not G33219;
	I31463<= not G33318;
	I31466<= not G33318;
	I31469<= not G33388;
	I31474<= not G33212;
	I31477<= not G33391;
	I31482<= not G33204;
	I31486<= not G33197;
	I31491<= not G33283;
	I31494<= not G33283;
	I31497<= not G33187;
	I31500<= not G33176;
	I31504<= not G33164;
	I31515<= not G33187;
	I31523<= not G33187;
	I31528<= not G33219;
	I31535<= not G33377;
	I31539<= not G33212;
	I31545<= not G33219;
	I31550<= not G33204;
	I31555<= not G33212;
	I31561<= not G33197;
	I31564<= not G33204;
	I31569<= not G33197;
	I31581<= not G33164;
	I31586<= not G33149;
	I31597<= not G33187;
	I31604<= not G33176;
	I31607<= not G33164;
	I31610<= not G33149;
	I31616<= not G33219;
	I31619<= not G33212;
	I31622<= not G33204;
	I31625<= not G33197;
	I31642<= not G33204;
	I31650<= not G33212;
	I31659<= not G33219;
	I31672<= not G33149;
	I31686<= not G33164;
	I31694<= not G33176;
	I31701<= not G33164;
	I31724<= not G33076;
	I31727<= not G33076;
	I31748<= not G33228;
	I31751<= not G33228;
	I31770<= not G33197;
	I31776<= not G33204;
	I31779<= not G33212;
	I31782<= not G33219;
	I31786<= not G33197;
	I31791<= not G33354;
	I31796<= not G33176;
	I31800<= not G33164;
	I31803<= not G33176;
	I31807<= not G33149;
	I31810<= not G33164;
	I31814<= not G33149;
	I31817<= not G33323;
	I31820<= not G33323;
	I31823<= not G33149;
	I31829<= not G33454;
	I31878<= not G33696;
	I32051<= not G33631;
	I32056<= not G33641;
	I32059<= not G33648;
	I32062<= not G33653;
	I32067<= not G33661;
	I32071<= not G33665;
	I32074<= not G33670;
	I32079<= not G33937;
	I32089<= not G33665;
	I32093<= not G33670;
	I32096<= not G33641;
	I32103<= not G33661;
	I32106<= not G33653;
	I32109<= not G33631;
	I32116<= not G33937;
	I32119<= not G33648;
	I32150<= not G33923;
	I32158<= not G33791;
	I32161<= not G33791;
	I32170<= not G33638;
	I32173<= not G33645;
	I32192<= not G33628;
	I32195<= not G33628;
	I32222<= not G34118;
	I32225<= not G34121;
	I32228<= not G34122;
	I32231<= not G34123;
	I32234<= not G34126;
	I32237<= not G34130;
	I32240<= not G34131;
	I32243<= not G34134;
	I32274<= not G34195;
	I32284<= not G34052;
	I32297<= not G34059;
	I32305<= not G34209;
	I32309<= not G34210;
	I32352<= not G34169;
	I32364<= not G34208;
	I32388<= not G34153;
	I32391<= not G34153;
	I32446<= not G34127;
	I32449<= not G34127;
	I32452<= not G34241;
	I32455<= not G34242;
	I32458<= not G34243;
	I32461<= not G34244;
	I32464<= not G34245;
	I32467<= not G34246;
	I32470<= not G34247;
	I32473<= not G34248;
	I32476<= not G34277;
	I32479<= not G34302;
	I32482<= not G34304;
	I32525<= not G34285;
	I32535<= not G34296;
	I32547<= not G34397;
	I32550<= not G34398;
	I32591<= not G34287;
	I32594<= not G34298;
	I32601<= not G34319;
	I32607<= not G34358;
	I32613<= not G34329;
	I32617<= not G34333;
	I32621<= not G34335;
	I32639<= not G34345;
	I32645<= not G34367;
	I32648<= not G34371;
	I32651<= not G34375;
	I32654<= not G34378;
	I32659<= not G34391;
	I32665<= not G34386;
	I32671<= not G34388;
	I32675<= not G34427;
	I32678<= not G34428;
	I32681<= not G34429;
	I32684<= not G34430;
	I32687<= not G34431;
	I32690<= not G34432;
	I32693<= not G34433;
	I32696<= not G34434;
	I32699<= not G34569;
	I32752<= not G34510;
	I32763<= not G34511;
	I32766<= not G34522;
	I32770<= not G34505;
	I32775<= not G34512;
	I32782<= not G34571;
	I32788<= not G34577;
	I32791<= not G34578;
	I32794<= not G34580;
	I32797<= not G34581;
	I32800<= not G34582;
	I32803<= not G34584;
	I32806<= not G34585;
	I32809<= not G34586;
	I32812<= not G34588;
	I32815<= not G34470;
	I32820<= not G34474;
	I32824<= not G34475;
	I32827<= not G34477;
	I32834<= not G34472;
	I32837<= not G34498;
	I32840<= not G34480;
	I32843<= not G34499;
	I32846<= not G34502;
	I32855<= not G34540;
	I32868<= not G34579;
	I32871<= not G34521;
	I32874<= not G34504;
	I32878<= not G34501;
	I32881<= not G34688;
	I32884<= not G34690;
	I32904<= not G34708;
	I32909<= not G34712;
	I32921<= not G34650;
	I32929<= not G34649;
	I32935<= not G34657;
	I32938<= not G34663;
	I32947<= not G34659;
	I32950<= not G34713;
	I32953<= not G34656;
	I32956<= not G34654;
	I32960<= not G34653;
	I32963<= not G34650;
	I32967<= not G34648;
	I32970<= not G34716;
	I32973<= not G34714;
	I32976<= not G34699;
	I32982<= not G34749;
	I32985<= not G34736;
	I32988<= not G34755;
	I32991<= not G34759;
	I32994<= not G34739;
	I32997<= not G34760;
	I33020<= not G34781;
	I33024<= not G34783;
	I33027<= not G34767;
	I33030<= not G34768;
	I33034<= not G34769;
	I33037<= not G34770;
	I33041<= not G34772;
	I33044<= not G34775;
	I33047<= not G34776;
	I33050<= not G34777;
	I33053<= not G34778;
	I33056<= not G34778;
	I33064<= not G34784;
	I33067<= not G34812;
	I33070<= not G34810;
	I33075<= not G34843;
	I33079<= not G34809;
	I33103<= not G34846;
	I33106<= not G34855;
	I33109<= not G34851;
	I33119<= not G34852;
	I33131<= not G34906;
	I33134<= not G34906;
	I33137<= not G34884;
	I33140<= not G34884;
	I33143<= not G34903;
	I33146<= not G34903;
	I33149<= not G34900;
	I33152<= not G34900;
	I33155<= not G34897;
	I33158<= not G34897;
	I33161<= not G34894;
	I33164<= not G34894;
	I33167<= not G34890;
	I33170<= not G34890;
	I33173<= not G34887;
	I33176<= not G34887;
	I33179<= not G34893;
	I33182<= not G34910;
	I33189<= not G34929;
	I33197<= not G34930;
	I33210<= not G34943;
	I33214<= not G34954;
	I33218<= not G34955;
	I33232<= not G34957;
	I33235<= not G34957;
	I33246<= not G34970;
	I33249<= not G34971;
	I33252<= not G34974;
	I33255<= not G34975;
	I33258<= not G34976;
	I33261<= not G34977;
	I33264<= not G34978;
	I33267<= not G34979;
	I33270<= not G34982;
	I33273<= not G34984;
	I33276<= not G34985;
	I33279<= not G34986;
	I33282<= not G34987;
	I33285<= not G34988;
	I33288<= not G34989;
	I33291<= not G34983;
	I33297<= not G35000;
	I33300<= not G35001;
	G7251<=G452 and G392;
	G7396<=G392 and G441;
	G7469<=G4382 and G4438;
	G7511<=G2145 and G2138 and G2130;
	G7520<=G2704 and G2697 and G2689;
	G7685<=G4382 and G4375;
	G7696<=G2955 and G2950;
	G7763<=G2965 and G2960;
	G7777<=G723 and G822 and G817;
	G7804<=G2975 and G2970;
	G7918<=G1205 and G1087;
	G7948<=G1548 and G1430;
	G8234<=G4515 and G4521;
	G8530<=G2902 and G2907;
	G8583<=G2917 and G2912;
	G8643<=G2927 and G2922;
	G8690<=G2941 and G2936;
	G8721<=G385 and G376 and G365;
	G9217<=G632 and G626;
	G9479<=G305 and G324;
	G9906<=G996 and G1157;
	G9967<=G1178 and G1157;
	G9968<=G1339 and G1500;
	G10034<=G1521 and G1500;
	G10290<=G4358 and G4349;
	G10476<=G7244 and G7259 and I13862;
	G10501<=G1233 and G9007;
	G10528<=G1576 and G9051;
	G10543<=G8238 and G437;
	G10565<=G8182 and G424;
	G10588<=G7004 and G5297;
	G10590<=G7246 and G7392 and I13937;
	G10616<=G7998 and G174;
	G10619<=G3080 and G7907;
	G10624<=G8387 and G3072;
	G10625<=G3431 and G7926;
	G10626<=G4057 and G7927;
	G10632<=G7475 and G7441 and G890;
	G10654<=G3085 and G8434;
	G10655<=G8440 and G3423;
	G10656<=G3782 and G7952;
	G10657<=G8451 and G4064;
	G10665<=G209 and G8292;
	G10674<=G6841 and G10200 and G2130;
	G10675<=G3436 and G8500;
	G10676<=G8506 and G3774;
	G10677<=G4141 and G7611;
	G10683<=G7289 and G4438;
	G10684<=G7998 and G411;
	G10704<=G2145 and G10200 and G2130;
	G10705<=G6850 and G10219 and G2689;
	G10706<=G3338 and G8691;
	G10707<=G3787 and G8561;
	G10719<=G6841 and G2138 and G2130;
	G10720<=G2704 and G10219 and G2689;
	G10721<=G3288 and G6875 and G3274 and G8481;
	G10724<=G3689 and G8728;
	G10732<=G6850 and G2697 and G2689;
	G10733<=G3639 and G6905 and G3625 and G8542;
	G10736<=G4040 and G8751;
	G10756<=G3990 and G6928 and G3976 and G8595;
	G10822<=G4264 and G8514;
	G10823<=G7704 and G5180 and G5188;
	G10827<=G8914 and G4258;
	G10828<=G6888 and G7640;
	G10829<=G7289 and G4375;
	G10838<=G7738 and G5527 and G5535;
	G10841<=G8509 and G8567;
	G10856<=G4269 and G8967;
	G10869<=G7766 and G5873 and G5881;
	G10873<=G3004 and G9015;
	G10874<=G7791 and G6219 and G6227;
	G10878<=G7858 and G1135;
	G10883<=G3355 and G9061;
	G10887<=G7812 and G6565 and G6573;
	G10890<=G7858 and G1105;
	G10896<=G1205 and G8654;
	G10898<=G3706 and G9100;
	G10902<=G7858 and G1129;
	G10917<=G9174 and G1087;
	G10921<=G1548 and G8685;
	G10925<=G7858 and G956;
	G10934<=G9197 and G7918;
	G10947<=G9200 and G1430;
	G10948<=G7880 and G1478;
	G10966<=G9226 and G7948;
	G10967<=G7880 and G1448;
	G10970<=G854 and G9582;
	G10998<=G8567 and G8509 and G8451 and G7650;
	G10999<=G7880 and G1472;
	G11003<=G7880 and G1300;
	G11010<=G4698 and G8933;
	G11016<=G4888 and G8984;
	G11018<=G7655 and G7643 and G7627;
	G11019<=G5092 and G9036;
	G11023<=G9669 and G5084;
	G11024<=G5436 and G9070;
	G11027<=G5097 and G9724;
	G11028<=G9730 and G5428;
	G11029<=G5782 and G9103;
	G11032<=G9354 and G7717;
	G11035<=G5441 and G9800;
	G11036<=G9806 and G5774;
	G11037<=G6128 and G9184;
	G11044<=G5343 and G10124;
	G11045<=G5787 and G9883;
	G11046<=G9889 and G6120;
	G11047<=G6474 and G9212;
	G11083<=G8836 and G802;
	G11111<=G5297 and G7004 and G5283 and G9780;
	G11114<=G5689 and G10160;
	G11115<=G6133 and G9954;
	G11116<=G9960 and G6466;
	G11123<=G5644 and G7028 and G5630 and G9864;
	G11126<=G6035 and G10185;
	G11127<=G6479 and G10022;
	G11139<=G5990 and G7051 and G5976 and G9935;
	G11142<=G6381 and G10207;
	G11144<=G239 and G8136 and G246 and I14198;
	G11160<=G6336 and G7074 and G6322 and G10003;
	G11163<=G6727 and G10224;
	G11166<=G8363 and G269 and G8296 and I14225;
	G11178<=G6682 and G7097 and G6668 and G10061;
	G11205<=G8217 and G8439;
	G11223<=G8281 and G8505;
	G11244<=G8346 and G8566;
	G11366<=G5016 and G10338;
	G11397<=G5360 and G7139;
	G11427<=G5706 and G7158;
	G11449<=G6052 and G7175;
	G11496<=G4382 and G7495;
	G11497<=G6398 and G7192;
	G11546<=G7289 and G4375;
	G11740<=G8769 and G703;
	G11890<=G7499 and G9155;
	G11893<=G1668 and G7268;
	G11915<=G1802 and G7315;
	G11916<=G2227 and G7328;
	G11937<=G1936 and G7362;
	G11939<=G2361 and G7380;
	G11956<=G2070 and G7411;
	G11960<=G2495 and G7424;
	G11967<=G311 and G7802;
	G11978<=G2629 and G7462;
	G12015<=G1002 and G7567;
	G12027<=G9499 and G9729;
	G12043<=G1345 and G7601;
	G12065<=G9557 and G9805;
	G12099<=G9619 and G9888;
	G12135<=G9684 and G9959;
	G12179<=G9745 and G10027;
	G12186<=G1178 and G7519;
	G12219<=G1189 and G7532;
	G12220<=G1521 and G7535;
	G12259<=G9480 and G640;
	G12284<=G1532 and G7557;
	G12527<=G8680 and G667;
	G12641<=G10295 and G3171 and G3179;
	G12687<=G9024 and G8977;
	G12692<=G10323 and G3522 and G3530;
	G12730<=G9024 and G4349;
	G12735<=G7121 and G3873 and G3881;
	G12761<=G969 and G7567;
	G12762<=G4358 and G8977;
	G12794<=G1008 and G7567;
	G12795<=G1312 and G7601;
	G12812<=G518 and G9158;
	G12817<=G1351 and G7601;
	G12920<=G1227 and G10960;
	G12924<=G1570 and G10980;
	G12931<=G392 and G11048;
	G12939<=G405 and G11048;
	G12953<=G411 and G11048;
	G12979<=G424 and G11048;
	G13019<=G194 and G11737;
	G13020<=G401 and G11048;
	G13025<=G8431 and G11026;
	G13029<=G8359 and G11030;
	G13030<=G429 and G11048;
	G13035<=G8497 and G11033;
	G13038<=G8509 and G11034;
	G13042<=G433 and G11048;
	G13046<=G6870 and G11270;
	G13047<=G8534 and G11042;
	G13048<=G8558 and G11043;
	G13059<=G6900 and G11303;
	G13060<=G8587 and G11110;
	G13063<=G8567 and G10808;
	G13080<=G6923 and G11357;
	G13081<=G8626 and G11122;
	G13156<=G10816 and G10812 and G10805;
	G13221<=G6946 and G11425;
	G13247<=G8964 and G11316;
	G13252<=G11561 and G11511 and G11469 and G699;
	G13265<=G9018 and G11493;
	G13277<=G3195 and G11432;
	G13282<=G3546 and G11480;
	G13287<=G1221 and G11472;
	G13290<=G3897 and G11534;
	G13294<=G1564 and G11513;
	G13299<=G437 and G11048;
	G13306<=G441 and G11048;
	G13313<=G475 and G11048;
	G13319<=G4076 and G8812 and G10658 and G8757;
	G13320<=G417 and G11048;
	G13321<=G847 and G11048;
	G13324<=G854 and G11326;
	G13333<=G4743 and G11755;
	G13345<=G4754 and G11773;
	G13349<=G4933 and G11780;
	G13383<=G4765 and G11797;
	G13384<=G4944 and G11804;
	G13393<=G703 and G11048;
	G13411<=G4955 and G11834;
	G13415<=G837 and G11048;
	G13436<=G9721 and G11811;
	G13461<=G2719 and G11819;
	G13473<=G9797 and G11841;
	G13491<=G6999 and G12160;
	G13492<=G9856 and G11865;
	G13493<=G9880 and G11866;
	G13497<=G2724 and G12155;
	G13507<=G7023 and G12198;
	G13508<=G9927 and G11888;
	G13509<=G9951 and G11889;
	G13523<=G7046 and G12246;
	G13524<=G9995 and G11910;
	G13525<=G10019 and G11911;
	G13541<=G7069 and G12308;
	G13542<=G10053 and G11927;
	G13564<=G4480 and G12820;
	G13566<=G7092 and G12358;
	G13567<=G10102 and G11948;
	G13604<=G4495 and G10487;
	G13632<=G10232 and G12228;
	G13633<=G4567 and G10509;
	G13656<=G278 and G11144;
	G13671<=G4498 and G10532;
	G13697<=G11166 and G8608;
	G13737<=G4501 and G10571;
	G13738<=G8880 and G10572;
	G13771<=G11441 and G11355 and G11302 and I16111;
	G13778<=G4540 and G10597;
	G13805<=G11489 and G11394 and G11356 and I16129;
	G13807<=G4504 and G10606;
	G13808<=G4543 and G10607;
	G13830<=G11543 and G11424 and G11395 and I16143;
	G13832<=G8880 and G10612;
	G13833<=G4546 and G10613;
	G13853<=G4549 and G10620;
	G13887<=G5204 and G12402;
	G13912<=G5551 and G12450;
	G13942<=G5897 and G12512;
	G13974<=G6243 and G12578;
	G13998<=G6589 and G12629;
	G14028<=G8673 and G11797;
	G14035<=G699 and G11048;
	G14061<=G8715 and G11834;
	G14097<=G878 and G10632;
	G14126<=G881 and G10632;
	G14148<=G884 and G10632;
	G14168<=G887 and G10632;
	G14180<=G872 and G10632;
	G14185<=G8686 and G11744;
	G14190<=G859 and G10632;
	G14193<=G7178 and G10590;
	G14202<=G869 and G10632;
	G14206<=G8655 and G11790;
	G14207<=G8639 and G11793;
	G14210<=G4392 and G10590;
	G14216<=G7631 and G10608;
	G14218<=G875 and G10632;
	G14220<=G8612 and G11820;
	G14221<=G8686 and G11823;
	G14222<=G8655 and G11826;
	G14233<=G8639 and G11855;
	G14256<=G2079 and G11872;
	G14257<=G8612 and G11878;
	G14261<=G4507 and G10738;
	G14295<=G1811 and G11894;
	G14296<=G2638 and G11897;
	G14316<=G2370 and G11920;
	G14438<=G1087 and G10726;
	G14496<=G12411 and G12244 and G12197 and I16618;
	G14506<=G1430 and G10755;
	G14528<=G12459 and G12306 and G12245 and I16646;
	G14537<=G10550 and G10529;
	G14555<=G12521 and G12356 and G12307 and I16671;
	G14565<=G11934 and G11952;
	G14566<=G10566 and G10551;
	G14567<=G10568 and G10552;
	G14581<=G12587 and G12428 and G12357 and I16695;
	G14585<=G1141 and G10905;
	G14586<=G11953 and G11970;
	G14587<=G10584 and G10567;
	G14588<=G11957 and G11974;
	G14589<=G10586 and G10569;
	G14608<=G12638 and G12476 and G12429 and I16721;
	G14610<=G1484 and G10935;
	G14612<=G11971 and G11993;
	G14613<=G10602 and G10585;
	G14614<=G11975 and G11997;
	G14615<=G10604 and G10587;
	G14641<=G11994 and G12020;
	G14643<=G11998 and G12023;
	G14644<=G10610 and G10605;
	G14654<=G7178 and G10476;
	G14680<=G12024 and G12053;
	G14681<=G4392 and G10476;
	G14708<=G74 and G12369;
	G14719<=G4392 and G10830;
	G14791<=G1146 and G10909;
	G14831<=G1152 and G10909;
	G14832<=G1489 and G10939;
	G14874<=G1099 and G10909;
	G14875<=G1495 and G10939;
	G14913<=G1442 and G10939;
	G15075<=G12850 and G12955;
	G15076<=G2130 and G12955;
	G15077<=G2138 and G12955;
	G15078<=G10361 and G12955;
	G15079<=G2151 and G12955;
	G15080<=G12855 and G12983;
	G15081<=G2689 and G12983;
	G15082<=G2697 and G12983;
	G15083<=G10362 and G12983;
	G15084<=G2710 and G12983;
	G15103<=G4180 and G14454;
	G15104<=G6955 and G14454;
	G15105<=G4235 and G14454;
	G15107<=G4258 and G14454;
	G15108<=G4264 and G14454;
	G15109<=G4269 and G14454;
	G15110<=G4245 and G14454;
	G15111<=G4281 and G14454;
	G15112<=G4284 and G14454;
	G15113<=G4291 and G14454;
	G15114<=G4239 and G14454;
	G15115<=G2946 and G14454;
	G15116<=G4297 and G14454;
	G15117<=G4300 and G14454;
	G15118<=G4253 and G14454;
	G15119<=G4249 and G14454;
	G15507<=G10970 and G13305;
	G15567<=G392 and G13312;
	G15574<=G4311 and G13202;
	G15589<=G411 and G13334;
	G15590<=G3139 and G13530;
	G15611<=G471 and G13437;
	G15612<=G3143 and G13530;
	G15613<=G3490 and G13555;
	G15631<=G168 and G13437;
	G15632<=G3494 and G13555;
	G15633<=G3841 and G13584;
	G15650<=G8362 and G13413;
	G15651<=G429 and G13414;
	G15652<=G174 and G13437;
	G15653<=G3119 and G13530;
	G15654<=G3845 and G13584;
	G15672<=G433 and G13458;
	G15673<=G182 and G13437;
	G15678<=G1094 and G13846;
	G15679<=G3470 and G13555;
	G15693<=G269 and G13474;
	G15694<=G457 and G13437;
	G15699<=G1437 and G13861;
	G15700<=G3089 and G13483;
	G15701<=G3821 and G13584;
	G15703<=G452 and G13437;
	G15704<=G3440 and G13504;
	G15706<=G13296 and G13484;
	G15707<=G4082 and G13506;
	G15711<=G460 and G13437;
	G15712<=G3791 and G13521;
	G15716<=G468 and G13437;
	G15722<=G464 and G13437;
	G15738<=G1111 and G13260;
	G15745<=G686 and G13223;
	G15749<=G1454 and G13273;
	G15757<=G3207 and G14066;
	G15779<=G13909 and G11214;
	G15783<=G3215 and G14098;
	G15784<=G3235 and G13977;
	G15785<=G3558 and G14107;
	G15786<=G13940 and G11233;
	G15793<=G3219 and G13873;
	G15794<=G3239 and G14008;
	G15795<=G3566 and G14130;
	G15796<=G3586 and G14015;
	G15797<=G3909 and G14139;
	G15804<=G3223 and G13889;
	G15805<=G3243 and G14041;
	G15807<=G3570 and G13898;
	G15808<=G3590 and G14048;
	G15809<=G3917 and G14154;
	G15810<=G3937 and G14055;
	G15812<=G3227 and G13915;
	G15813<=G3247 and G14069;
	G15814<=G3574 and G13920;
	G15815<=G3594 and G14075;
	G15817<=G3921 and G13929;
	G15818<=G3941 and G14082;
	G15819<=G3251 and G14101;
	G15820<=G3578 and G13955;
	G15821<=G3598 and G14110;
	G15822<=G3925 and G13960;
	G15823<=G3945 and G14116;
	G15836<=G3187 and G14104;
	G15837<=G3255 and G14127;
	G15838<=G3602 and G14133;
	G15839<=G3929 and G13990;
	G15840<=G3949 and G14142;
	G15841<=G4273 and G13868;
	G15847<=G3191 and G14005;
	G15848<=G3259 and G13892;
	G15849<=G3538 and G14136;
	G15850<=G3606 and G14151;
	G15851<=G3953 and G14157;
	G15852<=G13820 and G13223;
	G15856<=G9056 and G14223;
	G15857<=G3199 and G14038;
	G15858<=G3542 and G14045;
	G15859<=G3610 and G13923;
	G15860<=G3889 and G14160;
	G15861<=G3957 and G14170;
	G15863<=G13762 and G13223;
	G15870<=G3231 and G13948;
	G15871<=G3203 and G13951;
	G15872<=G9095 and G14234;
	G15873<=G3550 and G14072;
	G15874<=G3893 and G14079;
	G15875<=G3961 and G13963;
	G15876<=G13512 and G13223;
	G15880<=G3211 and G13980;
	G15881<=G3582 and G13983;
	G15882<=G3554 and G13986;
	G15883<=G9180 and G14258;
	G15884<=G3901 and G14113;
	G15902<=G441 and G13975;
	G15903<=G13796 and G13223;
	G15911<=G3111 and G13530;
	G15912<=G3562 and G14018;
	G15913<=G3933 and G14021;
	G15914<=G3905 and G14024;
	G15936<=G475 and G13999;
	G15937<=G11950 and G14387;
	G15966<=G3462 and G13555;
	G15967<=G3913 and G14058;
	G15978<=G246 and G14032;
	G15995<=G13314 and G1157 and G10666;
	G16023<=G3813 and G13584;
	G16025<=G446 and G14063;
	G16026<=G854 and G14065;
	G16047<=G13322 and G1500 and G10699;
	G16098<=G5148 and G14238;
	G16122<=G9491 and G14291;
	G16125<=G5152 and G14238;
	G16126<=G5495 and G14262;
	G16128<=G14333 and G14166;
	G16160<=G5499 and G14262;
	G16161<=G5841 and G14297;
	G16163<=G14254 and G14179;
	G16176<=G14596 and G11779;
	G16177<=G5128 and G14238;
	G16178<=G5845 and G14297;
	G16179<=G6187 and G14321;
	G16184<=G9285 and G14183;
	G16185<=G3263 and G14011;
	G16190<=G14626 and G11810;
	G16191<=G5475 and G14262;
	G16192<=G6191 and G14321;
	G16193<=G6533 and G14348;
	G16194<=G11547 and G6782 and G11640 and I17529;
	G16199<=G3614 and G14051;
	G16202<=G86 and G14197;
	G16203<=G5821 and G14297;
	G16204<=G6537 and G14348;
	G16205<=G11547 and G6782 and G11640 and I17542;
	G16207<=G9839 and G14204;
	G16208<=G3965 and G14085;
	G16211<=G5445 and G14215;
	G16212<=G6167 and G14321;
	G16213<=G6772 and G6782 and G11640 and I17552;
	G16221<=G5791 and G14231;
	G16222<=G6513 and G14348;
	G16224<=G14583 and G14232;
	G16233<=G6137 and G14251;
	G16234<=G6772 and G6782 and G11640 and I17575;
	G16243<=G6483 and G14275;
	G16244<=G11547 and G11592 and G6789 and I17585;
	G16245<=G14278 and G14708;
	G16279<=G4512 and G14424;
	G16283<=G11547 and G11592 and G6789 and I17606;
	G16303<=G4527 and G12921;
	G16324<=G13657 and G182;
	G16422<=G8216 and G13627;
	G16427<=G5216 and G14876;
	G16474<=G8280 and G13666;
	G16483<=G5224 and G14915;
	G16484<=G5244 and G14755;
	G16485<=G5563 and G14924;
	G16486<=G6772 and G11592 and G6789 and I17692;
	G16513<=G8345 and G13708;
	G16516<=G5228 and G14627;
	G16517<=G5248 and G14797;
	G16518<=G5571 and G14956;
	G16519<=G5591 and G14804;
	G16520<=G5909 and G14965;
	G16531<=G5232 and G14656;
	G16532<=G5252 and G14841;
	G16534<=G5575 and G14665;
	G16535<=G5595 and G14848;
	G16536<=G5917 and G14996;
	G16537<=G5937 and G14855;
	G16538<=G6255 and G15005;
	G16539<=G11547 and G6782 and G6789 and I17741;
	G16590<=G5236 and G14683;
	G16591<=G5256 and G14879;
	G16592<=G5579 and G14688;
	G16593<=G5599 and G14885;
	G16595<=G5921 and G14697;
	G16596<=G5941 and G14892;
	G16597<=G6263 and G15021;
	G16598<=G6283 and G14899;
	G16599<=G6601 and G15030;
	G16610<=G5260 and G14918;
	G16611<=G5583 and G14727;
	G16612<=G5603 and G14927;
	G16613<=G5925 and G14732;
	G16614<=G5945 and G14933;
	G16616<=G6267 and G14741;
	G16617<=G6287 and G14940;
	G16618<=G6609 and G15039;
	G16619<=G6629 and G14947;
	G16621<=G8278 and G13821;
	G16633<=G5196 and G14921;
	G16634<=G5264 and G14953;
	G16635<=G5607 and G14959;
	G16636<=G5929 and G14768;
	G16637<=G5949 and G14968;
	G16638<=G6271 and G14773;
	G16639<=G6291 and G14974;
	G16641<=G6613 and G14782;
	G16642<=G6633 and G14981;
	G16653<=G8343 and G13850;
	G16662<=G4552 and G14753;
	G16666<=G5200 and G14794;
	G16667<=G5268 and G14659;
	G16668<=G5543 and G14962;
	G16669<=G5611 and G14993;
	G16670<=G5953 and G14999;
	G16671<=G6275 and G14817;
	G16672<=G6295 and G15008;
	G16673<=G6617 and G14822;
	G16674<=G6637 and G15014;
	G16690<=G8399 and G13867;
	G16699<=G7134 and G12933;
	G16700<=G5208 and G14838;
	G16701<=G5547 and G14845;
	G16702<=G5615 and G14691;
	G16703<=G5889 and G15002;
	G16704<=G5957 and G15018;
	G16705<=G6299 and G15024;
	G16706<=G6621 and G14868;
	G16707<=G6641 and G15033;
	G16729<=G5240 and G14720;
	G16730<=G5212 and G14723;
	G16731<=G7153 and G12941;
	G16732<=G5555 and G14882;
	G16733<=G5893 and G14889;
	G16734<=G5961 and G14735;
	G16735<=G6235 and G15027;
	G16736<=G6303 and G15036;
	G16737<=G6645 and G15042;
	G16751<=G13155 and G13065;
	G16758<=G5220 and G14758;
	G16759<=G5587 and G14761;
	G16760<=G5559 and G14764;
	G16761<=G7170 and G12947;
	G16762<=G5901 and G14930;
	G16763<=G6239 and G14937;
	G16764<=G6307 and G14776;
	G16765<=G6581 and G15045;
	G16766<=G6649 and G12915;
	G16801<=G5120 and G14238;
	G16802<=G5567 and G14807;
	G16803<=G5933 and G14810;
	G16804<=G5905 and G14813;
	G16805<=G7187 and G12972;
	G16806<=G6247 and G14971;
	G16807<=G6585 and G14978;
	G16808<=G6653 and G14825;
	G16840<=G5467 and G14262;
	G16841<=G5913 and G14858;
	G16842<=G6279 and G14861;
	G16843<=G6251 and G14864;
	G16844<=G7212 and G13000;
	G16845<=G6593 and G15011;
	G16846<=G14034 and G12591 and G11185;
	G16855<=G4392 and G13107;
	G16868<=G5813 and G14297;
	G16869<=G6259 and G14902;
	G16870<=G6625 and G14905;
	G16871<=G6597 and G14908;
	G16884<=G6159 and G14321;
	G16885<=G6605 and G14950;
	G16896<=G262 and G13120;
	G16929<=G6505 and G14348;
	G16930<=G239 and G13132;
	G16957<=G13064 and G10418;
	G16965<=G269 and G13140;
	G16986<=G246 and G13142;
	G17057<=G446 and G13173;
	G17091<=G8659 and G12940;
	G17119<=G5272 and G14800;
	G17123<=G225 and G13209;
	G17133<=G10683 and G13222;
	G17134<=G5619 and G14851;
	G17138<=G255 and G13239;
	G17139<=G8635 and G12967;
	G17140<=G8616 and G12968;
	G17145<=G7469 and G13249;
	G17146<=G5965 and G14895;
	G17149<=G232 and G13255;
	G17150<=G8579 and G12995;
	G17151<=G8659 and G12996;
	G17152<=G8635 and G12997;
	G17153<=G6311 and G14943;
	G17156<=G305 and G13385;
	G17176<=G8616 and G13008;
	G17177<=G6657 and G14984;
	G17179<=G1041 and G13211;
	G17181<=G1945 and G13014;
	G17182<=G8579 and G13016;
	G17191<=G1384 and G13242;
	G17192<=G1677 and G13022;
	G17193<=G2504 and G13023;
	G17199<=G2236 and G13034;
	G17292<=G1075 and G13093;
	G17307<=G9498 and G14343;
	G17317<=G1079 and G13124;
	G17321<=G1418 and G13105;
	G17365<=G7650 and G13036;
	G17391<=G9556 and G14378;
	G17401<=G1083 and G13143;
	G17405<=G1422 and G13137;
	G17418<=G9618 and G14407;
	G17424<=G1426 and G13176;
	G17469<=G4076 and G13217;
	G17480<=G9683 and G14433;
	G17506<=G9744 and G14505;
	G17574<=G9554 and G14546;
	G17601<=G9616 and G14572;
	G17613<=G11547 and G11592 and G11640 and I18568;
	G17617<=G7885 and G13326;
	G17636<=G10829 and G13463;
	G17643<=G9681 and G14599;
	G17653<=G11547 and G11592 and G6789 and I18620;
	G17654<=G962 and G13284;
	G17655<=G7897 and G13342;
	G17671<=G7685 and G13485;
	G17682<=G9742 and G14637;
	G17690<=G11547 and G11592 and G11640 and I18671;
	G17692<=G1124 and G13307;
	G17693<=G1306 and G13291;
	G17719<=G9818 and G14675;
	G17724<=G11547 and G11592 and G11640 and I18713;
	G17725<=G11547 and G11592 and G6789 and I18716;
	G17726<=G1467 and G13315;
	G17747<=G6772 and G11592 and G11640 and I18740;
	G17752<=G7841 and G13174;
	G17753<=G13281 and G13175;
	G17766<=G6772 and G11592 and G11640 and I18762;
	G17767<=G6772 and G11592 and G6789 and I18765;
	G17768<=G13325 and G10741;
	G17769<=G1146 and G13188;
	G17770<=G7863 and G13189;
	G17771<=G13288 and G13190;
	G17780<=G6772 and G11592 and G11640 and I18782;
	G17781<=G6772 and G11592 and G6789 and I18785;
	G17783<=G7851 and G13110;
	G17784<=G1152 and G13215;
	G17785<=G13341 and G10762;
	G17786<=G1489 and G13216;
	G17793<=G6772 and G11592 and G6789 and I18803;
	G17809<=G7873 and G13125;
	G17810<=G1495 and G13246;
	G17817<=G11547 and G6782 and G11640 and I18819;
	G18103<=G401 and G17015;
	G18104<=G392 and G17015;
	G18105<=G417 and G17015;
	G18106<=G411 and G17015;
	G18107<=G429 and G17015;
	G18108<=G433 and G17015;
	G18109<=G437 and G17015;
	G18110<=G441 and G17015;
	G18111<=G174 and G17015;
	G18112<=G182 and G17015;
	G18113<=G405 and G17015;
	G18114<=G452 and G17015;
	G18115<=G460 and G17015;
	G18116<=G168 and G17015;
	G18117<=G464 and G17015;
	G18118<=G471 and G17015;
	G18119<=G475 and G17015;
	G18120<=G457 and G17015;
	G18121<=G424 and G17015;
	G18122<=G15052 and G17015;
	G18123<=G479 and G16886;
	G18124<=G102 and G16886;
	G18125<=G15053 and G16886;
	G18126<=G15054 and G16971;
	G18127<=G499 and G16971;
	G18128<=G504 and G16971;
	G18129<=G518 and G16971;
	G18130<=G528 and G16971;
	G18131<=G482 and G16971;
	G18132<=G513 and G16971;
	G18133<=G15055 and G17249;
	G18134<=G534 and G17249;
	G18135<=G136 and G17249;
	G18136<=G550 and G17249;
	G18137<=G538 and G17249;
	G18138<=G546 and G17249;
	G18139<=G542 and G17249;
	G18140<=G559 and G17533;
	G18141<=G568 and G17533;
	G18142<=G577 and G17533;
	G18143<=G586 and G17533;
	G18144<=G590 and G17533;
	G18145<=G582 and G17533;
	G18146<=G595 and G17533;
	G18147<=G599 and G17533;
	G18148<=G562 and G17533;
	G18149<=G608 and G17533;
	G18150<=G604 and G17533;
	G18151<=G617 and G17533;
	G18152<=G613 and G17533;
	G18153<=G626 and G17533;
	G18154<=G622 and G17533;
	G18155<=G15056 and G17533;
	G18156<=G572 and G17533;
	G18157<=G15057 and G17433;
	G18158<=G667 and G17433;
	G18159<=G671 and G17433;
	G18160<=G645 and G17433;
	G18161<=G691 and G17433;
	G18162<=G686 and G17433;
	G18163<=G79 and G17433;
	G18164<=G699 and G17433;
	G18165<=G650 and G17433;
	G18166<=G655 and G17433;
	G18167<=G718 and G17433;
	G18168<=G681 and G17433;
	G18169<=G676 and G17433;
	G18170<=G661 and G17433;
	G18171<=G728 and G17433;
	G18172<=G15058 and G17328;
	G18173<=G736 and G17328;
	G18174<=G739 and G17328;
	G18175<=G744 and G17328;
	G18176<=G732 and G17328;
	G18177<=G749 and G17328;
	G18178<=G758 and G17328;
	G18179<=G763 and G17328;
	G18180<=G767 and G17328;
	G18181<=G772 and G17328;
	G18182<=G776 and G17328;
	G18183<=G781 and G17328;
	G18184<=G785 and G17328;
	G18185<=G790 and G17328;
	G18186<=G753 and G17328;
	G18187<=G794 and G17328;
	G18188<=G807 and G17328;
	G18189<=G812 and G17821;
	G18190<=G822 and G17821;
	G18191<=G827 and G17821;
	G18192<=G817 and G17821;
	G18193<=G837 and G17821;
	G18194<=G843 and G17821;
	G18195<=G847 and G17821;
	G18196<=G703 and G17821;
	G18197<=G854 and G17821;
	G18198<=G15059 and G17821;
	G18199<=G832 and G17821;
	G18201<=G15061 and G15938;
	G18202<=G907 and G15938;
	G18203<=G911 and G15938;
	G18204<=G914 and G15938;
	G18205<=G904 and G15938;
	G18206<=G918 and G15938;
	G18207<=G925 and G15938;
	G18208<=G930 and G15938;
	G18209<=G921 and G15938;
	G18210<=G936 and G15938;
	G18211<=G15062 and G15979;
	G18212<=G947 and G15979;
	G18213<=G952 and G15979;
	G18214<=G939 and G15979;
	G18215<=G943 and G15979;
	G18216<=G967 and G15979;
	G18217<=G15063 and G16100;
	G18218<=G1008 and G16100;
	G18219<=G969 and G16100;
	G18220<=G1002 and G16100;
	G18221<=G1018 and G16100;
	G18222<=G1024 and G16100;
	G18223<=G1030 and G16100;
	G18224<=G1036 and G16100;
	G18225<=G1041 and G16100;
	G18226<=G15064 and G16129;
	G18227<=G1052 and G16129;
	G18228<=G1061 and G16129;
	G18229<=G1099 and G16326;
	G18230<=G1111 and G16326;
	G18231<=G1105 and G16326;
	G18232<=G1124 and G16326;
	G18233<=G1094 and G16326;
	G18234<=G1129 and G16326;
	G18235<=G1141 and G16326;
	G18236<=G15065 and G16326;
	G18237<=G1146 and G16326;
	G18238<=G1152 and G16326;
	G18239<=G1135 and G16326;
	G18240<=G15066 and G16431;
	G18241<=G1183 and G16431;
	G18242<=G962 and G16431;
	G18243<=G1189 and G16431;
	G18244<=G1171 and G16431;
	G18245<=G1193 and G16431;
	G18246<=G1199 and G16431;
	G18247<=G1178 and G16431;
	G18248<=G15067 and G16897;
	G18249<=G1216 and G16897;
	G18250<=G6821 and G16897;
	G18251<=G996 and G16897;
	G18252<=G990 and G16897;
	G18253<=G1211 and G16897;
	G18254<=G1236 and G16897;
	G18255<=G1087 and G16897;
	G18256<=G1242 and G16897;
	G18257<=G1205 and G16897;
	G18258<=G1221 and G16897;
	G18259<=G15068 and G16000;
	G18260<=G1252 and G16000;
	G18261<=G1256 and G16000;
	G18262<=G1259 and G16000;
	G18263<=G1249 and G16000;
	G18264<=G1263 and G16000;
	G18265<=G1270 and G16000;
	G18266<=G1274 and G16000;
	G18267<=G1266 and G16000;
	G18268<=G1280 and G16000;
	G18269<=G15069 and G16031;
	G18270<=G1291 and G16031;
	G18271<=G1296 and G16031;
	G18272<=G1283 and G16031;
	G18273<=G1287 and G16031;
	G18274<=G1311 and G16031;
	G18275<=G15070 and G16136;
	G18276<=G1351 and G16136;
	G18277<=G1312 and G16136;
	G18278<=G1345 and G16136;
	G18279<=G1361 and G16136;
	G18280<=G1367 and G16136;
	G18281<=G1373 and G16136;
	G18282<=G1379 and G16136;
	G18283<=G1384 and G16136;
	G18284<=G15071 and G16164;
	G18285<=G1395 and G16164;
	G18286<=G1404 and G16164;
	G18287<=G1442 and G16449;
	G18288<=G1454 and G16449;
	G18289<=G1448 and G16449;
	G18290<=G1467 and G16449;
	G18291<=G1437 and G16449;
	G18292<=G1472 and G16449;
	G18293<=G1484 and G16449;
	G18294<=G15072 and G16449;
	G18295<=G1489 and G16449;
	G18296<=G1495 and G16449;
	G18297<=G1478 and G16449;
	G18298<=G15073 and G16489;
	G18299<=G1526 and G16489;
	G18300<=G1306 and G16489;
	G18301<=G1532 and G16489;
	G18302<=G1514 and G16489;
	G18303<=G1536 and G16489;
	G18304<=G1542 and G16489;
	G18305<=G1521 and G16489;
	G18306<=G15074 and G16931;
	G18307<=G1559 and G16931;
	G18308<=G6832 and G16931;
	G18309<=G1339 and G16931;
	G18310<=G1333 and G16931;
	G18311<=G1554 and G16931;
	G18312<=G1579 and G16931;
	G18313<=G1430 and G16931;
	G18314<=G1585 and G16931;
	G18315<=G1548 and G16931;
	G18316<=G1564 and G16931;
	G18317<=G12846 and G17873;
	G18318<=G1604 and G17873;
	G18319<=G1600 and G17873;
	G18320<=G1616 and G17873;
	G18321<=G1620 and G17873;
	G18322<=G1608 and G17873;
	G18323<=G1632 and G17873;
	G18324<=G1644 and G17873;
	G18325<=G1624 and G17873;
	G18326<=G1664 and G17873;
	G18327<=G1636 and G17873;
	G18328<=G1657 and G17873;
	G18329<=G1612 and G17873;
	G18330<=G1668 and G17873;
	G18331<=G1682 and G17873;
	G18332<=G1677 and G17873;
	G18333<=G1691 and G17873;
	G18334<=G1696 and G17873;
	G18335<=G1687 and G17873;
	G18336<=G1700 and G17873;
	G18337<=G1706 and G17873;
	G18338<=G1710 and G17873;
	G18339<=G1714 and G17873;
	G18340<=G1720 and G17873;
	G18341<=G1648 and G17873;
	G18342<=G1592 and G17873;
	G18343<=G12847 and G17955;
	G18344<=G1740 and G17955;
	G18345<=G1736 and G17955;
	G18346<=G1752 and G17955;
	G18347<=G1756 and G17955;
	G18348<=G1744 and G17955;
	G18349<=G1768 and G17955;
	G18350<=G1779 and G17955;
	G18351<=G1760 and G17955;
	G18352<=G1798 and G17955;
	G18353<=G1772 and G17955;
	G18354<=G1792 and G17955;
	G18355<=G1748 and G17955;
	G18356<=G1802 and G17955;
	G18357<=G1816 and G17955;
	G18358<=G1811 and G17955;
	G18359<=G1825 and G17955;
	G18360<=G1830 and G17955;
	G18361<=G1821 and G17955;
	G18362<=G1834 and G17955;
	G18363<=G1840 and G17955;
	G18364<=G1844 and G17955;
	G18365<=G1848 and G17955;
	G18366<=G1854 and G17955;
	G18367<=G1783 and G17955;
	G18368<=G1728 and G17955;
	G18369<=G12848 and G15171;
	G18370<=G1874 and G15171;
	G18371<=G1870 and G15171;
	G18372<=G1886 and G15171;
	G18373<=G1890 and G15171;
	G18374<=G1878 and G15171;
	G18375<=G1902 and G15171;
	G18376<=G1913 and G15171;
	G18377<=G1894 and G15171;
	G18378<=G1932 and G15171;
	G18379<=G1906 and G15171;
	G18380<=G1926 and G15171;
	G18381<=G1882 and G15171;
	G18382<=G1936 and G15171;
	G18383<=G1950 and G15171;
	G18384<=G1945 and G15171;
	G18385<=G1959 and G15171;
	G18386<=G1964 and G15171;
	G18387<=G1955 and G15171;
	G18388<=G1968 and G15171;
	G18389<=G1974 and G15171;
	G18390<=G1978 and G15171;
	G18391<=G1982 and G15171;
	G18392<=G1988 and G15171;
	G18393<=G1917 and G15171;
	G18394<=G1862 and G15171;
	G18395<=G12849 and G15373;
	G18396<=G2008 and G15373;
	G18397<=G2004 and G15373;
	G18398<=G2020 and G15373;
	G18399<=G2024 and G15373;
	G18400<=G2012 and G15373;
	G18401<=G2036 and G15373;
	G18402<=G2047 and G15373;
	G18403<=G2028 and G15373;
	G18404<=G2066 and G15373;
	G18405<=G2040 and G15373;
	G18406<=G2060 and G15373;
	G18407<=G2016 and G15373;
	G18408<=G2070 and G15373;
	G18409<=G2084 and G15373;
	G18410<=G2079 and G15373;
	G18411<=G2093 and G15373;
	G18412<=G2098 and G15373;
	G18413<=G2089 and G15373;
	G18414<=G2102 and G15373;
	G18415<=G2108 and G15373;
	G18416<=G2112 and G15373;
	G18417<=G2116 and G15373;
	G18418<=G2122 and G15373;
	G18419<=G2051 and G15373;
	G18420<=G1996 and G15373;
	G18423<=G12851 and G18008;
	G18424<=G2165 and G18008;
	G18425<=G2161 and G18008;
	G18426<=G2177 and G18008;
	G18427<=G2181 and G18008;
	G18428<=G2169 and G18008;
	G18429<=G2193 and G18008;
	G18430<=G2204 and G18008;
	G18431<=G2185 and G18008;
	G18432<=G2223 and G18008;
	G18433<=G2197 and G18008;
	G18434<=G2217 and G18008;
	G18435<=G2173 and G18008;
	G18436<=G2227 and G18008;
	G18437<=G2241 and G18008;
	G18438<=G2236 and G18008;
	G18439<=G2250 and G18008;
	G18440<=G2255 and G18008;
	G18441<=G2246 and G18008;
	G18442<=G2259 and G18008;
	G18443<=G2265 and G18008;
	G18444<=G2269 and G18008;
	G18445<=G2273 and G18008;
	G18446<=G2279 and G18008;
	G18447<=G2208 and G18008;
	G18448<=G2153 and G18008;
	G18449<=G12852 and G15224;
	G18450<=G2299 and G15224;
	G18451<=G2295 and G15224;
	G18452<=G2311 and G15224;
	G18453<=G2315 and G15224;
	G18454<=G2303 and G15224;
	G18455<=G2327 and G15224;
	G18456<=G2338 and G15224;
	G18457<=G2319 and G15224;
	G18458<=G2357 and G15224;
	G18459<=G2331 and G15224;
	G18460<=G2351 and G15224;
	G18461<=G2307 and G15224;
	G18462<=G2361 and G15224;
	G18463<=G2375 and G15224;
	G18464<=G2370 and G15224;
	G18465<=G2384 and G15224;
	G18466<=G2389 and G15224;
	G18467<=G2380 and G15224;
	G18468<=G2393 and G15224;
	G18469<=G2399 and G15224;
	G18470<=G2403 and G15224;
	G18471<=G2407 and G15224;
	G18472<=G2413 and G15224;
	G18473<=G2342 and G15224;
	G18474<=G2287 and G15224;
	G18475<=G12853 and G15426;
	G18476<=G2433 and G15426;
	G18477<=G2429 and G15426;
	G18478<=G2445 and G15426;
	G18479<=G2449 and G15426;
	G18480<=G2437 and G15426;
	G18481<=G2461 and G15426;
	G18482<=G2472 and G15426;
	G18483<=G2453 and G15426;
	G18484<=G2491 and G15426;
	G18485<=G2465 and G15426;
	G18486<=G2485 and G15426;
	G18487<=G2441 and G15426;
	G18488<=G2495 and G15426;
	G18489<=G2509 and G15426;
	G18490<=G2504 and G15426;
	G18491<=G2518 and G15426;
	G18492<=G2523 and G15426;
	G18493<=G2514 and G15426;
	G18494<=G2527 and G15426;
	G18495<=G2533 and G15426;
	G18496<=G2537 and G15426;
	G18497<=G2541 and G15426;
	G18498<=G2547 and G15426;
	G18499<=G2476 and G15426;
	G18500<=G2421 and G15426;
	G18501<=G12854 and G15509;
	G18502<=G2567 and G15509;
	G18503<=G2563 and G15509;
	G18504<=G2579 and G15509;
	G18505<=G2583 and G15509;
	G18506<=G2571 and G15509;
	G18507<=G2595 and G15509;
	G18508<=G2606 and G15509;
	G18509<=G2587 and G15509;
	G18510<=G2625 and G15509;
	G18511<=G2599 and G15509;
	G18512<=G2619 and G15509;
	G18513<=G2575 and G15509;
	G18514<=G2629 and G15509;
	G18515<=G2643 and G15509;
	G18516<=G2638 and G15509;
	G18517<=G2652 and G15509;
	G18518<=G2657 and G15509;
	G18519<=G2648 and G15509;
	G18520<=G2661 and G15509;
	G18521<=G2667 and G15509;
	G18522<=G2671 and G15509;
	G18523<=G2675 and G15509;
	G18524<=G2681 and G15509;
	G18525<=G2610 and G15509;
	G18526<=G2555 and G15509;
	G18529<=G2712 and G15277;
	G18530<=G2715 and G15277;
	G18531<=G2719 and G15277;
	G18532<=G2724 and G15277;
	G18533<=G2729 and G15277;
	G18534<=G2735 and G15277;
	G18535<=G2741 and G15277;
	G18536<=G2748 and G15277;
	G18537<=G6856 and G15277;
	G18538<=G2759 and G15277;
	G18539<=G2763 and G15277;
	G18540<=G2775 and G15277;
	G18541<=G2767 and G15277;
	G18542<=G2787 and G15277;
	G18543<=G2779 and G15277;
	G18544<=G2791 and G15277;
	G18545<=G2783 and G15277;
	G18546<=G2795 and G15277;
	G18547<=G121 and G15277;
	G18548<=G2807 and G15277;
	G18549<=G2799 and G15277;
	G18550<=G2819 and G15277;
	G18551<=G2811 and G15277;
	G18552<=G2815 and G15277;
	G18553<=G2827 and G15277;
	G18554<=G2831 and G15277;
	G18555<=G2834 and G15277;
	G18556<=G2823 and G15277;
	G18557<=G2771 and G15277;
	G18558<=G2803 and G15277;
	G18559<=G12856 and G15277;
	G18560<=G2837 and G15277;
	G18561<=G2841 and G15277;
	G18563<=G2890 and G16349;
	G18564<=G2844 and G16349;
	G18565<=G2852 and G16349;
	G18566<=G2860 and G16349;
	G18567<=G2894 and G16349;
	G18568<=G37 and G16349;
	G18569<=G94 and G16349;
	G18570<=G2848 and G16349;
	G18571<=G2856 and G16349;
	G18572<=G2864 and G16349;
	G18573<=G2898 and G16349;
	G18574<=G2882 and G16349;
	G18575<=G2878 and G16349;
	G18576<=G2868 and G16349;
	G18577<=G2988 and G16349;
	G18578<=G2873 and G16349;
	G18579<=G2984 and G16349;
	G18580<=G2907 and G16349;
	G18581<=G2912 and G16349;
	G18582<=G2922 and G16349;
	G18583<=G2936 and G16349;
	G18584<=G2950 and G16349;
	G18585<=G2960 and G16349;
	G18586<=G2886 and G16349;
	G18587<=G2980 and G16349;
	G18588<=G2970 and G16349;
	G18589<=G2902 and G16349;
	G18590<=G2917 and G16349;
	G18591<=G2965 and G16349;
	G18592<=G2994 and G16349;
	G18593<=G2999 and G16349;
	G18594<=G12858 and G16349;
	G18595<=G2927 and G16349;
	G18596<=G2941 and G16349;
	G18597<=G2975 and G16349;
	G18598<=G3003 and G16349;
	G18599<=G2955 and G16349;
	G18600<=G3111 and G16987;
	G18601<=G3106 and G16987;
	G18602<=G3115 and G16987;
	G18603<=G3119 and G16987;
	G18604<=G3125 and G16987;
	G18605<=G3129 and G16987;
	G18606<=G3133 and G16987;
	G18607<=G3139 and G16987;
	G18608<=G15087 and G16987;
	G18609<=G3147 and G16987;
	G18610<=G15088 and G17059;
	G18611<=G15090 and G17200;
	G18612<=G3329 and G17200;
	G18613<=G3338 and G17200;
	G18614<=G3343 and G17200;
	G18615<=G3347 and G17200;
	G18616<=G6875 and G17200;
	G18617<=G3462 and G17062;
	G18618<=G3457 and G17062;
	G18619<=G3466 and G17062;
	G18620<=G3470 and G17062;
	G18621<=G3476 and G17062;
	G18622<=G3480 and G17062;
	G18623<=G3484 and G17062;
	G18624<=G3490 and G17062;
	G18625<=G15092 and G17062;
	G18626<=G3498 and G17062;
	G18627<=G15093 and G17093;
	G18628<=G15095 and G17226;
	G18629<=G3680 and G17226;
	G18630<=G3689 and G17226;
	G18631<=G3694 and G17226;
	G18632<=G3698 and G17226;
	G18633<=G6905 and G17226;
	G18634<=G3813 and G17096;
	G18635<=G3808 and G17096;
	G18636<=G3817 and G17096;
	G18637<=G3821 and G17096;
	G18638<=G3827 and G17096;
	G18639<=G3831 and G17096;
	G18640<=G3835 and G17096;
	G18641<=G3841 and G17096;
	G18642<=G15097 and G17096;
	G18643<=G3849 and G17096;
	G18644<=G15098 and G17125;
	G18645<=G15100 and G17271;
	G18646<=G4031 and G17271;
	G18647<=G4040 and G17271;
	G18648<=G4045 and G17271;
	G18649<=G4049 and G17271;
	G18650<=G6928 and G17271;
	G18651<=G15102 and G16249;
	G18652<=G4172 and G16249;
	G18653<=G4176 and G16249;
	G18654<=G4146 and G16249;
	G18655<=G15106 and G14454;
	G18656<=G15120 and G17128;
	G18657<=G4308 and G17128;
	G18658<=G15121 and G17183;
	G18659<=G4366 and G17183;
	G18662<=G15126 and G17367;
	G18663<=G4311 and G17367;
	G18664<=G4332 and G17367;
	G18665<=G4584 and G17367;
	G18666<=G4593 and G17367;
	G18667<=G4601 and G17367;
	G18668<=G4322 and G17367;
	G18669<=G4608 and G17367;
	G18670<=G4621 and G15758;
	G18671<=G4628 and G15758;
	G18672<=G15127 and G15758;
	G18673<=G4643 and G15758;
	G18674<=G4340 and G15758;
	G18675<=G4349 and G15758;
	G18676<=G4358 and G15758;
	G18677<=G4639 and G15758;
	G18678<=G66 and G15758;
	G18679<=G4633 and G15758;
	G18680<=G15128 and G15885;
	G18681<=G4653 and G15885;
	G18682<=G4646 and G15885;
	G18683<=G4674 and G15885;
	G18684<=G4681 and G15885;
	G18685<=G4688 and G15885;
	G18686<=G4659 and G15885;
	G18687<=G4664 and G15885;
	G18688<=G4704 and G16752;
	G18689<=G15129 and G16752;
	G18690<=G15130 and G16053;
	G18691<=G4727 and G16053;
	G18692<=G4732 and G16053;
	G18693<=G4717 and G16053;
	G18694<=G4722 and G16053;
	G18695<=G4737 and G16053;
	G18696<=G4741 and G16053;
	G18697<=G4749 and G16777;
	G18698<=G15131 and G16777;
	G18699<=G4760 and G16816;
	G18700<=G15132 and G16816;
	G18701<=G4771 and G16856;
	G18702<=G15133 and G16856;
	G18703<=G4776 and G16782;
	G18704<=G4793 and G16782;
	G18705<=G4801 and G16782;
	G18706<=G4785 and G16782;
	G18707<=G15134 and G16782;
	G18708<=G4818 and G16782;
	G18709<=G59 and G17302;
	G18710<=G15135 and G17302;
	G18711<=G15136 and G15915;
	G18712<=G4843 and G15915;
	G18713<=G4836 and G15915;
	G18714<=G4864 and G15915;
	G18715<=G4871 and G15915;
	G18716<=G4878 and G15915;
	G18717<=G4849 and G15915;
	G18718<=G4854 and G15915;
	G18719<=G4894 and G16795;
	G18720<=G15137 and G16795;
	G18721<=G15138 and G16077;
	G18722<=G4917 and G16077;
	G18723<=G4922 and G16077;
	G18724<=G4907 and G16077;
	G18725<=G4912 and G16077;
	G18726<=G4927 and G16077;
	G18727<=G4931 and G16077;
	G18728<=G4939 and G16821;
	G18729<=G15139 and G16821;
	G18730<=G4950 and G16861;
	G18731<=G15140 and G16861;
	G18732<=G4961 and G16877;
	G18733<=G15141 and G16877;
	G18734<=G4966 and G16826;
	G18735<=G4983 and G16826;
	G18736<=G4991 and G16826;
	G18737<=G4975 and G16826;
	G18738<=G15142 and G16826;
	G18739<=G5008 and G16826;
	G18740<=G4572 and G17384;
	G18741<=G15143 and G17384;
	G18742<=G5120 and G17847;
	G18743<=G5115 and G17847;
	G18744<=G5124 and G17847;
	G18745<=G5128 and G17847;
	G18746<=G5134 and G17847;
	G18747<=G5138 and G17847;
	G18748<=G5142 and G17847;
	G18749<=G5148 and G17847;
	G18750<=G15145 and G17847;
	G18751<=G5156 and G17847;
	G18752<=G15146 and G17926;
	G18753<=G15148 and G15595;
	G18754<=G5339 and G15595;
	G18755<=G5343 and G15595;
	G18756<=G5348 and G15595;
	G18757<=G5352 and G15595;
	G18758<=G7004 and G15595;
	G18759<=G5467 and G17929;
	G18760<=G5462 and G17929;
	G18761<=G5471 and G17929;
	G18762<=G5475 and G17929;
	G18763<=G5481 and G17929;
	G18764<=G5485 and G17929;
	G18765<=G5489 and G17929;
	G18766<=G5495 and G17929;
	G18767<=G15150 and G17929;
	G18768<=G5503 and G17929;
	G18769<=G15151 and G18062;
	G18770<=G15153 and G15615;
	G18771<=G5685 and G15615;
	G18772<=G5689 and G15615;
	G18773<=G5694 and G15615;
	G18774<=G5698 and G15615;
	G18775<=G7028 and G15615;
	G18776<=G5813 and G18065;
	G18777<=G5808 and G18065;
	G18778<=G5817 and G18065;
	G18779<=G5821 and G18065;
	G18780<=G5827 and G18065;
	G18781<=G5831 and G18065;
	G18782<=G5835 and G18065;
	G18783<=G5841 and G18065;
	G18784<=G15155 and G18065;
	G18785<=G5849 and G18065;
	G18786<=G15156 and G15345;
	G18787<=G15158 and G15634;
	G18788<=G6031 and G15634;
	G18789<=G6035 and G15634;
	G18790<=G6040 and G15634;
	G18791<=G6044 and G15634;
	G18792<=G7051 and G15634;
	G18793<=G6159 and G15348;
	G18794<=G6154 and G15348;
	G18795<=G6163 and G15348;
	G18796<=G6167 and G15348;
	G18797<=G6173 and G15348;
	G18798<=G6177 and G15348;
	G18799<=G6181 and G15348;
	G18800<=G6187 and G15348;
	G18801<=G15160 and G15348;
	G18802<=G6195 and G15348;
	G18803<=G15161 and G15480;
	G18804<=G15163 and G15656;
	G18805<=G6377 and G15656;
	G18806<=G6381 and G15656;
	G18807<=G6386 and G15656;
	G18808<=G6390 and G15656;
	G18809<=G7074 and G15656;
	G18810<=G6505 and G15483;
	G18811<=G6500 and G15483;
	G18812<=G6509 and G15483;
	G18813<=G6513 and G15483;
	G18814<=G6519 and G15483;
	G18815<=G6523 and G15483;
	G18816<=G6527 and G15483;
	G18817<=G6533 and G15483;
	G18818<=G15165 and G15483;
	G18819<=G6541 and G15483;
	G18820<=G15166 and G15563;
	G18821<=G15168 and G15680;
	G18822<=G6723 and G15680;
	G18823<=G6727 and G15680;
	G18824<=G6732 and G15680;
	G18825<=G6736 and G15680;
	G18826<=G7097 and G15680;
	G18890<=G10158 and G17625;
	G18893<=G16215 and G16030;
	G18906<=G13568 and G16264;
	G18909<=G16226 and G13570;
	G18910<=G16227 and G16075;
	G18933<=G16237 and G13597;
	G18934<=G3133 and G16096;
	G18935<=G4322 and G15574;
	G18943<=G269 and G16099;
	G18949<=G10183 and G17625;
	G18950<=G11193 and G16123;
	G18951<=G3484 and G16124;
	G18974<=G174 and G16127;
	G18981<=G11206 and G16158;
	G18982<=G3835 and G16159;
	G18987<=G182 and G16162;
	G18992<=G8341 and G16171;
	G18993<=G11224 and G16172;
	G19062<=G446 and G16180;
	G19069<=G8397 and G16186;
	G19139<=G452 and G16195;
	G19145<=G8450 and G16200;
	G19206<=G460 and G16206;
	G19207<=G7803 and G15992;
	G19266<=G246 and G16214;
	G19275<=G7823 and G16044;
	G19333<=G464 and G16223;
	G19350<=G15968 and G13505;
	G19354<=G471 and G16235;
	G19372<=G686 and G16289;
	G19383<=G16893 and G13223;
	G19384<=G667 and G16310;
	G19393<=G691 and G16325;
	G19461<=G11708 and G16846;
	G19462<=G7850 and G14182 and G14177 and G16646;
	G19487<=G499 and G16680;
	G19500<=G504 and G16712;
	G19516<=G7824 and G16097;
	G19521<=G513 and G16739;
	G19536<=G518 and G16768;
	G19540<=G1124 and G15904;
	G19545<=G3147 and G16769;
	G19556<=G11932 and G16809;
	G19560<=G15832 and G1157 and G10893;
	G19564<=G17175 and G13976;
	G19568<=G1467 and G15959;
	G19571<=G3498 and G16812;
	G19578<=G16183 and G11130;
	G19581<=G15843 and G1500 and G10918;
	G19585<=G17180 and G14004;
	G19588<=G3849 and G16853;
	G19594<=G11913 and G17268;
	G19596<=G1094 and G16681;
	G19601<=G16198 and G11149;
	G19610<=G1141 and G16069;
	G19613<=G1437 and G16713;
	G19631<=G1484 and G16093;
	G19637<=G5142 and G16958;
	G19651<=G1111 and G16119;
	G19655<=G2729 and G16966;
	G19656<=G2807 and G15844;
	G19660<=G12001 and G16968;
	G19661<=G5489 and G16969;
	G19671<=G1454 and G16155;
	G19674<=G2819 and G15867;
	G19680<=G12028 and G17013;
	G19681<=G5835 and G17014;
	G19684<=G2735 and G17297;
	G19691<=G9614 and G17085;
	G19692<=G12066 and G17086;
	G19693<=G6181 and G17087;
	G19715<=G9679 and G17120;
	G19716<=G12100 and G17121;
	G19717<=G6527 and G17122;
	G19735<=G9740 and G17135;
	G19736<=G12136 and G17136;
	G19740<=G2783 and G15907;
	G19746<=G9816 and G17147;
	G19749<=G732 and G16646;
	G19752<=G2771 and G15864;
	G19756<=G9899 and G17154;
	G19767<=G16810 and G14203;
	G19768<=G2803 and G15833;
	G19784<=G2775 and G15877;
	G19788<=G9983 and G17216;
	G19791<=G14253 and G17189;
	G19855<=G2787 and G15962;
	G19911<=G14707 and G17748;
	G19914<=G2815 and G15853;
	G19948<=G17515 and G16320;
	G20056<=G16291 and G9007 and G8954 and G8903;
	G20069<=G16312 and G9051 and G9011 and G8955;
	G20084<=G11591 and G16609;
	G20093<=G15372 and G14584;
	G20094<=G8872 and G16631;
	G20095<=G8873 and G16632;
	G20108<=G15508 and G11048;
	G20109<=G17954 and G17616;
	G20112<=G13540 and G16661;
	G20131<=G15170 and G14309;
	G20135<=G16258 and G16695;
	G20152<=G11545 and G16727;
	G20162<=G8737 and G16750;
	G20165<=G5156 and G17733;
	G20171<=G16479 and G10476;
	G20174<=G5503 and G17754;
	G20188<=G5849 and G17772;
	G20193<=G15578 and G17264;
	G20203<=G6195 and G17789;
	G20215<=G16479 and G10476;
	G20218<=G6541 and G17815;
	G20375<=G671 and G16846;
	G20559<=G336 and G15831;
	G20581<=G10801 and G15571;
	G20602<=G10803 and G15580;
	G20628<=G1046 and G15789;
	G20658<=G1389 and G15800;
	G20682<=G16238 and G4646;
	G20739<=G16259 and G4674;
	G20751<=G16260 and G4836;
	G20875<=G16281 and G4681;
	G20887<=G16282 and G4864;
	G20977<=G10123 and G17301;
	G21012<=G16304 and G4688;
	G21024<=G16306 and G4871;
	G21066<=G10043 and G17625;
	G21067<=G10085 and G17625;
	G21163<=G16321 and G4878;
	G21188<=G7666 and G15705;
	G21251<=G13969 and G17470;
	G21276<=G10157 and G17625;
	G21285<=G7857 and G16027;
	G21296<=G7879 and G16072;
	G21298<=G7697 and G15825;
	G21302<=G956 and G15731;
	G21303<=G10120 and G17625;
	G21332<=G996 and G15739;
	G21333<=G1300 and G15740;
	G21347<=G1339 and G15750;
	G21348<=G10121 and G17625;
	G21361<=G7869 and G16066;
	G21378<=G7887 and G16090;
	G21382<=G10086 and G17625;
	G21394<=G13335 and G15799;
	G21404<=G16069 and G13569;
	G21405<=G13377 and G15811;
	G21419<=G16681 and G13595;
	G21420<=G16093 and G13596;
	G21452<=G16119 and G13624;
	G21453<=G16713 and G13625;
	G21464<=G16181 and G10872;
	G21465<=G16155 and G13663;
	G21512<=G16225 and G10881;
	G21513<=G16196 and G10882;
	G21557<=G12980 and G15674;
	G21558<=G15904 and G13729;
	G21559<=G16236 and G10897;
	G21605<=G13005 and G15695;
	G21606<=G15959 and G13763;
	G21699<=G142 and G20283;
	G21700<=G150 and G20283;
	G21701<=G153 and G20283;
	G21702<=G157 and G20283;
	G21703<=G146 and G20283;
	G21704<=G164 and G20283;
	G21705<=G209 and G20283;
	G21706<=G222 and G20283;
	G21707<=G191 and G20283;
	G21708<=G15049 and G20283;
	G21709<=G283 and G20283;
	G21710<=G287 and G20283;
	G21711<=G291 and G20283;
	G21712<=G294 and G20283;
	G21713<=G298 and G20283;
	G21714<=G278 and G20283;
	G21715<=G160 and G20283;
	G21716<=G301 and G20283;
	G21717<=G15051 and G21037;
	G21718<=G370 and G21037;
	G21719<=G358 and G21037;
	G21720<=G376 and G21037;
	G21721<=G385 and G21037;
	G21728<=G3010 and G20330;
	G21729<=G3021 and G20330;
	G21730<=G3025 and G20330;
	G21731<=G3029 and G20330;
	G21732<=G3004 and G20330;
	G21733<=G3034 and G20330;
	G21734<=G3040 and G20330;
	G21735<=G3057 and G20330;
	G21736<=G3065 and G20330;
	G21737<=G3068 and G20330;
	G21738<=G3072 and G20330;
	G21739<=G3080 and G20330;
	G21740<=G3085 and G20330;
	G21741<=G15086 and G20330;
	G21742<=G3050 and G20330;
	G21743<=G3100 and G20330;
	G21744<=G3103 and G20330;
	G21745<=G3017 and G20330;
	G21746<=G3045 and G20330;
	G21747<=G3061 and G20330;
	G21748<=G15089 and G20785;
	G21749<=G3155 and G20785;
	G21750<=G3161 and G20785;
	G21751<=G3167 and G20785;
	G21752<=G3171 and G20785;
	G21753<=G3179 and G20785;
	G21754<=G3195 and G20785;
	G21755<=G3203 and G20785;
	G21756<=G3211 and G20785;
	G21757<=G3187 and G20785;
	G21758<=G3191 and G20785;
	G21759<=G3199 and G20785;
	G21760<=G3207 and G20785;
	G21761<=G3215 and G20785;
	G21762<=G3219 and G20785;
	G21763<=G3223 and G20785;
	G21764<=G3227 and G20785;
	G21765<=G3231 and G20785;
	G21766<=G3235 and G20785;
	G21767<=G3239 and G20785;
	G21768<=G3243 and G20785;
	G21769<=G3247 and G20785;
	G21770<=G3251 and G20785;
	G21771<=G3255 and G20785;
	G21772<=G3259 and G20785;
	G21773<=G3263 and G20785;
	G21774<=G3361 and G20391;
	G21775<=G3372 and G20391;
	G21776<=G3376 and G20391;
	G21777<=G3380 and G20391;
	G21778<=G3355 and G20391;
	G21779<=G3385 and G20391;
	G21780<=G3391 and G20391;
	G21781<=G3408 and G20391;
	G21782<=G3416 and G20391;
	G21783<=G3419 and G20391;
	G21784<=G3423 and G20391;
	G21785<=G3431 and G20391;
	G21786<=G3436 and G20391;
	G21787<=G15091 and G20391;
	G21788<=G3401 and G20391;
	G21789<=G3451 and G20391;
	G21790<=G3454 and G20391;
	G21791<=G3368 and G20391;
	G21792<=G3396 and G20391;
	G21793<=G3412 and G20391;
	G21794<=G15094 and G20924;
	G21795<=G3506 and G20924;
	G21796<=G3512 and G20924;
	G21797<=G3518 and G20924;
	G21798<=G3522 and G20924;
	G21799<=G3530 and G20924;
	G21800<=G3546 and G20924;
	G21801<=G3554 and G20924;
	G21802<=G3562 and G20924;
	G21803<=G3538 and G20924;
	G21804<=G3542 and G20924;
	G21805<=G3550 and G20924;
	G21806<=G3558 and G20924;
	G21807<=G3566 and G20924;
	G21808<=G3570 and G20924;
	G21809<=G3574 and G20924;
	G21810<=G3578 and G20924;
	G21811<=G3582 and G20924;
	G21812<=G3586 and G20924;
	G21813<=G3590 and G20924;
	G21814<=G3594 and G20924;
	G21815<=G3598 and G20924;
	G21816<=G3602 and G20924;
	G21817<=G3606 and G20924;
	G21818<=G3610 and G20924;
	G21819<=G3614 and G20924;
	G21820<=G3712 and G20453;
	G21821<=G3723 and G20453;
	G21822<=G3727 and G20453;
	G21823<=G3731 and G20453;
	G21824<=G3706 and G20453;
	G21825<=G3736 and G20453;
	G21826<=G3742 and G20453;
	G21827<=G3759 and G20453;
	G21828<=G3767 and G20453;
	G21829<=G3770 and G20453;
	G21830<=G3774 and G20453;
	G21831<=G3782 and G20453;
	G21832<=G3787 and G20453;
	G21833<=G15096 and G20453;
	G21834<=G3752 and G20453;
	G21835<=G3802 and G20453;
	G21836<=G3805 and G20453;
	G21837<=G3719 and G20453;
	G21838<=G3747 and G20453;
	G21839<=G3763 and G20453;
	G21840<=G15099 and G21070;
	G21841<=G3857 and G21070;
	G21842<=G3863 and G21070;
	G21843<=G3869 and G21070;
	G21844<=G3873 and G21070;
	G21845<=G3881 and G21070;
	G21846<=G3897 and G21070;
	G21847<=G3905 and G21070;
	G21848<=G3913 and G21070;
	G21849<=G3889 and G21070;
	G21850<=G3893 and G21070;
	G21851<=G3901 and G21070;
	G21852<=G3909 and G21070;
	G21853<=G3917 and G21070;
	G21854<=G3921 and G21070;
	G21855<=G3925 and G21070;
	G21856<=G3929 and G21070;
	G21857<=G3933 and G21070;
	G21858<=G3937 and G21070;
	G21859<=G3941 and G21070;
	G21860<=G3945 and G21070;
	G21861<=G3949 and G21070;
	G21862<=G3953 and G21070;
	G21863<=G3957 and G21070;
	G21864<=G3961 and G21070;
	G21865<=G3965 and G21070;
	G21866<=G4072 and G19801;
	G21867<=G4082 and G19801;
	G21868<=G4076 and G19801;
	G21869<=G4087 and G19801;
	G21870<=G4093 and G19801;
	G21871<=G4108 and G19801;
	G21872<=G4098 and G19801;
	G21873<=G6946 and G19801;
	G21874<=G4112 and G19801;
	G21875<=G4116 and G19801;
	G21876<=G4119 and G19801;
	G21877<=G6888 and G19801;
	G21878<=G4129 and G19801;
	G21879<=G4132 and G19801;
	G21880<=G4135 and G19801;
	G21881<=G4064 and G19801;
	G21882<=G4057 and G19801;
	G21883<=G4141 and G19801;
	G21884<=G4104 and G19801;
	G21885<=G4122 and G19801;
	G21886<=G4153 and G19801;
	G21887<=G15101 and G19801;
	G21888<=G4165 and G19801;
	G21889<=G4169 and G19801;
	G21890<=G4125 and G19801;
	G21906<=G5022 and G21468;
	G21907<=G5033 and G21468;
	G21908<=G5037 and G21468;
	G21909<=G5041 and G21468;
	G21910<=G5016 and G21468;
	G21911<=G5046 and G21468;
	G21912<=G5052 and G21468;
	G21913<=G5069 and G21468;
	G21914<=G5077 and G21468;
	G21915<=G5080 and G21468;
	G21916<=G5084 and G21468;
	G21917<=G5092 and G21468;
	G21918<=G5097 and G21468;
	G21919<=G15144 and G21468;
	G21920<=G5062 and G21468;
	G21921<=G5109 and G21468;
	G21922<=G5112 and G21468;
	G21923<=G5029 and G21468;
	G21924<=G5057 and G21468;
	G21925<=G5073 and G21468;
	G21926<=G15147 and G18997;
	G21927<=G5164 and G18997;
	G21928<=G5170 and G18997;
	G21929<=G5176 and G18997;
	G21930<=G5180 and G18997;
	G21931<=G5188 and G18997;
	G21932<=G5204 and G18997;
	G21933<=G5212 and G18997;
	G21934<=G5220 and G18997;
	G21935<=G5196 and G18997;
	G21936<=G5200 and G18997;
	G21937<=G5208 and G18997;
	G21938<=G5216 and G18997;
	G21939<=G5224 and G18997;
	G21940<=G5228 and G18997;
	G21941<=G5232 and G18997;
	G21942<=G5236 and G18997;
	G21943<=G5240 and G18997;
	G21944<=G5244 and G18997;
	G21945<=G5248 and G18997;
	G21946<=G5252 and G18997;
	G21947<=G5256 and G18997;
	G21948<=G5260 and G18997;
	G21949<=G5264 and G18997;
	G21950<=G5268 and G18997;
	G21951<=G5272 and G18997;
	G21952<=G5366 and G21514;
	G21953<=G5377 and G21514;
	G21954<=G5381 and G21514;
	G21955<=G5385 and G21514;
	G21956<=G5360 and G21514;
	G21957<=G5390 and G21514;
	G21958<=G5396 and G21514;
	G21959<=G5413 and G21514;
	G21960<=G5421 and G21514;
	G21961<=G5424 and G21514;
	G21962<=G5428 and G21514;
	G21963<=G5436 and G21514;
	G21964<=G5441 and G21514;
	G21965<=G15149 and G21514;
	G21966<=G5406 and G21514;
	G21967<=G5456 and G21514;
	G21968<=G5459 and G21514;
	G21969<=G5373 and G21514;
	G21970<=G5401 and G21514;
	G21971<=G5417 and G21514;
	G21972<=G15152 and G19074;
	G21973<=G5511 and G19074;
	G21974<=G5517 and G19074;
	G21975<=G5523 and G19074;
	G21976<=G5527 and G19074;
	G21977<=G5535 and G19074;
	G21978<=G5551 and G19074;
	G21979<=G5559 and G19074;
	G21980<=G5567 and G19074;
	G21981<=G5543 and G19074;
	G21982<=G5547 and G19074;
	G21983<=G5555 and G19074;
	G21984<=G5563 and G19074;
	G21985<=G5571 and G19074;
	G21986<=G5575 and G19074;
	G21987<=G5579 and G19074;
	G21988<=G5583 and G19074;
	G21989<=G5587 and G19074;
	G21990<=G5591 and G19074;
	G21991<=G5595 and G19074;
	G21992<=G5599 and G19074;
	G21993<=G5603 and G19074;
	G21994<=G5607 and G19074;
	G21995<=G5611 and G19074;
	G21996<=G5615 and G19074;
	G21997<=G5619 and G19074;
	G21998<=G5712 and G21562;
	G21999<=G5723 and G21562;
	G22000<=G5727 and G21562;
	G22001<=G5731 and G21562;
	G22002<=G5706 and G21562;
	G22003<=G5736 and G21562;
	G22004<=G5742 and G21562;
	G22005<=G5759 and G21562;
	G22006<=G5767 and G21562;
	G22007<=G5770 and G21562;
	G22008<=G5774 and G21562;
	G22009<=G5782 and G21562;
	G22010<=G5787 and G21562;
	G22011<=G15154 and G21562;
	G22012<=G5752 and G21562;
	G22013<=G5802 and G21562;
	G22014<=G5805 and G21562;
	G22015<=G5719 and G21562;
	G22016<=G5747 and G21562;
	G22017<=G5763 and G21562;
	G22018<=G15157 and G19147;
	G22019<=G5857 and G19147;
	G22020<=G5863 and G19147;
	G22021<=G5869 and G19147;
	G22022<=G5873 and G19147;
	G22023<=G5881 and G19147;
	G22024<=G5897 and G19147;
	G22025<=G5905 and G19147;
	G22026<=G5913 and G19147;
	G22027<=G5889 and G19147;
	G22028<=G5893 and G19147;
	G22029<=G5901 and G19147;
	G22030<=G5909 and G19147;
	G22031<=G5917 and G19147;
	G22032<=G5921 and G19147;
	G22033<=G5925 and G19147;
	G22034<=G5929 and G19147;
	G22035<=G5933 and G19147;
	G22036<=G5937 and G19147;
	G22037<=G5941 and G19147;
	G22038<=G5945 and G19147;
	G22039<=G5949 and G19147;
	G22040<=G5953 and G19147;
	G22041<=G5957 and G19147;
	G22042<=G5961 and G19147;
	G22043<=G5965 and G19147;
	G22044<=G6058 and G21611;
	G22045<=G6069 and G21611;
	G22046<=G6073 and G21611;
	G22047<=G6077 and G21611;
	G22048<=G6052 and G21611;
	G22049<=G6082 and G21611;
	G22050<=G6088 and G21611;
	G22051<=G6105 and G21611;
	G22052<=G6113 and G21611;
	G22053<=G6116 and G21611;
	G22054<=G6120 and G21611;
	G22055<=G6128 and G21611;
	G22056<=G6133 and G21611;
	G22057<=G15159 and G21611;
	G22058<=G6098 and G21611;
	G22059<=G6148 and G21611;
	G22060<=G6151 and G21611;
	G22061<=G6065 and G21611;
	G22062<=G6093 and G21611;
	G22063<=G6109 and G21611;
	G22064<=G15162 and G19210;
	G22065<=G6203 and G19210;
	G22066<=G6209 and G19210;
	G22067<=G6215 and G19210;
	G22068<=G6219 and G19210;
	G22069<=G6227 and G19210;
	G22070<=G6243 and G19210;
	G22071<=G6251 and G19210;
	G22072<=G6259 and G19210;
	G22073<=G6235 and G19210;
	G22074<=G6239 and G19210;
	G22075<=G6247 and G19210;
	G22076<=G6255 and G19210;
	G22077<=G6263 and G19210;
	G22078<=G6267 and G19210;
	G22079<=G6271 and G19210;
	G22080<=G6275 and G19210;
	G22081<=G6279 and G19210;
	G22082<=G6283 and G19210;
	G22083<=G6287 and G19210;
	G22084<=G6291 and G19210;
	G22085<=G6295 and G19210;
	G22086<=G6299 and G19210;
	G22087<=G6303 and G19210;
	G22088<=G6307 and G19210;
	G22089<=G6311 and G19210;
	G22090<=G6404 and G18833;
	G22091<=G6415 and G18833;
	G22092<=G6419 and G18833;
	G22093<=G6423 and G18833;
	G22094<=G6398 and G18833;
	G22095<=G6428 and G18833;
	G22096<=G6434 and G18833;
	G22097<=G6451 and G18833;
	G22098<=G6459 and G18833;
	G22099<=G6462 and G18833;
	G22100<=G6466 and G18833;
	G22101<=G6474 and G18833;
	G22102<=G6479 and G18833;
	G22103<=G15164 and G18833;
	G22104<=G6444 and G18833;
	G22105<=G6494 and G18833;
	G22106<=G6497 and G18833;
	G22107<=G6411 and G18833;
	G22108<=G6439 and G18833;
	G22109<=G6455 and G18833;
	G22110<=G15167 and G19277;
	G22111<=G6549 and G19277;
	G22112<=G6555 and G19277;
	G22113<=G6561 and G19277;
	G22114<=G6565 and G19277;
	G22115<=G6573 and G19277;
	G22116<=G6589 and G19277;
	G22117<=G6597 and G19277;
	G22118<=G6605 and G19277;
	G22119<=G6581 and G19277;
	G22120<=G6585 and G19277;
	G22121<=G6593 and G19277;
	G22122<=G6601 and G19277;
	G22123<=G6609 and G19277;
	G22124<=G6613 and G19277;
	G22125<=G6617 and G19277;
	G22126<=G6621 and G19277;
	G22127<=G6625 and G19277;
	G22128<=G6629 and G19277;
	G22129<=G6633 and G19277;
	G22130<=G6637 and G19277;
	G22131<=G6641 and G19277;
	G22132<=G6645 and G19277;
	G22133<=G6649 and G19277;
	G22134<=G6653 and G19277;
	G22135<=G6657 and G19277;
	G22142<=G7957 and G19140;
	G22143<=G19568 and G10971;
	G22145<=G14555 and G18832;
	G22149<=G14581 and G18880;
	G22157<=G14608 and G18892;
	G22158<=G13698 and G19609;
	G22160<=G8005 and G19795;
	G22161<=G13202 and G19071;
	G22165<=G15594 and G18903;
	G22172<=G8064 and G19857;
	G22191<=G8119 and G19875;
	G22193<=G19880 and G20682;
	G22208<=G19906 and G20739;
	G22209<=G19907 and G20751;
	G22216<=G13660 and G20000;
	G22218<=G19951 and G20875;
	G22219<=G19953 and G20887;
	G22298<=G19997 and G21012;
	G22299<=G19999 and G21024;
	G22307<=G20027 and G21163;
	G22308<=G1135 and G19738;
	G22309<=G1478 and G19751;
	G22310<=G19662 and G20235;
	G22316<=G2837 and G20270;
	G22329<=G11940 and G20329;
	G22340<=G19605 and G13522;
	G22342<=G9354 and G9285 and G21287;
	G22369<=G9354 and G7717 and G20783;
	G22384<=G9354 and G9285 and G20784;
	G22417<=G7753 and G9285 and G21186;
	G22432<=G9354 and G7717 and G21187;
	G22457<=G7753 and G7717 and G21288;
	G22472<=G7753 and G9285 and G21289;
	G22489<=G12954 and G19386;
	G22498<=G7753 and G7717 and G21334;
	G22515<=G12981 and G19395;
	G22518<=G12982 and G19398;
	G22525<=G13006 and G19411;
	G22534<=G8766 and G21389;
	G22538<=G14035 and G20248;
	G22588<=G79 and G20078;
	G22589<=G19267 and G19451;
	G22590<=G19274 and G19452;
	G22622<=G19336 and G19469;
	G22623<=G19337 and G19470;
	G22624<=G19344 and G19471;
	G22632<=G19356 and G19476;
	G22633<=G19359 and G19479;
	G22637<=G19363 and G19489;
	G22665<=G17174 and G20905;
	G22670<=G20114 and G9104;
	G22680<=G19530 and G7781;
	G22685<=G11891 and G20192;
	G22686<=G19335 and G19577;
	G22689<=G18918 and G9104;
	G22710<=G19358 and G19600;
	G22717<=G9291 and G20212;
	G22720<=G9253 and G20619;
	G22752<=G15792 and G19612;
	G22760<=G9360 and G20237;
	G22762<=G9305 and G20645;
	G22831<=G19441 and G19629;
	G22834<=G102 and G19630;
	G22835<=G15803 and G19633;
	G22843<=G9429 and G20272;
	G22846<=G9386 and G20676;
	G22848<=G19449 and G19649;
	G22849<=G1227 and G19653;
	G22851<=G496 and G19654;
	G22859<=G9456 and G20734;
	G22861<=G19792 and G19670;
	G22862<=G1570 and G19673;
	G22863<=G9547 and G20388;
	G22871<=G9523 and G20871;
	G22873<=G19854 and G19683;
	G22876<=G20136 and G9104;
	G22899<=G19486 and G19695;
	G22900<=G17137 and G19697;
	G22920<=G19764 and G19719;
	G22937<=G753 and G20540;
	G22938<=G19782 and G19739;
	G22939<=G9708 and G21062;
	G22942<=G9104 and G20219;
	G22982<=G19535 and G19747;
	G22990<=G19555 and G19760;
	G22991<=G645 and G20248;
	G22992<=G1227 and G19765;
	G23006<=G19575 and G19776;
	G23007<=G681 and G20248;
	G23008<=G1570 and G19783;
	G23009<=G20196 and G14219;
	G23023<=G650 and G20248;
	G23025<=G16021 and G19798;
	G23050<=G655 and G20248;
	G23056<=G16052 and G19860;
	G23062<=G718 and G20248;
	G23076<=G19128 and G9104;
	G23083<=G16076 and G19878;
	G23103<=G10143 and G20765;
	G23104<=G661 and G20248;
	G23121<=G19128 and G9104;
	G23130<=G728 and G20248;
	G23131<=G13919 and G19930;
	G23148<=G19128 and G9104;
	G23151<=G18994 and G7162;
	G23165<=G13954 and G19964;
	G23166<=G13959 and G19979;
	G23187<=G13989 and G20010;
	G23188<=G13994 and G20025;
	G23201<=G14027 and G20040;
	G23218<=G20200 and G16530;
	G23220<=G19417 and G20067;
	G23229<=G18994 and G4521;
	G23254<=G20056 and G20110;
	G23265<=G20069 and G20132;
	G23280<=G19417 and G20146;
	G23292<=G19879 and G16726;
	G23293<=G9104 and G19200;
	G23314<=G9104 and G19200;
	G23348<=G15570 and G21393;
	G23349<=G13662 and G20182;
	G23372<=G16448 and G20194;
	G23373<=G13699 and G20195;
	G23381<=G7239 and G21413;
	G23386<=G20034 and G20207;
	G23387<=G16506 and G20211;
	G23389<=G9072 and G19757;
	G23392<=G7247 and G21430;
	G23396<=G20051 and G20229;
	G23397<=G11154 and G20239;
	G23401<=G7262 and G21460;
	G23404<=G20063 and G20247;
	G23407<=G9295 and G20273;
	G23412<=G7297 and G21510;
	G23415<=G20077 and G20320;
	G23416<=G20082 and G20321;
	G23424<=G7345 and G21556;
	G23436<=G676 and G20375;
	G23439<=G13771 and G20452;
	G23451<=G13805 and G20510;
	G23471<=G20148 and G20523;
	G23474<=G13830 and G20533;
	G23475<=G19070 and G8971;
	G23484<=G20160 and G20541;
	G23497<=G20169 and G20569;
	G23498<=G20234 and G12998;
	G23513<=G19430 and G13007;
	G23514<=G20149 and G11829;
	G23531<=G10760 and G18930;
	G23532<=G19400 and G11852;
	G23533<=G19436 and G13015;
	G23540<=G16866 and G20622;
	G23551<=G10793 and G18948;
	G23553<=G19413 and G11875;
	G23554<=G20390 and G13024;
	G23564<=G16882 and G20648;
	G23572<=G20230 and G20656;
	G23577<=G19444 and G13033;
	G23581<=G20183 and G11900;
	G23599<=G19050 and G9104;
	G23606<=G16927 and G20679;
	G23618<=G19388 and G11917;
	G23619<=G19453 and G13045;
	G23639<=G19050 and G9104;
	G23646<=G16959 and G20737;
	G23657<=G19401 and G11941;
	G23658<=G14687 and G20852;
	G23675<=G19050 and G9104;
	G23682<=G16970 and G20874;
	G23690<=G14726 and G20978;
	G23691<=G14731 and G20993;
	G23708<=G19050 and G9104;
	G23724<=G14767 and G21123;
	G23725<=G14772 and G21138;
	G23742<=G19128 and G9104;
	G23754<=G14816 and G21189;
	G23755<=G14821 and G21204;
	G23774<=G14867 and G21252;
	G23775<=G14872 and G21267;
	G23779<=G1105 and G19355;
	G23799<=G14911 and G21279;
	G23801<=G1448 and G19362;
	G23802<=G9104 and G19050;
	G23811<=G4087 and G19364;
	G23828<=G9104 and G19128;
	G23836<=G4129 and G19495;
	G23837<=G21160 and G10804;
	G23854<=G4093 and G19506;
	G23855<=G4112 and G19455;
	G23856<=G4116 and G19483;
	G23857<=G19626 and G7908;
	G23872<=G19389 and G4157;
	G23873<=G21222 and G10815;
	G23884<=G4119 and G19510;
	G23885<=G4132 and G19513;
	G23900<=G1129 and G19408;
	G23901<=G19606 and G7963;
	G23917<=G1472 and G19428;
	G23919<=G4122 and G19546;
	G23920<=G4135 and G19549;
	G23921<=G19379 and G4146;
	G23957<=G4138 and G19589;
	G23958<=G9104 and G19200;
	G23990<=G19610 and G10951;
	G23991<=G19209 and G21428;
	G23996<=G19596 and G10951;
	G23998<=G19631 and G10971;
	G24001<=G19651 and G10951;
	G24002<=G19613 and G10971;
	G24004<=G37 and G21225;
	G24008<=G7909 and G19502;
	G24009<=G19671 and G10971;
	G24011<=G7939 and G19524;
	G24012<=G14496 and G21561;
	G24014<=G7933 and G19063;
	G24015<=G19540 and G10951;
	G24016<=G14528 and G21610;
	G24139<=G17619 and G21653;
	G24140<=G17663 and G21654;
	G24141<=G17657 and G21656;
	G24142<=G17700 and G21657;
	G24143<=G17694 and G21659;
	G24144<=G17727 and G21660;
	G24186<=G18102 and G22722;
	G24187<=G305 and G22722;
	G24188<=G316 and G22722;
	G24189<=G324 and G22722;
	G24190<=G329 and G22722;
	G24191<=G319 and G22722;
	G24192<=G311 and G22722;
	G24193<=G336 and G22722;
	G24194<=G106 and G22722;
	G24195<=G74 and G22722;
	G24196<=G333 and G22722;
	G24197<=G347 and G22722;
	G24198<=G351 and G22722;
	G24199<=G355 and G22722;
	G24217<=G18200 and G22594;
	G24218<=G872 and G22594;
	G24219<=G225 and G22594;
	G24220<=G255 and G22594;
	G24221<=G232 and G22594;
	G24222<=G262 and G22594;
	G24223<=G239 and G22594;
	G24224<=G269 and G22594;
	G24225<=G246 and G22594;
	G24226<=G446 and G22594;
	G24227<=G890 and G22594;
	G24228<=G862 and G22594;
	G24229<=G896 and G22594;
	G24230<=G901 and G22594;
	G24283<=G4411 and G22550;
	G24284<=G4375 and G22550;
	G24285<=G4388 and G22550;
	G24286<=G4405 and G22550;
	G24287<=G4401 and G22550;
	G24288<=G4417 and G22550;
	G24289<=G4427 and G22550;
	G24290<=G4430 and G22550;
	G24291<=G18660 and G22550;
	G24292<=G4443 and G22550;
	G24293<=G4438 and G22550;
	G24294<=G4452 and G22550;
	G24295<=G4434 and G22550;
	G24296<=G4382 and G22550;
	G24297<=G4455 and G22550;
	G24298<=G4392 and G22550;
	G24299<=G4456 and G22550;
	G24300<=G15123 and G22228;
	G24301<=G6961 and G22228;
	G24302<=G15124 and G22228;
	G24303<=G4369 and G22228;
	G24304<=G12875 and G22228;
	G24305<=G4477 and G22228;
	G24306<=G4483 and G22228;
	G24307<=G4486 and G22228;
	G24308<=G4489 and G22228;
	G24309<=G4480 and G22228;
	G24310<=G4495 and G22228;
	G24311<=G4498 and G22228;
	G24312<=G4501 and G22228;
	G24313<=G4504 and G22228;
	G24314<=G4515 and G22228;
	G24315<=G4521 and G22228;
	G24316<=G4527 and G22228;
	G24317<=G4534 and G22228;
	G24318<=G4555 and G22228;
	G24319<=G4561 and G22228;
	G24320<=G6973 and G22228;
	G24321<=G4558 and G22228;
	G24322<=G4423 and G22228;
	G24323<=G4546 and G22228;
	G24324<=G4540 and G22228;
	G24325<=G4543 and G22228;
	G24326<=G4552 and G22228;
	G24327<=G4549 and G22228;
	G24328<=G4567 and G22228;
	G24329<=G4462 and G22228;
	G24330<=G18661 and G22228;
	G24331<=G6977 and G22228;
	G24332<=G4459 and G22228;
	G24333<=G4512 and G22228;
	G24378<=G3106 and G22718;
	G24387<=G3457 and G22761;
	G24392<=G3115 and G23067;
	G24393<=G3808 and G22844;
	G24395<=G4704 and G22845;
	G24399<=G3133 and G23067;
	G24400<=G3466 and G23112;
	G24402<=G4749 and G22857;
	G24403<=G4894 and G22858;
	G24406<=G13623 and G22860;
	G24408<=G23989 and G18946;
	G24409<=G3484 and G23112;
	G24410<=G3817 and G23139;
	G24411<=G4584 and G22161;
	G24415<=G4760 and G22869;
	G24416<=G4939 and G22870;
	G24420<=G23997 and G18980;
	G24421<=G3835 and G23139;
	G24422<=G4771 and G22896;
	G24423<=G4950 and G22897;
	G24427<=G4961 and G22919;
	G24436<=G3125 and G23067;
	G24450<=G3129 and G23067;
	G24451<=G3476 and G23112;
	G24464<=G3480 and G23112;
	G24465<=G3827 and G23139;
	G24467<=G13761 and G23047;
	G24475<=G3831 and G23139;
	G24476<=G18879 and G22330;
	G24482<=G6875 and G23055;
	G24484<=G16288 and G23208;
	G24485<=G10710 and G22319;
	G24488<=G6905 and G23082;
	G24491<=G10727 and G22332;
	G24495<=G6928 and G23127;
	G24498<=G14036 and G23850;
	G24499<=G22217 and G19394;
	G24501<=G14000 and G23182;
	G24502<=G23428 and G13223;
	G24503<=G22225 and G19409;
	G24504<=G22226 and G19410;
	G24507<=G22304 and G19429;
	G24523<=G22318 and G19468;
	G24532<=G22331 and G19478;
	G24536<=G19516 and G22635;
	G24537<=G22626 and G10851;
	G24541<=G22626 and G10851;
	G24545<=G3333 and G23285;
	G24546<=G22447 and G19523;
	G24549<=G23162 and G20887;
	G24550<=G3684 and G23308;
	G24551<=G17148 and G23331;
	G24552<=G22487 and G19538;
	G24553<=G22983 and G19539;
	G24554<=G22490 and G19541;
	G24555<=G23184 and G21024;
	G24556<=G4035 and G23341;
	G24558<=G22516 and G19566;
	G24559<=G22993 and G19567;
	G24564<=G23198 and G21163;
	G24569<=G5115 and G23382;
	G24572<=G5462 and G23393;
	G24573<=G17198 and G23716;
	G24581<=G5124 and G23590;
	G24582<=G5808 and G23402;
	G24588<=G5142 and G23590;
	G24589<=G5471 and G23630;
	G24590<=G6154 and G23413;
	G24600<=G22591 and G19652;
	G24602<=G16507 and G22854;
	G24606<=G5489 and G23630;
	G24607<=G5817 and G23666;
	G24608<=G6500 and G23425;
	G24618<=G22625 and G19672;
	G24622<=G19856 and G22866;
	G24624<=G16524 and G22867;
	G24627<=G22763 and G19679;
	G24628<=G5835 and G23666;
	G24629<=G6163 and G23699;
	G24630<=G23255 and G14149;
	G24634<=G22634 and G19685;
	G24635<=G19874 and G22883;
	G24637<=G16586 and G22884;
	G24638<=G22763 and G19690;
	G24639<=G6181 and G23699;
	G24640<=G6509 and G23733;
	G24642<=G8290 and G22898;
	G24643<=G22636 and G19696;
	G24644<=G11714 and G22903;
	G24645<=G22639 and G19709;
	G24646<=G22640 and G19711;
	G24647<=G19903 and G22907;
	G24649<=G6527 and G23733;
	G24650<=G22641 and G19718;
	G24651<=G2741 and G23472;
	G24654<=G11735 and G22922;
	G24656<=G11736 and G22926;
	G24657<=G22644 and G19730;
	G24658<=G22645 and G19732;
	G24659<=G5134 and G23590;
	G24660<=G22648 and G19737;
	G24663<=G16621 and G22974;
	G24664<=G22652 and G19741;
	G24666<=G11753 and G22975;
	G24668<=G11754 and G22979;
	G24669<=G22653 and G19742;
	G24670<=G5138 and G23590;
	G24671<=G5481 and G23630;
	G24672<=G19534 and G22981;
	G24673<=G22659 and G19748;
	G24674<=G446 and G23496;
	G24675<=G17568 and G22342;
	G24676<=G2748 and G23782;
	G24679<=G13289 and G22985;
	G24680<=G16422 and G22986;
	G24681<=G16653 and G22988;
	G24682<=G22662 and G19754;
	G24684<=G11769 and G22989;
	G24686<=G5485 and G23630;
	G24687<=G5827 and G23666;
	G24688<=G22681 and G22663;
	G24698<=G22664 and G19761;
	G24700<=G645 and G23512;
	G24702<=G17464 and G22342;
	G24703<=G17592 and G22369;
	G24704<=G17593 and G22384;
	G24706<=G15910 and G22996;
	G24707<=G13295 and G22997;
	G24708<=G16474 and G22998;
	G24709<=G16690 and G23000;
	G24710<=G22679 and G19771;
	G24712<=G19592 and G23001;
	G24713<=G5831 and G23666;
	G24714<=G6173 and G23699;
	G24716<=G15935 and G23004;
	G24717<=G22684 and G19777;
	G24719<=G681 and G23530;
	G24721<=G17488 and G22369;
	G24722<=G17618 and G22417;
	G24723<=G17490 and G22384;
	G24724<=G17624 and G22432;
	G24725<=G19587 and G23012;
	G24726<=G15965 and G23015;
	G24727<=G13300 and G23016;
	G24728<=G16513 and G23017;
	G24729<=G22719 and G23018;
	G24730<=G6177 and G23699;
	G24731<=G6519 and G23733;
	G24743<=G22708 and G19789;
	G24745<=G650 and G23550;
	G24747<=G17510 and G22417;
	G24748<=G17656 and G22457;
	G24749<=G17511 and G22432;
	G24750<=G17662 and G22472;
	G24754<=G19604 and G23027;
	G24755<=G16022 and G23030;
	G24757<=G7004 and G23563;
	G24758<=G6523 and G23733;
	G24761<=G22751 and G19852;
	G24762<=G655 and G23573;
	G24763<=G17569 and G22457;
	G24764<=G17570 and G22472;
	G24765<=G17699 and G22498;
	G24769<=G19619 and G23058;
	G24771<=G7028 and G23605;
	G24772<=G16287 and G23061;
	G24773<=G22832 and G19872;
	G24774<=G718 and G23614;
	G24775<=G17594 and G22498;
	G24777<=G11345 and G23066;
	G24785<=G7051 and G23645;
	G24786<=G661 and G23654;
	G24788<=G11384 and G23111;
	G24790<=G7074 and G23681;
	G24794<=G11414 and G23138;
	G24796<=G7097 and G23714;
	G24797<=G22872 and G19960;
	G24803<=G22901 and G20005;
	G24812<=G19662 and G22192;
	G24817<=G22929 and G7235;
	G24820<=G13944 and G23978;
	G24822<=G3010 and G23534 and I24003;
	G24835<=G8720 and G23233;
	G24843<=G3010 and G23211 and I24015;
	G24846<=G3361 and G23555 and I24018;
	G24849<=G4165 and G22227;
	G24855<=G3050 and G23534 and I24027;
	G24858<=G3361 and G23223 and I24030;
	G24861<=G3712 and G23582 and I24033;
	G24864<=G11201 and G22305;
	G24865<=G11323 and G23253;
	G24872<=G23088 and G9104;
	G24881<=G3050 and G23211 and I24048;
	G24884<=G3401 and G23555 and I24051;
	G24887<=G3712 and G23239 and I24054;
	G24892<=G11559 and G23264;
	G24897<=G3401 and G23223 and I24064;
	G24900<=G3752 and G23582 and I24067;
	G24903<=G128 and G23889;
	G24904<=G11761 and G23279;
	G24908<=G3752 and G23239 and I24075;
	G24912<=G23687 and G20682;
	G24913<=G4821 and G23908;
	G24914<=G8721 and G23301;
	G24915<=G23087 and G20158;
	G24921<=G23721 and G20739;
	G24922<=G4831 and G23931;
	G24923<=G23129 and G20167;
	G24929<=G23751 and G20875;
	G24930<=G4826 and G23948;
	G24931<=G23153 and G20178;
	G24939<=G23771 and G21012;
	G24940<=G5011 and G23971;
	G24941<=G23171 and G20190;
	G24945<=G23183 and G20197;
	G24949<=G23796 and G20751;
	G24961<=G23193 and G20209;
	G24962<=G23194 and G20210;
	G24967<=G23197 and G20213;
	G24977<=G23209 and G20232;
	G24983<=G23217 and G20238;
	G24984<=G22929 and G12818;
	G24997<=G22929 and G10419;
	G24998<=G17412 and G23408;
	G25012<=G20644 and G23419;
	G25014<=G17474 and G23420;
	G25026<=G22929 and G10503;
	G25030<=G23251 and G20432;
	G25031<=G20675 and G23432;
	G25033<=G17500 and G23433;
	G25040<=G12738 and G23443;
	G25041<=G23261 and G20494;
	G25042<=G23262 and G20496;
	G25043<=G20733 and G23447;
	G25045<=G17525 and G23448;
	G25050<=G13056 and G22312;
	G25054<=G12778 and G23452;
	G25056<=G12779 and G23456;
	G25057<=G23275 and G20511;
	G25058<=G23276 and G20513;
	G25059<=G20870 and G23460;
	G25061<=G17586 and G23461;
	G25063<=G13078 and G22325;
	G25067<=G4722 and G22885;
	G25068<=G17574 and G23477;
	G25069<=G23296 and G20535;
	G25071<=G12804 and G23478;
	G25076<=G12805 and G23479;
	G25077<=G23297 and G20536;
	G25078<=G23298 and G20538;
	G25079<=G21011 and G23483;
	G25084<=G4737 and G22885;
	G25085<=G4912 and G22908;
	G25086<=G13941 and G23488;
	G25087<=G17307 and G23489;
	G25088<=G17601 and G23491;
	G25089<=G23317 and G20553;
	G25091<=G12830 and G23492;
	G25093<=G12831 and G23493;
	G25094<=G23318 and G20554;
	G25095<=G23319 and G20556;
	G25096<=G23778 and G20560;
	G25102<=G4727 and G22885;
	G25103<=G4927 and G22908;
	G25104<=G16800 and G23504;
	G25105<=G13973 and G23505;
	G25106<=G17391 and G23506;
	G25107<=G17643 and G23508;
	G25108<=G23345 and G20576;
	G25110<=G10427 and G23509;
	G25112<=G10428 and G23510;
	G25113<=G23346 and G20577;
	G25122<=G23374 and G20592;
	G25123<=G4732 and G22885;
	G25124<=G4917 and G22908;
	G25125<=G20187 and G23520;
	G25126<=G16839 and G23523;
	G25127<=G13997 and G23524;
	G25128<=G17418 and G23525;
	G25129<=G17682 and G23527;
	G25130<=G23358 and G20600;
	G25132<=G10497 and G23528;
	G25142<=G4717 and G22885;
	G25143<=G4922 and G22908;
	G25147<=G20202 and G23542;
	G25148<=G16867 and G23545;
	G25149<=G14030 and G23546;
	G25150<=G17480 and G23547;
	G25151<=G17719 and G23549;
	G25152<=G23383 and G20626;
	G25159<=G4907 and G22908;
	G25163<=G20217 and G23566;
	G25164<=G16883 and G23569;
	G25165<=G14062 and G23570;
	G25166<=G17506 and G23571;
	G25173<=G12234 and G23589;
	G25178<=G20241 and G23608;
	G25179<=G16928 and G23611;
	G25181<=G23405 and G20696;
	G25187<=G12296 and G23629;
	G25192<=G20276 and G23648;
	G25201<=G12346 and G23665;
	G25207<=G22513 and G10621;
	G25217<=G12418 and G23698;
	G25223<=G22523 and G10652;
	G25229<=G7636 and G22654;
	G25238<=G12466 and G23732;
	G25285<=G22152 and G13061;
	G25290<=G5022 and G22173 and I24482;
	G25323<=G6888 and G22359;
	G25328<=G5022 and G23764 and I24505;
	G25331<=G5366 and G22194 and I24508;
	G25357<=G23810 and G23786;
	G25366<=G7733 and G22406;
	G25367<=G6946 and G22407;
	G25368<=G6946 and G22408;
	G25371<=G5062 and G22173 and I24524;
	G25374<=G5366 and G23789 and I24527;
	G25377<=G5712 and G22210 and I24530;
	G25408<=G22682 and G9772;
	G25411<=G5062 and G23764 and I24546;
	G25414<=G5406 and G22194 and I24549;
	G25417<=G5712 and G23816 and I24552;
	G25420<=G6058 and G22220 and I24555;
	G25448<=G11202 and G22680;
	G25449<=G6946 and G22496;
	G25450<=G6888 and G22497;
	G25453<=G5406 and G23789 and I24576;
	G25456<=G5752 and G22210 and I24579;
	G25459<=G6058 and G23844 and I24582;
	G25462<=G6404 and G22300 and I24585;
	G25466<=G23574 and G21346;
	G25479<=G22646 and G9917;
	G25482<=G5752 and G23816 and I24597;
	G25485<=G6098 and G22220 and I24600;
	G25488<=G6404 and G23865 and I24603;
	G25491<=G23615 and G21355;
	G25502<=G6946 and G22527;
	G25503<=G6888 and G22529;
	G25507<=G6098 and G23844 and I24616;
	G25510<=G6444 and G22300 and I24619;
	G25518<=G6444 and G23865 and I24625;
	G25522<=G6888 and G22544;
	G25526<=G23720 and G21400;
	G25530<=G23750 and G21414;
	G25536<=G23770 and G21431;
	G25543<=G23795 and G21461;
	G25551<=G23822 and G21511;
	G25559<=G13004 and G22649;
	G25565<=G13013 and G22660;
	G25567<=I24674 and I24675;
	G25568<=I24679 and I24680;
	G25569<=I24684 and I24685;
	G25570<=I24689 and I24690;
	G25571<=I24694 and I24695;
	G25572<=I24699 and I24700;
	G25573<=I24704 and I24705;
	G25574<=I24709 and I24710;
	G25578<=G19402 and G24146;
	G25579<=G19422 and G24147;
	G25580<=G19268 and G24149;
	G25581<=G19338 and G24150;
	G25765<=G24989 and G24973;
	G25768<=G2912 and G24560;
	G25772<=G24944 and G24934;
	G25775<=G2922 and G24568;
	G25780<=G25532 and G25527;
	G25782<=G2936 and G24571;
	G25787<=G24792 and G20887;
	G25788<=G8010 and G24579;
	G25801<=G8097 and G24585;
	G25802<=G8106 and G24586;
	G25803<=G24798 and G21024;
	G25804<=G8069 and G24587;
	G25814<=G24760 and G13323;
	G25815<=G8155 and G24603;
	G25816<=G8164 and G24604;
	G25817<=G24807 and G21163;
	G25818<=G8124 and G24605;
	G25831<=G3151 and G24623;
	G25832<=G8219 and G24625;
	G25833<=G8228 and G24626;
	G25848<=G25539 and G18977;
	G25850<=G3502 and G24636;
	G25852<=G4593 and G24411;
	G25865<=G25545 and G18991;
	G25866<=G3853 and G24648;
	G25870<=G24840 and G16182;
	G25871<=G8334 and G24804;
	G25872<=G3119 and G24655;
	G25873<=G24854 and G16197;
	G25874<=G11118 and G24665;
	G25875<=G8390 and G24809;
	G25876<=G3470 and G24667;
	G25879<=G11135 and G24683;
	G25880<=G8443 and G24814;
	G25881<=G3821 and G24685;
	G25883<=G13728 and G24699;
	G25884<=G11153 and G24711;
	G25900<=G24390 and G19368;
	G25901<=G24853 and G16290;
	G25902<=G24398 and G19373;
	G25904<=G14001 and G24791;
	G25905<=G24879 and G16311;
	G25907<=G24799 and G22519;
	G25908<=G24782 and G22520;
	G25909<=G8745 and G24875;
	G25915<=G24926 and G9602;
	G25916<=G24432 and G19434;
	G25921<=G24936 and G9664;
	G25922<=G24959 and G20065;
	G25923<=G24443 and G19443;
	G25924<=G24976 and G16846;
	G25925<=G24990 and G23234;
	G25926<=G25005 and G24839;
	G25927<=G25004 and G20375;
	G25928<=G25022 and G23436;
	G25931<=G24574 and G19477;
	G25938<=G8997 and G24953;
	G25939<=G24583 and G19490;
	G25946<=G24496 and G19537;
	G25949<=G24701 and G19559;
	G25951<=G24500 and G19565;
	G25955<=G24720 and G19580;
	G25957<=G17190 and G24960;
	G25959<=G1648 and G24963;
	G25961<=G25199 and G20682;
	G25962<=G9258 and G24971;
	G25963<=G1657 and G24978;
	G25964<=G1783 and G24979;
	G25965<=G2208 and G24980;
	G25966<=G9364 and G24985;
	G25967<=G9373 and G24986;
	G25968<=G25215 and G20739;
	G25969<=G9310 and G24987;
	G25970<=G1792 and G24991;
	G25971<=G1917 and G24992;
	G25972<=G2217 and G24993;
	G25973<=G2342 and G24994;
	G25975<=G9434 and G24999;
	G25976<=G9443 and G25000;
	G25977<=G25236 and G20875;
	G25978<=G9391 and G25001;
	G25979<=G24517 and G19650;
	G25980<=G1926 and G25006;
	G25981<=G2051 and G25007;
	G25982<=G2351 and G25008;
	G25983<=G2476 and G25009;
	G25986<=G5160 and G25013;
	G25987<=G9501 and G25015;
	G25988<=G9510 and G25016;
	G25989<=G25258 and G21012;
	G25990<=G9461 and G25017;
	G25991<=G2060 and G25023;
	G25992<=G2485 and G25024;
	G25993<=G2610 and G25025;
	G26019<=G5507 and G25032;
	G26020<=G9559 and G25034;
	G26021<=G9568 and G25035;
	G26022<=G25271 and G20751;
	G26023<=G9528 and G25036;
	G26024<=G2619 and G25039;
	G26048<=G5853 and G25044;
	G26049<=G9621 and G25046;
	G26050<=G9630 and G25047;
	G26051<=G24896 and G14169;
	G26077<=G9607 and G25233;
	G26078<=G5128 and G25055;
	G26079<=G6199 and G25060;
	G26084<=G24926 and G9602;
	G26085<=G11906 and G25070;
	G26086<=G9672 and G25255;
	G26087<=G5475 and G25072;
	G26088<=G6545 and G25080;
	G26090<=G1624 and G25081;
	G26091<=G1691 and G25082;
	G26092<=G9766 and G25083;
	G26094<=G24936 and G9664;
	G26095<=G11923 and G25090;
	G26096<=G9733 and G25268;
	G26097<=G5821 and G25092;
	G26100<=G1677 and G25097;
	G26101<=G1760 and G25098;
	G26102<=G1825 and G25099;
	G26103<=G2185 and G25100;
	G26104<=G2250 and G25101;
	G26119<=G11944 and G25109;
	G26120<=G9809 and G25293;
	G26121<=G6167 and G25111;
	G26122<=G24557 and G19762;
	G26123<=G1696 and G25382;
	G26124<=G1811 and G25116;
	G26125<=G1894 and G25117;
	G26126<=G1959 and G25118;
	G26127<=G2236 and G25119;
	G26128<=G2319 and G25120;
	G26129<=G2384 and G25121;
	G26130<=G24890 and G19772;
	G26145<=G11962 and G25131;
	G26146<=G9892 and G25334;
	G26147<=G6513 and G25133;
	G26148<=G25357 and G11724 and G11709 and G11686;
	G26153<=G24565 and G19780;
	G26154<=G1830 and G25426;
	G26155<=G1945 and G25134;
	G26156<=G2028 and G25135;
	G26157<=G2093 and G25136;
	G26158<=G2255 and G25432;
	G26159<=G2370 and G25137;
	G26160<=G2453 and G25138;
	G26161<=G2518 and G25139;
	G26165<=G11980 and G25153;
	G26166<=G25357 and G11724 and G11709 and G7558;
	G26171<=G25357 and G6856 and G11709 and G11686;
	G26176<=G1964 and G25467;
	G26177<=G2079 and G25154;
	G26178<=G2389 and G25473;
	G26179<=G2504 and G25155;
	G26180<=G2587 and G25156;
	G26181<=G2652 and G25157;
	G26182<=G9978 and G25317;
	G26186<=G24580 and G23031;
	G26190<=G25357 and G11724 and G7586 and G11686;
	G26195<=G25357 and G6856 and G11709 and G7558;
	G26200<=G24688 and G10678 and G10658 and G10627;
	G26203<=G1632 and G25337;
	G26204<=G1720 and G25275;
	G26205<=G2098 and G25492;
	G26206<=G2523 and G25495;
	G26207<=G2638 and G25170;
	G26213<=G25357 and G11724 and G7586 and G7558;
	G26218<=G25357 and G6856 and G7586 and G11686;
	G26223<=G24688 and G10678 and G10658 and G8757;
	G26226<=G24688 and G8812 and G10658 and G10627;
	G26229<=G1724 and G25275;
	G26230<=G1768 and G25385;
	G26231<=G1854 and G25300;
	G26232<=G2193 and G25396;
	G26233<=G2279 and G25309;
	G26234<=G2657 and G25514;
	G26236<=G25357 and G6856 and G7586 and G7558;
	G26241<=G24688 and G10678 and G8778 and G10627;
	G26244<=G24688 and G8812 and G10658 and G8757;
	G26249<=G1858 and G25300;
	G26250<=G1902 and G25429;
	G26251<=G1988 and G25341;
	G26252<=G2283 and G25309;
	G26253<=G2327 and G25435;
	G26254<=G2413 and G25349;
	G26257<=G4253 and G25197;
	G26258<=G12875 and G25231;
	G26259<=G24430 and G25232;
	G26261<=G24688 and G10678 and G8778 and G8757;
	G26264<=G24688 and G8812 and G8778 and G10627;
	G26270<=G1700 and G25275;
	G26271<=G1992 and G25341;
	G26272<=G2036 and G25470;
	G26273<=G2122 and G25389;
	G26274<=G2130 and G25210;
	G26275<=G2417 and G25349;
	G26276<=G2461 and G25476;
	G26277<=G2547 and G25400;
	G26279<=G4249 and G25213;
	G26280<=G13051 and G25248;
	G26281<=G24688 and G8812 and G8778 and G8757;
	G26285<=G1834 and G25300;
	G26286<=G2126 and G25389;
	G26287<=G2138 and G25225;
	G26288<=G2259 and G25309;
	G26289<=G2551 and G25400;
	G26290<=G2595 and G25498;
	G26291<=G2681 and G25439;
	G26292<=G2689 and G25228;
	G26294<=G4245 and G25230;
	G26295<=G13070 and G25266;
	G26300<=G1968 and G25341;
	G26301<=G2145 and G25244;
	G26302<=G2393 and G25349;
	G26303<=G2685 and G25439;
	G26304<=G2697 and G25246;
	G26306<=G13087 and G25286;
	G26307<=G13070 and G25288;
	G26308<=G6961 and G25289;
	G26310<=G2102 and G25389;
	G26311<=G2527 and G25400;
	G26312<=G2704 and G25264;
	G26313<=G12645 and G25326;
	G26323<=G10262 and G25273;
	G26324<=G2661 and G25439;
	G26325<=G12644 and G25370;
	G26336<=G10307 and G25480;
	G26339<=G225 and G24836;
	G26341<=G24746 and G20105;
	G26345<=G13051 and G25505;
	G26347<=G262 and G24850;
	G26350<=G13087 and G25517;
	G26351<=G239 and G24869;
	G26356<=G15581 and G25523;
	G26357<=G22547 and G25525;
	G26358<=G19522 and G25528;
	G26360<=G10589 and G25533;
	G26362<=G19557 and G25538;
	G26378<=G19576 and G25544;
	G26379<=G19904 and G25546;
	G26380<=G19572 and G25547;
	G26381<=G4456 and G25548;
	G26387<=G24813 and G20231;
	G26388<=G19595 and G25552;
	G26389<=G19949 and G25553;
	G26390<=G4423 and G25554;
	G26391<=G19593 and G25555;
	G26393<=G19467 and G25558;
	G26394<=G22530 and G25560;
	G26395<=G22547 and G25561;
	G26397<=G19475 and G25563;
	G26398<=G24946 and G10474;
	G26399<=G15572 and G25566;
	G26423<=G19488 and G24356;
	G26484<=G24946 and G8841;
	G26485<=G24968 and G10502;
	G26486<=G4423 and G24358;
	G26487<=G15702 and G24359;
	G26511<=G19265 and G24364;
	G26513<=G19501 and G24365;
	G26514<=G7400 and G25564;
	G26516<=G24968 and G8876;
	G26517<=G15708 and G24367;
	G26541<=G319 and G24375;
	G26542<=G13102 and G24376;
	G26543<=G12910 and G24377;
	G26544<=G7446 and G24357;
	G26547<=G13283 and G25027;
	G26571<=G10472 and G24386;
	G26572<=G7443 and G24439;
	G26602<=G7487 and G24453;
	G26604<=G13248 and G25051;
	G26606<=G1018 and G24510;
	G26610<=G14198 and G24405;
	G26611<=G24935 and G20580;
	G26612<=G901 and G24407;
	G26613<=G1361 and G24518;
	G26629<=G14173 and G24418;
	G26630<=G7592 and G24419;
	G26633<=G24964 and G20616;
	G26635<=G25321 and G20617;
	G26650<=G10796 and G24424;
	G26651<=G22707 and G24425;
	G26652<=G10799 and G24426;
	G26670<=G13385 and G24428;
	G26671<=G316 and G24429;
	G26684<=G25407 and G20673;
	G26689<=G15754 and G24431;
	G26711<=G25446 and G20713;
	G26712<=G24508 and G24463;
	G26713<=G25447 and G20714;
	G26719<=G10709 and G24438;
	G26749<=G24494 and G23578;
	G26750<=G24514 and G24474;
	G26753<=G16024 and G24452;
	G26778<=G25501 and G20923;
	G26779<=G24497 and G23620;
	G26780<=G4098 and G24437;
	G26783<=G25037 and G21048;
	G26799<=G25247 and G21068;
	G26808<=G25521 and G21185;
	G26815<=G4108 and G24528;
	G26819<=G106 and G24490;
	G26821<=G24821 and G13103;
	G26822<=G24841 and G13116;
	G26823<=G24401 and G13106;
	G26826<=G24907 and G15747;
	G26828<=G24919 and G15756;
	G26829<=G2844 and G24505;
	G26833<=G2852 and G24509;
	G26838<=G2860 and G24515;
	G26839<=G2988 and G24516;
	G26842<=G2894 and G24522;
	G26844<=G25261 and G21418;
	G26845<=G24391 and G21426;
	G26846<=G37 and G24524;
	G26847<=G2873 and G24525;
	G26848<=G2950 and G24526;
	G26849<=G2994 and G24527;
	G26852<=G24975 and G24958;
	G26853<=G94 and G24533;
	G26854<=G2868 and G24534;
	G26855<=G2960 and G24535;
	G26857<=G25062 and G25049;
	G26858<=G2970 and G24540;
	G26861<=G25021 and G25003;
	G26863<=G24974 and G24957;
	G26864<=G2907 and G24548;
	G26871<=G25038 and G25020;
	G26977<=G23032 and G26261 and G26424 and G25550;
	G26994<=G23032 and G26226 and G26424 and G25557;
	G27020<=G4601 and G25852;
	G27025<=G26334 and G7917;
	G27028<=G26342 and G1157;
	G27029<=G26327 and G11031;
	G27030<=G26343 and G7947;
	G27032<=G7704 and G5180 and G5188 and G26200;
	G27033<=G25767 and G19273;
	G27034<=G26328 and G8609;
	G27035<=G26348 and G1500;
	G27036<=G26329 and G11038;
	G27039<=G7738 and G5527 and G5535 and G26223;
	G27040<=G7812 and G6565 and G6573 and G26226;
	G27041<=G8519 and G26330;
	G27042<=G25774 and G19343;
	G27043<=G26335 and G8632;
	G27044<=G7766 and G5873 and G5881 and G26241;
	G27045<=G10295 and G3171 and G3179 and G26244;
	G27050<=G25789 and G22338;
	G27057<=G7791 and G6219 and G6227 and G26261;
	G27058<=G10323 and G3522 and G3530 and G26264;
	G27073<=G7121 and G3873 and G3881 and G26281;
	G27083<=G25819 and G22456;
	G27085<=G25835 and G22494;
	G27086<=G25836 and G22495;
	G27087<=G13872 and G26284;
	G27090<=G25997 and G16423;
	G27094<=G25997 and G16472;
	G27095<=G25997 and G16473;
	G27096<=G26026 and G16475;
	G27097<=G25867 and G22526;
	G27098<=G25868 and G22528;
	G27099<=G14094 and G26352;
	G27103<=G25997 and G16509;
	G27104<=G25997 and G16510;
	G27105<=G26026 and G16511;
	G27106<=G26026 and G16512;
	G27107<=G26055 and G16514;
	G27113<=G25997 and G16522;
	G27114<=G25997 and G16523;
	G27115<=G26026 and G16526;
	G27116<=G26026 and G16527;
	G27117<=G26055 and G16528;
	G27118<=G26055 and G16529;
	G27119<=G25877 and G22542;
	G27120<=G25878 and G22543;
	G27121<=G136 and G26326;
	G27127<=G25997 and G16582;
	G27128<=G25997 and G16583;
	G27129<=G26026 and G16584;
	G27130<=G26026 and G16585;
	G27131<=G26055 and G16588;
	G27132<=G26055 and G16589;
	G27134<=G25997 and G16602;
	G27136<=G26026 and G16605;
	G27137<=G26026 and G16606;
	G27138<=G26055 and G16607;
	G27139<=G26055 and G16608;
	G27140<=G25885 and G22593;
	G27145<=G14121 and G26382;
	G27146<=G26148 and G8187 and G1648;
	G27148<=G25997 and G16622;
	G27149<=G25997 and G16623;
	G27151<=G26026 and G16626;
	G27153<=G26055 and G16629;
	G27154<=G26055 and G16630;
	G27158<=G26609 and G16645;
	G27160<=G14163 and G26340;
	G27161<=G26166 and G8241 and G1783;
	G27162<=G26171 and G8259 and G2208;
	G27177<=G25997 and G16651;
	G27178<=G25997 and G16652;
	G27180<=G26026 and G16654;
	G27181<=G26026 and G16655;
	G27183<=G26055 and G16658;
	G27184<=G26628 and G13756;
	G27185<=G26190 and G8302 and G1917;
	G27186<=G26195 and G8316 and G2342;
	G27201<=G25997 and G16685;
	G27202<=G25997 and G13876;
	G27203<=G26026 and G16688;
	G27204<=G26026 and G16689;
	G27206<=G26055 and G16691;
	G27207<=G26055 and G16692;
	G27208<=G9037 and G26598;
	G27209<=G26213 and G8365 and G2051;
	G27210<=G26218 and G8373 and G2476;
	G27211<=G25997 and G16716;
	G27212<=G25997 and G16717;
	G27213<=G26026 and G16721;
	G27214<=G26026 and G13901;
	G27215<=G26055 and G16724;
	G27216<=G26055 and G16725;
	G27217<=G26236 and G8418 and G2610;
	G27218<=G25997 and G16740;
	G27219<=G26026 and G16742;
	G27220<=G26026 and G16743;
	G27221<=G26055 and G16747;
	G27222<=G26055 and G13932;
	G27227<=G26026 and G16771;
	G27228<=G26055 and G16773;
	G27229<=G26055 and G16774;
	G27230<=G25906 and G19558;
	G27234<=G26055 and G16814;
	G27235<=G25910 and G19579;
	G27246<=G26690 and G26673;
	G27247<=G2759 and G26745;
	G27249<=G25929 and G19678;
	G27251<=G26721 and G26694;
	G27252<=G26733 and G26703;
	G27254<=G25935 and G19688;
	G27255<=G25936 and G19689;
	G27256<=G25937 and G19698;
	G27259<=G26755 and G26725;
	G27260<=G26766 and G26737;
	G27262<=G25997 and G17092;
	G27263<=G25940 and G19713;
	G27264<=G25941 and G19714;
	G27265<=G26785 and G26759;
	G27266<=G26789 and G26770;
	G27267<=G26026 and G17124;
	G27268<=G25942 and G19733;
	G27269<=G25943 and G19734;
	G27270<=G26805 and G26793;
	G27272<=G26055 and G17144;
	G27275<=G25945 and G19745;
	G27276<=G9750 and G26607;
	G27277<=G26359 and G14191;
	G27280<=G9825 and G26614;
	G27281<=G9830 and G26615;
	G27284<=G9908 and G26631;
	G27285<=G9912 and G26632;
	G27286<=G6856 and G26634;
	G27287<=G26545 and G23011;
	G27288<=G26515 and G23013;
	G27291<=G11969 and G26653;
	G27292<=G1714 and G26654;
	G27293<=G9972 and G26655;
	G27294<=G9975 and G26656;
	G27298<=G26573 and G23026;
	G27299<=G26546 and G23028;
	G27300<=G12370 and G26672;
	G27301<=G11992 and G26679;
	G27302<=G1848 and G26680;
	G27303<=G11996 and G26681;
	G27304<=G2273 and G26682;
	G27305<=G10041 and G26683;
	G27309<=G26603 and G23057;
	G27310<=G26574 and G23059;
	G27311<=G12431 and G26693;
	G27312<=G12019 and G26700;
	G27313<=G1982 and G26701;
	G27314<=G12436 and G26702;
	G27315<=G12022 and G26709;
	G27316<=G2407 and G26710;
	G27323<=G26268 and G23086;
	G27324<=G10150 and G26720;
	G27325<=G12478 and G26724;
	G27326<=G12048 and G26731;
	G27327<=G2116 and G26732;
	G27328<=G12482 and G26736;
	G27329<=G12052 and G26743;
	G27330<=G2541 and G26744;
	G27331<=G10177 and G26754;
	G27332<=G12538 and G26758;
	G27333<=G10180 and G26765;
	G27334<=G12539 and G26769;
	G27335<=G12087 and G26776;
	G27336<=G2675 and G26777;
	G27339<=G26400 and G17308;
	G27340<=G10199 and G26784;
	G27341<=G10203 and G26788;
	G27342<=G12592 and G26792;
	G27346<=G26400 and G17389;
	G27347<=G26400 and G17390;
	G27348<=G26488 and G17392;
	G27350<=G10217 and G26803;
	G27351<=G10218 and G26804;
	G27357<=G26400 and G17414;
	G27358<=G26400 and G17415;
	G27359<=G26488 and G17416;
	G27360<=G26488 and G17417;
	G27361<=G26519 and G17419;
	G27362<=G26080 and G20036;
	G27363<=G10231 and G26812;
	G27369<=G25894 and G25324;
	G27370<=G26400 and G17472;
	G27371<=G26400 and G17473;
	G27372<=G26488 and G17476;
	G27373<=G26488 and G17477;
	G27374<=G26519 and G17478;
	G27375<=G26519 and G17479;
	G27376<=G26549 and G17481;
	G27378<=G26089 and G20052;
	G27384<=G26400 and G17496;
	G27385<=G26400 and G17497;
	G27386<=G26488 and G17498;
	G27387<=G26488 and G17499;
	G27388<=G26519 and G17502;
	G27389<=G26519 and G17503;
	G27390<=G26549 and G17504;
	G27391<=G26549 and G17505;
	G27392<=G26576 and G17507;
	G27393<=G26099 and G20066;
	G27395<=G8046 and G26314 and G9187 and G9077;
	G27404<=G26400 and G17518;
	G27406<=G26488 and G17521;
	G27407<=G26488 and G17522;
	G27408<=G26519 and G17523;
	G27409<=G26519 and G17524;
	G27410<=G26549 and G17527;
	G27411<=G26549 and G17528;
	G27412<=G26576 and G17529;
	G27413<=G26576 and G17530;
	G27414<=G255 and G26827;
	G27416<=G8046 and G26314 and G9187 and G504;
	G27421<=G8038 and G26314 and G9187 and G9077;
	G27427<=G26400 and G17575;
	G27428<=G26400 and G17576;
	G27430<=G26488 and G17579;
	G27432<=G26519 and G17582;
	G27433<=G26519 and G17583;
	G27434<=G26549 and G17584;
	G27435<=G26549 and G17585;
	G27436<=G26576 and G17588;
	G27437<=G26576 and G17589;
	G27439<=G232 and G26831;
	G27440<=G8046 and G26314 and G518 and G504;
	G27445<=G8038 and G26314 and G9187 and G504;
	G27451<=G26400 and G17599;
	G27452<=G26400 and G17600;
	G27454<=G26488 and G17602;
	G27455<=G26488 and G17603;
	G27457<=G26519 and G17606;
	G27459<=G26549 and G17609;
	G27460<=G26549 and G17610;
	G27461<=G26576 and G17611;
	G27462<=G26576 and G17612;
	G27467<=G269 and G26832;
	G27469<=G8046 and G26314 and G518 and G9077;
	G27474<=G8038 and G26314 and G518 and G504;
	G27480<=G26400 and G17638;
	G27481<=G26400 and G14630;
	G27482<=G26488 and G17641;
	G27483<=G26488 and G17642;
	G27485<=G26519 and G17644;
	G27486<=G26519 and G17645;
	G27488<=G26549 and G17648;
	G27490<=G26576 and G17651;
	G27491<=G26576 and G17652;
	G27493<=G246 and G26837;
	G27494<=G8038 and G26314 and G518 and G9077;
	G27500<=G26400 and G17672;
	G27501<=G26400 and G17673;
	G27502<=G26488 and G17677;
	G27503<=G26488 and G14668;
	G27504<=G26519 and G17680;
	G27505<=G26519 and G17681;
	G27507<=G26549 and G17683;
	G27508<=G26549 and G17684;
	G27510<=G26576 and G17687;
	G27517<=G26400 and G17707;
	G27518<=G26488 and G17709;
	G27519<=G26488 and G17710;
	G27520<=G26519 and G17714;
	G27521<=G26519 and G14700;
	G27522<=G26549 and G17717;
	G27523<=G26549 and G17718;
	G27525<=G26576 and G17720;
	G27526<=G26576 and G17721;
	G27534<=G26488 and G17735;
	G27535<=G26519 and G17737;
	G27536<=G26519 and G17738;
	G27537<=G26549 and G17742;
	G27538<=G26549 and G14744;
	G27539<=G26576 and G17745;
	G27540<=G26576 and G17746;
	G27541<=G26278 and G23334;
	G27545<=G26519 and G17756;
	G27546<=G26549 and G17758;
	G27547<=G26549 and G17759;
	G27548<=G26576 and G17763;
	G27549<=G26576 and G14785;
	G27553<=G26293 and G23353;
	G27557<=G26549 and G17774;
	G27558<=G26576 and G17776;
	G27559<=G26576 and G17777;
	G27560<=G26299 and G20191;
	G27564<=G26305 and G23378;
	G27568<=G26576 and G17791;
	G27588<=G26690 and G26673;
	G27594<=G26721 and G26694;
	G27595<=G26733 and G26703;
	G27598<=G25899 and G10475;
	G27599<=G26337 and G20033;
	G27600<=G26755 and G26725;
	G27601<=G26766 and G26737;
	G27602<=G23032 and G26244 and G26424 and G24966;
	G27612<=G25887 and G8844;
	G27614<=G26785 and G26759;
	G27615<=G26789 and G26770;
	G27616<=G26349 and G20449;
	G27617<=G23032 and G26264 and G26424 and G24982;
	G27627<=G13266 and G25790;
	G27628<=G26400 and G18061;
	G27633<=G13076 and G25766;
	G27634<=G26805 and G26793;
	G27635<=G23032 and G26281 and G26424 and G24996;
	G27645<=G26488 and G15344;
	G27646<=G13094 and G25773;
	G27648<=G25882 and G8974;
	G27649<=G10820 and G25820;
	G27650<=G26519 and G15479;
	G27651<=G22448 and G25781;
	G27653<=G26549 and G15562;
	G27658<=G22491 and G25786;
	G27660<=G24688 and G26424 and G22763;
	G27661<=G26576 and G15568;
	G27664<=G1024 and G25911;
	G27665<=G26872 and G23519;
	G27666<=G26865 and G23521;
	G27667<=G26361 and G20601;
	G27668<=G1367 and G25917;
	G27669<=G26840 and G13278;
	G27673<=G25769 and G23541;
	G27674<=G26873 and G23543;
	G27676<=G26377 and G20627;
	G27677<=G13021 and G25888;
	G27678<=G947 and G25830;
	G27682<=G25777 and G23565;
	G27683<=G25770 and G23567;
	G27684<=G26386 and G20657;
	G27685<=G13032 and G25895;
	G27686<=G1291 and G25849;
	G27690<=G25784 and G23607;
	G27691<=G25778 and G23609;
	G27692<=G26392 and G20697;
	G27696<=G25800 and G23647;
	G27697<=G25785 and G23649;
	G27699<=G26396 and G20766;
	G27700<=G22342 and G25182 and G26424 and G26148;
	G27710<=G26422 and G20904;
	G27711<=G22369 and G25193 and G26424 and G26166;
	G27714<=G22384 and G25195 and G26424 and G26171;
	G27723<=G26512 and G21049;
	G27724<=G22417 and G25208 and G26424 and G26190;
	G27727<=G22432 and G25211 and G26424 and G26195;
	G27759<=G22457 and G25224 and G26424 and G26213;
	G27762<=G22472 and G25226 and G26424 and G26218;
	G27765<=G4146 and G25886;
	G27817<=G22498 and G25245 and G26424 and G26236;
	G27820<=G7670 and G25932;
	G27821<=G7680 and G25892;
	G27822<=G4157 and G25893;
	G27932<=G25944 and G19369;
	G27957<=G25947 and G15995;
	G27958<=G25950 and G22449;
	G27959<=G25948 and G19374;
	G27962<=G25954 and G19597;
	G27963<=G25952 and G16047;
	G27964<=G25956 and G22492;
	G27965<=G25834 and G13117;
	G27968<=G25958 and G19614;
	G27981<=G26751 and G23924;
	G27988<=G26781 and G23941;
	G27992<=G26800 and G23964;
	G27995<=G26809 and G23985;
	G27997<=G26813 and G23995;
	G27999<=G23032 and G26200 and G26424 and G25529;
	G28010<=G23032 and G26223 and G26424 and G25535;
	G28020<=G23032 and G26241 and G26424 and G25542;
	G28035<=G24103 and I26530 and I26531;
	G28107<=G27970 and G18874;
	G28108<=G7975 and G27237;
	G28110<=G27974 and G18886;
	G28111<=G27343 and G22716;
	G28112<=G27352 and G26162;
	G28113<=G8016 and G27242;
	G28114<=G25869 and G27051;
	G28115<=G27354 and G22759;
	G28116<=G27366 and G26183;
	G28117<=G8075 and G27245;
	G28124<=G27368 and G22842;
	G28125<=G27381 and G26209;
	G28130<=G27353 and G23063;
	G28133<=G27367 and G23108;
	G28136<=G27382 and G23135;
	G28139<=G27337 and G26054;
	G28141<=G10831 and G11797 and G11261 and G27163;
	G28143<=G27344 and G26083;
	G28144<=G4608 and G27020;
	G28148<=G27355 and G26093;
	G28150<=G10862 and G11834 and G11283 and G27187;
	G28151<=G8426 and G27295;
	G28152<=G26297 and G27279;
	G28153<=G26424 and G22763 and G27031;
	G28154<=G8492 and G27306;
	G28158<=G26424 and G22763 and G27037;
	G28159<=G8553 and G27317;
	G28160<=G26309 and G27463;
	G28164<=G8651 and G27528;
	G28165<=G27018 and G22455;
	G28171<=G27016 and G19385;
	G28178<=G27019 and G19397;
	G28182<=G8770 and G27349;
	G28183<=G27024 and G19421;
	G28185<=G27026 and G19435;
	G28192<=G8891 and G27415;
	G28193<=G8851 and G27629;
	G28197<=G27647 and G11344;
	G28198<=G26649 and G27492;
	G28199<=G27479 and G16684;
	G28200<=G27652 and G11383;
	G28201<=G27499 and G16720;
	G28202<=G27659 and G11413;
	G28204<=G26098 and G27654;
	G28205<=G27516 and G16746;
	G28210<=G9229 and G27554;
	G28213<=G27720 and G23380;
	G28214<=G27731 and G26625;
	G28215<=G9264 and G27565;
	G28217<=G27733 and G23391;
	G28218<=G27768 and G26645;
	G28219<=G9316 and G27573;
	G28223<=G27338 and G17194;
	G28224<=G27163 and G22763 and G27064;
	G28225<=G27770 and G23400;
	G28226<=G27825 and G26667;
	G28227<=G9397 and G27583;
	G28228<=G27126 and G19636;
	G28229<=G27345 and G17213;
	G28231<=G27187 and G22763 and G27074;
	G28232<=G27732 and G23586;
	G28233<=G27827 and G23411;
	G28234<=G27877 and G26686;
	G28235<=G9467 and G27592;
	G28236<=G8515 and G27971;
	G28237<=G9492 and G27597;
	G28238<=G27133 and G19658;
	G28239<=G27135 and G19659;
	G28240<=G27356 and G17239;
	G28242<=G27769 and G23626;
	G28243<=G27879 and G23423;
	G28244<=G27926 and G26715;
	G28245<=G11367 and G27975;
	G28246<=G8572 and G27976;
	G28247<=G27147 and G19675;
	G28248<=G27150 and G19676;
	G28249<=G27152 and G19677;
	G28251<=G27826 and G23662;
	G28252<=G27159 and G19682;
	G28253<=G23719 and G27700;
	G28254<=G7268 and G1668 and G27395;
	G28255<=G8515 and G27983;
	G28256<=G11398 and G27984;
	G28257<=G27179 and G19686;
	G28258<=G27182 and G19687;
	G28260<=G27703 and G26518;
	G28261<=G27878 and G23695;
	G28263<=G23747 and G27711;
	G28264<=G7315 and G1802 and G27416;
	G28265<=G11367 and G27989;
	G28266<=G23748 and G27714;
	G28267<=G7328 and G2227 and G27421;
	G28268<=G8572 and G27990;
	G28269<=G27205 and G19712;
	G28272<=G27721 and G26548;
	G28273<=G27927 and G23729;
	G28280<=G23761 and G27724;
	G28281<=G7362 and G1936 and G27440;
	G28282<=G23762 and G27727;
	G28283<=G7380 and G2361 and G27445;
	G28284<=G11398 and G27994;
	G28285<=G9657 and G27717;
	G28289<=G27734 and G26575;
	G28290<=G23780 and G27759;
	G28291<=G7411 and G2070 and G27469;
	G28292<=G23781 and G27762;
	G28293<=G7424 and G2495 and G27474;
	G28299<=G9716 and G27670;
	G28300<=G27771 and G26605;
	G28301<=G27224 and G19750;
	G28302<=G23809 and G27817;
	G28303<=G7462 and G2629 and G27494;
	G28304<=G27226 and G19753;
	G28311<=G9792 and G27679;
	G28312<=G27828 and G26608;
	G28313<=G27231 and G19766;
	G28314<=G27552 and G14205;
	G28315<=G27232 and G19769;
	G28318<=G27233 and G19770;
	G28324<=G9875 and G27687;
	G28327<=G27365 and G19785;
	G28330<=G27238 and G19786;
	G28333<=G27239 and G19787;
	G28339<=G9946 and G27693;
	G28341<=G27240 and G19790;
	G28343<=G27380 and G19799;
	G28346<=G27243 and G19800;
	G28352<=G10014 and G27705;
	G28360<=G27401 and G19861;
	G28415<=G27250 and G19963;
	G28426<=G27257 and G20006;
	G28427<=G27258 and G20008;
	G28439<=G27273 and G10233;
	G28440<=G27274 and G20059;
	G28442<=G27278 and G20072;
	G28451<=G27283 and G20090;
	G28453<=G27582 and G10233;
	G28454<=G26976 and G12233;
	G28455<=G27289 and G20103;
	G28456<=G27290 and G20104;
	G28458<=G27187 and G12730 and G20887 and I26948;
	G28466<=G27960 and G17637;
	G28467<=G26993 and G12295;
	G28471<=G27187 and G12762 and G21024 and I26960;
	G28477<=G27966 and G17676;
	G28478<=G27007 and G12345;
	G28484<=G27187 and G10290 and G21163 and I26972;
	G28488<=G27969 and G17713;
	G28489<=G27010 and G12417;
	G28494<=G27973 and G17741;
	G28495<=G27012 and G12465;
	G28499<=G27982 and G17762;
	G28523<=G27704 and G15585;
	G28524<=G6821 and G27084;
	G28528<=G27187 and G12730;
	G28530<=G27383 and G20240;
	G28531<=G27722 and G15608;
	G28532<=G27394 and G20265;
	G28535<=G11981 and G27088;
	G28537<=G6832 and G27089;
	G28539<=G27187 and G12762;
	G28541<=G27403 and G20274;
	G28542<=G27405 and G20275;
	G28543<=G27735 and G15628;
	G28547<=G6821 and G27091;
	G28550<=G12009 and G27092;
	G28553<=G27187 and G10290;
	G28554<=G27426 and G20372;
	G28555<=G27429 and G20373;
	G28556<=G27431 and G20374;
	G28557<=G27772 and G15647;
	G28558<=G7301 and G27046;
	G28563<=G11981 and G27100;
	G28567<=G6832 and G27101;
	G28569<=G27453 and G20433;
	G28570<=G27456 and G20434;
	G28571<=G27458 and G20435;
	G28572<=G27829 and G15669;
	G28573<=G7349 and G27059;
	G28583<=G12009 and G27112;
	G28585<=G27063 and G10530;
	G28586<=G27484 and G20497;
	G28587<=G27487 and G20498;
	G28588<=G27489 and G20499;
	G28597<=G27515 and G20508;
	G28599<=G27027 and G8922;
	G28601<=G27506 and G20514;
	G28602<=G27509 and G20515;
	G28612<=G27524 and G20539;
	G28616<=G27532 and G20551;
	G28617<=G27533 and G20552;
	G28624<=G22357 and G27009;
	G28626<=G27542 and G20573;
	G28627<=G27543 and G20574;
	G28630<=G27544 and G20575;
	G28637<=G22399 and G27011;
	G28638<=G27551 and G20583;
	G28639<=G27767 and G20597;
	G28642<=G27555 and G20598;
	G28645<=G27556 and G20599;
	G28652<=G27282 and G10288;
	G28653<=G7544 and G27014;
	G28654<=G1030 and G27108;
	G28655<=G27561 and G20603;
	G28657<=G27562 and G20606;
	G28658<=G27563 and G20611;
	G28660<=G27824 and G20623;
	G28663<=G27566 and G20624;
	G28666<=G27567 and G20625;
	G28672<=G7577 and G27017;
	G28673<=G1373 and G27122;
	G28674<=G27569 and G20629;
	G28676<=G27570 and G20632;
	G28677<=G27571 and G20635;
	G28679<=G27572 and G20638;
	G28683<=G27876 and G20649;
	G28686<=G27574 and G20650;
	G28689<=G27575 and G20651;
	G28692<=G27578 and G20661;
	G28694<=G27579 and G20664;
	G28695<=G27580 and G20666;
	G28697<=G27581 and G20669;
	G28703<=G27925 and G20680;
	G28706<=G27584 and G20681;
	G28710<=G27589 and G20703;
	G28712<=G27590 and G20708;
	G28714<=G27591 and G20711;
	G28722<=G27955 and G20738;
	G28725<=G27596 and G20779;
	G28739<=G21434 and G26424 and G25274 and G27395;
	G28761<=G21434 and G26424 and G25299 and G27416;
	G28768<=G21434 and G26424 and G25308 and G27421;
	G28789<=G21434 and G26424 and G25340 and G27440;
	G28799<=G21434 and G26424 and G25348 and G27445;
	G28812<=G26972 and G13037;
	G28813<=G4104 and G27038;
	G28833<=G21434 and G26424 and G25388 and G27469;
	G28846<=G21434 and G26424 and G25399 and G27474;
	G28880<=G21434 and G26424 and G25438 and G27494;
	G28889<=G17292 and G25169 and G26424 and G27395;
	G28919<=G27663 and G21295;
	G28924<=G17317 and G25183 and G26424 and G27416;
	G28939<=G17321 and G25184 and G26424 and G27421;
	G28959<=G17401 and G25194 and G26424 and G27440;
	G28970<=G17405 and G25196 and G26424 and G27445;
	G28982<=G27163 and G12687 and G20682 and I27349;
	G28991<=G14438 and G25209 and G26424 and G27469;
	G28998<=G17424 and G25212 and G26424 and G27474;
	G29008<=G27163 and G12730 and G20739 and I27364;
	G29029<=G14506 and G25227 and G26424 and G27494;
	G29036<=G27163 and G12762 and G20875 and I27381;
	G29073<=G27163 and G10290 and G21012 and I27409;
	G29110<=G27187 and G12687 and G20751 and I27429;
	G29178<=G27163 and G12687;
	G29182<=G27163 and G12730;
	G29188<=G27163 and G12762;
	G29192<=G27163 and G10290;
	G29199<=G27187 and G12687;
	G29201<=G24081 and I27503 and I27504;
	G29202<=G24088 and I27508 and I27509;
	G29203<=G24095 and I27513 and I27514;
	G29204<=G24110 and I27518 and I27519;
	G29205<=G24117 and I27523 and I27524;
	G29206<=G24124 and I27528 and I27529;
	G29207<=G24131 and I27533 and I27534;
	G29208<=G24138 and I27538 and I27539;
	G29314<=G29005 and G22144;
	G29315<=G29188 and G7051 and G5990;
	G29316<=G28528 and G6875 and G3288;
	G29320<=G29068 and G22147;
	G29321<=G29033 and G22148;
	G29322<=G29192 and G7074 and G6336;
	G29323<=G28539 and G6905 and G3639;
	G29324<=G29078 and G18883;
	G29326<=G29105 and G22155;
	G29327<=G29070 and G22156;
	G29328<=G28553 and G6928 and G3990;
	G29329<=G7995 and G28353;
	G29330<=G29114 and G18894;
	G29331<=G29143 and G22169;
	G29332<=G29107 and G22170;
	G29334<=G29148 and G18908;
	G29336<=G4704 and G28363;
	G29337<=G29166 and G22180;
	G29338<=G29145 and G22181;
	G29344<=G29168 and G18932;
	G29345<=G4749 and G28376;
	G29346<=G4894 and G28381;
	G29347<=G29176 and G22201;
	G29349<=G4760 and G28391;
	G29350<=G4939 and G28395;
	G29351<=G4771 and G28406;
	G29352<=G4950 and G28410;
	G29354<=G4961 and G28421;
	G29360<=G27364 and G28294;
	G29362<=G27379 and G28307;
	G29363<=G8458 and G28444;
	G29364<=G27400 and G28321;
	G29367<=G8575 and G28325;
	G29369<=G28209 and G22341;
	G29375<=G13946 and G28370;
	G29376<=G14002 and G28504;
	G29377<=G28132 and G19387;
	G29378<=G28137 and G22493;
	G29380<=G28134 and G19396;
	G29381<=G28135 and G19399;
	G29382<=G26424 and G22763 and G28172;
	G29383<=G28138 and G19412;
	G29384<=G26424 and G22763 and G28179;
	G29475<=G14033 and G28500;
	G29477<=G14090 and G28441;
	G29494<=G9073 and G28479;
	G29509<=G1600 and G28755;
	G29510<=G28856 and G22342;
	G29511<=G1736 and G28783;
	G29512<=G2161 and G28793;
	G29513<=G28448 and G14095;
	G29514<=G1608 and G28780;
	G29515<=G28888 and G22342;
	G29516<=G28895 and G22369;
	G29517<=G1870 and G28827;
	G29518<=G28906 and G22384;
	G29519<=G2295 and G28840;
	G29521<=G1744 and G28824;
	G29522<=G28923 and G22369;
	G29523<=G28930 and G22417;
	G29524<=G2004 and G28864;
	G29525<=G2169 and G28837;
	G29526<=G28938 and G22384;
	G29527<=G28945 and G22432;
	G29528<=G2429 and G28874;
	G29530<=G1612 and G28820;
	G29531<=G1664 and G28559;
	G29532<=G1878 and G28861;
	G29533<=G28958 and G22417;
	G29534<=G28965 and G22457;
	G29535<=G2303 and G28871;
	G29536<=G28969 and G22432;
	G29537<=G28976 and G22472;
	G29538<=G2563 and G28914;
	G29547<=G1748 and G28857;
	G29548<=G1798 and G28575;
	G29549<=G2012 and G28900;
	G29550<=G28990 and G22457;
	G29551<=G2173 and G28867;
	G29552<=G2223 and G28579;
	G29553<=G2437 and G28911;
	G29554<=G28997 and G22472;
	G29555<=G29004 and G22498;
	G29563<=G1616 and G28853;
	G29564<=G1882 and G28896;
	G29565<=G1932 and G28590;
	G29566<=G2307 and G28907;
	G29567<=G2357 and G28593;
	G29568<=G2571 and G28950;
	G29569<=G29028 and G22498;
	G29570<=G2763 and G28598;
	G29571<=G28452 and G11762;
	G29572<=G1620 and G28885;
	G29573<=G1752 and G28892;
	G29574<=G2016 and G28931;
	G29575<=G2066 and G28604;
	G29576<=G2177 and G28903;
	G29577<=G2441 and G28946;
	G29578<=G2491 and G28606;
	G29579<=G28457 and G7964;
	G29580<=G28519 and G14186;
	G29581<=G28462 and G11796;
	G29582<=G27766 and G28608;
	G29584<=G1706 and G29018;
	G29585<=G1756 and G28920;
	G29586<=G1886 and G28927;
	G29587<=G2181 and G28935;
	G29588<=G2311 and G28942;
	G29589<=G2575 and G28977;
	G29590<=G2625 and G28615;
	G29591<=G28552 and G11346;
	G29592<=G28469 and G11832;
	G29593<=G28470 and G7985;
	G29594<=G28529 and G14192;
	G29595<=G28475 and G11833;
	G29596<=G27823 and G28620;
	G29598<=G28823 and G22342;
	G29599<=G1710 and G29018;
	G29600<=G1840 and G29049;
	G29601<=G1890 and G28955;
	G29602<=G2020 and G28962;
	G29603<=G2265 and G29060;
	G29604<=G2315 and G28966;
	G29605<=G2445 and G28973;
	G29606<=G28480 and G8011;
	G29607<=G28509 and G14208;
	G29608<=G28568 and G11385;
	G29609<=G28482 and G11861;
	G29610<=G28483 and G8026;
	G29611<=G28540 and G14209;
	G29612<=G27875 and G28633;
	G29613<=G28208 and G19763;
	G29614<=G28860 and G22369;
	G29615<=G1844 and G29049;
	G29616<=G1974 and G29085;
	G29617<=G2024 and G28987;
	G29618<=G28870 and G22384;
	G29619<=G2269 and G29060;
	G29620<=G2399 and G29097;
	G29621<=G2449 and G28994;
	G29622<=G2579 and G29001;
	G29623<=G28496 and G11563;
	G29624<=G28491 and G8070;
	G29625<=G28514 and G14226;
	G29626<=G28584 and G11415;
	G29627<=G28493 and G11884;
	G29628<=G27924 and G28648;
	G29629<=G28211 and G19779;
	G29630<=G28212 and G19781;
	G29631<=G1682 and G28656;
	G29632<=G28899 and G22417;
	G29633<=G1978 and G29085;
	G29634<=G2108 and G29121;
	G29635<=G28910 and G22432;
	G29636<=G2403 and G29097;
	G29637<=G2533 and G29134;
	G29638<=G2583 and G29025;
	G29639<=G28510 and G11618;
	G29640<=G28498 and G8125;
	G29641<=G28520 and G14237;
	G29642<=G27954 and G28669;
	G29644<=G28216 and G19794;
	G29645<=G1714 and G29018;
	G29646<=G1816 and G28675;
	G29647<=G28934 and G22457;
	G29648<=G2112 and G29121;
	G29649<=G2241 and G28678;
	G29650<=G28949 and G22472;
	G29651<=G2537 and G29134;
	G29652<=G2667 and G29157;
	G29656<=G28515 and G11666;
	G29661<=G1687 and G29015;
	G29662<=G1848 and G29049;
	G29663<=G1950 and G28693;
	G29664<=G2273 and G29060;
	G29665<=G2375 and G28696;
	G29666<=G28980 and G22498;
	G29667<=G2671 and G29157;
	G29668<=G28527 and G14255;
	G29683<=G1821 and G29046;
	G29684<=G1982 and G29085;
	G29685<=G2084 and G28711;
	G29686<=G2246 and G29057;
	G29687<=G2407 and G29097;
	G29688<=G2509 and G28713;
	G29693<=G28207 and G10233;
	G29708<=G1955 and G29082;
	G29709<=G2116 and G29121;
	G29710<=G2380 and G29094;
	G29711<=G2541 and G29134;
	G29712<=G2643 and G28726;
	G29718<=G28512 and G11136;
	G29731<=G2089 and G29118;
	G29732<=G2514 and G29131;
	G29733<=G2675 and G29157;
	G29736<=G28522 and G10233;
	G29740<=G2648 and G29154;
	G29742<=G28288 and G10233;
	G29743<=G28206 and G10233;
	G29746<=G28279 and G20037;
	G29747<=G28286 and G23196;
	G29749<=G28295 and G23214;
	G29750<=G28296 and G23215;
	G29751<=G28297 and G23216;
	G29752<=G28516 and G10233;
	G29757<=G28305 and G23221;
	G29758<=G28306 and G23222;
	G29759<=G28308 and G23226;
	G29760<=G28309 and G23227;
	G29761<=G28310 and G23228;
	G29762<=G28298 and G10233;
	G29766<=G28316 and G23235;
	G29767<=G28317 and G23236;
	G29769<=G28319 and G23237;
	G29770<=G28320 and G23238;
	G29771<=G28322 and G23242;
	G29772<=G28323 and G23243;
	G29773<=G28203 and G10233;
	G29774<=G28287 and G10233;
	G29782<=G28328 and G23245;
	G29783<=G28329 and G23246;
	G29784<=G28331 and G23247;
	G29785<=G28332 and G23248;
	G29787<=G28334 and G23249;
	G29788<=G28335 and G23250;
	G29789<=G28270 and G10233;
	G29794<=G28342 and G23256;
	G29795<=G28344 and G23257;
	G29796<=G28345 and G23258;
	G29797<=G28347 and G23259;
	G29798<=G28348 and G23260;
	G29799<=G28271 and G10233;
	G29803<=G28414 and G26836;
	G29804<=G1592 and G29014;
	G29805<=G28357 and G23270;
	G29806<=G28358 and G23271;
	G29807<=G28359 and G23272;
	G29808<=G28361 and G23273;
	G29809<=G28362 and G23274;
	G29810<=G28259 and G11317;
	G29834<=G28368 and G23278;
	G29835<=G28326 and G24866;
	G29836<=G28425 and G26841;
	G29837<=G28369 and G20144;
	G29838<=G1636 and G29044;
	G29839<=G1728 and G29045;
	G29840<=G2153 and G29056;
	G29841<=G28371 and G23283;
	G29842<=G28372 and G23284;
	G29843<=G28373 and G23289;
	G29844<=G28374 and G23290;
	G29845<=G28375 and G23291;
	G29850<=G28340 and G24893;
	G29851<=G1668 and G29079;
	G29852<=G1772 and G29080;
	G29853<=G1862 and G29081;
	G29854<=G2197 and G29092;
	G29855<=G2287 and G29093;
	G29856<=G28385 and G23303;
	G29857<=G28386 and G23304;
	G29858<=G28387 and G23306;
	G29859<=G28388 and G23307;
	G29860<=G28389 and G23312;
	G29861<=G28390 and G23313;
	G29865<=G1802 and G29115;
	G29866<=G1906 and G29116;
	G29867<=G1996 and G29117;
	G29868<=G2227 and G29128;
	G29869<=G2331 and G29129;
	G29870<=G2421 and G29130;
	G29871<=G28400 and G23332;
	G29872<=G28401 and G23333;
	G29874<=G28402 and G23336;
	G29875<=G28403 and G23337;
	G29876<=G28404 and G23339;
	G29877<=G28405 and G23340;
	G29880<=G1936 and G29149;
	G29881<=G2040 and G29150;
	G29882<=G2361 and G29151;
	G29883<=G2465 and G29152;
	G29884<=G2555 and G29153;
	G29885<=G28416 and G23350;
	G29887<=G28417 and G23351;
	G29888<=G28418 and G23352;
	G29890<=G28419 and G23355;
	G29891<=G28420 and G23356;
	G29894<=G2070 and G29169;
	G29895<=G2495 and G29170;
	G29896<=G2599 and G29171;
	G29899<=G28428 and G23375;
	G29901<=G28429 and G23376;
	G29902<=G28430 and G23377;
	G29907<=G2629 and G29177;
	G29909<=G28435 and G23388;
	G29924<=G13031 and G29190;
	G29926<=G1604 and G28736;
	G29937<=G13044 and G29196;
	G29938<=G23552 and G28889;
	G29940<=G1740 and G28758;
	G29943<=G2165 and G28765;
	G29949<=G23575 and G28924;
	G29951<=G1874 and G28786;
	G29952<=G23576 and G28939;
	G29954<=G2299 and G28796;
	G29959<=G28953 and G12823;
	G29962<=G23616 and G28959;
	G29964<=G2008 and G28830;
	G29966<=G23617 and G28970;
	G29968<=G2433 and G28843;
	G29969<=G28121 and G20509;
	G29973<=G28981 and G9206;
	G29974<=G29173 and G12914;
	G29975<=G28986 and G10420;
	G29979<=G23655 and G28991;
	G29982<=G23656 and G28998;
	G29984<=G2567 and G28877;
	G29985<=G28127 and G20532;
	G29986<=G28468 and G23473;
	G29987<=G29197 and G26424 and G22763;
	G29988<=G29187 and G12235;
	G29989<=G29006 and G10489;
	G29990<=G29007 and G9239;
	G29991<=G29179 and G12922;
	G29992<=G29012 and G10490;
	G30000<=G23685 and G29029;
	G30001<=G28490 and G23486;
	G30002<=G28481 and G23487;
	G30003<=G28149 and G9021;
	G30004<=G28521 and G25837;
	G30005<=G28230 and G24394;
	G30006<=G29032 and G9259;
	G30007<=G29141 and G12929;
	G30008<=G29191 and G12297;
	G30009<=G29034 and G10518;
	G30010<=G29035 and G9274;
	G30011<=G29183 and G12930;
	G30015<=G29040 and G10519;
	G30023<=G28508 and G20570;
	G30024<=G28497 and G23501;
	G30025<=G28492 and G23502;
	G30026<=G28476 and G25064;
	G30027<=G29104 and G12550;
	G30028<=G29069 and G9311;
	G30029<=G29164 and G12936;
	G30030<=G29198 and G12347;
	G30031<=G29071 and G10540;
	G30032<=G29072 and G9326;
	G30033<=G29189 and G12937;
	G30034<=G29077 and G10541;
	G30035<=G22539 and G28120;
	G30041<=G28511 and G23518;
	G30042<=G29142 and G12601;
	G30043<=G29106 and G9392;
	G30044<=G29174 and G12944;
	G30045<=G29200 and G12419;
	G30046<=G29108 and G10564;
	G30047<=G29109 and G9407;
	G30048<=G29193 and G12945;
	G30049<=G13114 and G28167;
	G30050<=G22545 and G28126;
	G30051<=G28513 and G20604;
	G30056<=G29165 and G12659;
	G30057<=G29144 and G9462;
	G30058<=G29180 and G12950;
	G30059<=G28106 and G12467;
	G30060<=G29146 and G10581;
	G30061<=G1036 and G28188;
	G30062<=G13129 and G28174;
	G30064<=G28517 and G20630;
	G30066<=G28518 and G20636;
	G30069<=G29175 and G12708;
	G30070<=G29167 and G9529;
	G30071<=G29184 and G12975;
	G30073<=G1379 and G28194;
	G30075<=G28525 and G20662;
	G30078<=G28526 and G20667;
	G30080<=G28121 and G20674;
	G30082<=G29181 and G12752;
	G30083<=G28533 and G20698;
	G30084<=G28534 and G20700;
	G30086<=G28536 and G20704;
	G30089<=G28538 and G20709;
	G30091<=G28127 and G20716;
	G30094<=G28544 and G20767;
	G30095<=G28545 and G20768;
	G30096<=G28546 and G20770;
	G30098<=G28548 and G20774;
	G30099<=G28549 and G20776;
	G30101<=G28551 and G20780;
	G30107<=G28560 and G20909;
	G30108<=G28561 and G20910;
	G30109<=G28562 and G20912;
	G30110<=G28564 and G20916;
	G30111<=G28565 and G20917;
	G30112<=G28566 and G20919;
	G30118<=G28574 and G21050;
	G30120<=G28576 and G21051;
	G30121<=G28577 and G21052;
	G30122<=G28578 and G21054;
	G30124<=G28580 and G21055;
	G30125<=G28581 and G21056;
	G30126<=G28582 and G21058;
	G30131<=G28589 and G21178;
	G30133<=G28591 and G21179;
	G30135<=G28592 and G21180;
	G30137<=G28594 and G21181;
	G30138<=G28595 and G21182;
	G30139<=G28596 and G21184;
	G30140<=G28600 and G23749;
	G30145<=G28603 and G21247;
	G30149<=G28605 and G21248;
	G30151<=G28607 and G21249;
	G30152<=G28609 and G23767;
	G30153<=G28610 and G23768;
	G30154<=G28611 and G23769;
	G30158<=G28613 and G21274;
	G30161<=G28614 and G21275;
	G30164<=G28618 and G23787;
	G30165<=G28619 and G23788;
	G30166<=G28621 and G23792;
	G30167<=G28622 and G23793;
	G30168<=G28623 and G23794;
	G30172<=G28625 and G21286;
	G30173<=G28118 and G13082;
	G30174<=G28628 and G23812;
	G30175<=G28629 and G23813;
	G30177<=G28631 and G23814;
	G30178<=G28632 and G23815;
	G30179<=G28634 and G23819;
	G30180<=G28635 and G23820;
	G30181<=G28636 and G23821;
	G30185<=G28640 and G23838;
	G30186<=G28641 and G23839;
	G30187<=G28643 and G23840;
	G30188<=G28644 and G23841;
	G30190<=G28646 and G23842;
	G30191<=G28647 and G23843;
	G30192<=G28649 and G23847;
	G30193<=G28650 and G23848;
	G30194<=G28651 and G23849;
	G30196<=G28659 and G23858;
	G30197<=G28661 and G23859;
	G30198<=G28662 and G23860;
	G30199<=G28664 and G23861;
	G30200<=G28665 and G23862;
	G30202<=G28667 and G23863;
	G30203<=G28668 and G23864;
	G30204<=G28670 and G23868;
	G30205<=G28671 and G23869;
	G30207<=G28680 and G23874;
	G30208<=G28681 and G23875;
	G30209<=G28682 and G23876;
	G30210<=G28684 and G23877;
	G30211<=G28685 and G23878;
	G30212<=G28687 and G23879;
	G30213<=G28688 and G23880;
	G30215<=G28690 and G23881;
	G30216<=G28691 and G23882;
	G30219<=G28698 and G23887;
	G30220<=G28699 and G23888;
	G30221<=G28700 and G23893;
	G30222<=G28701 and G23894;
	G30223<=G28702 and G23895;
	G30224<=G28704 and G23896;
	G30225<=G28705 and G23897;
	G30226<=G28707 and G23898;
	G30227<=G28708 and G23899;
	G30228<=G28715 and G23903;
	G30229<=G28716 and G23904;
	G30230<=G28717 and G23906;
	G30231<=G28718 and G23907;
	G30232<=G28719 and G23912;
	G30233<=G28720 and G23913;
	G30234<=G28721 and G23914;
	G30235<=G28723 and G23915;
	G30236<=G28724 and G23916;
	G30238<=G28727 and G23922;
	G30239<=G28728 and G23923;
	G30241<=G28729 and G23926;
	G30242<=G28730 and G23927;
	G30243<=G28731 and G23929;
	G30244<=G28732 and G23930;
	G30245<=G28733 and G23935;
	G30246<=G28734 and G23936;
	G30247<=G28735 and G23937;
	G30248<=G28743 and G23938;
	G30250<=G28744 and G23939;
	G30251<=G28745 and G23940;
	G30253<=G28746 and G23943;
	G30254<=G28747 and G23944;
	G30255<=G28748 and G23946;
	G30256<=G28749 and G23947;
	G30257<=G28750 and G23952;
	G30258<=G28751 and G23953;
	G30261<=G28772 and G23961;
	G30263<=G28773 and G23962;
	G30264<=G28774 and G23963;
	G30266<=G28775 and G23966;
	G30267<=G28776 and G23967;
	G30268<=G28777 and G23969;
	G30269<=G28778 and G23970;
	G30272<=G28814 and G23982;
	G30274<=G28815 and G23983;
	G30275<=G28816 and G23984;
	G30277<=G28817 and G23987;
	G30278<=G28818 and G23988;
	G30281<=G28850 and G23992;
	G30283<=G28851 and G23993;
	G30284<=G28852 and G23994;
	G30289<=G28884 and G24000;
	G30308<=G29178 and G7004 and G5297;
	G30315<=G29182 and G7028 and G5644;
	G30316<=G29199 and G7097 and G6682;
	G30564<=G21358 and G29385;
	G30566<=G26247 and G29507;
	G30576<=G18898 and G29800;
	G30577<=G26267 and G29679;
	G30583<=G19666 and G29355;
	G30589<=G18898 and G29811;
	G30590<=G18911 and G29812;
	G30592<=G30270 and G18929;
	G30594<=G18898 and G29846;
	G30595<=G18911 and G29847;
	G30596<=G30279 and G18947;
	G30598<=G18898 and G29862;
	G30599<=G18911 and G29863;
	G30600<=G30287 and G18975;
	G30604<=G18911 and G29878;
	G30607<=G30291 and G18989;
	G30612<=G26338 and G29597;
	G30614<=G20154 and G29814;
	G30670<=G11330 and G29359;
	G30671<=G29319 and G22317;
	G30673<=G20175 and G29814;
	G30730<=G26346 and G29778;
	G30731<=G11374 and G29361;
	G30735<=G29814 and G22319;
	G30825<=G29814 and G22332;
	G30914<=G29873 and G20887;
	G30915<=G29886 and G24778;
	G30918<=G8681 and G29707;
	G30919<=G29898 and G23286;
	G30920<=G29889 and G21024;
	G30921<=G29900 and G24789;
	G30925<=G29908 and G23309;
	G30926<=G29903 and G21163;
	G30927<=G29910 and G24795;
	G30930<=G29915 and G23342;
	G30935<=G8808 and G29745;
	G30936<=G8830 and G29916;
	G30937<=G22626 and G29814;
	G30982<=G8895 and G29933;
	G31015<=G29476 and G22758;
	G31016<=G29478 and G22840;
	G31017<=G29479 and G22841;
	G31018<=G29480 and G22855;
	G31019<=G29481 and G22856;
	G31021<=G26025 and G29814;
	G31066<=G29483 and G22865;
	G31067<=G29484 and G22868;
	G31069<=G29793 and G14150;
	G31070<=G29814 and G25985;
	G31115<=G29487 and G22882;
	G31118<=G29490 and G22906;
	G31120<=G1700 and G29976;
	G31122<=G12144 and G29993;
	G31123<=G1834 and G29994;
	G31124<=G2259 and G29997;
	G31125<=G29502 and G22973;
	G31128<=G12187 and G30016;
	G31129<=G1968 and G30017;
	G31130<=G12191 and G30019;
	G31131<=G2393 and G30020;
	G31132<=G29504 and G22987;
	G31139<=G12221 and G30036;
	G31140<=G2102 and G30037;
	G31141<=G12224 and G30038;
	G31142<=G2527 and G30039;
	G31143<=G29506 and G22999;
	G31145<=G9970 and G30052;
	G31146<=G12285 and G30053;
	G31147<=G12286 and G30054;
	G31148<=G2661 and G30055;
	G31149<=G29508 and G23021;
	G31150<=G1682 and G30063;
	G31151<=G10037 and G30065;
	G31152<=G10039 and G30067;
	G31153<=G12336 and G30068;
	G31154<=G19128 and G29814;
	G31166<=G1816 and G30074;
	G31167<=G10080 and G30076;
	G31168<=G2241 and G30077;
	G31169<=G10083 and G30079;
	G31170<=G19128 and G29814;
	G31182<=G30240 and G20682;
	G31183<=G30249 and G25174;
	G31184<=G1950 and G30085;
	G31185<=G10114 and G30087;
	G31186<=G2375 and G30088;
	G31187<=G10118 and G30090;
	G31188<=G20028 and G29653;
	G31194<=G19128 and G29814;
	G31206<=G30260 and G23890;
	G31207<=G30252 and G20739;
	G31208<=G30262 and G25188;
	G31209<=G2084 and G30097;
	G31210<=G2509 and G30100;
	G31211<=G10156 and G30102;
	G31212<=G20028 and G29669;
	G31218<=G30271 and G23909;
	G31219<=G30265 and G20875;
	G31220<=G30273 and G25202;
	G31222<=G2643 and G30113;
	G31223<=G20028 and G29689;
	G31224<=G30280 and G23932;
	G31225<=G30276 and G21012;
	G31226<=G30282 and G25218;
	G31228<=G20028 and G29713;
	G31229<=G30288 and G23949;
	G31230<=G30285 and G20751;
	G31231<=G30290 and G25239;
	G31232<=G30294 and G23972;
	G31237<=G29366 and G25325;
	G31238<=G29583 and G20053;
	G31240<=G14793 and G30206;
	G31242<=G29373 and G25409;
	G31252<=G29643 and G20101;
	G31261<=G14754 and G30259;
	G31266<=G30129 and G27742;
	G31270<=G29692 and G23282;
	G31271<=G29706 and G23300;
	G31272<=G30117 and G27742;
	G31273<=G30143 and G27779;
	G31275<=G30147 and G27800;
	G31278<=G29716 and G23302;
	G31280<=G29717 and G23305;
	G31281<=G30106 and G27742;
	G31282<=G30130 and G27779;
	G31283<=G30156 and G27837;
	G31285<=G30134 and G27800;
	G31286<=G30159 and G27858;
	G31290<=G29734 and G23335;
	G31292<=G29735 and G23338;
	G31296<=G30119 and G27779;
	G31297<=G30144 and G27837;
	G31298<=G30169 and G27886;
	G31299<=G30123 and G27800;
	G31300<=G30148 and G27858;
	G31301<=G30170 and G27907;
	G31305<=G29741 and G23354;
	G31309<=G30132 and G27837;
	G31310<=G30157 and G27886;
	G31312<=G30136 and G27858;
	G31313<=G30160 and G27907;
	G31314<=G30183 and G27937;
	G31321<=G30146 and G27886;
	G31323<=G30150 and G27907;
	G31324<=G30171 and G27937;
	G31327<=G19200 and G29814;
	G31374<=G29748 and G23390;
	G31376<=G24952 and G29814;
	G31467<=G30162 and G27937;
	G31470<=G29753 and G23398;
	G31471<=G29754 and G23399;
	G31475<=G29756 and G23406;
	G31477<=G29763 and G23409;
	G31478<=G29764 and G23410;
	G31480<=G1644 and G30296;
	G31481<=G29768 and G23417;
	G31484<=G29775 and G23418;
	G31485<=G29776 and G23421;
	G31486<=G29777 and G23422;
	G31488<=G1779 and G30302;
	G31489<=G2204 and G30305;
	G31490<=G29786 and G23429;
	G31492<=G29790 and G23431;
	G31493<=G29791 and G23434;
	G31494<=G29792 and G23435;
	G31495<=G1913 and G30309;
	G31496<=G2338 and G30312;
	G31497<=G20041 and G29930;
	G31499<=G29801 and G23446;
	G31500<=G29802 and G23449;
	G31501<=G2047 and G29310;
	G31502<=G2472 and G29311;
	G31503<=G20041 and G29945;
	G31504<=G29370 and G10553;
	G31505<=G30195 and G24379;
	G31508<=G29813 and G23459;
	G31513<=G2606 and G29318;
	G31514<=G20041 and G29956;
	G31516<=G29848 and G23476;
	G31517<=G29849 and G23482;
	G31518<=G20041 and G29970;
	G31519<=G29864 and G23490;
	G31520<=G29879 and G23507;
	G31523<=G7528 and G29333;
	G31524<=G29897 and G20593;
	G31525<=G29892 and G23526;
	G31526<=G22521 and G29342;
	G31527<=G7553 and G29343;
	G31528<=G19050 and G29814;
	G31540<=G29904 and G23548;
	G31541<=G22536 and G29348;
	G31542<=G19050 and G29814;
	G31554<=G19050 and G29814;
	G31566<=G19050 and G29814;
	G31579<=G19128 and G29814;
	G31654<=G29325 and G13062;
	G31672<=G29814 and G19050;
	G31707<=G30081 and G23886;
	G31710<=G29814 and G19128;
	G31744<=G30092 and G23902;
	G31746<=G30093 and G23905;
	G31750<=G30103 and G23925;
	G31752<=G30104 and G23928;
	G31756<=G30114 and G23942;
	G31758<=G30115 and G23945;
	G31759<=G21291 and G29385;
	G31763<=G30127 and G23965;
	G31765<=G30128 and G23968;
	G31769<=G30141 and G23986;
	G31776<=G21329 and G29385;
	G31777<=G21343 and G29385;
	G31778<=G21369 and G29385;
	G31780<=G30163 and G23999;
	G31784<=G30176 and G24003;
	G31786<=G30189 and G24010;
	G31787<=G21281 and G29385;
	G31788<=G21352 and G29385;
	G31789<=G30201 and G24013;
	G31790<=G21299 and G29385;
	G31792<=G30214 and G24017;
	G31933<=G939 and G30735;
	G31934<=G31670 and G18827;
	G31936<=G31213 and G24005;
	G31940<=G943 and G30735;
	G31941<=G1283 and G30825;
	G31943<=G4717 and G30614;
	G31944<=G31745 and G22146;
	G31948<=G30670 and G18884;
	G31949<=G1287 and G30825;
	G31959<=G4907 and G30673;
	G31960<=G31749 and G22153;
	G31961<=G31751 and G22154;
	G31962<=G8033 and G31013;
	G31963<=G30731 and G18895;
	G31966<=G31754 and G22166;
	G31967<=G31755 and G22167;
	G31968<=G31757 and G22168;
	G31969<=G31189 and G22139;
	G31974<=G31760 and G22176;
	G31975<=G31761 and G22177;
	G31976<=G31762 and G22178;
	G31977<=G31764 and G22179;
	G31985<=G4722 and G30614;
	G31986<=G31766 and G22197;
	G31987<=G31767 and G22198;
	G31988<=G31768 and G22199;
	G31989<=G31770 and G22200;
	G31990<=G31772 and G18945;
	G31991<=G4912 and G30673;
	G31992<=G31773 and G22213;
	G31993<=G31774 and G22214;
	G31994<=G31775 and G22215;
	G31995<=G28274 and G30569;
	G31996<=G31779 and G18979;
	G32008<=G31781 and G22223;
	G32009<=G31782 and G22224;
	G32010<=G31785 and G22303;
	G32011<=G8287 and G31134;
	G32012<=G8297 and G31233;
	G32013<=G8673 and G30614;
	G32014<=G8715 and G30673;
	G32016<=G8522 and G31138;
	G32018<=G4146 and G30937;
	G32019<=G30579 and G22358;
	G32020<=G4157 and G30937;
	G32028<=G30569 and G29339;
	G32029<=G31318 and G16482;
	G32030<=G4172 and G30937;
	G32031<=G31372 and G13464;
	G32032<=G31373 and G16515;
	G32034<=G14124 and G31239;
	G32035<=G4176 and G30937;
	G32036<=G31469 and G13486;
	G32039<=G31476 and G20070;
	G32040<=G14122 and G31243;
	G32041<=G13913 and G31262;
	G32042<=G27244 and G31070;
	G32043<=G31482 and G16173;
	G32044<=G31483 and G20085;
	G32045<=G31491 and G16187;
	G32046<=G10925 and G30735;
	G32047<=G27248 and G31070;
	G32048<=G31498 and G13869;
	G32049<=G10902 and G30735;
	G32050<=G11003 and G30825;
	G32051<=G31506 and G10831;
	G32052<=G31507 and G13885;
	G32053<=G14176 and G31509;
	G32054<=G10890 and G30735;
	G32055<=G10999 and G30825;
	G32056<=G27271 and G31021;
	G32067<=G4727 and G30614;
	G32068<=G31515 and G10862;
	G32069<=G10878 and G30735;
	G32070<=G10967 and G30825;
	G32071<=G27236 and G31070;
	G32082<=G4917 and G30673;
	G32083<=G947 and G30735;
	G32084<=G10948 and G30825;
	G32085<=G27253 and G31021;
	G32086<=G7597 and G30735;
	G32087<=G1291 and G30825;
	G32088<=G27241 and G31070;
	G32089<=G27261 and G31021;
	G32095<=G7619 and G30825;
	G32096<=G31601 and G29893;
	G32097<=G25960 and G31021;
	G32098<=G4732 and G30614;
	G32103<=G31609 and G29905;
	G32104<=G31616 and G29906;
	G32105<=G4922 and G30673;
	G32106<=G31601 and G29911;
	G32107<=G31624 and G29912;
	G32108<=G31631 and G29913;
	G32109<=G31609 and G29920;
	G32110<=G31639 and G29921;
	G32111<=G31616 and G29922;
	G32112<=G31646 and G29923;
	G32113<=G31601 and G29925;
	G32114<=G31624 and G29927;
	G32115<=G31631 and G29928;
	G32116<=G31658 and G29929;
	G32119<=G31609 and G29939;
	G32120<=G31639 and G29941;
	G32121<=G31616 and G29942;
	G32122<=G31646 and G29944;
	G32126<=G31601 and G29948;
	G32127<=G31624 and G29950;
	G32128<=G31631 and G29953;
	G32129<=G31658 and G29955;
	G32139<=G31601 and G29960;
	G32140<=G31609 and G29961;
	G32141<=G31639 and G29963;
	G32142<=G31616 and G29965;
	G32143<=G31646 and G29967;
	G32145<=G31609 and G29977;
	G32146<=G31624 and G29978;
	G32147<=G31616 and G29980;
	G32148<=G31631 and G29981;
	G32149<=G31658 and G29983;
	G32150<=G31624 and G29995;
	G32151<=G31639 and G29996;
	G32152<=G31631 and G29998;
	G32153<=G31646 and G29999;
	G32154<=G31277 and G14184;
	G32156<=G31639 and G30018;
	G32157<=G31646 and G30021;
	G32158<=G31658 and G30022;
	G32159<=G31658 and G30040;
	G32160<=G31001 and G22995;
	G32161<=G3151 and G31154;
	G32162<=G31002 and G23014;
	G32163<=G3502 and G31170;
	G32164<=G30733 and G25171;
	G32165<=G31669 and G27742;
	G32166<=G31007 and G23029;
	G32167<=G3853 and G31194;
	G32168<=G30597 and G25185;
	G32169<=G31014 and G23046;
	G32170<=G31671 and G27779;
	G32171<=G31706 and G27800;
	G32172<=G2767 and G31608;
	G32173<=G160 and G31134;
	G32174<=G31708 and G27837;
	G32175<=G31709 and G27858;
	G32176<=G2779 and G31623;
	G32177<=G30608 and G25214;
	G32178<=G31747 and G27886;
	G32179<=G31748 and G27907;
	G32180<=G2791 and G31638;
	G32181<=G31020 and G19912;
	G32182<=G31753 and G27937;
	G32183<=G2795 and G31653;
	G32184<=G30611 and G25249;
	G32187<=G30672 and G25287;
	G32188<=G27586 and G31376;
	G32189<=G30824 and G25369;
	G32190<=G142 and G31233;
	G32191<=G27593 and G31376;
	G32193<=G30732 and G25410;
	G32194<=G30601 and G28436;
	G32195<=G30734 and G25451;
	G32196<=G27587 and G31376;
	G32197<=G31144 and G20088;
	G32198<=G4253 and G31327;
	G32199<=G30916 and G25506;
	G32200<=G27468 and G31376;
	G32203<=G4249 and G31327;
	G32204<=G4245 and G31327;
	G32205<=G30922 and G28463;
	G32206<=G30609 and G25524;
	G32207<=G31221 and G23323;
	G32224<=G4300 and G31327;
	G32232<=G31241 and G20266;
	G32234<=G31601 and G30292;
	G32241<=G31244 and G20323;
	G32242<=G31245 and G20324;
	G32244<=G31609 and G30297;
	G32246<=G31246 and G20326;
	G32248<=G31616 and G30299;
	G32254<=G31247 and G20379;
	G32255<=G31248 and G20381;
	G32256<=G31249 and G20382;
	G32258<=G31624 and G30303;
	G32260<=G31250 and G20385;
	G32261<=G31251 and G20386;
	G32263<=G31631 and G30306;
	G32265<=G2799 and G30567;
	G32269<=G31253 and G20443;
	G32270<=G31254 and G20444;
	G32272<=G31639 and G30310;
	G32273<=G31255 and G20446;
	G32274<=G31256 and G20447;
	G32276<=G31646 and G30313;
	G32278<=G2811 and G30572;
	G32281<=G31257 and G20500;
	G32282<=G31258 and G20503;
	G32283<=G31259 and G20506;
	G32284<=G31260 and G20507;
	G32286<=G31658 and G29312;
	G32287<=G2823 and G30578;
	G32290<=G31267 and G20525;
	G32291<=G31268 and G20527;
	G32292<=G31269 and G20530;
	G32293<=G2827 and G30593;
	G32295<=G27931 and G31376;
	G32300<=G31274 and G20544;
	G32301<=G31276 and G20547;
	G32302<=G31279 and G23485;
	G32303<=G27550 and G31376;
	G32304<=G31284 and G20564;
	G32305<=G31287 and G20567;
	G32306<=G31289 and G23499;
	G32307<=G31291 and G23500;
	G32308<=G31293 and G23503;
	G32309<=G5160 and G31528;
	G32310<=G27577 and G31376;
	G32311<=G31295 and G20582;
	G32312<=G31302 and G20591;
	G32313<=G31303 and G23515;
	G32314<=G31304 and G23516;
	G32315<=G31306 and G23517;
	G32316<=G31307 and G23522;
	G32317<=G5507 and G31542;
	G32321<=G27613 and G31376;
	G32322<=G31308 and G20605;
	G32323<=G31311 and G20610;
	G32324<=G31315 and G23537;
	G32325<=G31316 and G23538;
	G32326<=G31317 and G23539;
	G32327<=G31319 and G23544;
	G32328<=G5853 and G31554;
	G32330<=G31320 and G20631;
	G32331<=G31322 and G20637;
	G32332<=G31325 and G23558;
	G32333<=G31326 and G23559;
	G32334<=G31375 and G23568;
	G32335<=G6199 and G31566;
	G32336<=G31596 and G11842;
	G32337<=G31465 and G20663;
	G32338<=G31466 and G20668;
	G32339<=G31474 and G20672;
	G32340<=G31468 and G23585;
	G32341<=G31472 and G23610;
	G32342<=G6545 and G31579;
	G32343<=G31473 and G20710;
	G32345<=G2138 and G31672;
	G32348<=G2145 and G31672;
	G32350<=G2697 and G31710;
	G32356<=G2704 and G31710;
	G32369<=G2130 and G31672;
	G32376<=G2689 and G31710;
	G32396<=G4698 and G30983;
	G32397<=G31068 and G15830;
	G32400<=G4743 and G30989;
	G32401<=G31116 and G13432;
	G32402<=G4888 and G30990;
	G32403<=G31117 and G15842;
	G32409<=G4754 and G30996;
	G32410<=G4933 and G30997;
	G32411<=G31119 and G13469;
	G32412<=G4765 and G30998;
	G32413<=G31121 and G19518;
	G32414<=G4944 and G30999;
	G32418<=G31126 and G16239;
	G32419<=G4955 and G31000;
	G32420<=G31127 and G19533;
	G32425<=G31668 and G21604;
	G32428<=G31133 and G16261;
	G33071<=G31591 and G32404;
	G33073<=G32386 and G18828;
	G33074<=G32387 and G18830;
	G33081<=G32388 and G18875;
	G33082<=G32389 and G18877;
	G33086<=G32390 and G18887;
	G33087<=G32391 and G18888;
	G33091<=G32392 and G18897;
	G33099<=G32395 and G18944;
	G33101<=G32398 and G18976;
	G33102<=G32399 and G18978;
	G33104<=G26296 and G32137;
	G33105<=G26298 and G32138;
	G33106<=G32408 and G18990;
	G33110<=G32404 and G32415;
	G33111<=G24005 and G32421;
	G33113<=G31964 and G22339;
	G33114<=G22139 and G31945;
	G33121<=G8748 and G32212;
	G33122<=G8859 and G32192;
	G33124<=G8945 and G32296;
	G33126<=G9044 and G32201;
	G33186<=G32037 and G22830;
	G33233<=G32094 and G23005;
	G33237<=G32394 and G25198;
	G33239<=G32117 and G19902;
	G33241<=G32173 and G23128;
	G33242<=G32123 and G19931;
	G33243<=G32124 and G19947;
	G33244<=G32190 and G23152;
	G33245<=G32125 and G19961;
	G33247<=G32130 and G19980;
	G33248<=G32131 and G19996;
	G33249<=G32144 and G20026;
	G33252<=G32155 and G20064;
	G33263<=G32393 and G25481;
	G33264<=G31965 and G21306;
	G33269<=G31970 and G15582;
	G33304<=G32427 and G31971;
	G33305<=G31935 and G17811;
	G33311<=G31942 and G12925;
	G33322<=G32202 and G20450;
	G33327<=G32208 and G20561;
	G33328<=G32209 and G20584;
	G33329<=G32210 and G20585;
	G33330<=G32211 and G20588;
	G33331<=G32216 and G20607;
	G33332<=G32217 and G20608;
	G33333<=G32218 and G20612;
	G33334<=G32219 and G20613;
	G33338<=G32220 and G20633;
	G33339<=G32221 and G20634;
	G33340<=G32222 and G20639;
	G33341<=G32223 and G20640;
	G33342<=G32226 and G20660;
	G33343<=G32227 and G20665;
	G33344<=G32228 and G20670;
	G33345<=G32229 and G20671;
	G33349<=G32233 and G20699;
	G33350<=G32235 and G20702;
	G33351<=G32236 and G20707;
	G33352<=G32237 and G20712;
	G33353<=G32240 and G20732;
	G33355<=G32243 and G20769;
	G33356<=G32245 and G20772;
	G33357<=G32247 and G20775;
	G33358<=G32249 and G20778;
	G33359<=G32252 and G20853;
	G33360<=G32253 and G20869;
	G33361<=G32257 and G20911;
	G33362<=G32259 and G20914;
	G33363<=G32262 and G20918;
	G33364<=G32264 and G20921;
	G33365<=G32267 and G20994;
	G33366<=G32268 and G21010;
	G33367<=G32271 and G21053;
	G33368<=G32275 and G21057;
	G33369<=G32277 and G21060;
	G33370<=G32279 and G21139;
	G33371<=G32280 and G21155;
	G33372<=G32285 and G21183;
	G33373<=G32288 and G21205;
	G33374<=G32289 and G21221;
	G33376<=G32294 and G21268;
	G33379<=G30984 and G32364;
	G33381<=G11842 and G32318;
	G33392<=G32344 and G21362;
	G33399<=G32346 and G21379;
	G33400<=G32347 and G21380;
	G33401<=G32349 and G21381;
	G33402<=G32351 and G21395;
	G33403<=G32352 and G21396;
	G33404<=G32353 and G21397;
	G33405<=G32354 and G21398;
	G33406<=G32355 and G21399;
	G33407<=G32357 and G21406;
	G33408<=G32358 and G21407;
	G33409<=G32359 and G21408;
	G33410<=G32360 and G21409;
	G33411<=G32361 and G21410;
	G33412<=G32362 and G21411;
	G33414<=G32367 and G21421;
	G33415<=G32368 and G21422;
	G33416<=G32370 and G21423;
	G33417<=G32371 and G21424;
	G33418<=G32372 and G21425;
	G33420<=G32373 and G21454;
	G33421<=G32374 and G21455;
	G33422<=G32375 and G21456;
	G33423<=G32225 and G29657;
	G33425<=G32380 and G21466;
	G33428<=G32230 and G29672;
	G33429<=G32231 and G29676;
	G33431<=G32364 and G32377;
	G33433<=G32238 and G29694;
	G33434<=G32239 and G29702;
	G33440<=G32250 and G29719;
	G33441<=G32251 and G29722;
	G33446<=G32385 and G21607;
	G33450<=G32266 and G29737;
	G33461<=G32463 and I31001 and I31002;
	G33462<=G32470 and I31006 and I31007;
	G33463<=G32477 and I31011 and I31012;
	G33464<=G32484 and I31016 and I31017;
	G33465<=G32491 and I31021 and I31022;
	G33466<=G32498 and I31026 and I31027;
	G33467<=G32505 and I31031 and I31032;
	G33468<=G32512 and I31036 and I31037;
	G33469<=G32519 and I31041 and I31042;
	G33470<=G32528 and I31046 and I31047;
	G33471<=G32535 and I31051 and I31052;
	G33472<=G32542 and I31056 and I31057;
	G33473<=G32549 and I31061 and I31062;
	G33474<=G32556 and I31066 and I31067;
	G33475<=G32563 and I31071 and I31072;
	G33476<=G32570 and I31076 and I31077;
	G33477<=G32577 and I31081 and I31082;
	G33478<=G32584 and I31086 and I31087;
	G33479<=G32593 and I31091 and I31092;
	G33480<=G32600 and I31096 and I31097;
	G33481<=G32607 and I31101 and I31102;
	G33482<=G32614 and I31106 and I31107;
	G33483<=G32621 and I31111 and I31112;
	G33484<=G32628 and I31116 and I31117;
	G33485<=G32635 and I31121 and I31122;
	G33486<=G32642 and I31126 and I31127;
	G33487<=G32649 and I31131 and I31132;
	G33488<=G32658 and I31136 and I31137;
	G33489<=G32665 and I31141 and I31142;
	G33490<=G32672 and I31146 and I31147;
	G33491<=G32679 and I31151 and I31152;
	G33492<=G32686 and I31156 and I31157;
	G33493<=G32693 and I31161 and I31162;
	G33494<=G32700 and I31166 and I31167;
	G33495<=G32707 and I31171 and I31172;
	G33496<=G32714 and I31176 and I31177;
	G33497<=G32723 and I31181 and I31182;
	G33498<=G32730 and I31186 and I31187;
	G33499<=G32737 and I31191 and I31192;
	G33500<=G32744 and I31196 and I31197;
	G33501<=G32751 and I31201 and I31202;
	G33502<=G32758 and I31206 and I31207;
	G33503<=G32765 and I31211 and I31212;
	G33504<=G32772 and I31216 and I31217;
	G33505<=G32779 and I31221 and I31222;
	G33506<=G32788 and I31226 and I31227;
	G33507<=G32795 and I31231 and I31232;
	G33508<=G32802 and I31236 and I31237;
	G33509<=G32809 and I31241 and I31242;
	G33510<=G32816 and I31246 and I31247;
	G33511<=G32823 and I31251 and I31252;
	G33512<=G32830 and I31256 and I31257;
	G33513<=G32837 and I31261 and I31262;
	G33514<=G32844 and I31266 and I31267;
	G33515<=G32853 and I31271 and I31272;
	G33516<=G32860 and I31276 and I31277;
	G33517<=G32867 and I31281 and I31282;
	G33518<=G32874 and I31286 and I31287;
	G33519<=G32881 and I31291 and I31292;
	G33520<=G32888 and I31296 and I31297;
	G33521<=G32895 and I31301 and I31302;
	G33522<=G32902 and I31306 and I31307;
	G33523<=G32909 and I31311 and I31312;
	G33524<=G32918 and I31316 and I31317;
	G33525<=G32925 and I31321 and I31322;
	G33526<=G32932 and I31326 and I31327;
	G33527<=G32939 and I31331 and I31332;
	G33528<=G32946 and I31336 and I31337;
	G33529<=G32953 and I31341 and I31342;
	G33530<=G32960 and I31346 and I31347;
	G33531<=G32967 and I31351 and I31352;
	G33532<=G32974 and I31356 and I31357;
	G33639<=G33386 and G18829;
	G33640<=G33387 and G18831;
	G33646<=G33389 and G18876;
	G33647<=G33390 and G18878;
	G33652<=G33393 and G18889;
	G33657<=G30991 and G33443;
	G33674<=G33164 and G10710 and G22319;
	G33675<=G33164 and G10727 and G22332;
	G33676<=G33125 and G7970;
	G33677<=G33443 and G31937;
	G33678<=G33149 and G10710 and G22319;
	G33680<=G33128 and G4688;
	G33681<=G33129 and G7991;
	G33683<=G33149 and G10727 and G22332;
	G33684<=G33139 and G13565;
	G33687<=G33132 and G4878;
	G33689<=G33144 and G11006;
	G33690<=G33146 and G16280;
	G33693<=G33145 and G13594;
	G33697<=G33160 and G13330;
	G33700<=G33148 and G11012;
	G33701<=G33162 and G16305;
	G33704<=G33176 and G10710 and G22319;
	G33707<=G33174 and G13346;
	G33710<=G14037 and G33246;
	G33711<=G33176 and G10727 and G22332;
	G33715<=G33135 and G19416;
	G33717<=G14092 and G33306;
	G33718<=G33147 and G19432;
	G33719<=G33141 and G19433;
	G33720<=G33161 and G19439;
	G33721<=G33163 and G19440;
	G33722<=G33175 and G19445;
	G33723<=G14091 and G33299;
	G33724<=G14145 and G33258;
	G33725<=G22626 and G10851 and G33176;
	G33727<=G33115 and G19499;
	G33728<=G22626 and G10851 and G33187;
	G33730<=G7202 and G4621 and G33127 and G4633;
	G33731<=G33116 and G19520;
	G33734<=G7806 and G33136 and I31593;
	G33735<=G33118 and G19553;
	G33742<=G7828 and G33142 and I31600;
	G33743<=G33119 and G19574;
	G33758<=G33133 and G20269;
	G33759<=G33123 and G22847;
	G33760<=G33143 and G20328;
	G33784<=G33107 and G20531;
	G33785<=G33100 and G20550;
	G33786<=G33130 and G20572;
	G33787<=G33103 and G20595;
	G33789<=G33159 and G23022;
	G33790<=G33108 and G20643;
	G33795<=G33138 and G20782;
	G33796<=G33117 and G25267;
	G33798<=G33227 and G20058;
	G33801<=G33437 and G25327;
	G33802<=G33097 and G14545;
	G33803<=G33231 and G20071;
	G33805<=G33232 and G20079;
	G33807<=G33112 and G25452;
	G33808<=G33109 and G22161;
	G33809<=G33432 and G30184;
	G33810<=G33427 and G12768;
	G33811<=G33439 and G17573;
	G33812<=G23088 and G33187 and G9104;
	G33814<=G33098 and G28144;
	G33815<=G33449 and G12911;
	G33816<=G33234 and G20096;
	G33817<=G33235 and G20102;
	G33818<=G33236 and G20113;
	G33819<=G23088 and G33176 and G9104;
	G33820<=G33075 and G26830;
	G33821<=G33238 and G20153;
	G33822<=G33385 and G20157;
	G33828<=G33090 and G24411;
	G33829<=G33240 and G20164;
	G33830<=G33382 and G20166;
	G33831<=G23088 and G33149 and G9104;
	G33832<=G33088 and G27991;
	G33833<=G33093 and G25852;
	G33834<=G33095 and G29172;
	G33835<=G4340 and G33413;
	G33836<=G33096 and G27020;
	G33837<=G33251 and G20233;
	G33840<=G33253 and G20267;
	G33841<=G33254 and G20268;
	G33842<=G33255 and G20322;
	G33843<=G33256 and G20325;
	G33844<=G33257 and G20327;
	G33846<=G33259 and G20380;
	G33847<=G33260 and G20383;
	G33848<=G33261 and G20384;
	G33849<=G33262 and G20387;
	G33855<=G33265 and G20441;
	G33856<=G33266 and G20442;
	G33857<=G33267 and G20445;
	G33858<=G33268 and G20448;
	G33859<=G33426 and G10531;
	G33860<=G33270 and G20501;
	G33861<=G33271 and G20502;
	G33862<=G33272 and G20504;
	G33863<=G33273 and G20505;
	G33864<=G33274 and G20524;
	G33865<=G33275 and G20526;
	G33866<=G33276 and G20528;
	G33867<=G33277 and G20529;
	G33868<=G33278 and G20542;
	G33869<=G33279 and G20543;
	G33870<=G33280 and G20545;
	G33871<=G33281 and G20546;
	G33872<=G33282 and G20548;
	G33873<=G33291 and G20549;
	G33876<=G33286 and G20562;
	G33877<=G33287 and G20563;
	G33878<=G33288 and G20565;
	G33879<=G33289 and G20566;
	G33880<=G33290 and G20568;
	G33881<=G33292 and G20586;
	G33882<=G33293 and G20587;
	G33883<=G33294 and G20589;
	G33884<=G33295 and G20590;
	G33885<=G33296 and G20609;
	G33886<=G33297 and G20614;
	G33887<=G33298 and G20615;
	G33889<=G33303 and G20641;
	G33890<=G33310 and G20659;
	G33892<=G33312 and G20701;
	G33893<=G33313 and G20706;
	G33896<=G33314 and G20771;
	G33897<=G33315 and G20777;
	G33898<=G33419 and G15655;
	G33899<=G32132 and G33335;
	G33900<=G33316 and G20913;
	G33901<=G33317 and G20920;
	G33902<=G33085 and G13202;
	G33903<=G33447 and G19146;
	G33904<=G33321 and G21059;
	G33905<=G33089 and G15574;
	G33906<=G33084 and G22311;
	G33907<=G23088 and G33219 and G9104;
	G33908<=G33092 and G18935;
	G33909<=G33131 and G10708;
	G33910<=G33134 and G7836;
	G33911<=G33137 and G10725;
	G33913<=G23088 and G33204 and G9104;
	G33915<=G33140 and G7846;
	G33919<=G33438 and G10795;
	G33921<=G33187 and G9104 and G19200;
	G33922<=G33448 and G7202;
	G33924<=G33335 and G33346;
	G33927<=G33094 and G21412;
	G33941<=G33380 and G21560;
	G33942<=G33383 and G21608;
	G33943<=G33384 and G21609;
	G34045<=G33766 and G22942;
	G34050<=G33772 and G22942;
	G34054<=G33778 and G22942;
	G34061<=G33800 and G23076;
	G34063<=G33806 and G23121;
	G34065<=G33813 and G23148;
	G34066<=G33730 and G19352;
	G34069<=G8774 and G33797;
	G34071<=G8854 and G33799;
	G34072<=G33839 and G24872;
	G34073<=G8948 and G33823;
	G34074<=G33685 and G19498;
	G34075<=G33692 and G19517;
	G34076<=G33694 and G19519;
	G34077<=G22957 and G9104 and G33736;
	G34078<=G33699 and G19531;
	G34079<=G33703 and G19532;
	G34080<=G22957 and G9104 and G33750;
	G34081<=G33706 and G19552;
	G34082<=G33709 and G19554;
	G34083<=G33714 and G19573;
	G34084<=G9214 and G33851;
	G34085<=G33761 and G9104 and G18957;
	G34086<=G20114 and G33766 and G9104;
	G34087<=G33766 and G9104 and G18957;
	G34088<=G33736 and G9104 and G18957;
	G34089<=G22957 and G9104 and G33744;
	G34091<=G22957 and G9104 and G33761;
	G34092<=G33750 and G9104 and G18957;
	G34093<=G20114 and G33755 and G9104;
	G34096<=G22957 and G9104 and G33772;
	G34097<=G33772 and G9104 and G18957;
	G34098<=G33744 and G9104 and G18957;
	G34102<=G33912 and G23599;
	G34104<=G33916 and G23639;
	G34105<=G33778 and G9104 and G18957;
	G34106<=G33917 and G23675;
	G34108<=G22957 and G9104 and G33766;
	G34109<=G33918 and G23708;
	G34110<=G33732 and G22935;
	G34111<=G33733 and G22936;
	G34112<=G22957 and G9104 and G33778;
	G34113<=G33734 and G19744;
	G34114<=G33920 and G23742;
	G34115<=G20516 and G9104 and G33750;
	G34116<=G33933 and G25140;
	G34117<=G33742 and G19755;
	G34119<=G20516 and G9104 and G33755;
	G34120<=G33930 and G25158;
	G34133<=G33845 and G23958;
	G34135<=G33926 and G23802;
	G34136<=G33850 and G23293;
	G34137<=G33928 and G23802;
	G34138<=G33929 and G23828;
	G34139<=G33827 and G23314;
	G34140<=G33931 and G23802;
	G34141<=G33932 and G23828;
	G34143<=G33934 and G23828;
	G34146<=G33788 and G20091;
	G34157<=G33794 and G20159;
	G34169<=G33804 and G31227;
	G34171<=G33925 and G24360;
	G34173<=G33679 and G24368;
	G34178<=G33712 and G24361;
	G34179<=G33686 and G24372;
	G34180<=G33716 and G24373;
	G34182<=G33691 and G24384;
	G34183<=G33695 and G24385;
	G34184<=G33698 and G24388;
	G34185<=G33702 and G24389;
	G34186<=G33705 and G24396;
	G34187<=G33708 and G24397;
	G34191<=G33713 and G24404;
	G34196<=G33682 and G24485;
	G34198<=G33688 and G24491;
	G34203<=G33726 and G24537;
	G34205<=G33729 and G24541;
	G34211<=G33891 and G21349;
	G34212<=G33761 and G22689;
	G34213<=G33766 and G22689;
	G34214<=G33772 and G22689;
	G34215<=G33778 and G22670;
	G34216<=G33778 and G22689;
	G34217<=G33736 and G22876;
	G34218<=G33744 and G22670;
	G34219<=G33736 and G22942;
	G34223<=G33744 and G22876;
	G34224<=G33736 and G22670;
	G34225<=G33744 and G22942;
	G34226<=G33914 and G21467;
	G34228<=G33750 and G22942;
	G34230<=G33761 and G22942;
	G34279<=G34231 and G19208;
	G34281<=G34043 and G19276;
	G34284<=G34046 and G19351;
	G34287<=G11370 and G34124;
	G34291<=G34055 and G19366;
	G34295<=G34057 and G19370;
	G34298<=G8679 and G34132;
	G34301<=G34064 and G19415;
	G34309<=G13947 and G34147;
	G34310<=G14003 and G34162;
	G34319<=G9535 and G34156;
	G34322<=G14188 and G34174;
	G34324<=G14064 and G34161;
	G34329<=G14511 and G34181;
	G34333<=G9984 and G34192;
	G34334<=G34090 and G19865;
	G34335<=G8461 and G34197;
	G34337<=G34095 and G19881;
	G34338<=G34099 and G19905;
	G34340<=G34100 and G19950;
	G34341<=G34101 and G19952;
	G34342<=G34103 and G19998;
	G34344<=G34107 and G20038;
	G34348<=G34125 and G20128;
	G34363<=G34148 and G20389;
	G34364<=G34048 and G24366;
	G34365<=G34149 and G20451;
	G34367<=G7404 and G34042;
	G34370<=G34067 and G10554;
	G34371<=G7450 and G34044;
	G34375<=G13077 and G34049;
	G34378<=G13095 and G34053;
	G34380<=G34158 and G20571;
	G34381<=G34166 and G20594;
	G34382<=G34167 and G20618;
	G34385<=G34168 and G20642;
	G34386<=G10800 and G34060;
	G34388<=G10802 and G34062;
	G34389<=G34170 and G20715;
	G34390<=G34172 and G21069;
	G34393<=G34189 and G21304;
	G34394<=G34190 and G21305;
	G34395<=G34193 and G21336;
	G34396<=G34194 and G21337;
	G34397<=G7673 and G34068;
	G34398<=G7684 and G34070;
	G34401<=G34199 and G21383;
	G34410<=G34204 and G21427;
	G34413<=G34094 and G22670;
	G34414<=G34206 and G21457;
	G34415<=G34207 and G21458;
	G34470<=G7834 and G34325;
	G34474<=G20083 and G34326;
	G34475<=G27450 and G34327;
	G34476<=G34399 and G18891;
	G34477<=G26344 and G34328;
	G34478<=G34402 and G18904;
	G34479<=G34403 and G18905;
	G34481<=G34404 and G18916;
	G34482<=G34405 and G18917;
	G34483<=G34406 and G18938;
	G34484<=G34407 and G18939;
	G34485<=G34411 and G18952;
	G34486<=G34412 and G18953;
	G34487<=G34416 and G18983;
	G34488<=G34417 and G18988;
	G34489<=G34421 and G19068;
	G34492<=G34272 and G33430;
	G34493<=G34273 and G19360;
	G34495<=G34274 and G19365;
	G34497<=G34275 and G33072;
	G34498<=G13888 and G34336;
	G34499<=G31288 and G34339;
	G34500<=G34276 and G30568;
	G34502<=G26363 and G34343;
	G34503<=G34278 and G19437;
	G34506<=G8833 and G34354;
	G34507<=G34280 and G19454;
	G34508<=G34282 and G19472;
	G34509<=G34283 and G19473;
	G34513<=G9003 and G34346;
	G34514<=G34286 and G19480;
	G34515<=G34288 and G19491;
	G34516<=G34289 and G19492;
	G34517<=G34290 and G19493;
	G34518<=G34292 and G19503;
	G34519<=G34293 and G19504;
	G34520<=G34294 and G19505;
	G34523<=G9162 and G34351;
	G34524<=G9083 and G34359;
	G34525<=G34297 and G19528;
	G34526<=G34300 and G19569;
	G34527<=G34303 and G19603;
	G34528<=G34305 and G19617;
	G34529<=G34306 and G19634;
	G34532<=G34314 and G19710;
	G34533<=G34318 and G19731;
	G34534<=G34321 and G19743;
	G34538<=G34330 and G20054;
	G34541<=G34331 and G20087;
	G34542<=G34332 and G20089;
	G34554<=G34347 and G20495;
	G34555<=G34349 and G20512;
	G34556<=G34350 and G20537;
	G34557<=G34352 and G20555;
	G34558<=G34353 and G20578;
	G34560<=G34366 and G17366;
	G34561<=G34368 and G17410;
	G34562<=G34369 and G17411;
	G34563<=G34372 and G17465;
	G34564<=G34373 and G17466;
	G34565<=G34374 and G17471;
	G34566<=G34376 and G17489;
	G34567<=G34377 and G17491;
	G34568<=G34379 and G17512;
	G34571<=G27225 and G34299;
	G34572<=G34387 and G33326;
	G34577<=G24577 and G34307;
	G34578<=G24578 and G34308;
	G34580<=G29539 and G34311;
	G34581<=G22864 and G34312;
	G34582<=G7764 and G34313;
	G34584<=G24653 and G34315;
	G34585<=G24705 and G34316;
	G34586<=G11025 and G34317;
	G34588<=G26082 and G34323;
	G34655<=G34573 and G18885;
	G34658<=G34574 and G18896;
	G34661<=G34575 and G18907;
	G34662<=G34576 and G18931;
	G34665<=G34583 and G19067;
	G34666<=G34587 and G19144;
	G34667<=G34471 and G33424;
	G34678<=G34490 and G19431;
	G34679<=G14093 and G34539;
	G34681<=G34491 and G19438;
	G34684<=G14178 and G34545;
	G34685<=G14164 and G34550;
	G34686<=G34494 and G19494;
	G34687<=G14181 and G34543;
	G34694<=G34530 and G19885;
	G34696<=G34531 and G20004;
	G34700<=G34535 and G20129;
	G34701<=G34536 and G20179;
	G34702<=G34537 and G20208;
	G34706<=G34496 and G10570;
	G34707<=G34544 and G20579;
	G34709<=G34549 and G17242;
	G34710<=G34553 and G20903;
	G34715<=G34570 and G33375;
	G34738<=G34660 and G33442;
	G34740<=G34664 and G19414;
	G34741<=G8899 and G34697;
	G34742<=G9000 and G34698;
	G34743<=G8951 and G34703;
	G34744<=G34668 and G19481;
	G34745<=G34669 and G19482;
	G34746<=G34670 and G19526;
	G34747<=G34671 and G19527;
	G34748<=G34672 and G19529;
	G34750<=G34673 and G19542;
	G34751<=G34674 and G19543;
	G34752<=G34675 and G19544;
	G34753<=G34676 and G19586;
	G34754<=G34677 and G19602;
	G34756<=G34680 and G19618;
	G34757<=G34682 and G19635;
	G34758<=G34683 and G19657;
	G34763<=G34689 and G19915;
	G34764<=G34691 and G20009;
	G34765<=G34692 and G20057;
	G34771<=G34693 and G20147;
	G34774<=G34695 and G20180;
	G34782<=G34711 and G33888;
	G34811<=G14165 and G34766;
	G34841<=G34761 and G20080;
	G34842<=G34762 and G20168;
	G34857<=G16540 and G34813;
	G34858<=G16540 and G34816;
	G34859<=G16540 and G34820;
	G34860<=G16540 and G34823;
	G34861<=G16540 and G34827;
	G34862<=G16540 and G34830;
	G34863<=G16540 and G34833;
	G34865<=G16540 and G34836;
	G34866<=G34819 and G20106;
	G34867<=G34826 and G20145;
	G34868<=G34813 and G19866;
	G34869<=G34816 and G19869;
	G34870<=G34820 and G19882;
	G34871<=G34823 and G19908;
	G34872<=G34827 and G19954;
	G34873<=G34830 and G20046;
	G34874<=G34833 and G20060;
	G34875<=G34836 and G20073;
	G34876<=G34844 and G20534;
	G34909<=G34856 and G20130;
	G34948<=G16540 and G34935;
	G34953<=G34935 and G19957;
	G34955<=G34931 and G34320;
	G34961<=G34944 and G23019;
	G34962<=G34945 and G23020;
	G34963<=G34946 and G23041;
	G34964<=G34947 and G23060;
	G34965<=G34949 and G23084;
	G34966<=G34950 and G23170;
	G34967<=G34951 and G23189;
	G34968<=G34952 and G23203;
	G34969<=G34960 and G19570;
	G34999<=G34998 and G23085;
	I13862<=G7232 and G7219 and G7258;
	I13937<=G7340 and G7293 and G7261;
	I14198<=G225 and G8237 and G232 and G8180;
	I14225<=G8457 and G255 and G8406 and G262;
	I16111<=G8691 and G11409 and G11381;
	I16129<=G8728 and G11443 and G11411;
	I16143<=G8751 and G11491 and G11445;
	I16618<=G10124 and G12341 and G12293;
	I16646<=G10160 and G12413 and G12343;
	I16671<=G10185 and G12461 and G12415;
	I16695<=G10207 and G12523 and G12463;
	I16721<=G10224 and G12589 and G12525;
	I17529<=G13156 and G11450 and G6756;
	I17542<=G13156 and G6767 and G6756;
	I17552<=G13156 and G11450 and G11498;
	I17575<=G13156 and G11450 and G6756;
	I17585<=G14988 and G11450 and G11498;
	I17606<=G14988 and G11450 and G6756;
	I17692<=G14988 and G11450 and G6756;
	I17741<=G14988 and G11450 and G11498;
	I18568<=G13156 and G11450 and G11498;
	I18620<=G13156 and G11450 and G11498;
	I18671<=G13156 and G11450 and G6756;
	I18713<=G13156 and G6767 and G6756;
	I18716<=G13156 and G11450 and G6756;
	I18740<=G13156 and G11450 and G11498;
	I18762<=G13156 and G6767 and G11498;
	I18765<=G13156 and G11450 and G11498;
	I18782<=G13156 and G11450 and G6756;
	I18785<=G13156 and G6767 and G11498;
	I18803<=G13156 and G11450 and G6756;
	I18819<=G13156 and G11450 and G11498;
	I24003<=G8097 and G8334 and G3045;
	I24015<=G8334 and G7975 and G3045;
	I24018<=G8155 and G8390 and G3396;
	I24027<=G3029 and G3034 and G8426;
	I24030<=G8390 and G8016 and G3396;
	I24033<=G8219 and G8443 and G3747;
	I24048<=G3034 and G3040 and G8426;
	I24051<=G3380 and G3385 and G8492;
	I24054<=G8443 and G8075 and G3747;
	I24064<=G3385 and G3391 and G8492;
	I24067<=G3731 and G3736 and G8553;
	I24075<=G3736 and G3742 and G8553;
	I24482<=G9364 and G9607 and G5057;
	I24505<=G9607 and G9229 and G5057;
	I24508<=G9434 and G9672 and G5401;
	I24524<=G5041 and G5046 and G9716;
	I24527<=G9672 and G9264 and G5401;
	I24530<=G9501 and G9733 and G5747;
	I24546<=G5046 and G5052 and G9716;
	I24549<=G5385 and G5390 and G9792;
	I24552<=G9733 and G9316 and G5747;
	I24555<=G9559 and G9809 and G6093;
	I24576<=G5390 and G5396 and G9792;
	I24579<=G5731 and G5736 and G9875;
	I24582<=G9809 and G9397 and G6093;
	I24585<=G9621 and G9892 and G6439;
	I24597<=G5736 and G5742 and G9875;
	I24600<=G6077 and G6082 and G9946;
	I24603<=G9892 and G9467 and G6439;
	I24616<=G6082 and G6088 and G9946;
	I24619<=G6423 and G6428 and G10014;
	I24625<=G6428 and G6434 and G10014;
	I24674<=G19919 and G24019 and G24020 and G24021;
	I24675<=G24022 and G24023 and G24024 and G24025;
	I24679<=G19968 and G24026 and G24027 and G24028;
	I24680<=G24029 and G24030 and G24031 and G24032;
	I24684<=G20014 and G24033 and G24034 and G24035;
	I24685<=G24036 and G24037 and G24038 and G24039;
	I24689<=G20841 and G24040 and G24041 and G24042;
	I24690<=G24043 and G24044 and G24045 and G24046;
	I24694<=G20982 and G24047 and G24048 and G24049;
	I24695<=G24050 and G24051 and G24052 and G24053;
	I24699<=G21127 and G24054 and G24055 and G24056;
	I24700<=G24057 and G24058 and G24059 and G24060;
	I24704<=G21193 and G24061 and G24062 and G24063;
	I24705<=G24064 and G24065 and G24066 and G24067;
	I24709<=G21256 and G24068 and G24069 and G24070;
	I24710<=G24071 and G24072 and G24073 and G24074;
	I26530<=G26365 and G24096 and G24097 and G24098;
	I26531<=G24099 and G24100 and G24101 and G24102;
	I26948<=G24981 and G26424 and G22698;
	I26960<=G24995 and G26424 and G22698;
	I26972<=G25011 and G26424 and G22698;
	I27349<=G25534 and G26424 and G22698;
	I27364<=G25541 and G26424 and G22698;
	I27381<=G25549 and G26424 and G22698;
	I27409<=G25556 and G26424 and G22698;
	I27429<=G25562 and G26424 and G22698;
	I27503<=G19890 and G24075 and G24076 and G28032;
	I27504<=G24077 and G24078 and G24079 and G24080;
	I27508<=G19935 and G24082 and G24083 and G28033;
	I27509<=G24084 and G24085 and G24086 and G24087;
	I27513<=G19984 and G24089 and G24090 and G28034;
	I27514<=G24091 and G24092 and G24093 and G24094;
	I27518<=G20720 and G24104 and G24105 and G24106;
	I27519<=G28036 and G24107 and G24108 and G24109;
	I27523<=G20857 and G24111 and G24112 and G24113;
	I27524<=G28037 and G24114 and G24115 and G24116;
	I27528<=G20998 and G24118 and G24119 and G24120;
	I27529<=G28038 and G24121 and G24122 and G24123;
	I27533<=G21143 and G24125 and G24126 and G24127;
	I27534<=G28039 and G24128 and G24129 and G24130;
	I27538<=G21209 and G24132 and G24133 and G24134;
	I27539<=G28040 and G24135 and G24136 and G24137;
	I31001<=G29385 and G32456 and G32457 and G32458;
	I31002<=G32459 and G32460 and G32461 and G32462;
	I31006<=G31376 and G31796 and G32464 and G32465;
	I31007<=G32466 and G32467 and G32468 and G32469;
	I31011<=G30735 and G31797 and G32471 and G32472;
	I31012<=G32473 and G32474 and G32475 and G32476;
	I31016<=G30825 and G31798 and G32478 and G32479;
	I31017<=G32480 and G32481 and G32482 and G32483;
	I31021<=G31070 and G31799 and G32485 and G32486;
	I31022<=G32487 and G32488 and G32489 and G32490;
	I31026<=G31194 and G31800 and G32492 and G32493;
	I31027<=G32494 and G32495 and G32496 and G32497;
	I31031<=G30614 and G31801 and G32499 and G32500;
	I31032<=G32501 and G32502 and G32503 and G32504;
	I31036<=G30673 and G31802 and G32506 and G32507;
	I31037<=G32508 and G32509 and G32510 and G32511;
	I31041<=G31566 and G31803 and G32513 and G32514;
	I31042<=G32515 and G32516 and G32517 and G32518;
	I31046<=G29385 and G32521 and G32522 and G32523;
	I31047<=G32524 and G32525 and G32526 and G32527;
	I31051<=G31376 and G31804 and G32529 and G32530;
	I31052<=G32531 and G32532 and G32533 and G32534;
	I31056<=G30735 and G31805 and G32536 and G32537;
	I31057<=G32538 and G32539 and G32540 and G32541;
	I31061<=G30825 and G31806 and G32543 and G32544;
	I31062<=G32545 and G32546 and G32547 and G32548;
	I31066<=G31070 and G31807 and G32550 and G32551;
	I31067<=G32552 and G32553 and G32554 and G32555;
	I31071<=G31170 and G31808 and G32557 and G32558;
	I31072<=G32559 and G32560 and G32561 and G32562;
	I31076<=G30614 and G31809 and G32564 and G32565;
	I31077<=G32566 and G32567 and G32568 and G32569;
	I31081<=G30673 and G31810 and G32571 and G32572;
	I31082<=G32573 and G32574 and G32575 and G32576;
	I31086<=G31554 and G31811 and G32578 and G32579;
	I31087<=G32580 and G32581 and G32582 and G32583;
	I31091<=G29385 and G32586 and G32587 and G32588;
	I31092<=G32589 and G32590 and G32591 and G32592;
	I31096<=G31376 and G31812 and G32594 and G32595;
	I31097<=G32596 and G32597 and G32598 and G32599;
	I31101<=G30735 and G31813 and G32601 and G32602;
	I31102<=G32603 and G32604 and G32605 and G32606;
	I31106<=G30825 and G31814 and G32608 and G32609;
	I31107<=G32610 and G32611 and G32612 and G32613;
	I31111<=G31070 and G31815 and G32615 and G32616;
	I31112<=G32617 and G32618 and G32619 and G32620;
	I31116<=G31154 and G31816 and G32622 and G32623;
	I31117<=G32624 and G32625 and G32626 and G32627;
	I31121<=G30614 and G31817 and G32629 and G32630;
	I31122<=G32631 and G32632 and G32633 and G32634;
	I31126<=G30673 and G31818 and G32636 and G32637;
	I31127<=G32638 and G32639 and G32640 and G32641;
	I31131<=G31542 and G31819 and G32643 and G32644;
	I31132<=G32645 and G32646 and G32647 and G32648;
	I31136<=G29385 and G32651 and G32652 and G32653;
	I31137<=G32654 and G32655 and G32656 and G32657;
	I31141<=G31376 and G31820 and G32659 and G32660;
	I31142<=G32661 and G32662 and G32663 and G32664;
	I31146<=G30735 and G31821 and G32666 and G32667;
	I31147<=G32668 and G32669 and G32670 and G32671;
	I31151<=G30825 and G31822 and G32673 and G32674;
	I31152<=G32675 and G32676 and G32677 and G32678;
	I31156<=G31070 and G31823 and G32680 and G32681;
	I31157<=G32682 and G32683 and G32684 and G32685;
	I31161<=G30614 and G31824 and G32687 and G32688;
	I31162<=G32689 and G32690 and G32691 and G32692;
	I31166<=G30673 and G31825 and G32694 and G32695;
	I31167<=G32696 and G32697 and G32698 and G32699;
	I31171<=G31528 and G31826 and G32701 and G32702;
	I31172<=G32703 and G32704 and G32705 and G32706;
	I31176<=G31579 and G31827 and G32708 and G32709;
	I31177<=G32710 and G32711 and G32712 and G32713;
	I31181<=G29385 and G32716 and G32717 and G32718;
	I31182<=G32719 and G32720 and G32721 and G32722;
	I31186<=G31376 and G31828 and G32724 and G32725;
	I31187<=G32726 and G32727 and G32728 and G32729;
	I31191<=G30735 and G31829 and G32731 and G32732;
	I31192<=G32733 and G32734 and G32735 and G32736;
	I31196<=G30825 and G31830 and G32738 and G32739;
	I31197<=G32740 and G32741 and G32742 and G32743;
	I31201<=G31672 and G31831 and G32745 and G32746;
	I31202<=G32747 and G32748 and G32749 and G32750;
	I31206<=G31710 and G31832 and G32752 and G32753;
	I31207<=G32754 and G32755 and G32756 and G32757;
	I31211<=G31021 and G31833 and G32759 and G32760;
	I31212<=G32761 and G32762 and G32763 and G32764;
	I31216<=G30937 and G31834 and G32766 and G32767;
	I31217<=G32768 and G32769 and G32770 and G32771;
	I31221<=G31327 and G31835 and G32773 and G32774;
	I31222<=G32775 and G32776 and G32777 and G32778;
	I31226<=G29385 and G32781 and G32782 and G32783;
	I31227<=G32784 and G32785 and G32786 and G32787;
	I31231<=G31376 and G31836 and G32789 and G32790;
	I31232<=G32791 and G32792 and G32793 and G32794;
	I31236<=G30735 and G31837 and G32796 and G32797;
	I31237<=G32798 and G32799 and G32800 and G32801;
	I31241<=G30825 and G31838 and G32803 and G32804;
	I31242<=G32805 and G32806 and G32807 and G32808;
	I31246<=G31672 and G31839 and G32810 and G32811;
	I31247<=G32812 and G32813 and G32814 and G32815;
	I31251<=G31710 and G31840 and G32817 and G32818;
	I31252<=G32819 and G32820 and G32821 and G32822;
	I31256<=G31021 and G31841 and G32824 and G32825;
	I31257<=G32826 and G32827 and G32828 and G32829;
	I31261<=G30937 and G31842 and G32831 and G32832;
	I31262<=G32833 and G32834 and G32835 and G32836;
	I31266<=G31327 and G31843 and G32838 and G32839;
	I31267<=G32840 and G32841 and G32842 and G32843;
	I31271<=G29385 and G32846 and G32847 and G32848;
	I31272<=G32849 and G32850 and G32851 and G32852;
	I31276<=G31376 and G31844 and G32854 and G32855;
	I31277<=G32856 and G32857 and G32858 and G32859;
	I31281<=G30735 and G31845 and G32861 and G32862;
	I31282<=G32863 and G32864 and G32865 and G32866;
	I31286<=G30825 and G31846 and G32868 and G32869;
	I31287<=G32870 and G32871 and G32872 and G32873;
	I31291<=G31021 and G31847 and G32875 and G32876;
	I31292<=G32877 and G32878 and G32879 and G32880;
	I31296<=G30937 and G31848 and G32882 and G32883;
	I31297<=G32884 and G32885 and G32886 and G32887;
	I31301<=G31327 and G31849 and G32889 and G32890;
	I31302<=G32891 and G32892 and G32893 and G32894;
	I31306<=G30614 and G31850 and G32896 and G32897;
	I31307<=G32898 and G32899 and G32900 and G32901;
	I31311<=G30673 and G31851 and G32903 and G32904;
	I31312<=G32905 and G32906 and G32907 and G32908;
	I31316<=G29385 and G32911 and G32912 and G32913;
	I31317<=G32914 and G32915 and G32916 and G32917;
	I31321<=G31376 and G31852 and G32919 and G32920;
	I31322<=G32921 and G32922 and G32923 and G32924;
	I31326<=G30735 and G31853 and G32926 and G32927;
	I31327<=G32928 and G32929 and G32930 and G32931;
	I31331<=G30825 and G31854 and G32933 and G32934;
	I31332<=G32935 and G32936 and G32937 and G32938;
	I31336<=G31672 and G31855 and G32940 and G32941;
	I31337<=G32942 and G32943 and G32944 and G32945;
	I31341<=G31710 and G31856 and G32947 and G32948;
	I31342<=G32949 and G32950 and G32951 and G32952;
	I31346<=G31021 and G31857 and G32954 and G32955;
	I31347<=G32956 and G32957 and G32958 and G32959;
	I31351<=G30937 and G31858 and G32961 and G32962;
	I31352<=G32963 and G32964 and G32965 and G32966;
	I31356<=G31327 and G31859 and G32968 and G32969;
	I31357<=G32970 and G32971 and G32972 and G32973;
	I31593<=G31003 and G8350 and G7788;
	I31600<=G31009 and G8400 and G7809;
	G7133<= not (I11825 and I11826);
	G7150<= not (G5016 and G5062);
	G7167<= not (G5360 and G5406);
	G7184<= not (G5706 and G5752);
	G7201<= not (I11865 and I11866);
	G7209<= not (G6052 and G6098);
	G7223<= not (I11878 and I11879);
	G7227<= not (G4584 and G4593);
	G7228<= not (G6398 and G6444);
	G7442<= not (G896 and G890);
	G7549<= not (G1018 and G1030);
	G7582<= not (G1361 and G1373);
	G7598<= not (I12075 and I12076);
	G7611<= not (G4057 and G4064);
	G7620<= not (I12097 and I12098);
	G7690<= not (G4669 and G4659 and G4653);
	G7701<= not (G4859 and G4849 and G4843);
	G7803<= not (I12204 and I12205);
	G7823<= not (I12218 and I12219);
	G7836<= not (G4653 and G4688);
	G7846<= not (G4843 and G4878);
	G7850<= not (G554 and G807);
	G7857<= not (I12241 and I12242);
	G7869<= not (I12252 and I12253);
	G7879<= not (I12262 and I12263);
	G7885<= not (I12270 and I12271);
	G7887<= not (I12278 and I12279);
	G7897<= not (I12288 and I12289);
	G8010<= not (I12345 and I12346);
	G8069<= not (I12373 and I12374);
	G8105<= not (G3068 and G3072);
	G8124<= not (I12402 and I12403);
	G8163<= not (G3419 and G3423);
	G8227<= not (G3770 and G3774);
	G8238<= not (I12469 and I12470);
	G8292<= not (G218 and G215);
	G8347<= not (G4358 and G4349 and G4340);
	G8359<= not (I12545 and I12546);
	G8434<= not (G3080 and G3072);
	G8500<= not (G3431 and G3423);
	G8561<= not (G3782 and G3774);
	G8609<= not (G1171 and G1157);
	G8632<= not (G1514 and G1500);
	G8678<= not (G376 and G358);
	G8691<= not (G3267 and G3310 and G3281 and G3303);
	G8728<= not (G3618 and G3661 and G3632 and G3654);
	G8737<= not (I12729 and I12730);
	G8751<= not (G3969 and G4012 and G3983 and G4005);
	G8769<= not (G691 and G714);
	G8803<= not (G128 and G4646);
	G8806<= not (G358 and G370 and G376 and G385);
	G8829<= not (G5011 and G4836);
	G8847<= not (G4831 and G4681);
	G8871<= not (I12841 and I12842);
	G8873<= not (I12849 and I12850);
	G8889<= not (G3684 and G4871);
	G8913<= not (I12877 and I12878);
	G8967<= not (G4264 and G4258);
	G9092<= not (G3004 and G3050);
	G9177<= not (G3355 and G3401);
	G9203<= not (G3706 and G3752);
	G9246<= not (G847 and G812);
	G9258<= not (I13044 and I13045);
	G9295<= not (I13066 and I13067);
	G9310<= not (I13078 and I13079);
	G9334<= not (G827 and G832);
	G9372<= not (G5080 and G5084);
	G9391<= not (I13110 and I13111);
	G9442<= not (G5424 and G5428);
	G9461<= not (I13140 and I13141);
	G9485<= not (G1657 and G1624);
	G9509<= not (G5770 and G5774);
	G9528<= not (I13183 and I13184);
	G9538<= not (G1792 and G1760);
	G9543<= not (G2217 and G2185);
	G9567<= not (G6116 and G6120);
	G9591<= not (G1926 and G1894);
	G9595<= not (G2351 and G2319);
	G9629<= not (G6462 and G6466);
	G9645<= not (G2060 and G2028);
	G9654<= not (G2485 and G2453);
	G9663<= not (G128 and G4646);
	G9705<= not (G2619 and G2587);
	G9715<= not (G5011 and G4836);
	G9724<= not (G5092 and G5084);
	G9750<= not (I13335 and I13336);
	G9775<= not (G4831 and G4681);
	G9800<= not (G5436 and G5428);
	G9823<= not (I13383 and I13384);
	G9825<= not (I13391 and I13392);
	G9830<= not (I13402 and I13403);
	G9852<= not (G3684 and G4871);
	G9883<= not (G5782 and G5774);
	G9904<= not (I13443 and I13444);
	G9908<= not (I13453 and I13454);
	G9912<= not (I13463 and I13464);
	G9954<= not (G6128 and G6120);
	G9966<= not (I13498 and I13499);
	G9972<= not (I13510 and I13511);
	G9975<= not (I13519 and I13520);
	G10022<= not (G6474 and G6466);
	G10041<= not (I13565 and I13566);
	G10124<= not (G5276 and G5320 and G5290 and G5313);
	G10160<= not (G5623 and G5666 and G5637 and G5659);
	G10185<= not (G5969 and G6012 and G5983 and G6005);
	G10207<= not (G6315 and G6358 and G6329 and G6351);
	G10224<= not (G6661 and G6704 and G6675 and G6697);
	G10307<= not (I13730 and I13731);
	G10336<= not (I13750 and I13751);
	G10472<= not (I13851 and I13852);
	G10511<= not (G4628 and G7202 and G4621);
	G10515<= not (G10337 and G5022);
	G10520<= not (G7195 and G7115);
	G10529<= not (G1592 and G7308);
	G10537<= not (G7138 and G5366);
	G10550<= not (G7268 and G7308);
	G10551<= not (G1728 and G7356);
	G10552<= not (G2153 and G7374);
	G10556<= not (G7971 and G8133);
	G10561<= not (G7157 and G5712);
	G10566<= not (G7315 and G7356);
	G10567<= not (G1862 and G7405);
	G10568<= not (G7328 and G7374);
	G10569<= not (G2287 and G7418);
	G10573<= not (G7992 and G8179);
	G10578<= not (G7174 and G6058);
	G10583<= not (G7475 and G862);
	G10584<= not (G7362 and G7405);
	G10585<= not (G1996 and G7451);
	G10586<= not (G7380 and G7418);
	G10587<= not (G2421 and G7456);
	G10598<= not (G7191 and G6404);
	G10601<= not (G896 and G7397);
	G10602<= not (G7411 and G7451);
	G10603<= not (G10077 and G9751);
	G10604<= not (G7424 and G7456);
	G10605<= not (G2555 and G7490);
	G10609<= not (G10111 and G9826);
	G10610<= not (G7462 and G7490);
	G10611<= not (G10115 and G9831);
	G10614<= not (G9024 and G8977 and G8928);
	G10617<= not (G10151 and G9909);
	G10618<= not (G10153 and G9913);
	G10622<= not (G10178 and G9973);
	G10623<= not (G10181 and G9976);
	G10653<= not (G10204 and G10042);
	G10726<= not (G7304 and G7661 and G979 and G1061);
	G10737<= not (G6961 and G9848);
	G10738<= not (G6961 and G10308);
	G10754<= not (G7936 and G7913 and G8411);
	G10755<= not (G7352 and G7675 and G1322 and G1404);
	G10759<= not (G7537 and G324);
	G10775<= not (G7960 and G7943 and G8470);
	G10796<= not (G7537 and G7523);
	G10820<= not (G9985 and G9920 and G9843);
	G10905<= not (G1116 and G7304);
	G10909<= not (G7304 and G1116);
	G10916<= not (G1146 and G7854);
	G10928<= not (G8181 and G8137 and G417);
	G10929<= not (G1099 and G7854);
	G10935<= not (G1459 and G7352);
	G10939<= not (G7352 and G1459);
	G10946<= not (G1489 and G7876);
	G10951<= not (G7845 and G7868);
	G10961<= not (G1442 and G7876);
	G10971<= not (G7867 and G7886);
	G11002<= not (G7475 and G862);
	G11020<= not (G9187 and G9040);
	G11117<= not (G8087 and G8186 and G8239);
	G11118<= not (I14170 and I14171);
	G11130<= not (G1221 and G7918);
	G11134<= not (G8138 and G8240 and G8301);
	G11135<= not (I14186 and I14187);
	G11149<= not (G1564 and G7948);
	G11153<= not (I14205 and I14206);
	G11154<= not (I14212 and I14213);
	G11155<= not (G4776 and G7892 and G9030);
	G11169<= not (I14229 and I14230);
	G11172<= not (G8478 and G3096);
	G11173<= not (G4966 and G7898 and G9064);
	G11189<= not (I14248 and I14249);
	G11190<= not (G8539 and G3447);
	G11193<= not (I14258 and I14259);
	G11200<= not (G8592 and G3798);
	G11206<= not (I14276 and I14277);
	G11224<= not (I14290 and I14291);
	G11245<= not (G7636 and G7733 and G7697);
	G11251<= not (G8438 and G3092);
	G11279<= not (G8504 and G3443);
	G11292<= not (I14331 and I14332);
	G11302<= not (G9496 and G3281);
	G11312<= not (G8565 and G3794);
	G11320<= not (G4633 and G4621 and G7202);
	G11323<= not (I14351 and I14352);
	G11326<= not (G8993 and G376 and G365 and G370);
	G11330<= not (G9483 and G1193);
	G11350<= not (I14369 and I14370);
	G11355<= not (G9551 and G3310);
	G11356<= not (G9552 and G3632);
	G11374<= not (G9536 and G1536);
	G11381<= not (G9660 and G3274);
	G11382<= not (G8644 and G6895 and G8663);
	G11389<= not (I14399 and I14400);
	G11394<= not (G9600 and G3661);
	G11395<= not (G9601 and G3983);
	G11396<= not (G8713 and G4688);
	G11405<= not (G2741 and G2735 and G6856 and G2748);
	G11409<= not (G9842 and G3298);
	G11410<= not (G6875 and G6895 and G8696);
	G11411<= not (G9713 and G3625);
	G11412<= not (G8666 and G6918 and G8697);
	G11419<= not (I14428 and I14429);
	G11424<= not (G9662 and G4012);
	G11426<= not (G8742 and G4878);
	G11432<= not (G10295 and G8864);
	G11441<= not (G9599 and G3267);
	G11442<= not (G8644 and G3288 and G3343);
	G11443<= not (G9916 and G3649);
	G11444<= not (G6905 and G6918 and G8733);
	G11445<= not (G9771 and G3976);
	G11446<= not (G8700 and G6941 and G8734);
	G11479<= not (G6875 and G3288 and G3347);
	G11480<= not (G10323 and G8906);
	G11489<= not (G9661 and G3618);
	G11490<= not (G8666 and G3639 and G3694);
	G11491<= not (G9982 and G4000);
	G11492<= not (G6928 and G6941 and G8756);
	G11511<= not (I14481 and I14482);
	G11533<= not (G6905 and G3639 and G3698);
	G11534<= not (G7121 and G8958);
	G11543<= not (G9714 and G3969);
	G11544<= not (G8700 and G3990 and G4045);
	G11545<= not (I14498 and I14499);
	G11559<= not (I14509 and I14510);
	G11561<= not (I14517 and I14518);
	G11590<= not (G6928 and G3990 and G4049);
	G11591<= not (I14531 and I14532);
	G11639<= not (G8933 and G4722);
	G11674<= not (G8676 and G4674);
	G11675<= not (G8984 and G4912);
	G11676<= not (G358 and G8944 and G376 and G385);
	G11679<= not (G8836 and G802);
	G11707<= not (G8718 and G4864);
	G11708<= not (G10147 and G10110);
	G11761<= not (I14610 and I14611);
	G11858<= not (G9014 and G3010);
	G11881<= not (G9060 and G3361);
	G11892<= not (G7777 and G9086);
	G11903<= not (G9099 and G3712);
	G11906<= not (I14713 and I14714);
	G11914<= not (G8187 and G1648);
	G11923<= not (I14734 and I14735);
	G11933<= not (G837 and G9334 and G7197);
	G11934<= not (G8139 and G8187);
	G11936<= not (G8241 and G1783);
	G11938<= not (G8259 and G2208);
	G11944<= not (I14765 and I14766);
	G11951<= not (G9166 and G847 and G703);
	G11952<= not (G1624 and G8187);
	G11953<= not (G8195 and G8241);
	G11955<= not (G8302 and G1917);
	G11957<= not (G8205 and G8259);
	G11959<= not (G8316 and G2342);
	G11961<= not (G9777 and G5105);
	G11962<= not (I14789 and I14790);
	G11968<= not (G837 and G9334 and G9086);
	G11969<= not (G7252 and G1636);
	G11970<= not (G1760 and G8241);
	G11971<= not (G8249 and G8302);
	G11973<= not (G8365 and G2051);
	G11974<= not (G2185 and G8259);
	G11975<= not (G8267 and G8316);
	G11977<= not (G8373 and G2476);
	G11979<= not (G9861 and G5452);
	G11980<= not (I14817 and I14818);
	G11990<= not (G9166 and G703);
	G11992<= not (G7275 and G1772);
	G11993<= not (G1894 and G8302);
	G11994<= not (G8310 and G8365);
	G11996<= not (G7280 and G2197);
	G11997<= not (G2319 and G8316);
	G11998<= not (G8324 and G8373);
	G12000<= not (G8418 and G2610);
	G12001<= not (I14854 and I14855);
	G12008<= not (G9932 and G5798);
	G12014<= not (G7197 and G703);
	G12016<= not (G1648 and G8093);
	G12019<= not (G7322 and G1906);
	G12020<= not (G2028 and G8365);
	G12022<= not (G7335 and G2331);
	G12023<= not (G2453 and G8373);
	G12024<= not (G8381 and G8418);
	G12028<= not (I14884 and I14885);
	G12035<= not (G10000 and G6144);
	G12042<= not (G9086 and G703);
	G12044<= not (G1657 and G8139);
	G12045<= not (G1783 and G8146);
	G12048<= not (G7369 and G2040);
	G12049<= not (G2208 and G8150);
	G12052<= not (G7387 and G2465);
	G12053<= not (G2587 and G8418);
	G12066<= not (I14924 and I14925);
	G12073<= not (G10058 and G6490);
	G12078<= not (G8187 and G8093);
	G12079<= not (G1792 and G8195);
	G12080<= not (G1917 and G8201);
	G12083<= not (G2217 and G8205);
	G12084<= not (G2342 and G8211);
	G12087<= not (G7431 and G2599);
	G12100<= not (I14956 and I14957);
	G12111<= not (G847 and G9166);
	G12112<= not (G8139 and G1624);
	G12114<= not (G8241 and G8146);
	G12115<= not (G1926 and G8249);
	G12116<= not (G2051 and G8255);
	G12118<= not (G8259 and G8150);
	G12119<= not (G2351 and G8267);
	G12120<= not (G2476 and G8273);
	G12124<= not (G8741 and G4674);
	G12125<= not (G9728 and G5101);
	G12136<= not (I14992 and I14993);
	G12144<= not (I15003 and I15004);
	G12145<= not (G8195 and G1760);
	G12147<= not (G8302 and G8201);
	G12148<= not (G2060 and G8310);
	G12149<= not (G8205 and G2185);
	G12151<= not (G8316 and G8211);
	G12152<= not (G2485 and G8324);
	G12153<= not (G2610 and G8330);
	G12155<= not (G7753 and G7717);
	G12159<= not (G8765 and G4864);
	G12169<= not (G9804 and G5448);
	G12185<= not (G9905 and G799);
	G12187<= not (I15042 and I15043);
	G12188<= not (G8249 and G1894);
	G12190<= not (G8365 and G8255);
	G12191<= not (I15052 and I15053);
	G12192<= not (G8267 and G2319);
	G12194<= not (G8373 and G8273);
	G12195<= not (G2619 and G8381);
	G12196<= not (G8764 and G4688);
	G12197<= not (G7296 and G5290);
	G12207<= not (G9887 and G5794);
	G12221<= not (I15079 and I15080);
	G12222<= not (G8310 and G2028);
	G12224<= not (I15088 and I15089);
	G12225<= not (G8324 and G2453);
	G12227<= not (G8418 and G8330);
	G12232<= not (G8804 and G4878);
	G12239<= not (I15106 and I15107);
	G12244<= not (G7343 and G5320);
	G12245<= not (G7344 and G5637);
	G12255<= not (G9958 and G6140);
	G12285<= not (I15122 and I15123);
	G12286<= not (I15129 and I15130);
	G12287<= not (G8381 and G2587);
	G12289<= not (G9978 and G9766 and G9708);
	G12292<= not (G4698 and G8933);
	G12293<= not (G7436 and G5283);
	G12294<= not (G10044 and G7018 and G10090);
	G12301<= not (I15148 and I15149);
	G12306<= not (G7394 and G5666);
	G12307<= not (G7395 and G5983);
	G12317<= not (G10026 and G6486);
	G12323<= not (G9480 and G640);
	G12332<= not (I15167 and I15168);
	G12336<= not (I15175 and I15176);
	G12340<= not (G4888 and G8984);
	G12341<= not (G7512 and G5308);
	G12342<= not (G7004 and G7018 and G10129);
	G12343<= not (G7470 and G5630);
	G12344<= not (G10093 and G7041 and G10130);
	G12351<= not (I15194 and I15195);
	G12356<= not (G7438 and G6012);
	G12357<= not (G7439 and G6329);
	G12369<= not (G9049 and G637);
	G12370<= not (I15213 and I15214);
	G12402<= not (G7704 and G10266);
	G12411<= not (G7393 and G5276);
	G12412<= not (G10044 and G5297 and G5348);
	G12413<= not (G7521 and G5654);
	G12414<= not (G7028 and G7041 and G10165);
	G12415<= not (G7496 and G5976);
	G12416<= not (G10133 and G7064 and G10166);
	G12423<= not (I15242 and I15243);
	G12428<= not (G7472 and G6358);
	G12429<= not (G7473 and G6675);
	G12431<= not (I15254 and I15255);
	G12436<= not (I15263 and I15264);
	G12449<= not (G7004 and G5297 and G5352);
	G12450<= not (G7738 and G10281);
	G12459<= not (G7437 and G5623);
	G12460<= not (G10093 and G5644 and G5694);
	G12461<= not (G7536 and G6000);
	G12462<= not (G7051 and G7064 and G10190);
	G12463<= not (G7513 and G6322);
	G12464<= not (G10169 and G7087 and G10191);
	G12471<= not (I15288 and I15289);
	G12476<= not (G7498 and G6704);
	G12478<= not (I15299 and I15300);
	G12482<= not (I15307 and I15308);
	G12491<= not (G7285 and G4462 and G6961);
	G12511<= not (G7028 and G5644 and G5698);
	G12512<= not (G7766 and G10312);
	G12521<= not (G7471 and G5969);
	G12522<= not (G10133 and G5990 and G6040);
	G12523<= not (G7563 and G6346);
	G12524<= not (G7074 and G7087 and G10212);
	G12525<= not (G7522 and G6668);
	G12526<= not (G10194 and G7110 and G10213);
	G12538<= not (I15334 and I15335);
	G12539<= not (I15341 and I15342);
	G12577<= not (G7051 and G5990 and G6044);
	G12578<= not (G7791 and G10341);
	G12587<= not (G7497 and G6315);
	G12588<= not (G10169 and G6336 and G6386);
	G12589<= not (G7591 and G6692);
	G12590<= not (G7097 and G7110 and G10229);
	G12592<= not (I15364 and I15365);
	G12628<= not (G7074 and G6336 and G6390);
	G12629<= not (G7812 and G7142);
	G12638<= not (G7514 and G6661);
	G12639<= not (G10194 and G6682 and G6732);
	G12644<= not (G10233 and G4531);
	G12686<= not (G7097 and G6682 and G6736);
	G12767<= not (G4467 and G6961);
	G12796<= not (G4467 and G6961);
	G12797<= not (G10275 and G7655 and G7643 and G7627);
	G12819<= not (G9848 and G6961);
	G12822<= not (G6978 and G7236 and G7224 and G7163);
	G12910<= not (G11002 and G10601);
	G12915<= not (G12806 and G12632);
	G12933<= not (G7150 and G10515);
	G12941<= not (G7167 and G10537);
	G12947<= not (G7184 and G10561);
	G12969<= not (G4388 and G7178 and G10476);
	G12971<= not (G9024 and G8977 and G10664);
	G12972<= not (G7209 and G10578);
	G12999<= not (G4392 and G10476 and G4401);
	G13000<= not (G7228 and G10598);
	G13040<= not (G5196 and G12002 and G5308 and G9780);
	G13043<= not (G10521 and G969);
	G13050<= not (G5543 and G12029 and G5654 and G9864);
	G13057<= not (G969 and G11294);
	G13058<= not (G10544 and G1312);
	G13066<= not (G4430 and G7178 and G10590);
	G13067<= not (G5240 and G12059 and G5331 and G9780);
	G13069<= not (G5889 and G12067 and G6000 and G9935);
	G13079<= not (G1312 and G11336);
	G13083<= not (G4392 and G10590 and G4434);
	G13084<= not (G5587 and G12093 and G5677 and G9864);
	G13086<= not (G6235 and G12101 and G6346 and G10003);
	G13092<= not (G1061 and G10761);
	G13093<= not (G10649 and G7661 and G979 and G1061);
	G13097<= not (G5204 and G12002 and G5339 and G9780);
	G13098<= not (G5933 and G12129 and G6023 and G9935);
	G13100<= not (G6581 and G12137 and G6692 and G10061);
	G13102<= not (G7523 and G10759);
	G13104<= not (G1404 and G10794);
	G13105<= not (G10671 and G7675 and G1322 and G1404);
	G13108<= not (G5551 and G12029 and G5685 and G9864);
	G13109<= not (G6279 and G12173 and G6369 and G10003);
	G13115<= not (G1008 and G11786 and G11294);
	G13118<= not (G5897 and G12067 and G6031 and G9935);
	G13119<= not (G6625 and G12211 and G6715 and G10061);
	G13121<= not (G11117 and G8411);
	G13124<= not (G10666 and G7661 and G979 and G1061);
	G13130<= not (G1351 and G11815 and G11336);
	G13131<= not (G6243 and G12101 and G6377 and G10003);
	G13134<= not (G11134 and G8470);
	G13137<= not (G10699 and G7675 and G1322 and G1404);
	G13139<= not (G6589 and G12137 and G6723 and G10061);
	G13143<= not (G10695 and G7661 and G979 and G1061);
	G13176<= not (G10715 and G7675 and G1322 and G1404);
	G13210<= not (G7479 and G10521);
	G13217<= not (G4082 and G10808);
	G13240<= not (G1046 and G10521);
	G13241<= not (G7503 and G10544);
	G13248<= not (G9985 and G12399 and G9843);
	G13256<= not (G11846 and G11294 and G11812);
	G13257<= not (G1389 and G10544);
	G13260<= not (G1116 and G10666);
	G13264<= not (G11869 and G11336 and G11849);
	G13266<= not (G12440 and G9920 and G9843);
	G13273<= not (G1459 and G10699);
	G13281<= not (G10916 and G1099);
	G13283<= not (G12440 and G12399 and G9843);
	G13284<= not (G10695 and G1157);
	G13288<= not (G10946 and G1442);
	G13291<= not (G10715 and G1500);
	G13307<= not (G1116 and G10695);
	G13315<= not (G1459 and G10715);
	G13330<= not (G4664 and G11006);
	G13346<= not (G4854 and G11012);
	G13432<= not (G4793 and G10831);
	G13459<= not (G7479 and G11294 and G11846);
	G13462<= not (G12449 and G12412 and G12342 and G12294);
	G13464<= not (G10831 and G4793 and G4776);
	G13469<= not (G4983 and G10862);
	G13475<= not (G1008 and G11294 and G11786);
	G13476<= not (G7503 and G11336 and G11869);
	G13478<= not (G12511 and G12460 and G12414 and G12344);
	G13479<= not (G12686 and G12639 and G12590 and G12526);
	G13486<= not (G10862 and G4983 and G4966);
	G13495<= not (G1008 and G11786 and G7972);
	G13496<= not (G1351 and G11336 and G11815);
	G13498<= not (G12577 and G12522 and G12462 and G12416);
	G13499<= not (G11479 and G11442 and G11410 and G11382);
	G13511<= not (G182 and G174 and G203 and G12812);
	G13513<= not (G1351 and G11815 and G8002);
	G13515<= not (G12628 and G12588 and G12524 and G12464);
	G13516<= not (G11533 and G11490 and G11444 and G11412);
	G13527<= not (G182 and G168 and G203 and G12812);
	G13528<= not (G11294 and G7549 and G1008);
	G13529<= not (G11590 and G11544 and G11492 and G11446);
	G13544<= not (G7972 and G10521 and G7549 and G1008);
	G13551<= not (G11812 and G7479 and G7903 and G10521);
	G13554<= not (G11336 and G7582 and G1351);
	G13573<= not (G8002 and G10544 and G7582 and G1351);
	G13580<= not (G11849 and G7503 and G7922 and G10544);
	G13600<= not (G3021 and G11039);
	G13627<= not (G11172 and G8388);
	G13628<= not (G3372 and G11107);
	G13634<= not (G11797 and G11261);
	G13666<= not (G11190 and G8441);
	G13667<= not (G3723 and G11119);
	G13672<= not (G8933 and G11261);
	G13676<= not (G11834 and G11283);
	G13708<= not (G11200 and G8507);
	G13709<= not (G11755 and G11261);
	G13712<= not (G8984 and G11283);
	G13727<= not (G174 and G203 and G168 and G12812);
	G13739<= not (G11773 and G11261);
	G13742<= not (G11780 and G11283);
	G13756<= not (G203 and G12812);
	G13764<= not (G11252 and G3072);
	G13779<= not (G11804 and G11283);
	G13795<= not (G11216 and G401);
	G13797<= not (G8102 and G11273);
	G13798<= not (G11280 and G3423);
	G13821<= not (G11251 and G8340);
	G13822<= not (G8160 and G11306);
	G13823<= not (G11313 and G3774);
	G13834<= not (G4754 and G11773);
	G13846<= not (G1116 and G10649);
	G13850<= not (G11279 and G8396);
	G13851<= not (G8224 and G11360);
	G13854<= not (G4765 and G11797);
	G13855<= not (G4944 and G11804);
	G13861<= not (G1459 and G10671);
	G13866<= not (G3239 and G11194 and G3321 and G11519);
	G13867<= not (G11312 and G8449);
	G13870<= not (G11773 and G4732);
	G13871<= not (G4955 and G11834);
	G13873<= not (G11566 and G11729);
	G13882<= not (G3590 and G11207 and G3672 and G11576);
	G13884<= not (G11797 and G4727);
	G13886<= not (G11804 and G4922);
	G13889<= not (G11566 and G11435);
	G13892<= not (G11653 and G11473);
	G13896<= not (G3227 and G11194 and G3281 and G11350);
	G13897<= not (G3211 and G11217 and G3329 and G11519);
	G13898<= not (G11621 and G11747);
	G13907<= not (G3941 and G11225 and G4023 and G11631);
	G13909<= not (G11396 and G8847 and G11674 and G8803);
	G13911<= not (G11834 and G4917);
	G13915<= not (G11566 and G11473);
	G13918<= not (G3259 and G11217 and G3267 and G11350);
	G13920<= not (G11621 and G11483);
	G13923<= not (G11692 and G11527);
	G13927<= not (G3578 and G11207 and G3632 and G11389);
	G13928<= not (G3562 and G11238 and G3680 and G11576);
	G13929<= not (G11669 and G11763);
	G13940<= not (G11426 and G8889 and G11707 and G8829);
	G13945<= not (G691 and G11740);
	G13948<= not (G11610 and G8864);
	G13951<= not (G10295 and G11729);
	G13955<= not (G11621 and G11527);
	G13958<= not (G3610 and G11238 and G3618 and G11389);
	G13960<= not (G11669 and G11537);
	G13963<= not (G11715 and G11584);
	G13967<= not (G3929 and G11225 and G3983 and G11419);
	G13968<= not (G3913 and G11255 and G4031 and G11631);
	G13977<= not (G11610 and G11729);
	G13980<= not (G10295 and G11435);
	G13983<= not (G11658 and G8906);
	G13986<= not (G10323 and G11747);
	G13990<= not (G11669 and G11584);
	G13993<= not (G3961 and G11255 and G3969 and G11419);
	G14005<= not (G11514 and G11729);
	G14008<= not (G11610 and G11435);
	G14011<= not (G10295 and G11473);
	G14014<= not (G3199 and G11217 and G3298 and G11519);
	G14015<= not (G11658 and G11747);
	G14018<= not (G10323 and G11483);
	G14021<= not (G11697 and G8958);
	G14024<= not (G7121 and G11763);
	G14038<= not (G11514 and G11435);
	G14041<= not (G11610 and G11473);
	G14045<= not (G11571 and G11747);
	G14048<= not (G11658 and G11483);
	G14051<= not (G10323 and G11527);
	G14054<= not (G3550 and G11238 and G3649 and G11576);
	G14055<= not (G11697 and G11763);
	G14058<= not (G7121 and G11537);
	G14066<= not (G11514 and G11473);
	G14069<= not (G11653 and G8864);
	G14072<= not (G11571 and G11483);
	G14075<= not (G11658 and G11527);
	G14079<= not (G11626 and G11763);
	G14082<= not (G11697 and G11537);
	G14085<= not (G7121 and G11584);
	G14088<= not (G3901 and G11255 and G4000 and G11631);
	G14089<= not (G11755 and G4717);
	G14098<= not (G11566 and G8864);
	G14101<= not (G11653 and G11729);
	G14104<= not (G11514 and G8864);
	G14107<= not (G11571 and G11527);
	G14110<= not (G11692 and G8906);
	G14113<= not (G11626 and G11537);
	G14116<= not (G11697 and G11584);
	G14120<= not (G11780 and G4907);
	G14123<= not (G10685 and G10928);
	G14127<= not (G11653 and G11435);
	G14130<= not (G11621 and G8906);
	G14133<= not (G11692 and G11747);
	G14136<= not (G11571 and G8906);
	G14139<= not (G11626 and G11584);
	G14142<= not (G11715 and G8958);
	G14146<= not (G11020 and G691);
	G14151<= not (G11692 and G11483);
	G14154<= not (G11669 and G8958);
	G14157<= not (G11715 and G11763);
	G14160<= not (G11626 and G8958);
	G14170<= not (G11715 and G11537);
	G14177<= not (G11741 and G11721 and G753);
	G14223<= not (G9092 and G11858);
	G14234<= not (G9177 and G11881);
	G14254<= not (G11968 and G11933 and G11951);
	G14258<= not (G9203 and G11903);
	G14279<= not (G12111 and G9246);
	G14317<= not (G5033 and G11862);
	G14333<= not (G12042 and G12014 and G11990 and G11892);
	G14343<= not (G11961 and G9670);
	G14344<= not (G5377 and G11885);
	G14378<= not (G11979 and G9731);
	G14379<= not (G5723 and G11907);
	G14407<= not (G12008 and G9807);
	G14408<= not (G6069 and G11924);
	G14422<= not (G3187 and G11194 and G3298 and G8481);
	G14433<= not (G12035 and G9890);
	G14434<= not (G6415 and G11945);
	G14452<= not (G3538 and G11207 and G3649 and G8542);
	G14489<= not (G12126 and G5084);
	G14505<= not (G12073 and G9961);
	G14517<= not (G3231 and G11217 and G3321 and G8481);
	G14519<= not (G3889 and G11225 and G4000 and G8595);
	G14520<= not (G9369 and G12163);
	G14521<= not (G12170 and G5428);
	G14542<= not (G3582 and G11238 and G3672 and G8542);
	G14546<= not (G12125 and G9613);
	G14547<= not (G9439 and G12201);
	G14548<= not (G12208 and G5774);
	G14569<= not (G3195 and G11194 and G3329 and G8481);
	G14570<= not (G3933 and G11255 and G4023 and G8595);
	G14572<= not (G12169 and G9678);
	G14573<= not (G9506 and G12249);
	G14574<= not (G12256 and G6120);
	G14590<= not (G3546 and G11207 and G3680 and G8542);
	G14596<= not (G12196 and G9775 and G12124 and G9663);
	G14598<= not (G5248 and G12002 and G5331 and G12497);
	G14599<= not (G12207 and G9739);
	G14600<= not (G9564 and G12311);
	G14601<= not (G12318 and G6466);
	G14625<= not (G3897 and G11225 and G4031 and G8595);
	G14626<= not (G12232 and G9852 and G12159 and G9715);
	G14627<= not (G12553 and G12772);
	G14636<= not (G5595 and G12029 and G5677 and G12563);
	G14637<= not (G12255 and G9815);
	G14638<= not (G9626 and G12361);
	G14655<= not (G4743 and G11755);
	G14656<= not (G12553 and G12405);
	G14659<= not (G12646 and G12443);
	G14663<= not (G5236 and G12002 and G5290 and G12239);
	G14664<= not (G5220 and G12059 and G5339 and G12497);
	G14665<= not (G12604 and G12798);
	G14674<= not (G5941 and G12067 and G6023 and G12614);
	G14675<= not (G12317 and G9898);
	G14677<= not (I16779 and I16780);
	G14682<= not (G4933 and G11780);
	G14683<= not (G12553 and G12443);
	G14686<= not (G5268 and G12059 and G5276 and G12239);
	G14688<= not (G12604 and G12453);
	G14691<= not (G12695 and G12505);
	G14695<= not (G5583 and G12029 and G5637 and G12301);
	G14696<= not (G5567 and G12093 and G5685 and G12563);
	G14697<= not (G12662 and G12824);
	G14706<= not (G6287 and G12101 and G6369 and G12672);
	G14720<= not (G12593 and G10266);
	G14723<= not (G7704 and G12772);
	G14727<= not (G12604 and G12505);
	G14730<= not (G5615 and G12093 and G5623 and G12301);
	G14732<= not (G12662 and G12515);
	G14735<= not (G12739 and G12571);
	G14739<= not (G5929 and G12067 and G5983 and G12351);
	G14740<= not (G5913 and G12129 and G6031 and G12614);
	G14741<= not (G12711 and G10421);
	G14750<= not (G6633 and G12137 and G6715 and G12721);
	G14755<= not (G12593 and G12772);
	G14758<= not (G7704 and G12405);
	G14761<= not (G12651 and G10281);
	G14764<= not (G7738 and G12798);
	G14768<= not (G12662 and G12571);
	G14771<= not (G5961 and G12129 and G5969 and G12351);
	G14773<= not (G12711 and G12581);
	G14776<= not (G12780 and G12622);
	G14780<= not (G6275 and G12101 and G6329 and G12423);
	G14781<= not (G6259 and G12173 and G6377 and G12672);
	G14782<= not (G12755 and G10491);
	G14794<= not (G12492 and G12772);
	G14797<= not (G12593 and G12405);
	G14800<= not (G7704 and G12443);
	G14803<= not (G5208 and G12059 and G5308 and G12497);
	G14804<= not (G12651 and G12798);
	G14807<= not (G7738 and G12453);
	G14810<= not (G12700 and G10312);
	G14813<= not (G7766 and G12824);
	G14817<= not (G12711 and G12622);
	G14820<= not (G6307 and G12173 and G6315 and G12423);
	G14822<= not (G12755 and G12632);
	G14825<= not (G12806 and G12680);
	G14829<= not (G6621 and G12137 and G6675 and G12471);
	G14830<= not (G6605 and G12211 and G6723 and G12721);
	G14838<= not (G12492 and G12405);
	G14841<= not (G12593 and G12443);
	G14845<= not (G12558 and G12798);
	G14848<= not (G12651 and G12453);
	G14851<= not (G7738 and G12505);
	G14854<= not (G5555 and G12093 and G5654 and G12563);
	G14855<= not (G12700 and G12824);
	G14858<= not (G7766 and G12515);
	G14861<= not (G12744 and G10341);
	G14864<= not (G7791 and G10421);
	G14868<= not (G12755 and G12680);
	G14871<= not (G6653 and G12211 and G6661 and G12471);
	G14876<= not (G12492 and G12443);
	G14879<= not (G12646 and G10266);
	G14882<= not (G12558 and G12453);
	G14885<= not (G12651 and G12505);
	G14889<= not (G12609 and G12824);
	G14892<= not (G12700 and G12515);
	G14895<= not (G7766 and G12571);
	G14898<= not (G5901 and G12129 and G6000 and G12614);
	G14899<= not (G12744 and G10421);
	G14902<= not (G7791 and G12581);
	G14905<= not (G12785 and G7142);
	G14908<= not (G7812 and G10491);
	G14915<= not (G12553 and G10266);
	G14918<= not (G12646 and G12772);
	G14921<= not (G12492 and G10266);
	G14924<= not (G12558 and G12505);
	G14927<= not (G12695 and G10281);
	G14930<= not (G12609 and G12515);
	G14933<= not (G12700 and G12571);
	G14937<= not (G12667 and G10421);
	G14940<= not (G12744 and G12581);
	G14943<= not (G7791 and G12622);
	G14946<= not (G6247 and G12173 and G6346 and G12672);
	G14947<= not (G12785 and G10491);
	G14950<= not (G7812 and G12632);
	G14953<= not (G12646 and G12405);
	G14956<= not (G12604 and G10281);
	G14959<= not (G12695 and G12798);
	G14962<= not (G12558 and G10281);
	G14965<= not (G12609 and G12571);
	G14968<= not (G12739 and G10312);
	G14971<= not (G12667 and G12581);
	G14974<= not (G12744 and G12622);
	G14978<= not (G12716 and G10491);
	G14981<= not (G12785 and G12632);
	G14984<= not (G7812 and G12680);
	G14987<= not (G6593 and G12211 and G6692 and G12721);
	G14993<= not (G12695 and G12453);
	G14996<= not (G12662 and G10312);
	G14999<= not (G12739 and G12824);
	G15002<= not (G12609 and G10312);
	G15005<= not (G12667 and G12622);
	G15008<= not (G12780 and G10341);
	G15011<= not (G12716 and G12632);
	G15014<= not (G12785 and G12680);
	G15018<= not (G12739 and G12515);
	G15021<= not (G12711 and G10341);
	G15024<= not (G12780 and G10421);
	G15027<= not (G12667 and G10341);
	G15030<= not (G12716 and G12680);
	G15033<= not (G12806 and G7142);
	G15036<= not (G12780 and G12581);
	G15039<= not (G12755 and G7142);
	G15042<= not (G12806 and G10491);
	G15045<= not (G12716 and G7142);
	G15572<= not (G12969 and G7219);
	G15581<= not (G7232 and G12999);
	G15591<= not (G4332 and G4322 and G13202);
	G15674<= not (G921 and G13110);
	G15695<= not (G1266 and G13125);
	G15702<= not (G13066 and G7293);
	G15708<= not (G7340 and G13083);
	G15709<= not (G5224 and G14399 and G5327 and G9780);
	G15710<= not (G319 and G13385);
	G15713<= not (G5571 and G14425 and G5673 and G9864);
	G15715<= not (G336 and G305 and G13385);
	G15717<= not (G10754 and G13092);
	G15719<= not (G5256 and G14490 and G5335 and G9780);
	G15720<= not (G5917 and G14497 and G6019 and G9935);
	G15721<= not (G7564 and G311 and G13385);
	G15723<= not (G10775 and G13104);
	G15725<= not (G5603 and G14522 and G5681 and G9864);
	G15726<= not (G6263 and G14529 and G6365 and G10003);
	G15728<= not (G5200 and G14399 and G5313 and G9780);
	G15729<= not (G5949 and G14549 and G6027 and G9935);
	G15730<= not (G6609 and G14556 and G6711 and G10061);
	G15734<= not (G5228 and G12059 and G5290 and G14631);
	G15735<= not (G5547 and G14425 and G5659 and G9864);
	G15736<= not (G6295 and G14575 and G6373 and G10003);
	G15737<= not (G13240 and G13115 and G7903 and G13210);
	G15741<= not (G5244 and G14490 and G5320 and G14631);
	G15742<= not (G5575 and G12093 and G5637 and G14669);
	G15743<= not (G5893 and G14497 and G6005 and G9935);
	G15744<= not (G6641 and G14602 and G6719 and G10061);
	G15748<= not (G13257 and G13130 and G7922 and G13241);
	G15751<= not (G5591 and G14522 and G5666 and G14669);
	G15752<= not (G5921 and G12129 and G5983 and G14701);
	G15753<= not (G6239 and G14529 and G6351 and G10003);
	G15780<= not (G5937 and G14549 and G6012 and G14701);
	G15781<= not (G6267 and G12173 and G6329 and G14745);
	G15782<= not (G6585 and G14556 and G6697 and G10061);
	G15787<= not (G6283 and G14575 and G6358 and G14745);
	G15788<= not (G6613 and G12211 and G6675 and G14786);
	G15798<= not (G6629 and G14602 and G6704 and G14786);
	G15829<= not (G4112 and G13831);
	G15832<= not (G7903 and G7479 and G13256);
	G15833<= not (G14714 and G12378 and G12337);
	G15843<= not (G7922 and G7503 and G13264);
	G15844<= not (G14714 and G9340 and G12378);
	G15853<= not (G14714 and G9417 and G12337);
	G15864<= not (G14833 and G12543 and G12487);
	G15867<= not (G14714 and G9417 and G9340);
	G15877<= not (G14833 and G9340 and G12543);
	G15904<= not (I17380 and I17381);
	G15907<= not (G14833 and G9417 and G12487);
	G15959<= not (I17405 and I17406);
	G15962<= not (G14833 and G9417 and G9340);
	G16069<= not (I17447 and I17448);
	G16093<= not (I17461 and I17462);
	G16097<= not (G13319 and G10998);
	G16119<= not (I17475 and I17476);
	G16155<= not (I17495 and I17496);
	G16181<= not (G13475 and G13495 and G13057 and G13459);
	G16196<= not (G13496 and G13513 and G13079 and G13476);
	G16225<= not (G13544 and G13528 and G13043);
	G16236<= not (G13573 and G13554 and G13058);
	G16238<= not (G4698 and G13883 and G12054);
	G16259<= not (G4743 and G13908 and G12054);
	G16260<= not (G4888 and G13910 and G12088);
	G16264<= not (G518 and G9158 and G13223);
	G16275<= not (G9291 and G13480);
	G16278<= not (G8102 and G8057 and G13664);
	G16281<= not (G4754 and G13937 and G12054);
	G16282<= not (G4933 and G13939 and G12088);
	G16291<= not (G13551 and G13545);
	G16296<= not (G9360 and G13501);
	G16299<= not (G8160 and G8112 and G13706);
	G16304<= not (G4765 and G13970 and G12054);
	G16306<= not (G4944 and G13971 and G12088);
	G16312<= not (G13580 and G13574);
	G16316<= not (G9429 and G13518);
	G16319<= not (G8224 and G8170 and G13736);
	G16321<= not (G4955 and G13996 and G12088);
	G16507<= not (G13797 and G13764);
	G16524<= not (G13822 and G13798);
	G16586<= not (G13851 and G13823);
	G16604<= not (G3251 and G11194 and G3267 and G13877);
	G16625<= not (G3203 and G13700 and G3274 and G11519);
	G16628<= not (G3602 and G11207 and G3618 and G13902);
	G16657<= not (G3554 and G13730 and G3625 and G11576);
	G16660<= not (G3953 and G11225 and G3969 and G13933);
	G16663<= not (G13854 and G13834 and G14655 and G12292);
	G16681<= not (I17884 and I17885);
	G16687<= not (G3255 and G13700 and G3325 and G11519);
	G16694<= not (G3905 and G13772 and G3976 and G11631);
	G16696<= not (G13871 and G13855 and G14682 and G12340);
	G16713<= not (I17924 and I17925);
	G16719<= not (G3243 and G13700 and G3310 and G11350);
	G16723<= not (G3606 and G13730 and G3676 and G11576);
	G16728<= not (G13884 and G13870 and G14089 and G11639);
	G16741<= not (G3207 and G13765 and G3303 and G11519);
	G16745<= not (G3594 and G13730 and G3661 and G11389);
	G16749<= not (G3957 and G13772 and G4027 and G11631);
	G16757<= not (G13911 and G13886 and G14120 and G11675);
	G16770<= not (G3263 and G13765 and G3274 and G8481);
	G16772<= not (G3558 and G13799 and G3654 and G11576);
	G16776<= not (G3945 and G13772 and G4012 and G11419);
	G16813<= not (G3614 and G13799 and G3625 and G8542);
	G16815<= not (G3909 and G13824 and G4005 and G11631);
	G16854<= not (G3965 and G13824 and G3976 and G8595);
	G16875<= not (G3223 and G13765 and G3317 and G11519);
	G16893<= not (G10685 and G13252 and G703);
	G16925<= not (G3574 and G13799 and G3668 and G11576);
	G16956<= not (G3925 and G13824 and G4019 and G11631);
	G17137<= not (G13727 and G13511 and G13527);
	G17217<= not (G7239 and G14194);
	G17220<= not (G9369 and G9298 and G14376);
	G17225<= not (G8612 and G14367);
	G17243<= not (G7247 and G14212);
	G17246<= not (G9439 and G9379 and G14405);
	G17287<= not (G7262 and G14228);
	G17290<= not (G9506 and G9449 and G14431);
	G17297<= not (G2729 and G14291);
	G17312<= not (G7297 and G14248);
	G17315<= not (G9564 and G9516 and G14503);
	G17363<= not (G8635 and G14367);
	G17364<= not (G8639 and G14367);
	G17396<= not (G7345 and G14272);
	G17399<= not (G9626 and G9574 and G14535);
	G17412<= not (G14520 and G14489);
	G17468<= not (G3215 and G13700 and G3317 and G8481);
	G17474<= not (G14547 and G14521);
	G17492<= not (G8655 and G14367);
	G17493<= not (G8659 and G14367);
	G17495<= not (G3566 and G13730 and G3668 and G8542);
	G17500<= not (G14573 and G14548);
	G17513<= not (G3247 and G13765 and G3325 and G8481);
	G17514<= not (G3917 and G13772 and G4019 and G8595);
	G17520<= not (G5260 and G12002 and G5276 and G14631);
	G17525<= not (G14600 and G14574);
	G17568<= not (I18486 and I18487);
	G17571<= not (G8579 and G14367);
	G17572<= not (G3598 and G13799 and G3676 and G8542);
	G17578<= not (G5212 and G14399 and G5283 and G12497);
	G17581<= not (G5607 and G12029 and G5623 and G14669);
	G17586<= not (G14638 and G14601);
	G17592<= not (I18530 and I18531);
	G17593<= not (I18537 and I18538);
	G17595<= not (G8616 and G14367);
	G17596<= not (G8686 and G14367);
	G17597<= not (G3191 and G13700 and G3303 and G8481);
	G17598<= not (G3949 and G13824 and G4027 and G8595);
	G17605<= not (G5559 and G14425 and G5630 and G12563);
	G17608<= not (G5953 and G12067 and G5969 and G14701);
	G17618<= not (I18580 and I18581);
	G17624<= not (I18588 and I18589);
	G17634<= not (G3219 and G11217 and G3281 and G13877);
	G17635<= not (G3542 and G13730 and G3654 and G8542);
	G17640<= not (G5264 and G14399 and G5335 and G12497);
	G17647<= not (G5905 and G14497 and G5976 and G12614);
	G17650<= not (G6299 and G12101 and G6315 and G14745);
	G17656<= not (I18626 and I18627);
	G17662<= not (I18634 and I18635);
	G17668<= not (G3235 and G13765 and G3310 and G13877);
	G17669<= not (G3570 and G11238 and G3632 and G13902);
	G17670<= not (G3893 and G13772 and G4005 and G8595);
	G17675<= not (G5252 and G14399 and G5320 and G12239);
	G17679<= not (G5611 and G14425 and G5681 and G12563);
	G17686<= not (G6251 and G14529 and G6322 and G12672);
	G17689<= not (G6645 and G12137 and G6661 and G14786);
	G17699<= not (I18681 and I18682);
	G17705<= not (G3586 and G13799 and G3661 and G13902);
	G17706<= not (G3921 and G11255 and G3983 and G13933);
	G17708<= not (G5216 and G14490 and G5313 and G12497);
	G17712<= not (G5599 and G14425 and G5666 and G12301);
	G17716<= not (G5957 and G14497 and G6027 and G12614);
	G17723<= not (G6597 and G14556 and G6668 and G12721);
	G17732<= not (G3937 and G13824 and G4012 and G13933);
	G17734<= not (G5272 and G14490 and G5283 and G9780);
	G17736<= not (G5563 and G14522 and G5659 and G12563);
	G17740<= not (G5945 and G14497 and G6012 and G12351);
	G17744<= not (G6303 and G14529 and G6373 and G12672);
	G17748<= not (G562 and G14708 and G12323);
	G17755<= not (G5619 and G14522 and G5630 and G9864);
	G17757<= not (G5909 and G14549 and G6005 and G12614);
	G17761<= not (G6291 and G14529 and G6358 and G12423);
	G17765<= not (G6649 and G14556 and G6719 and G12721);
	G17773<= not (G5965 and G14549 and G5976 and G9935);
	G17775<= not (G6255 and G14575 and G6351 and G12672);
	G17779<= not (G6637 and G14556 and G6704 and G12471);
	G17788<= not (G5232 and G14490 and G5327 and G12497);
	G17790<= not (G6311 and G14575 and G6322 and G10003);
	G17792<= not (G6601 and G14602 and G6697 and G12721);
	G17814<= not (G5579 and G14522 and G5673 and G12563);
	G17816<= not (G6657 and G14602 and G6668 and G10061);
	G17820<= not (G5925 and G14549 and G6019 and G12614);
	G17846<= not (G6271 and G14575 and G6365 and G12672);
	G17872<= not (G6617 and G14602 and G6711 and G12721);
	G19265<= not (G15721 and G15715 and G13091 and G15710);
	G19335<= not (G15717 and G1056);
	G19358<= not (G15723 and G1399);
	G19442<= not (G11431 and G17794);
	G19450<= not (G11471 and G17794);
	G19455<= not (G15969 and G10841 and G7781);
	G19466<= not (G11562 and G17794);
	G19474<= not (G11609 and G17794);
	G19483<= not (G15969 and G10841 and G10922);
	G19495<= not (G15969 and G10841 and G7781);
	G19506<= not (G4087 and G15825);
	G19510<= not (G15969 and G10841 and G10899);
	G19513<= not (G15969 and G10841 and G10922);
	G19530<= not (G15829 and G10841);
	G19546<= not (G15969 and G10841 and G10884);
	G19549<= not (G15969 and G10841 and G10899);
	G19589<= not (G15969 and G10841 and G10884);
	G19597<= not (G1199 and G15995);
	G19611<= not (G1070 and G1199 and G15995);
	G19614<= not (G1542 and G16047);
	G19632<= not (G1413 and G1542 and G16047);
	G19764<= not (I20166 and I20167);
	G19782<= not (I20188 and I20189);
	G19792<= not (I20204 and I20205);
	G19795<= not (G13600 and G16275);
	G19854<= not (I20222 and I20223);
	G19856<= not (G13626 and G16278 and G8105);
	G19857<= not (G13628 and G16296);
	G19874<= not (G13665 and G16299 and G8163);
	G19875<= not (G13667 and G16316);
	G19886<= not (G11403 and G17794);
	G19903<= not (G13707 and G16319 and G8227);
	G19913<= not (G11430 and G17794);
	G19916<= not (G3029 and G16313);
	G19962<= not (G11470 and G17794);
	G19965<= not (G3380 and G16424);
	G20007<= not (G11512 and G17794);
	G20011<= not (G3731 and G16476);
	G20039<= not (G11250 and G17794);
	G20055<= not (G11269 and G17794);
	G20068<= not (G11293 and G17794);
	G20076<= not (G13795 and G16521);
	G20081<= not (G11325 and G17794);
	G20092<= not (G11373 and G17794);
	G20107<= not (G11404 and G17794);
	G20111<= not (G17513 and G14517 and G17468 and G14422);
	G20133<= not (G17668 and G17634 and G17597 and G14569);
	G20134<= not (G17572 and G14542 and G17495 and G14452);
	G20150<= not (G17705 and G17669 and G17635 and G14590);
	G20151<= not (G17598 and G14570 and G17514 and G14519);
	G20161<= not (G17732 and G17706 and G17670 and G14625);
	G20163<= not (G16663 and G13938);
	G20170<= not (G16741 and G13897 and G16687 and G13866);
	G20172<= not (G16876 and G8131);
	G20173<= not (G16696 and G13972);
	G20181<= not (G13252 and G16846);
	G20184<= not (G16770 and G13918 and G16719 and G13896);
	G20185<= not (G16772 and G13928 and G16723 and G13882);
	G20186<= not (G16926 and G8177);
	G20198<= not (G16813 and G13958 and G16745 and G13927);
	G20199<= not (G16815 and G13968 and G16749 and G13907);
	G20200<= not (I20461 and I20462);
	G20201<= not (I20468 and I20469);
	G20214<= not (G16854 and G13993 and G16776 and G13967);
	G20216<= not (I20487 and I20488);
	G20236<= not (G16875 and G14014 and G16625 and G16604);
	G20248<= not (G17056 and G14146 and G14123);
	G20271<= not (G16925 and G14054 and G16657 and G16628);
	G20371<= not (G16956 and G14088 and G16694 and G16660);
	G20619<= not (G14317 and G17217);
	G20644<= not (G14342 and G17220 and G9372);
	G20645<= not (G14344 and G17243);
	G20675<= not (G14377 and G17246 and G9442);
	G20676<= not (G14379 and G17287);
	G20733<= not (G14406 and G17290 and G9509);
	G20734<= not (G14408 and G17312);
	G20783<= not (G14616 and G17225);
	G20784<= not (G14616 and G17595);
	G20838<= not (G5041 and G17284);
	G20870<= not (G14432 and G17315 and G9567);
	G20871<= not (G14434 and G17396);
	G20979<= not (G5385 and G17309);
	G21011<= not (G14504 and G17399 and G9629);
	G21124<= not (G5731 and G17393);
	G21186<= not (G14616 and G17363);
	G21187<= not (G14616 and G17364);
	G21190<= not (G6077 and G17420);
	G21253<= not (G6423 and G17482);
	G21272<= not (G11268 and G17157);
	G21283<= not (G11291 and G17157);
	G21287<= not (G14616 and G17571);
	G21288<= not (G14616 and G17492);
	G21289<= not (G14616 and G17493);
	G21294<= not (G11324 and G17157);
	G21301<= not (G11371 and G17157);
	G21307<= not (G15719 and G13067 and G15709 and G13040);
	G21330<= not (G11401 and G17157);
	G21331<= not (G11402 and G17157);
	G21334<= not (G14616 and G17596);
	G21338<= not (G15741 and G15734 and G15728 and G13097);
	G21339<= not (G15725 and G13084 and G15713 and G13050);
	G21344<= not (G11428 and G17157);
	G21345<= not (G11429 and G17157);
	G21350<= not (G15751 and G15742 and G15735 and G13108);
	G21351<= not (G15729 and G13098 and G15720 and G13069);
	G21353<= not (G11467 and G17157);
	G21354<= not (G11468 and G17157);
	G21356<= not (G15780 and G15752 and G15743 and G13118);
	G21357<= not (G15736 and G13109 and G15726 and G13086);
	G21359<= not (G11509 and G17157);
	G21360<= not (G11510 and G17157);
	G21363<= not (G17708 and G14664 and G17640 and G14598);
	G21364<= not (G15787 and G15781 and G15753 and G13131);
	G21365<= not (G15744 and G13119 and G15730 and G13100);
	G21377<= not (G11560 and G17157);
	G21384<= not (G17734 and G14686 and G17675 and G14663);
	G21385<= not (G17736 and G14696 and G17679 and G14636);
	G21386<= not (G15798 and G15788 and G15782 and G13139);
	G21388<= not (G11608 and G17157);
	G21401<= not (G17755 and G14730 and G17712 and G14695);
	G21402<= not (G17757 and G14740 and G17716 and G14674);
	G21403<= not (G11652 and G17157);
	G21415<= not (G17773 and G14771 and G17740 and G14739);
	G21416<= not (G17775 and G14781 and G17744 and G14706);
	G21417<= not (G11677 and G17157);
	G21429<= not (G17788 and G14803 and G17578 and G17520);
	G21432<= not (G17790 and G14820 and G17761 and G14780);
	G21433<= not (G17792 and G14830 and G17765 and G14750);
	G21459<= not (G17814 and G14854 and G17605 and G17581);
	G21462<= not (G17816 and G14871 and G17779 and G14829);
	G21509<= not (G17820 and G14898 and G17647 and G17608);
	G21555<= not (G17846 and G14946 and G17686 and G17650);
	G21603<= not (G17872 and G14987 and G17723 and G17689);
	G22306<= not (G4584 and G4616 and G13202 and G19071);
	G22312<= not (G907 and G19063);
	G22325<= not (G1252 and G19140);
	G22638<= not (G18957 and G2886);
	G22642<= not (G7870 and G19560);
	G22643<= not (G20136 and G18954);
	G22650<= not (G7888 and G19581);
	G22651<= not (G20114 and G2873);
	G22661<= not (G20136 and G94);
	G22663<= not (I21977 and I21978);
	G22666<= not (G18957 and G2878);
	G22668<= not (G20219 and G2912);
	G22681<= not (I21993 and I21994);
	G22687<= not (G19560 and G7870);
	G22688<= not (G20219 and G2936);
	G22709<= not (G1193 and G19611);
	G22711<= not (G19581 and G7888);
	G22712<= not (G18957 and G2864);
	G22713<= not (G20114 and G2890);
	G22715<= not (G20114 and G2999);
	G22753<= not (G1536 and G19632);
	G22754<= not (G20114 and G19376);
	G22755<= not (G20136 and G18984);
	G22757<= not (G20114 and G7891);
	G22833<= not (G1193 and G19560 and G10666);
	G22836<= not (G18918 and G2852);
	G22837<= not (G20219 and G2907);
	G22838<= not (G20219 and G2960);
	G22839<= not (G20114 and G2988);
	G22850<= not (G1536 and G19581 and G10699);
	G22852<= not (G18957 and G2856);
	G22853<= not (G20219 and G2922);
	G22864<= not (G7780 and G21156);
	G22874<= not (G18918 and G2844);
	G22875<= not (G20516 and G2980);
	G22885<= not (G9104 and G20154);
	G22902<= not (G18957 and G2848);
	G22908<= not (G9104 and G20175);
	G22921<= not (G20219 and G2950);
	G22940<= not (G18918 and G2860);
	G22941<= not (G20219 and G2970);
	G22984<= not (G20114 and G2868);
	G23010<= not (G20516 and G2984);
	G23047<= not (G482 and G20000);
	G23067<= not (G20887 and G10721);
	G23105<= not (G8097 and G19887);
	G23112<= not (G21024 and G10733);
	G23132<= not (G8155 and G19932);
	G23139<= not (G21163 and G10756);
	G23167<= not (G8219 and G19981);
	G23195<= not (G20136 and G37);
	G23210<= not (G18957 and G2882);
	G23266<= not (G18918 and G2894);
	G23281<= not (G18957 and G2898);
	G23286<= not (G6875 and G20887);
	G23309<= not (G6905 and G21024);
	G23324<= not (G703 and G20181);
	G23342<= not (G6928 and G21163);
	G23357<= not (G20201 and G11231);
	G23379<= not (G20216 and G11248);
	G23428<= not (G13945 and G20522);
	G23552<= not (I22684 and I22685);
	G23575<= not (I22711 and I22712);
	G23576<= not (I22718 and I22719);
	G23590<= not (G20682 and G11111);
	G23616<= not (I22754 and I22755);
	G23617<= not (I22761 and I22762);
	G23623<= not (G9364 and G20717);
	G23630<= not (G20739 and G11123);
	G23655<= not (I22793 and I22794);
	G23656<= not (I22800 and I22801);
	G23659<= not (G9434 and G20854);
	G23666<= not (G20875 and G11139);
	G23685<= not (I22823 and I22824);
	G23692<= not (G9501 and G20995);
	G23699<= not (G21012 and G11160);
	G23719<= not (I22845 and I22846);
	G23726<= not (G9559 and G21140);
	G23733<= not (G20751 and G11178);
	G23747<= not (I22865 and I22866);
	G23748<= not (I22872 and I22873);
	G23756<= not (G9621 and G21206);
	G23761<= not (I22893 and I22894);
	G23762<= not (I22900 and I22901);
	G23778<= not (I22922 and I22923);
	G23780<= not (I22930 and I22931);
	G23781<= not (I22937 and I22938);
	G23782<= not (G2741 and G21062);
	G23786<= not (I22945 and I22946);
	G23809<= not (I22966 and I22967);
	G23810<= not (I22973 and I22974);
	G23850<= not (G12185 and G19462);
	G23890<= not (G7004 and G20682);
	G23909<= not (G7028 and G20739);
	G23932<= not (G7051 and G20875);
	G23949<= not (G7074 and G21012);
	G23972<= not (G7097 and G20751);
	G23975<= not (I23119 and I23120);
	G23978<= not (G572 and G21389 and G12323);
	G24362<= not (G21370 and G22136);
	G24369<= not (I23586 and I23587);
	G24380<= not (I23601 and I23602);
	G24528<= not (G4098 and G22654);
	G24544<= not (G22666 and G22661 and G22651);
	G24547<= not (G22638 and G22643 and G22754);
	G24566<= not (G22755 and G22713);
	G24567<= not (G22957 and G2917);
	G24570<= not (G22957 and G2941);
	G24574<= not (G22709 and G22687);
	G24576<= not (G22957 and G2902);
	G24583<= not (G22753 and G22711);
	G24584<= not (G22852 and G22836 and G22715);
	G24591<= not (G22833 and G22642);
	G24601<= not (G22957 and G2965);
	G24609<= not (G22850 and G22650);
	G24620<= not (G22902 and G22874);
	G24621<= not (G22957 and G2927);
	G24652<= not (G22712 and G22940 and G22757);
	G24661<= not (G23210 and G23195 and G22984);
	G24662<= not (G22957 and G2955);
	G24677<= not (G22957 and G2975);
	G24678<= not (G22994 and G23010);
	G24760<= not (I23918 and I23919);
	G24776<= not (G3040 and G23052);
	G24787<= not (G3391 and G23079);
	G24792<= not (I23950 and I23951);
	G24793<= not (G3742 and G23124);
	G24798<= not (I23962 and I23963);
	G24802<= not (I23970 and I23971);
	G24804<= not (G19916 and G23105);
	G24807<= not (I23979 and I23980);
	G24808<= not (I23986 and I23987);
	G24809<= not (G19965 and G23132);
	G24814<= not (G20011 and G23167);
	G24880<= not (G23281 and G23266 and G22839);
	G24890<= not (G13852 and G22929);
	G24905<= not (G534 and G23088);
	G24906<= not (G8743 and G23088);
	G24916<= not (G19450 and G23154);
	G24917<= not (G19913 and G23172);
	G24918<= not (G136 and G23088);
	G24924<= not (G20007 and G23172);
	G24925<= not (G20092 and G23154);
	G24926<= not (G20172 and G20163 and G23357 and G13995);
	G24932<= not (G19886 and G23172);
	G24933<= not (G19466 and G23154);
	G24934<= not (G21283 and G23462);
	G24936<= not (G20186 and G20173 and G23379 and G14029);
	G24942<= not (G20039 and G23172);
	G24943<= not (G20068 and G23172);
	G24944<= not (G21354 and G23363);
	G24950<= not (G19442 and G23154);
	G24951<= not (G199 and G23088);
	G24957<= not (G21359 and G23462);
	G24958<= not (G21330 and G23462);
	G24972<= not (G19962 and G23172);
	G24973<= not (G21272 and G23462);
	G24974<= not (G21301 and G23363);
	G24975<= not (G21388 and G23363);
	G24988<= not (G546 and G23088);
	G24989<= not (G21345 and G23363);
	G25002<= not (G19474 and G23154);
	G25003<= not (G21353 and G23462);
	G25018<= not (G20107 and G23154);
	G25019<= not (G20055 and G23172);
	G25020<= not (G21377 and G23462);
	G25021<= not (G21417 and G23363);
	G25038<= not (G21331 and G23363);
	G25048<= not (G542 and G23088);
	G25049<= not (G21344 and G23462);
	G25062<= not (G21403 and G23363);
	G25172<= not (G5052 and G23560);
	G25186<= not (G5396 and G23602);
	G25199<= not (I24364 and I24365);
	G25200<= not (G5742 and G23642);
	G25215<= not (I24384 and I24385);
	G25216<= not (G6088 and G23678);
	G25233<= not (G20838 and G23623);
	G25236<= not (I24415 and I24416);
	G25237<= not (G6434 and G23711);
	G25255<= not (G20979 and G23659);
	G25258<= not (I24439 and I24440);
	G25268<= not (G21124 and G23692);
	G25271<= not (I24462 and I24463);
	G25275<= not (G22342 and G11991);
	G25293<= not (G21190 and G23726);
	G25300<= not (G22369 and G12018);
	G25309<= not (G22384 and G12021);
	G25334<= not (G21253 and G23756);
	G25337<= not (G22342 and G1648 and G8187);
	G25341<= not (G22417 and G12047);
	G25349<= not (G22432 and G12051);
	G25381<= not (G538 and G23088);
	G25382<= not (G12333 and G22342);
	G25385<= not (G22369 and G1783 and G8241);
	G25389<= not (G22457 and G12082);
	G25396<= not (G22384 and G2208 and G8259);
	G25400<= not (G22472 and G12086);
	G25425<= not (G20081 and G23172);
	G25426<= not (G12371 and G22369);
	G25429<= not (G22417 and G1917 and G8302);
	G25432<= not (G12374 and G22384);
	G25435<= not (G22432 and G2342 and G8316);
	G25439<= not (G22498 and G12122);
	G25467<= not (G12432 and G22417);
	G25470<= not (G22457 and G2051 and G8365);
	G25473<= not (G12437 and G22432);
	G25476<= not (G22472 and G2476 and G8373);
	G25492<= not (G12479 and G22457);
	G25495<= not (G12483 and G22472);
	G25498<= not (G22498 and G2610 and G8418);
	G25514<= not (G12540 and G22498);
	G25527<= not (G21294 and G23462);
	G25531<= not (G22763 and G2868);
	G25532<= not (G21360 and G23363);
	G25537<= not (G22763 and G2873);
	G25779<= not (G19694 and G24362);
	G25888<= not (G914 and G24439);
	G25895<= not (G1259 and G24453);
	G25953<= not (G22756 and G24570 and G22688);
	G25974<= not (G24576 and G22837);
	G25984<= not (G24567 and G22668);
	G25985<= not (G24631 and G23956);
	G25995<= not (G24621 and G22853);
	G25996<= not (G24601 and G22838);
	G26025<= not (G22405 and G24631);
	G26052<= not (G22714 and G24662 and G22921);
	G26053<= not (G22875 and G24677 and G22941);
	G26208<= not (G7975 and G24751);
	G26235<= not (G8016 and G24766);
	G26248<= not (I25220 and I25221);
	G26255<= not (G8075 and G24779);
	G26269<= not (I25243 and I25244);
	G26352<= not (G744 and G24875 and G11679);
	G26382<= not (G577 and G24953 and G12323);
	G26666<= not (G9229 and G25144);
	G26685<= not (G9264 and G25160);
	G26714<= not (G9316 and G25175);
	G26745<= not (G6856 and G25317);
	G26752<= not (G9397 and G25189);
	G26782<= not (G9467 and G25203);
	G27141<= not (I25846 and I25847);
	G27223<= not (I25908 and I25909);
	G27273<= not (G10504 and G26131 and G26105);
	G27282<= not (G11192 and G26269 and G26248 and G479);
	G27295<= not (G24776 and G26208);
	G27306<= not (G24787 and G26235);
	G27317<= not (G24793 and G26255);
	G27365<= not (I26050 and I26051);
	G27377<= not (G10685 and G25930);
	G27380<= not (I26071 and I26072);
	G27401<= not (I26094 and I26095);
	G27463<= not (G287 and G26330 and G23204);
	G27468<= not (G24951 and G24932 and G24925 and G26852);
	G27550<= not (G24943 and G25772);
	G27577<= not (G25019 and G25002 and G24988 and G25765);
	G27582<= not (G10857 and G26131 and G26105);
	G27586<= not (G24924 and G24916 and G24905 and G26863);
	G27587<= not (G24917 and G25018 and G24918 and G26857);
	G27593<= not (G24972 and G24950 and G24906 and G26861);
	G27613<= not (G24942 and G24933 and G25048 and G26871);
	G27654<= not (G164 and G26598 and G23042);
	G27670<= not (G25172 and G26666);
	G27679<= not (G25186 and G26685);
	G27687<= not (G25200 and G26714);
	G27693<= not (G25216 and G26752);
	G27705<= not (G25237 and G26782);
	G27738<= not (G21228 and G25243 and G26424 and G26148);
	G27767<= not (I26367 and I26368);
	G27775<= not (G21228 and G25262 and G26424 and G26166);
	G27796<= not (G21228 and G25263 and G26424 and G26171);
	G27824<= not (I26394 and I26395);
	G27833<= not (G21228 and G25282 and G26424 and G26190);
	G27854<= not (G21228 and G25283 and G26424 and G26195);
	G27876<= not (I26418 and I26419);
	G27882<= not (G21228 and G25307 and G26424 and G26213);
	G27903<= not (G21228 and G25316 and G26424 and G26218);
	G27925<= not (I26439 and I26440);
	G27931<= not (G25425 and G25381 and G25780);
	G27933<= not (G21228 and G25356 and G26424 and G26236);
	G27955<= not (I26460 and I26461);
	G28109<= not (G27051 and G25783);
	G28131<= not (G27051 and G25838);
	G28167<= not (G925 and G27046);
	G28174<= not (G1270 and G27059);
	G28203<= not (G12546 and G27985 and G27977);
	G28206<= not (G12546 and G26105 and G27985);
	G28207<= not (G12546 and G26131 and G27977);
	G28259<= not (G10504 and G26987 and G26973);
	G28270<= not (G10504 and G26105 and G26987);
	G28271<= not (G10533 and G27004 and G26990);
	G28287<= not (G10504 and G26131 and G26973);
	G28288<= not (G10533 and G26105 and G27004);
	G28298<= not (G10533 and G26131 and G26990);
	G28336<= not (G27064 and G24756 and G27163 and G19644);
	G28349<= not (G27074 and G24770 and G27187 and G19644);
	G28363<= not (G27064 and G13593);
	G28376<= not (G27064 and G13620);
	G28381<= not (G27074 and G13621);
	G28391<= not (G27064 and G13637);
	G28395<= not (G27074 and G13655);
	G28406<= not (G27064 and G13675);
	G28410<= not (G27074 and G13679);
	G28421<= not (G27074 and G13715);
	G28448<= not (G23975 and G27377);
	G28500<= not (G590 and G27629 and G12323);
	G28504<= not (G758 and G27528 and G11679);
	G28512<= not (G10857 and G27155 and G27142);
	G28516<= not (G10857 and G26105 and G27155);
	G28522<= not (G10857 and G26131 and G27142);
	G28736<= not (G27742 and G7308 and G7252);
	G28755<= not (G27742 and G7268 and G1592);
	G28758<= not (G27779 and G7356 and G7275);
	G28765<= not (G27800 and G7374 and G7280);
	G28780<= not (G27742 and G7308 and G1636);
	G28783<= not (G27779 and G7315 and G1728);
	G28786<= not (G27837 and G7405 and G7322);
	G28793<= not (G27800 and G7328 and G2153);
	G28796<= not (G27858 and G7418 and G7335);
	G28820<= not (G27742 and G1668 and G1592);
	G28823<= not (G27738 and G14565);
	G28824<= not (G27779 and G7356 and G1772);
	G28827<= not (G27837 and G7362 and G1862);
	G28830<= not (G27886 and G7451 and G7369);
	G28837<= not (G27800 and G7374 and G2197);
	G28840<= not (G27858 and G7380 and G2287);
	G28843<= not (G27907 and G7456 and G7387);
	G28853<= not (G27742 and G1636 and G7252);
	G28856<= not (G27738 and G8093);
	G28857<= not (G27779 and G1802 and G1728);
	G28860<= not (G27775 and G14586);
	G28861<= not (G27837 and G7405 and G1906);
	G28864<= not (G27886 and G7411 and G1996);
	G28867<= not (G27800 and G2227 and G2153);
	G28870<= not (G27796 and G14588);
	G28871<= not (G27858 and G7418 and G2331);
	G28874<= not (G27907 and G7424 and G2421);
	G28877<= not (G27937 and G7490 and G7431);
	G28885<= not (G27742 and G1668 and G7268);
	G28888<= not (G27738 and G8139);
	G28892<= not (G27779 and G1772 and G7275);
	G28895<= not (G27775 and G8146);
	G28896<= not (G27837 and G1936 and G1862);
	G28899<= not (G27833 and G14612);
	G28900<= not (G27886 and G7451 and G2040);
	G28903<= not (G27800 and G2197 and G7280);
	G28906<= not (G27796 and G8150);
	G28907<= not (G27858 and G2361 and G2287);
	G28910<= not (G27854 and G14614);
	G28911<= not (G27907 and G7456 and G2465);
	G28914<= not (G27937 and G7462 and G2555);
	G28920<= not (G27779 and G1802 and G7315);
	G28923<= not (G27775 and G8195);
	G28927<= not (G27837 and G1906 and G7322);
	G28930<= not (G27833 and G8201);
	G28931<= not (G27886 and G2070 and G1996);
	G28934<= not (G27882 and G14641);
	G28935<= not (G27800 and G2227 and G7328);
	G28938<= not (G27796 and G8205);
	G28942<= not (G27858 and G2331 and G7335);
	G28945<= not (G27854 and G8211);
	G28946<= not (G27907 and G2495 and G2421);
	G28949<= not (G27903 and G14643);
	G28950<= not (G27937 and G7490 and G2599);
	G28955<= not (G27837 and G1936 and G7362);
	G28958<= not (G27833 and G8249);
	G28962<= not (G27886 and G2040 and G7369);
	G28965<= not (G27882 and G8255);
	G28966<= not (G27858 and G2361 and G7380);
	G28969<= not (G27854 and G8267);
	G28973<= not (G27907 and G2465 and G7387);
	G28976<= not (G27903 and G8273);
	G28977<= not (G27937 and G2629 and G2555);
	G28980<= not (G27933 and G14680);
	G28987<= not (G27886 and G2070 and G7411);
	G28990<= not (G27882 and G8310);
	G28994<= not (G27907 and G2495 and G7424);
	G28997<= not (G27903 and G8324);
	G29001<= not (G27937 and G2599 and G7431);
	G29004<= not (G27933 and G8330);
	G29015<= not (G27742 and G9586);
	G29018<= not (G9586 and G27742);
	G29025<= not (G27937 and G2629 and G7462);
	G29028<= not (G27933 and G8381);
	G29046<= not (G27779 and G9640);
	G29049<= not (G9640 and G27779);
	G29057<= not (G27800 and G9649);
	G29060<= not (G9649 and G27800);
	G29082<= not (G27837 and G9694);
	G29085<= not (G9694 and G27837);
	G29094<= not (G27858 and G9700);
	G29097<= not (G9700 and G27858);
	G29118<= not (G27886 and G9755);
	G29121<= not (G9755 and G27886);
	G29131<= not (G27907 and G9762);
	G29134<= not (G9762 and G27907);
	G29154<= not (G27937 and G9835);
	G29157<= not (G9835 and G27937);
	G29186<= not (G27051 and G4507);
	G29335<= not (G25540 and G28131);
	G29355<= not (G24383 and G28109);
	G29540<= not (G28336 and G13464);
	G29556<= not (G28349 and G13486);
	G29657<= not (G28363 and G13634);
	G29660<= not (G28448 and G9582);
	G29672<= not (G28376 and G13672);
	G29676<= not (G28381 and G13676);
	G29679<= not (G153 and G28353 and G23042);
	G29694<= not (G28391 and G13709);
	G29702<= not (G28395 and G13712);
	G29719<= not (G28406 and G13739);
	G29722<= not (G28410 and G13742);
	G29737<= not (G28421 and G13779);
	G29778<= not (G294 and G28444 and G23204);
	G30573<= not (G29355 and G19666);
	G30580<= not (G29335 and G19666);
	G31003<= not (G27163 and G29497 and G19644);
	G31009<= not (G27187 and G29503 and G19644);
	G31262<= not (G767 and G29916 and G11679);
	G31509<= not (G599 and G29933 and G12323);
	G31669<= not (I29254 and I29255);
	G31671<= not (I29262 and I29263);
	G31706<= not (I29270 and I29271);
	G31708<= not (I29278 and I29279);
	G31709<= not (I29285 and I29286);
	G31747<= not (I29296 and I29297);
	G31748<= not (I29303 and I29304);
	G31753<= not (I29314 and I29315);
	G31950<= not (G7285 and G30573);
	G31971<= not (G30573 and G10511);
	G31978<= not (G30580 and G15591);
	G31997<= not (G22306 and G30580);
	G32057<= not (G31003 and G13297);
	G32072<= not (G31009 and G13301);
	G33083<= not (G7805 and G32118);
	G33299<= not (G608 and G32296 and G12323);
	G33306<= not (G776 and G32212 and G11679);
	G33394<= not (G10159 and G4474 and G32426);
	G33669<= not (G33378 and G862);
	G33679<= not (G33394 and G10737 and G10308);
	G33838<= not (G33083 and G4369);
	G33925<= not (G33394 and G4462 and G4467);
	G33930<= not (G33394 and G12767 and G9848);
	G33933<= not (G33394 and G12491 and G12819 and G12796);
	G34048<= not (G33669 and G10583 and G7442);
	G34051<= not (I31973 and I31974);
	G34056<= not (I31984 and I31985);
	G34162<= not (G785 and G33823 and G11679);
	G34174<= not (G617 and G33851 and G12323);
	G34220<= not (I32186 and I32187);
	G34227<= not (I32203 and I32204);
	G34422<= not (I32432 and I32433);
	G34424<= not (I32440 and I32441);
	G34469<= not (I32517 and I32518);
	G34545<= not (G11679 and G794 and G34354);
	G34550<= not (G626 and G34359 and G12323);
	G34650<= not (I32757 and I32758);
	I11824<= not (G4593 and G4601);
	I11825<= not (G4593 and I11824);
	I11826<= not (G4601 and I11824);
	I11864<= not (G4434 and G4401);
	I11865<= not (G4434 and I11864);
	I11866<= not (G4401 and I11864);
	I11877<= not (G4388 and G4430);
	I11878<= not (G4388 and I11877);
	I11879<= not (G4430 and I11877);
	I12074<= not (G996 and G979);
	I12075<= not (G996 and I12074);
	I12076<= not (G979 and I12074);
	I12096<= not (G1339 and G1322);
	I12097<= not (G1339 and I12096);
	I12098<= not (G1322 and I12096);
	I12203<= not (G1094 and G1135);
	I12204<= not (G1094 and I12203);
	I12205<= not (G1135 and I12203);
	I12217<= not (G1437 and G1478);
	I12218<= not (G1437 and I12217);
	I12219<= not (G1478 and I12217);
	I12240<= not (G1111 and G1105);
	I12241<= not (G1111 and I12240);
	I12242<= not (G1105 and I12240);
	I12251<= not (G1124 and G1129);
	I12252<= not (G1124 and I12251);
	I12253<= not (G1129 and I12251);
	I12261<= not (G1454 and G1448);
	I12262<= not (G1454 and I12261);
	I12263<= not (G1448 and I12261);
	I12269<= not (G1141 and G956);
	I12270<= not (G1141 and I12269);
	I12271<= not (G956 and I12269);
	I12277<= not (G1467 and G1472);
	I12278<= not (G1467 and I12277);
	I12279<= not (G1472 and I12277);
	I12287<= not (G1484 and G1300);
	I12288<= not (G1484 and I12287);
	I12289<= not (G1300 and I12287);
	I12344<= not (G3106 and G3111);
	I12345<= not (G3106 and I12344);
	I12346<= not (G3111 and I12344);
	I12372<= not (G3457 and G3462);
	I12373<= not (G3457 and I12372);
	I12374<= not (G3462 and I12372);
	I12401<= not (G3808 and G3813);
	I12402<= not (G3808 and I12401);
	I12403<= not (G3813 and I12401);
	I12468<= not (G405 and G392);
	I12469<= not (G405 and I12468);
	I12470<= not (G392 and I12468);
	I12544<= not (G191 and G194);
	I12545<= not (G191 and I12544);
	I12546<= not (G194 and I12544);
	I12728<= not (G4291 and G4287);
	I12729<= not (G4291 and I12728);
	I12730<= not (G4287 and I12728);
	I12840<= not (G4222 and G4235);
	I12841<= not (G4222 and I12840);
	I12842<= not (G4235 and I12840);
	I12848<= not (G4281 and G4277);
	I12849<= not (G4281 and I12848);
	I12850<= not (G4277 and I12848);
	I12876<= not (G4200 and G4180);
	I12877<= not (G4200 and I12876);
	I12878<= not (G4180 and I12876);
	I13043<= not (G5115 and G5120);
	I13044<= not (G5115 and I13043);
	I13045<= not (G5120 and I13043);
	I13065<= not (G4308 and G4304);
	I13066<= not (G4308 and I13065);
	I13067<= not (G4304 and I13065);
	I13077<= not (G5462 and G5467);
	I13078<= not (G5462 and I13077);
	I13079<= not (G5467 and I13077);
	I13109<= not (G5808 and G5813);
	I13110<= not (G5808 and I13109);
	I13111<= not (G5813 and I13109);
	I13139<= not (G6154 and G6159);
	I13140<= not (G6154 and I13139);
	I13141<= not (G6159 and I13139);
	I13182<= not (G6500 and G6505);
	I13183<= not (G6500 and I13182);
	I13184<= not (G6505 and I13182);
	I13334<= not (G1687 and G1691);
	I13335<= not (G1687 and I13334);
	I13336<= not (G1691 and I13334);
	I13382<= not (G269 and G246);
	I13383<= not (G269 and I13382);
	I13384<= not (G246 and I13382);
	I13390<= not (G1821 and G1825);
	I13391<= not (G1821 and I13390);
	I13392<= not (G1825 and I13390);
	I13401<= not (G2246 and G2250);
	I13402<= not (G2246 and I13401);
	I13403<= not (G2250 and I13401);
	I13442<= not (G262 and G239);
	I13443<= not (G262 and I13442);
	I13444<= not (G239 and I13442);
	I13452<= not (G1955 and G1959);
	I13453<= not (G1955 and I13452);
	I13454<= not (G1959 and I13452);
	I13462<= not (G2380 and G2384);
	I13463<= not (G2380 and I13462);
	I13464<= not (G2384 and I13462);
	I13497<= not (G255 and G232);
	I13498<= not (G255 and I13497);
	I13499<= not (G232 and I13497);
	I13509<= not (G2089 and G2093);
	I13510<= not (G2089 and I13509);
	I13511<= not (G2093 and I13509);
	I13518<= not (G2514 and G2518);
	I13519<= not (G2514 and I13518);
	I13520<= not (G2518 and I13518);
	I13564<= not (G2648 and G2652);
	I13565<= not (G2648 and I13564);
	I13566<= not (G2652 and I13564);
	I13729<= not (G4534 and G4537);
	I13730<= not (G4534 and I13729);
	I13731<= not (G4537 and I13729);
	I13749<= not (G4608 and G4584);
	I13750<= not (G4608 and I13749);
	I13751<= not (G4584 and I13749);
	I13850<= not (G862 and G7397);
	I13851<= not (G862 and I13850);
	I13852<= not (G7397 and I13850);
	I14169<= not (G8389 and G3119);
	I14170<= not (G8389 and I14169);
	I14171<= not (G3119 and I14169);
	I14185<= not (G8442 and G3470);
	I14186<= not (G8442 and I14185);
	I14187<= not (G3470 and I14185);
	I14204<= not (G8508 and G3821);
	I14205<= not (G8508 and I14204);
	I14206<= not (G3821 and I14204);
	I14211<= not (G9252 and G9295);
	I14212<= not (G9252 and I14211);
	I14213<= not (G9295 and I14211);
	I14228<= not (G979 and G8055);
	I14229<= not (G979 and I14228);
	I14230<= not (G8055 and I14228);
	I14247<= not (G1322 and G8091);
	I14248<= not (G1322 and I14247);
	I14249<= not (G8091 and I14247);
	I14257<= not (G8154 and G3133);
	I14258<= not (G8154 and I14257);
	I14259<= not (G3133 and I14257);
	I14275<= not (G8218 and G3484);
	I14276<= not (G8218 and I14275);
	I14277<= not (G3484 and I14275);
	I14289<= not (G8282 and G3835);
	I14290<= not (G8282 and I14289);
	I14291<= not (G3835 and I14289);
	I14330<= not (G225 and G9966);
	I14331<= not (G225 and I14330);
	I14332<= not (G9966 and I14330);
	I14350<= not (G8890 and G8848);
	I14351<= not (G8890 and I14350);
	I14352<= not (G8848 and I14350);
	I14368<= not (G8481 and G3303);
	I14369<= not (G8481 and I14368);
	I14370<= not (G3303 and I14368);
	I14398<= not (G8542 and G3654);
	I14399<= not (G8542 and I14398);
	I14400<= not (G3654 and I14398);
	I14427<= not (G8595 and G4005);
	I14428<= not (G8595 and I14427);
	I14429<= not (G4005 and I14427);
	I14480<= not (G10074 and G655);
	I14481<= not (G10074 and I14480);
	I14482<= not (G655 and I14480);
	I14497<= not (G9020 and G8737);
	I14498<= not (G9020 and I14497);
	I14499<= not (G8737 and I14497);
	I14508<= not (G370 and G8721);
	I14509<= not (G370 and I14508);
	I14510<= not (G8721 and I14508);
	I14516<= not (G10147 and G661);
	I14517<= not (G10147 and I14516);
	I14518<= not (G661 and I14516);
	I14530<= not (G8840 and G8873);
	I14531<= not (G8840 and I14530);
	I14532<= not (G8873 and I14530);
	I14609<= not (G8993 and G8678);
	I14610<= not (G8993 and I14609);
	I14611<= not (G8678 and I14609);
	I14712<= not (G9671 and G5128);
	I14713<= not (G9671 and I14712);
	I14714<= not (G5128 and I14712);
	I14733<= not (G9732 and G5475);
	I14734<= not (G9732 and I14733);
	I14735<= not (G5475 and I14733);
	I14764<= not (G9808 and G5821);
	I14765<= not (G9808 and I14764);
	I14766<= not (G5821 and I14764);
	I14788<= not (G9891 and G6167);
	I14789<= not (G9891 and I14788);
	I14790<= not (G6167 and I14788);
	I14816<= not (G9962 and G6513);
	I14817<= not (G9962 and I14816);
	I14818<= not (G6513 and I14816);
	I14853<= not (G9433 and G5142);
	I14854<= not (G9433 and I14853);
	I14855<= not (G5142 and I14853);
	I14883<= not (G9500 and G5489);
	I14884<= not (G9500 and I14883);
	I14885<= not (G5489 and I14883);
	I14923<= not (G9558 and G5835);
	I14924<= not (G9558 and I14923);
	I14925<= not (G5835 and I14923);
	I14955<= not (G9620 and G6181);
	I14956<= not (G9620 and I14955);
	I14957<= not (G6181 and I14955);
	I14991<= not (G9685 and G6527);
	I14992<= not (G9685 and I14991);
	I14993<= not (G6527 and I14991);
	I15002<= not (G9691 and G1700);
	I15003<= not (G9691 and I15002);
	I15004<= not (G1700 and I15002);
	I15041<= not (G9752 and G1834);
	I15042<= not (G9752 and I15041);
	I15043<= not (G1834 and I15041);
	I15051<= not (G9759 and G2259);
	I15052<= not (G9759 and I15051);
	I15053<= not (G2259 and I15051);
	I15078<= not (G9827 and G1968);
	I15079<= not (G9827 and I15078);
	I15080<= not (G1968 and I15078);
	I15087<= not (G9832 and G2393);
	I15088<= not (G9832 and I15087);
	I15089<= not (G2393 and I15087);
	I15105<= not (G9780 and G5313);
	I15106<= not (G9780 and I15105);
	I15107<= not (G5313 and I15105);
	I15121<= not (G9910 and G2102);
	I15122<= not (G9910 and I15121);
	I15123<= not (G2102 and I15121);
	I15128<= not (G9914 and G2527);
	I15129<= not (G9914 and I15128);
	I15130<= not (G2527 and I15128);
	I15147<= not (G9864 and G5659);
	I15148<= not (G9864 and I15147);
	I15149<= not (G5659 and I15147);
	I15166<= not (G9904 and G9823);
	I15167<= not (G9904 and I15166);
	I15168<= not (G9823 and I15166);
	I15174<= not (G9977 and G2661);
	I15175<= not (G9977 and I15174);
	I15176<= not (G2661 and I15174);
	I15193<= not (G9935 and G6005);
	I15194<= not (G9935 and I15193);
	I15195<= not (G6005 and I15193);
	I15212<= not (G10035 and G1714);
	I15213<= not (G10035 and I15212);
	I15214<= not (G1714 and I15212);
	I15241<= not (G10003 and G6351);
	I15242<= not (G10003 and I15241);
	I15243<= not (G6351 and I15241);
	I15253<= not (G10078 and G1848);
	I15254<= not (G10078 and I15253);
	I15255<= not (G1848 and I15253);
	I15262<= not (G10081 and G2273);
	I15263<= not (G10081 and I15262);
	I15264<= not (G2273 and I15262);
	I15287<= not (G10061 and G6697);
	I15288<= not (G10061 and I15287);
	I15289<= not (G6697 and I15287);
	I15298<= not (G10112 and G1982);
	I15299<= not (G10112 and I15298);
	I15300<= not (G1982 and I15298);
	I15306<= not (G10116 and G2407);
	I15307<= not (G10116 and I15306);
	I15308<= not (G2407 and I15306);
	I15333<= not (G10152 and G2116);
	I15334<= not (G10152 and I15333);
	I15335<= not (G2116 and I15333);
	I15340<= not (G10154 and G2541);
	I15341<= not (G10154 and I15340);
	I15342<= not (G2541 and I15340);
	I15363<= not (G10182 and G2675);
	I15364<= not (G10182 and I15363);
	I15365<= not (G2675 and I15363);
	I16778<= not (G11292 and G12332);
	I16779<= not (G11292 and I16778);
	I16780<= not (G12332 and I16778);
	I17379<= not (G13336 and G1129);
	I17380<= not (G13336 and I17379);
	I17381<= not (G1129 and I17379);
	I17404<= not (G13378 and G1472);
	I17405<= not (G13378 and I17404);
	I17406<= not (G1472 and I17404);
	I17446<= not (G13336 and G956);
	I17447<= not (G13336 and I17446);
	I17448<= not (G956 and I17446);
	I17460<= not (G13378 and G1300);
	I17461<= not (G13378 and I17460);
	I17462<= not (G1300 and I17460);
	I17474<= not (G13336 and G1105);
	I17475<= not (G13336 and I17474);
	I17476<= not (G1105 and I17474);
	I17494<= not (G13378 and G1448);
	I17495<= not (G13378 and I17494);
	I17496<= not (G1448 and I17494);
	I17883<= not (G13336 and G1135);
	I17884<= not (G13336 and I17883);
	I17885<= not (G1135 and I17883);
	I17923<= not (G13378 and G1478);
	I17924<= not (G13378 and I17923);
	I17925<= not (G1478 and I17923);
	I18485<= not (G1677 and G14611);
	I18486<= not (G1677 and I18485);
	I18487<= not (G14611 and I18485);
	I18529<= not (G1811 and G14640);
	I18530<= not (G1811 and I18529);
	I18531<= not (G14640 and I18529);
	I18536<= not (G2236 and G14642);
	I18537<= not (G2236 and I18536);
	I18538<= not (G14642 and I18536);
	I18579<= not (G1945 and G14678);
	I18580<= not (G1945 and I18579);
	I18581<= not (G14678 and I18579);
	I18587<= not (G2370 and G14679);
	I18588<= not (G2370 and I18587);
	I18589<= not (G14679 and I18587);
	I18625<= not (G2079 and G14712);
	I18626<= not (G2079 and I18625);
	I18627<= not (G14712 and I18625);
	I18633<= not (G2504 and G14713);
	I18634<= not (G2504 and I18633);
	I18635<= not (G14713 and I18633);
	I18680<= not (G2638 and G14752);
	I18681<= not (G2638 and I18680);
	I18682<= not (G14752 and I18680);
	I20165<= not (G16246 and G990);
	I20166<= not (G16246 and I20165);
	I20167<= not (G990 and I20165);
	I20187<= not (G16272 and G1333);
	I20188<= not (G16272 and I20187);
	I20189<= not (G1333 and I20187);
	I20203<= not (G16246 and G11147);
	I20204<= not (G16246 and I20203);
	I20205<= not (G11147 and I20203);
	I20221<= not (G16272 and G11170);
	I20222<= not (G16272 and I20221);
	I20223<= not (G11170 and I20221);
	I20460<= not (G17515 and G14187);
	I20461<= not (G17515 and I20460);
	I20462<= not (G14187 and I20460);
	I20467<= not (G16663 and G16728);
	I20468<= not (G16663 and I20467);
	I20469<= not (G16728 and I20467);
	I20486<= not (G16696 and G16757);
	I20487<= not (G16696 and I20486);
	I20488<= not (G16757 and I20486);
	I21976<= not (G7680 and G19620);
	I21977<= not (G7680 and I21976);
	I21978<= not (G19620 and I21976);
	I21992<= not (G7670 and G19638);
	I21993<= not (G7670 and I21992);
	I21994<= not (G19638 and I21992);
	I22683<= not (G11893 and G21434);
	I22684<= not (G11893 and I22683);
	I22685<= not (G21434 and I22683);
	I22710<= not (G11915 and G21434);
	I22711<= not (G11915 and I22710);
	I22712<= not (G21434 and I22710);
	I22717<= not (G11916 and G21434);
	I22718<= not (G11916 and I22717);
	I22719<= not (G21434 and I22717);
	I22753<= not (G11937 and G21434);
	I22754<= not (G11937 and I22753);
	I22755<= not (G21434 and I22753);
	I22760<= not (G11939 and G21434);
	I22761<= not (G11939 and I22760);
	I22762<= not (G21434 and I22760);
	I22792<= not (G11956 and G21434);
	I22793<= not (G11956 and I22792);
	I22794<= not (G21434 and I22792);
	I22799<= not (G11960 and G21434);
	I22800<= not (G11960 and I22799);
	I22801<= not (G21434 and I22799);
	I22822<= not (G11978 and G21434);
	I22823<= not (G11978 and I22822);
	I22824<= not (G21434 and I22822);
	I22844<= not (G12113 and G21228);
	I22845<= not (G12113 and I22844);
	I22846<= not (G21228 and I22844);
	I22864<= not (G12146 and G21228);
	I22865<= not (G12146 and I22864);
	I22866<= not (G21228 and I22864);
	I22871<= not (G12150 and G21228);
	I22872<= not (G12150 and I22871);
	I22873<= not (G21228 and I22871);
	I22892<= not (G12189 and G21228);
	I22893<= not (G12189 and I22892);
	I22894<= not (G21228 and I22892);
	I22899<= not (G12193 and G21228);
	I22900<= not (G12193 and I22899);
	I22901<= not (G21228 and I22899);
	I22921<= not (G14677 and G21284);
	I22922<= not (G14677 and I22921);
	I22923<= not (G21284 and I22921);
	I22929<= not (G12223 and G21228);
	I22930<= not (G12223 and I22929);
	I22931<= not (G21228 and I22929);
	I22936<= not (G12226 and G21228);
	I22937<= not (G12226 and I22936);
	I22938<= not (G21228 and I22936);
	I22944<= not (G9492 and G19620);
	I22945<= not (G9492 and I22944);
	I22946<= not (G19620 and I22944);
	I22965<= not (G12288 and G21228);
	I22966<= not (G12288 and I22965);
	I22967<= not (G21228 and I22965);
	I22972<= not (G9657 and G19638);
	I22973<= not (G9657 and I22972);
	I22974<= not (G19638 and I22972);
	I23118<= not (G20076 and G417);
	I23119<= not (G20076 and I23118);
	I23120<= not (G417 and I23118);
	I23585<= not (G22409 and G4332);
	I23586<= not (G22409 and I23585);
	I23587<= not (G4332 and I23585);
	I23600<= not (G22360 and G4322);
	I23601<= not (G22360 and I23600);
	I23602<= not (G4322 and I23600);
	I23917<= not (G23975 and G9333);
	I23918<= not (G23975 and I23917);
	I23919<= not (G9333 and I23917);
	I23949<= not (G23162 and G13603);
	I23950<= not (G23162 and I23949);
	I23951<= not (G13603 and I23949);
	I23961<= not (G23184 and G13631);
	I23962<= not (G23184 and I23961);
	I23963<= not (G13631 and I23961);
	I23969<= not (G22202 and G490);
	I23970<= not (G22202 and I23969);
	I23971<= not (G490 and I23969);
	I23978<= not (G23198 and G13670);
	I23979<= not (G23198 and I23978);
	I23980<= not (G13670 and I23978);
	I23985<= not (G22182 and G482);
	I23986<= not (G22182 and I23985);
	I23987<= not (G482 and I23985);
	I24363<= not (G23687 and G14320);
	I24364<= not (G23687 and I24363);
	I24365<= not (G14320 and I24363);
	I24383<= not (G23721 and G14347);
	I24384<= not (G23721 and I24383);
	I24385<= not (G14347 and I24383);
	I24414<= not (G23751 and G14382);
	I24415<= not (G23751 and I24414);
	I24416<= not (G14382 and I24414);
	I24438<= not (G23771 and G14411);
	I24439<= not (G23771 and I24438);
	I24440<= not (G14411 and I24438);
	I24461<= not (G23796 and G14437);
	I24462<= not (G23796 and I24461);
	I24463<= not (G14437 and I24461);
	I25219<= not (G482 and G24718);
	I25220<= not (G482 and I25219);
	I25221<= not (G24718 and I25219);
	I25242<= not (G490 and G24744);
	I25243<= not (G490 and I25242);
	I25244<= not (G24744 and I25242);
	I25845<= not (G26212 and G24799);
	I25846<= not (G26212 and I25845);
	I25847<= not (G24799 and I25845);
	I25907<= not (G26256 and G24782);
	I25908<= not (G26256 and I25907);
	I25909<= not (G24782 and I25907);
	I26049<= not (G25997 and G13500);
	I26050<= not (G25997 and I26049);
	I26051<= not (G13500 and I26049);
	I26070<= not (G26026 and G13517);
	I26071<= not (G26026 and I26070);
	I26072<= not (G13517 and I26070);
	I26093<= not (G26055 and G13539);
	I26094<= not (G26055 and I26093);
	I26095<= not (G13539 and I26093);
	I26366<= not (G26400 and G14211);
	I26367<= not (G26400 and I26366);
	I26368<= not (G14211 and I26366);
	I26393<= not (G26488 and G14227);
	I26394<= not (G26488 and I26393);
	I26395<= not (G14227 and I26393);
	I26417<= not (G26519 and G14247);
	I26418<= not (G26519 and I26417);
	I26419<= not (G14247 and I26417);
	I26438<= not (G26549 and G14271);
	I26439<= not (G26549 and I26438);
	I26440<= not (G14271 and I26438);
	I26459<= not (G26576 and G14306);
	I26460<= not (G26576 and I26459);
	I26461<= not (G14306 and I26459);
	I29253<= not (G29482 and G12017);
	I29254<= not (G29482 and I29253);
	I29255<= not (G12017 and I29253);
	I29261<= not (G29485 and G12046);
	I29262<= not (G29485 and I29261);
	I29263<= not (G12046 and I29261);
	I29269<= not (G29486 and G12050);
	I29270<= not (G29486 and I29269);
	I29271<= not (G12050 and I29269);
	I29277<= not (G29488 and G12081);
	I29278<= not (G29488 and I29277);
	I29279<= not (G12081 and I29277);
	I29284<= not (G29489 and G12085);
	I29285<= not (G29489 and I29284);
	I29286<= not (G12085 and I29284);
	I29295<= not (G29495 and G12117);
	I29296<= not (G29495 and I29295);
	I29297<= not (G12117 and I29295);
	I29302<= not (G29496 and G12121);
	I29303<= not (G29496 and I29302);
	I29304<= not (G12121 and I29302);
	I29313<= not (G29501 and G12154);
	I29314<= not (G29501 and I29313);
	I29315<= not (G12154 and I29313);
	I31972<= not (G33641 and G33631);
	I31973<= not (G33641 and I31972);
	I31974<= not (G33631 and I31972);
	I31983<= not (G33653 and G33648);
	I31984<= not (G33653 and I31983);
	I31985<= not (G33648 and I31983);
	I32185<= not (G33665 and G33661);
	I32186<= not (G33665 and I32185);
	I32187<= not (G33661 and I32185);
	I32202<= not (G33937 and G33670);
	I32203<= not (G33937 and I32202);
	I32204<= not (G33670 and I32202);
	I32431<= not (G34056 and G34051);
	I32432<= not (G34056 and I32431);
	I32433<= not (G34051 and I32431);
	I32439<= not (G34227 and G34220);
	I32440<= not (G34227 and I32439);
	I32441<= not (G34220 and I32439);
	I32516<= not (G34424 and G34422);
	I32517<= not (G34424 and I32516);
	I32518<= not (G34422 and I32516);
	I32756<= not (G34469 and G25779);
	I32757<= not (G34469 and I32756);
	I32758<= not (G25779 and I32756);
	G7404<=G933 or G939;
	G7450<=G1277 or G1283;
	G7673<=G4153 or G4172;
	G7684<=G4072 or G4176;
	G7764<=G2999 or G2932;
	G7834<=G2886 or G2946;
	G7932<=G4072 or G4153;
	G8417<=G1056 or G1116 or I12583;
	G8461<=G301 or G534;
	G8476<=G1399 or G1459 or I12611;
	G8679<=G222 or G199;
	G8790<=I12782 or I12783;
	G8863<=G1644 or G1664;
	G8904<=G1779 or G1798;
	G8905<=G2204 or G2223;
	G8921<=I12902 or I12903;
	G8956<=G1913 or G1932;
	G8957<=G2338 or G2357;
	G9012<=G2047 or G2066;
	G9013<=G2472 or G2491;
	G9055<=G2606 or G2625;
	G9483<=G1008 or G969;
	G9535<=G209 or G538;
	G9536<=G1351 or G1312;
	G9984<=G4300 or G4242;
	G10589<=G7223 or G7201;
	G10800<=G7517 or G952;
	G10802<=G7533 or G1296;
	G11025<=G2980 or G7831;
	G11370<=G8807 or G550;
	G11372<=G490 or G482 or G8038;
	G11380<=G8583 or G8530;
	G11737<=G8359 or G8292;
	G12768<=G7785 or G7202;
	G12832<=G10347 or G10348;
	G12911<=G10278 or G12768;
	G12925<=G8928 or G10511;
	G12954<=G12186 or G9906;
	G12981<=G12219 or G9967;
	G12982<=G12220 or G9968;
	G13006<=G12284 or G10034;
	G13077<=G11330 or G943;
	G13091<=G329 or G319 or G10796;
	G13095<=G11374 or G1287;
	G13155<=G11496 or G11546;
	G13211<=G11294 or G7567;
	G13242<=G11336 or G7601;
	G13289<=G10619 or G10624;
	G13295<=G10625 or G10655;
	G13296<=G10626 or G10657;
	G13300<=G10656 or G10676;
	G13385<=G11967 or G9479;
	G13526<=G209 or G10685 or G301;
	G13540<=G10822 or G10827;
	G13543<=G10543 or G10565;
	G13570<=G9223 or G11130;
	G13597<=G9247 or G11149;
	G13623<=G482 or G12527;
	G13657<=G7251 or G10616;
	G13660<=G8183 or G12527;
	G13662<=G10896 or G10917;
	G13699<=G10921 or G10947;
	G13728<=G6804 or G12527;
	G13761<=G490 or G12527;
	G13762<=G499 or G12527;
	G13794<=G7396 or G10684;
	G13820<=G11184 or G9187 or G12527;
	G13858<=G209 or G10685;
	G13888<=G2941 or G11691;
	G13914<=G8643 or G11380;
	G13938<=G11213 or G11191;
	G13941<=G11019 or G11023;
	G13969<=G11448 or G8913;
	G13972<=G11232 or G11203;
	G13973<=G11024 or G11028;
	G13997<=G11029 or G11036;
	G14030<=G11037 or G11046;
	G14044<=G10776 or G8703;
	G14062<=G11047 or G11116;
	G14078<=G10776 or G8703;
	G14119<=G10776 or G8703;
	G14182<=G11741 or G11721 or G753;
	G14187<=G8871 or G11771;
	G14309<=G10320 or G11048;
	G14387<=G9086 or G11048;
	G14511<=G10685 or G546;
	G14583<=G10685 or G542;
	G14844<=G10776 or G8703;
	G14888<=G10776 or G8703;
	G14936<=G10776 or G8703;
	G14977<=G10776 or G8703;
	G15017<=G10776 or G8703;
	G15124<=G13605 or G4581;
	G15125<=G10363 or G13605;
	G15582<=G8977 or G12925;
	G15727<=G13383 or G13345 or G13333 or G11010;
	G15732<=G13411 or G13384 or G13349 or G11016;
	G15789<=G10819 or G13211;
	G15792<=G12920 or G10501;
	G15800<=G10821 or G13242;
	G15803<=G12924 or G10528;
	G15910<=G13025 or G10654;
	G15935<=G13029 or G10665;
	G15965<=G13035 or G10675;
	G15968<=G13038 or G10677;
	G16021<=G13047 or G10706;
	G16022<=G13048 or G10707;
	G16052<=G13060 or G10724;
	G16076<=G13081 or G10736;
	G16173<=G8796 or G13464;
	G16187<=G8822 or G13486;
	G16239<=G7892 or G13432;
	G16258<=G13247 or G10856;
	G16261<=G7898 or G13469;
	G16430<=G182 or G13657;
	G16448<=G13287 or G10934;
	G16506<=G13294 or G10966;
	G16800<=G13436 or G11027;
	G16810<=G13461 or G11032;
	G16811<=G8690 or G13914;
	G16839<=G13473 or G11035;
	G16866<=G13492 or G11044;
	G16867<=G13493 or G11045;
	G16876<=G14028 or G11773 or G11755;
	G16882<=G13508 or G11114;
	G16883<=G13509 or G11115;
	G16926<=G14061 or G11804 or G11780;
	G16927<=G13524 or G11126;
	G16928<=G13525 or G11127;
	G16959<=G13542 or G11142;
	G16970<=G13567 or G11163;
	G17264<=G7118 or G14309;
	G17268<=G9220 or G14387;
	G17464<=G14334 or G14313 or G11935 or I18385;
	G17488<=G14361 or G14335 or G11954 or I18417;
	G17490<=G14364 or G14337 or G11958 or I18421;
	G17510<=G14393 or G14362 or G11972 or I18449;
	G17511<=G14396 or G14365 or G11976 or I18452;
	G17569<=G14416 or G14394 or G11995 or I18492;
	G17570<=G14419 or G14397 or G11999 or I18495;
	G17594<=G14450 or G14420 or G12025 or I18543;
	G18879<=G17365 or G14423;
	G18994<=G16303 or G13632;
	G19267<=G17752 or G17768;
	G19274<=G17753 or G14791;
	G19336<=G17769 or G14831;
	G19337<=G17770 or G17785;
	G19344<=G17771 or G14832;
	G19356<=G17784 or G14874;
	G19359<=G17786 or G14875;
	G19363<=G17810 or G14913;
	G19441<=G15507 or G12931;
	G19449<=G15567 or G12939;
	G19467<=G16896 or G14097;
	G19475<=G16930 or G14126;
	G19486<=G15589 or G12979;
	G19488<=G16965 or G14148;
	G19501<=G16986 or G14168;
	G19522<=G17057 or G14180;
	G19525<=G7696 or G16811;
	G19534<=G15650 or G13019;
	G19535<=G15651 or G13020;
	G19555<=G15672 or G13030;
	G19557<=G17123 or G14190;
	G19572<=G17133 or G14193;
	G19575<=G15693 or G13042;
	G19576<=G17138 or G14202;
	G19587<=G15700 or G13046;
	G19593<=G17145 or G14210;
	G19595<=G17149 or G14218;
	G19604<=G15704 or G13059;
	G19605<=G15707 or G13063;
	G19619<=G15712 or G13080;
	G19879<=G15841 or G13265;
	G19904<=G17636 or G14654;
	G19949<=G17671 or G14681;
	G20034<=G15902 or G13299;
	G20051<=G15936 or G13306;
	G20063<=G15978 or G13313;
	G20077<=G16025 or G13320;
	G20082<=G16026 or G13321;
	G20083<=G2902 or G17058;
	G20148<=G16128 or G13393;
	G20160<=G16163 or G13415;
	G20169<=G16184 or G13460;
	G20187<=G16202 or G13491;
	G20196<=G16207 or G13497;
	G20202<=G16211 or G13507;
	G20217<=G16221 or G13523;
	G20241<=G16233 or G13541;
	G20276<=G16243 or G13566;
	G20522<=G691 or G16893;
	G20905<=G7216 or G17264;
	G21891<=G19948 or G15103;
	G21892<=G19788 or G15104;
	G21893<=G20094 or G18655;
	G21894<=G20112 or G15107;
	G21895<=G20135 or G15108;
	G21896<=G20084 or G15110;
	G21897<=G20095 or G15111;
	G21898<=G20152 or G15112;
	G21899<=G20162 or G15113;
	G21900<=G20977 or G15114;
	G21901<=G21251 or G15115;
	G22152<=G21188 or G17469;
	G22217<=G21302 or G17617;
	G22225<=G21332 or G17654;
	G22226<=G21333 or G17655;
	G22304<=G21347 or G17693;
	G22318<=G21394 or G17783;
	G22331<=G21405 or G17809;
	G22447<=G21464 or G12761;
	G22487<=G21512 or G12794;
	G22490<=G21513 or G12795;
	G22516<=G21559 or G12817;
	G22530<=G16751 or G20171;
	G22531<=G20773 or G20922;
	G22547<=G16855 or G20215;
	G22585<=G20915 or G21061;
	G22591<=G18893 or G18909;
	G22625<=G18910 or G18933;
	G22634<=G18934 or G15590;
	G22636<=G18943 or G15611;
	G22639<=G18950 or G15612;
	G22640<=G18951 or G15613;
	G22641<=G18974 or G15631;
	G22644<=G18981 or G15632;
	G22645<=G18982 or G15633;
	G22648<=G18987 or G15652;
	G22652<=G18992 or G15653;
	G22653<=G18993 or G15654;
	G22659<=G19062 or G15673;
	G22662<=G19069 or G15679;
	G22664<=G19139 or G15694;
	G22669<=G7763 or G19525;
	G22679<=G19145 or G15701;
	G22684<=G19206 or G15703;
	G22707<=G20559 or G17156;
	G22708<=G19266 or G15711;
	G22751<=G19333 or G15716;
	G22832<=G19354 or G15722;
	G22872<=G19372 or G19383;
	G22901<=G19384 or G15745;
	G23087<=G19487 or G15852;
	G23129<=G19500 or G15863;
	G23153<=G19521 or G15876;
	G23162<=G20184 or G20170 or I22267;
	G23171<=G19536 or G15903;
	G23183<=G19545 or G15911;
	G23184<=G20198 or G20185 or I22280;
	G23193<=G19556 or G15937;
	G23194<=G19564 or G19578;
	G23197<=G19571 or G15966;
	G23198<=G20214 or G20199 or I22298;
	G23209<=G19585 or G19601;
	G23217<=G19588 or G16023;
	G23251<=G19637 or G16098;
	G23255<=G19655 or G16122;
	G23261<=G19660 or G16125;
	G23262<=G19661 or G16126;
	G23275<=G19680 or G16160;
	G23276<=G19681 or G16161;
	G23296<=G19691 or G16177;
	G23297<=G19692 or G16178;
	G23298<=G19693 or G16179;
	G23317<=G19715 or G16191;
	G23318<=G19716 or G16192;
	G23319<=G19717 or G16193;
	G23345<=G19735 or G16203;
	G23346<=G19736 or G16204;
	G23358<=G19746 or G16212;
	G23374<=G19767 or G13514;
	G23383<=G19756 or G16222;
	G23405<=G19791 or G16245;
	G23574<=G20093 or G20108;
	G23615<=G20109 or G20131;
	G23687<=G21384 or G21363 or I22830;
	G23716<=G9194 or G20905;
	G23720<=G20165 or G16801;
	G23721<=G21401 or G21385 or I22852;
	G23750<=G20174 or G16840;
	G23751<=G21415 or G21402 or I22880;
	G23770<=G20188 or G16868;
	G23771<=G21432 or G21416 or I22912;
	G23795<=G20203 or G16884;
	G23796<=G21462 or G21433 or I22958;
	G23822<=G20218 or G16929;
	G23825<=G20705 or G20781;
	G23989<=G20581 or G17179;
	G23997<=G20602 or G17191;
	G24151<=G18088 or G21661;
	G24200<=G22831 or G18103;
	G24201<=G22848 or G18104;
	G24202<=G22899 or G18106;
	G24203<=G22982 or G18107;
	G24204<=G22990 or G18108;
	G24205<=G23006 or G18109;
	G24206<=G23386 or G18110;
	G24207<=G23396 or G18119;
	G24208<=G23404 or G18121;
	G24209<=G23415 or G18122;
	G24210<=G22900 or G18125;
	G24211<=G23572 or G18138;
	G24212<=G23280 or G18155;
	G24213<=G23220 or G18186;
	G24214<=G23471 or G18195;
	G24215<=G23484 or G18196;
	G24216<=G23416 or G18197;
	G24231<=G22589 or G18201;
	G24232<=G22686 or G18228;
	G24233<=G22590 or G18236;
	G24234<=G22622 or G18237;
	G24235<=G22632 or G18238;
	G24236<=G22489 or G18241;
	G24237<=G22515 or G18242;
	G24238<=G23254 or G18248;
	G24239<=G22752 or G18250;
	G24240<=G22861 or G18251;
	G24241<=G22920 or G18252;
	G24242<=G22834 or G18253;
	G24243<=G22992 or G18254;
	G24244<=G23349 or G18255;
	G24245<=G22849 or G18256;
	G24246<=G23372 or G18257;
	G24247<=G22623 or G18259;
	G24248<=G22710 or G18286;
	G24249<=G22624 or G18294;
	G24250<=G22633 or G18295;
	G24251<=G22637 or G18296;
	G24252<=G22518 or G18299;
	G24253<=G22525 or G18300;
	G24254<=G23265 or G18306;
	G24255<=G22835 or G18308;
	G24256<=G22873 or G18309;
	G24257<=G22938 or G18310;
	G24258<=G22851 or G18311;
	G24259<=G23008 or G18312;
	G24260<=G23373 or G18313;
	G24261<=G22862 or G18314;
	G24262<=G23387 or G18315;
	G24263<=G23497 or G18529;
	G24264<=G22310 or G18559;
	G24265<=G22316 or G18560;
	G24266<=G22329 or G18561;
	G24267<=G23439 or G18611;
	G24268<=G23025 or G18612;
	G24269<=G23131 or G18613;
	G24270<=G23165 or G18614;
	G24271<=G23451 or G18628;
	G24272<=G23056 or G18629;
	G24273<=G23166 or G18630;
	G24274<=G23187 or G18631;
	G24275<=G23474 or G18645;
	G24276<=G23083 or G18646;
	G24277<=G23188 or G18647;
	G24278<=G23201 or G18648;
	G24279<=G23218 or G15105;
	G24280<=G23292 or G15109;
	G24281<=G23397 or G18656;
	G24282<=G23407 or G18657;
	G24334<=G23991 or G18676;
	G24335<=G22165 or G18678;
	G24336<=G24012 or G18753;
	G24337<=G23540 or G18754;
	G24338<=G23658 or G18755;
	G24339<=G23690 or G18756;
	G24340<=G24016 or G18770;
	G24341<=G23564 or G18771;
	G24342<=G23691 or G18772;
	G24343<=G23724 or G18773;
	G24344<=G22145 or G18787;
	G24345<=G23606 or G18788;
	G24346<=G23725 or G18789;
	G24347<=G23754 or G18790;
	G24348<=G22149 or G18804;
	G24349<=G23646 or G18805;
	G24350<=G23755 or G18806;
	G24351<=G23774 or G18807;
	G24352<=G22157 or G18821;
	G24353<=G23682 or G18822;
	G24354<=G23775 or G18823;
	G24355<=G23799 or G18824;
	G24363<=G7831 or G22138;
	G24374<=G19345 or G24004;
	G24390<=G23779 or G21285;
	G24398<=G23801 or G21296;
	G24401<=G23811 or G21298;
	G24430<=G23151 or G8234;
	G24432<=G23900 or G21361;
	G24433<=G10878 or G22400;
	G24443<=G23917 or G21378;
	G24444<=G10890 or G22400;
	G24447<=G10948 or G22450;
	G24457<=G10902 or G22400;
	G24460<=G10967 or G22450;
	G24468<=G10925 or G22400;
	G24471<=G10999 or G22450;
	G24478<=G11003 or G22450;
	G24496<=G24008 or G21557;
	G24500<=G24011 or G21605;
	G24510<=G22488 or G7567;
	G24517<=G22158 or G18906;
	G24518<=G22517 or G7601;
	G24557<=G22308 or G19207;
	G24561<=I23755 or I23756;
	G24565<=G22309 or G19275;
	G24577<=G2856 or G22531;
	G24578<=G2882 or G23825;
	G24580<=G22340 or G13096;
	G24641<=G22151 or G22159;
	G24653<=G2848 or G22585;
	G24705<=G2890 or G23267;
	G24715<=G22189 or G22207;
	G24746<=G22588 or G19461;
	G24782<=G23857 or G23872;
	G24799<=G23901 or G23921;
	G24813<=G22685 or G19594;
	G24821<=G21404 or G23990;
	G24840<=G21419 or G23996;
	G24841<=G21420 or G23998;
	G24842<=G7804 or G22669;
	G24853<=G21452 or G24001;
	G24854<=G21453 or G24002;
	G24879<=G21465 or G24009;
	G24896<=G22863 or G19684;
	G24907<=G21558 or G24015;
	G24919<=G21606 or G22143;
	G24935<=G22937 or G19749;
	G24946<=G22360 or G22409 or G8130;
	G24952<=G21326 or G21340 or I24117;
	G24965<=G22667 or G23825;
	G24968<=G22360 or G22409 or G23389;
	G25010<=G23267 or G2932;
	G25037<=G23103 or G19911;
	G25261<=G23348 or G20193;
	G25539<=G23531 or G20628;
	G25545<=G23551 or G20658;
	G25575<=G24139 or G24140;
	G25576<=G24141 or G24142;
	G25577<=G24143 or G24144;
	G25582<=G21662 or G24152;
	G25583<=G21666 or G24153;
	G25584<=G21670 or G24154;
	G25585<=G21674 or G24155;
	G25586<=G21678 or G24156;
	G25587<=G21682 or G24157;
	G25588<=G21686 or G24158;
	G25589<=G21690 or G24159;
	G25590<=G21694 or G24160;
	G25591<=G24642 or G21705;
	G25592<=G24672 or G21706;
	G25593<=G24716 or G21707;
	G25594<=G24772 or G21708;
	G25595<=G24835 or G21717;
	G25596<=G24865 or G21718;
	G25597<=G24892 or G21719;
	G25598<=G24904 or G21720;
	G25599<=G24914 or G21721;
	G25600<=G24650 or G18111;
	G25601<=G24660 or G18112;
	G25602<=G24673 or G18113;
	G25603<=G24698 or G18114;
	G25604<=G24717 or G18115;
	G25605<=G24743 or G18116;
	G25606<=G24761 or G18117;
	G25607<=G24773 or G18118;
	G25608<=G24643 or G18120;
	G25609<=G24915 or G18126;
	G25610<=G24923 or G18127;
	G25611<=G24931 or G18128;
	G25612<=G24941 or G18132;
	G25613<=G25181 or G18140;
	G25614<=G24797 or G18161;
	G25615<=G24803 or G18162;
	G25616<=G25096 or G18172;
	G25617<=G25466 or G18189;
	G25618<=G25491 or G18192;
	G25619<=G24961 or G18193;
	G25621<=G24523 or G18205;
	G25622<=G24546 or G18217;
	G25623<=G24552 or G18219;
	G25624<=G24408 or G18224;
	G25625<=G24553 or G18226;
	G25626<=G24499 or G18235;
	G25627<=G24503 or G18247;
	G25628<=G24600 or G18249;
	G25629<=G24962 or G18258;
	G25630<=G24532 or G18263;
	G25631<=G24554 or G18275;
	G25632<=G24558 or G18277;
	G25633<=G24420 or G18282;
	G25634<=G24559 or G18284;
	G25635<=G24504 or G18293;
	G25636<=G24507 or G18305;
	G25637<=G24618 or G18307;
	G25638<=G24977 or G18316;
	G25639<=G25122 or G18530;
	G25643<=G24602 or G21736;
	G25644<=G24622 or G21737;
	G25645<=G24679 or G21738;
	G25646<=G24706 or G21739;
	G25647<=G24725 or G21740;
	G25648<=G24644 or G21741;
	G25649<=G24654 or G21742;
	G25650<=G24663 or G21743;
	G25651<=G24680 or G21744;
	G25652<=G24777 or G21747;
	G25653<=G24664 or G18602;
	G25654<=G24634 or G18606;
	G25655<=G24645 or G18607;
	G25656<=G24945 or G18609;
	G25657<=G24624 or G21782;
	G25658<=G24635 or G21783;
	G25659<=G24707 or G21784;
	G25660<=G24726 or G21785;
	G25661<=G24754 or G21786;
	G25662<=G24656 or G21787;
	G25663<=G24666 or G21788;
	G25664<=G24681 or G21789;
	G25665<=G24708 or G21790;
	G25666<=G24788 or G21793;
	G25667<=G24682 or G18619;
	G25668<=G24646 or G18623;
	G25669<=G24657 or G18624;
	G25670<=G24967 or G18626;
	G25671<=G24637 or G21828;
	G25672<=G24647 or G21829;
	G25673<=G24727 or G21830;
	G25674<=G24755 or G21831;
	G25675<=G24769 or G21832;
	G25676<=G24668 or G21833;
	G25677<=G24684 or G21834;
	G25678<=G24709 or G21835;
	G25679<=G24728 or G21836;
	G25680<=G24794 or G21839;
	G25681<=G24710 or G18636;
	G25682<=G24658 or G18640;
	G25683<=G24669 or G18641;
	G25684<=G24983 or G18643;
	G25685<=G24476 or G21866;
	G25686<=G24712 or G21881;
	G25687<=G24729 or G21882;
	G25688<=G24812 or G21887;
	G25689<=G24849 or G21888;
	G25690<=G24864 or G21889;
	G25691<=G24536 or G21890;
	G25693<=G24627 or G18707;
	G25694<=G24638 or G18738;
	G25695<=G24998 or G21914;
	G25696<=G25012 or G21915;
	G25697<=G25086 or G21916;
	G25698<=G25104 or G21917;
	G25699<=G25125 or G21918;
	G25700<=G25040 or G21919;
	G25701<=G25054 or G21920;
	G25702<=G25068 or G21921;
	G25703<=G25087 or G21922;
	G25704<=G25173 or G21925;
	G25705<=G25069 or G18744;
	G25706<=G25030 or G18748;
	G25707<=G25041 or G18749;
	G25708<=G25526 or G18751;
	G25709<=G25014 or G21960;
	G25710<=G25031 or G21961;
	G25711<=G25105 or G21962;
	G25712<=G25126 or G21963;
	G25713<=G25147 or G21964;
	G25714<=G25056 or G21965;
	G25715<=G25071 or G21966;
	G25716<=G25088 or G21967;
	G25717<=G25106 or G21968;
	G25718<=G25187 or G21971;
	G25719<=G25089 or G18761;
	G25720<=G25042 or G18765;
	G25721<=G25057 or G18766;
	G25722<=G25530 or G18768;
	G25723<=G25033 or G22006;
	G25724<=G25043 or G22007;
	G25725<=G25127 or G22008;
	G25726<=G25148 or G22009;
	G25727<=G25163 or G22010;
	G25728<=G25076 or G22011;
	G25729<=G25091 or G22012;
	G25730<=G25107 or G22013;
	G25731<=G25128 or G22014;
	G25732<=G25201 or G22017;
	G25733<=G25108 or G18778;
	G25734<=G25058 or G18782;
	G25735<=G25077 or G18783;
	G25736<=G25536 or G18785;
	G25737<=G25045 or G22052;
	G25738<=G25059 or G22053;
	G25739<=G25149 or G22054;
	G25740<=G25164 or G22055;
	G25741<=G25178 or G22056;
	G25742<=G25093 or G22057;
	G25743<=G25110 or G22058;
	G25744<=G25129 or G22059;
	G25745<=G25150 or G22060;
	G25746<=G25217 or G22063;
	G25747<=G25130 or G18795;
	G25748<=G25078 or G18799;
	G25749<=G25094 or G18800;
	G25750<=G25543 or G18802;
	G25751<=G25061 or G22098;
	G25752<=G25079 or G22099;
	G25753<=G25165 or G22100;
	G25754<=G25179 or G22101;
	G25755<=G25192 or G22102;
	G25756<=G25112 or G22103;
	G25757<=G25132 or G22104;
	G25758<=G25151 or G22105;
	G25759<=G25166 or G22106;
	G25760<=G25238 or G22109;
	G25761<=G25152 or G18812;
	G25762<=G25095 or G18816;
	G25763<=G25113 or G18817;
	G25764<=G25551 or G18819;
	G25767<=G25207 or G12015;
	G25774<=G25223 or G12043;
	G25789<=G25285 or G14543;
	G25791<=G25411 or G25371 or G25328 or G25290;
	G25805<=G25453 or G25414 or G25374 or G25331;
	G25819<=G25323 or G23836;
	G25821<=G25482 or G25456 or G25417 or G25377;
	G25834<=G25366 or G23854;
	G25835<=G25367 or G23855;
	G25836<=G25368 or G23856;
	G25839<=G25507 or G25485 or G25459 or G25420;
	G25856<=G25518 or G25510 or G25488 or G25462;
	G25867<=G25449 or G23884;
	G25868<=G25450 or G23885;
	G25877<=G25502 or G23919;
	G25878<=G25503 or G23920;
	G25885<=G25522 or G23957;
	G25894<=G24817 or G23229;
	G25906<=G25559 or G24014;
	G25910<=G25565 or G22142;
	G25911<=G22514 or G24510;
	G25917<=G22524 or G24518;
	G25929<=G24395 or G22193;
	G25935<=G24402 or G22208;
	G25936<=G24403 or G22209;
	G25937<=G24406 or G22216;
	G25940<=G24415 or G22218;
	G25941<=G24416 or G22219;
	G25942<=G24422 or G22298;
	G25943<=G24423 or G22299;
	G25945<=G24427 or G22307;
	G25960<=G24566 or G24678;
	G26080<=G19393 or G24502;
	G26082<=G2898 or G24561;
	G26089<=G24501 or G22534;
	G26099<=G24506 or G22538;
	G26278<=G24545 or G24549;
	G26293<=G24550 or G24555;
	G26299<=G24551 or G22665;
	G26305<=G24556 or G24564;
	G26327<=G8462 or G24591;
	G26328<=G1183 or G24591;
	G26329<=G8526 or G24609;
	G26334<=G1171 or G24591;
	G26335<=G1526 or G24609;
	G26342<=G8407 or G24591;
	G26343<=G1514 or G24609;
	G26344<=G2927 or G25010;
	G26348<=G8466 or G24609;
	G26349<=G24630 or G13409;
	G26359<=G24651 or G22939;
	G26361<=G24674 or G22991;
	G26363<=G2965 or G24965;
	G26365<=G25504 or G25141;
	G26377<=G24700 or G23007;
	G26386<=G24719 or G23023;
	G26392<=G24745 or G23050;
	G26396<=G24762 or G23062;
	G26422<=G24774 or G23104;
	G26512<=G24786 or G23130;
	G26616<=G24881 or G24855 or G24843 or G24822;
	G26636<=G24897 or G24884 or G24858 or G24846;
	G26657<=G24908 or G24900 or G24887 or G24861;
	G26673<=G24433 or G10674;
	G26690<=G10776 or G24433;
	G26694<=G24444 or G10704;
	G26703<=G24447 or G10705;
	G26721<=G10776 or G24444;
	G26725<=G24457 or G10719;
	G26733<=G10776 or G24447;
	G26737<=G24460 or G10720;
	G26751<=G24903 or G24912;
	G26755<=G10776 or G24457;
	G26759<=G24468 or G7511;
	G26766<=G10776 or G24460;
	G26770<=G24471 or G10732;
	G26781<=G24913 or G24921;
	G26785<=G10776 or G24468;
	G26789<=G10776 or G24471;
	G26793<=G24478 or G7520;
	G26800<=G24922 or G24929;
	G26805<=G10776 or G24478;
	G26809<=G24930 or G24939;
	G26813<=G24940 or G24949;
	G26866<=G20204 or G20242 or G24363;
	G26874<=I25612 or I25613;
	G26875<=G21652 or G25575;
	G26876<=G21655 or G25576;
	G26877<=G21658 or G25577;
	G26878<=G25578 or G25579;
	G26879<=G25580 or G25581;
	G26880<=G26610 or G24186;
	G26881<=G26629 or G24187;
	G26882<=G26650 or G24188;
	G26883<=G26670 or G24189;
	G26884<=G26511 or G24190;
	G26885<=G26541 or G24191;
	G26886<=G26651 or G24192;
	G26887<=G26542 or G24193;
	G26888<=G26671 or G24194;
	G26889<=G26689 or G24195;
	G26890<=G26630 or G24196;
	G26891<=G26652 or G24197;
	G26892<=G26719 or G24198;
	G26893<=G26753 or G24199;
	G26894<=G25979 or G18129;
	G26895<=G26783 or G18148;
	G26896<=G26341 or G18171;
	G26897<=G26611 or G18176;
	G26898<=G26387 or G18194;
	G26899<=G26844 or G18199;
	G26900<=G26819 or G24217;
	G26901<=G26362 or G24218;
	G26902<=G26378 or G24219;
	G26903<=G26388 or G24220;
	G26904<=G26393 or G24221;
	G26905<=G26397 or G24222;
	G26906<=G26423 or G24223;
	G26907<=G26513 or G24224;
	G26908<=G26358 or G24225;
	G26909<=G26543 or G24227;
	G26910<=G26571 or G24228;
	G26911<=G26612 or G24230;
	G26912<=G25946 or G18209;
	G26913<=G25848 or G18225;
	G26914<=G25949 or G18227;
	G26915<=G25900 or G18230;
	G26916<=G25916 or G18232;
	G26917<=G26122 or G18233;
	G26918<=G25931 or G18243;
	G26919<=G25951 or G18267;
	G26920<=G25865 or G18283;
	G26921<=G25955 or G18285;
	G26922<=G25902 or G18288;
	G26923<=G25923 or G18290;
	G26924<=G26153 or G18291;
	G26925<=G25939 or G18301;
	G26926<=G26633 or G18531;
	G26927<=G26711 or G18539;
	G26928<=G26713 or G18541;
	G26929<=G26635 or G18543;
	G26930<=G26799 or G18544;
	G26931<=G26778 or G18547;
	G26932<=G26684 or G18549;
	G26933<=G26808 or G18551;
	G26934<=G26845 or G18556;
	G26938<=G26186 or G21883;
	G26939<=G25907 or G21884;
	G26940<=G25908 or G21886;
	G26944<=G26130 or G18658;
	G26945<=G26379 or G24283;
	G26946<=G26389 or G24284;
	G26947<=G26394 or G24285;
	G26948<=G26399 or G24286;
	G26949<=G26356 or G24287;
	G26950<=G26357 or G24288;
	G26951<=G26390 or G24289;
	G26952<=G26360 or G24290;
	G26953<=G26486 or G24291;
	G26954<=G26380 or G24292;
	G26955<=G26391 or G24293;
	G26956<=G26487 or G24294;
	G26957<=G26517 or G24295;
	G26958<=G26395 or G24297;
	G26959<=G26381 or G24299;
	G26960<=G26258 or G24304;
	G26961<=G26280 or G24306;
	G26962<=G26295 or G24307;
	G26963<=G26306 or G24308;
	G26964<=G26259 or G24316;
	G26965<=G26336 or G24317;
	G26966<=G26345 or G24318;
	G26967<=G26350 or G24319;
	G26968<=G26307 or G24321;
	G26969<=G26313 or G24329;
	G26970<=G26308 or G24332;
	G26971<=G26325 or G24333;
	G26972<=G26780 or G25229;
	G27008<=G26866 or G21370 or I25736;
	G27016<=G26821 or G14585;
	G27019<=G26822 or G14610;
	G27024<=G26826 or G17692;
	G27026<=G26828 or G17726;
	G27031<=G26213 or G26190 or G26166 or G26148;
	G27037<=G26236 or G26218 or G26195 or G26171;
	G27108<=G22522 or G25911;
	G27122<=G22537 or G25917;
	G27126<=G24378 or G25787;
	G27133<=G25788 or G24392;
	G27135<=G24387 or G25803;
	G27147<=G25802 or G24399;
	G27150<=G25804 or G24400;
	G27152<=G24393 or G25817;
	G27159<=G25814 or G12953;
	G27179<=G25816 or G24409;
	G27182<=G25818 or G24410;
	G27205<=G25833 or G24421;
	G27224<=G25870 or G15678;
	G27225<=G2975 or G26364;
	G27226<=G25872 or G24436;
	G27231<=G25873 or G15699;
	G27232<=G25874 or G24450;
	G27233<=G25876 or G24451;
	G27236<=G24620 or G25974;
	G27238<=G25879 or G24464;
	G27239<=G25881 or G24465;
	G27240<=G25883 or G24467;
	G27241<=G24584 or G25984;
	G27243<=G25884 or G24475;
	G27244<=G24652 or G25995;
	G27248<=G24880 or G25953;
	G27250<=G25901 or G15738;
	G27253<=G24661 or G26052;
	G27257<=G25904 or G24498;
	G27258<=G25905 or G15749;
	G27261<=G24544 or G25996;
	G27271<=G24547 or G26053;
	G27274<=G15779 or G25915;
	G27278<=G15786 or G25921;
	G27283<=G25922 or G25924;
	G27289<=G25925 or G25927;
	G27290<=G25926 or G25928;
	G27383<=G24569 or G25961;
	G27394<=G25957 or G24573;
	G27403<=G25962 or G24581;
	G27405<=G24572 or G25968;
	G27426<=G25967 or G24588;
	G27429<=G25969 or G24589;
	G27431<=G24582 or G25977;
	G27450<=G2917 or G26483;
	G27453<=G25976 or G24606;
	G27456<=G25978 or G24607;
	G27458<=G24590 or G25989;
	G27484<=G25988 or G24628;
	G27487<=G25990 or G24629;
	G27489<=G24608 or G26022;
	G27506<=G26021 or G24639;
	G27509<=G26023 or G24640;
	G27515<=G26051 or G13431;
	G27524<=G26050 or G24649;
	G27532<=G16176 or G26084;
	G27533<=G26078 or G24659;
	G27542<=G16190 or G26094;
	G27543<=G26085 or G24670;
	G27544<=G26087 or G24671;
	G27551<=G26091 or G24675;
	G27552<=G26092 or G24676;
	G27555<=G26095 or G24686;
	G27556<=G26097 or G24687;
	G27561<=G26100 or G24702;
	G27562<=G26102 or G24703;
	G27563<=G26104 or G24704;
	G27566<=G26119 or G24713;
	G27567<=G26121 or G24714;
	G27569<=G26124 or G24721;
	G27570<=G26126 or G24722;
	G27571<=G26127 or G24723;
	G27572<=G26129 or G24724;
	G27574<=G26145 or G24730;
	G27575<=G26147 or G24731;
	G27578<=G26155 or G24747;
	G27579<=G26157 or G24748;
	G27580<=G26159 or G24749;
	G27581<=G26161 or G24750;
	G27584<=G26165 or G24758;
	G27589<=G26177 or G24763;
	G27590<=G26179 or G24764;
	G27591<=G26181 or G24765;
	G27596<=G26207 or G24775;
	G27663<=G26323 or G24820;
	G27742<=G17292 or G26673;
	G27779<=G17317 or G26694;
	G27800<=G17321 or G26703;
	G27837<=G17401 or G26725;
	G27858<=G17405 or G26737;
	G27886<=G14438 or G26759;
	G27907<=G17424 or G26770;
	G27937<=G14506 or G26793;
	G27970<=G26514 or G25050;
	G27972<=G26131 or G26105;
	G27974<=G26544 or G25063;
	G27980<=G26105 or G26131;
	G28030<=G24018 or G26874;
	G28041<=G24145 or G26878;
	G28042<=G24148 or G26879;
	G28043<=G27323 or G21714;
	G28044<=G27256 or G18130;
	G28045<=G27378 or G18141;
	G28046<=G27667 or G18157;
	G28047<=G27676 or G18160;
	G28048<=G27362 or G18163;
	G28049<=G27684 or G18164;
	G28050<=G27692 or G18165;
	G28051<=G27699 or G18166;
	G28052<=G27710 or G18167;
	G28053<=G27393 or G18168;
	G28054<=G27723 or G18170;
	G28055<=G27560 or G18190;
	G28056<=G27230 or G18210;
	G28057<=G27033 or G18218;
	G28058<=G27235 or G18268;
	G28059<=G27042 or G18276;
	G28060<=G27616 or G18532;
	G28061<=G27287 or G21735;
	G28062<=G27288 or G21746;
	G28063<=G27541 or G21773;
	G28064<=G27298 or G21781;
	G28065<=G27299 or G21792;
	G28066<=G27553 or G21819;
	G28067<=G27309 or G21827;
	G28068<=G27310 or G21838;
	G28069<=G27564 or G21865;
	G28070<=G27050 or G21867;
	G28071<=G27085 or G21873;
	G28072<=G27086 or G21874;
	G28073<=G27097 or G21875;
	G28074<=G27119 or G21876;
	G28075<=G27083 or G21877;
	G28076<=G27098 or G21878;
	G28077<=G27120 or G21879;
	G28078<=G27140 or G21880;
	G28082<=G27369 or G24315;
	G28083<=G27249 or G18689;
	G28084<=G27254 or G18698;
	G28085<=G27263 or G18700;
	G28086<=G27268 or G18702;
	G28087<=G27255 or G18720;
	G28088<=G27264 or G18729;
	G28089<=G27269 or G18731;
	G28090<=G27275 or G18733;
	G28091<=G27665 or G21913;
	G28092<=G27666 or G21924;
	G28093<=G27981 or G21951;
	G28094<=G27673 or G21959;
	G28095<=G27674 or G21970;
	G28096<=G27988 or G21997;
	G28097<=G27682 or G22005;
	G28098<=G27683 or G22016;
	G28099<=G27992 or G22043;
	G28100<=G27690 or G22051;
	G28101<=G27691 or G22062;
	G28102<=G27995 or G22089;
	G28103<=G27696 or G22097;
	G28104<=G27697 or G22108;
	G28105<=G27997 or G22135;
	G28118<=G27821 or G26815;
	G28132<=G27932 or G27957;
	G28134<=G27958 or G27962;
	G28135<=G27959 or G27963;
	G28138<=G27964 or G27968;
	G28140<=I26643 or I26644;
	G28172<=G27469 or G27440 or G27416 or G27395;
	G28179<=G27494 or G27474 or G27445 or G27421;
	G28180<=G20242 or G27511;
	G28186<=G27209 or G27185 or G27161 or G27146;
	G28188<=G22535 or G27108;
	G28191<=G27217 or G27210 or G27186 or G27162;
	G28194<=G22540 or G27122;
	G28208<=G27025 or G27028;
	G28209<=G27223 or G27141;
	G28211<=G27029 or G27034;
	G28212<=G27030 or G27035;
	G28216<=G27036 or G27043;
	G28220<=G23495 or I26741 or I26742;
	G28230<=G27669 or G14261;
	G28279<=G27087 or G25909;
	G28286<=G27090 or G15757;
	G28295<=G27094 or G15783;
	G28296<=G27095 or G15784;
	G28297<=G27096 or G15785;
	G28305<=G27103 or G15793;
	G28306<=G27104 or G15794;
	G28308<=G27105 or G15795;
	G28309<=G27106 or G15796;
	G28310<=G27107 or G15797;
	G28316<=G27113 or G15804;
	G28317<=G27114 or G15805;
	G28319<=G27115 or G15807;
	G28320<=G27116 or G15808;
	G28322<=G27117 or G15809;
	G28323<=G27118 or G15810;
	G28328<=G27127 or G15812;
	G28329<=G27128 or G15813;
	G28331<=G27129 or G15814;
	G28332<=G27130 or G15815;
	G28334<=G27131 or G15817;
	G28335<=G27132 or G15818;
	G28342<=G27134 or G15819;
	G28344<=G27136 or G15820;
	G28345<=G27137 or G15821;
	G28347<=G27138 or G15822;
	G28348<=G27139 or G15823;
	G28357<=G27148 or G15836;
	G28358<=G27149 or G15837;
	G28359<=G27151 or G15838;
	G28361<=G27153 or G15839;
	G28362<=G27154 or G15840;
	G28368<=G27158 or G27184;
	G28369<=G27160 or G25938;
	G28371<=G27177 or G15847;
	G28372<=G27178 or G15848;
	G28373<=G27180 or G15849;
	G28374<=G27181 or G15850;
	G28375<=G27183 or G15851;
	G28385<=G27201 or G15857;
	G28386<=G27202 or G13277;
	G28387<=G27203 or G15858;
	G28388<=G27204 or G15859;
	G28389<=G27206 or G15860;
	G28390<=G27207 or G15861;
	G28400<=G27211 or G15870;
	G28401<=G27212 or G15871;
	G28402<=G27213 or G15873;
	G28403<=G27214 or G13282;
	G28404<=G27215 or G15874;
	G28405<=G27216 or G15875;
	G28416<=G27218 or G15880;
	G28417<=G27219 or G15881;
	G28418<=G27220 or G15882;
	G28419<=G27221 or G15884;
	G28420<=G27222 or G13290;
	G28428<=G27227 or G15912;
	G28429<=G27228 or G15913;
	G28430<=G27229 or G15914;
	G28435<=G27234 or G15967;
	G28490<=G27262 or G16185;
	G28497<=G27267 or G16199;
	G28511<=G27272 or G16208;
	G28513<=G27276 or G26123;
	G28517<=G27280 or G26154;
	G28518<=G27281 or G26158;
	G28525<=G27284 or G26176;
	G28526<=G27285 or G26178;
	G28527<=G27286 or G26182;
	G28533<=G27291 or G26203;
	G28534<=G27292 or G26204;
	G28536<=G27293 or G26205;
	G28538<=G27294 or G26206;
	G28544<=G27300 or G26229;
	G28545<=G27301 or G26230;
	G28546<=G27302 or G26231;
	G28548<=G27303 or G26232;
	G28549<=G27304 or G26233;
	G28551<=G27305 or G26234;
	G28560<=G27311 or G26249;
	G28561<=G27312 or G26250;
	G28562<=G27313 or G26251;
	G28564<=G27314 or G26252;
	G28565<=G27315 or G26253;
	G28566<=G27316 or G26254;
	G28574<=G27324 or G26270;
	G28576<=G27325 or G26271;
	G28577<=G27326 or G26272;
	G28578<=G27327 or G26273;
	G28580<=G27328 or G26275;
	G28581<=G27329 or G26276;
	G28582<=G27330 or G26277;
	G28589<=G27331 or G26285;
	G28591<=G27332 or G26286;
	G28592<=G27333 or G26288;
	G28594<=G27334 or G26289;
	G28595<=G27335 or G26290;
	G28596<=G27336 or G26291;
	G28600<=G27339 or G16427;
	G28603<=G27340 or G26300;
	G28605<=G27341 or G26302;
	G28607<=G27342 or G26303;
	G28609<=G27346 or G16483;
	G28610<=G27347 or G16484;
	G28611<=G27348 or G16485;
	G28613<=G27350 or G26310;
	G28614<=G27351 or G26311;
	G28618<=G27357 or G16516;
	G28619<=G27358 or G16517;
	G28621<=G27359 or G16518;
	G28622<=G27360 or G16519;
	G28623<=G27361 or G16520;
	G28625<=G27363 or G26324;
	G28628<=G27370 or G16531;
	G28629<=G27371 or G16532;
	G28631<=G27372 or G16534;
	G28632<=G27373 or G16535;
	G28634<=G27374 or G16536;
	G28635<=G27375 or G16537;
	G28636<=G27376 or G16538;
	G28640<=G27384 or G16590;
	G28641<=G27385 or G16591;
	G28643<=G27386 or G16592;
	G28644<=G27387 or G16593;
	G28646<=G27388 or G16595;
	G28647<=G27389 or G16596;
	G28649<=G27390 or G16597;
	G28650<=G27391 or G16598;
	G28651<=G27392 or G16599;
	G28659<=G27404 or G16610;
	G28661<=G27406 or G16611;
	G28662<=G27407 or G16612;
	G28664<=G27408 or G16613;
	G28665<=G27409 or G16614;
	G28667<=G27410 or G16616;
	G28668<=G27411 or G16617;
	G28670<=G27412 or G16618;
	G28671<=G27413 or G16619;
	G28680<=G27427 or G16633;
	G28681<=G27428 or G16634;
	G28682<=G27430 or G16635;
	G28684<=G27432 or G16636;
	G28685<=G27433 or G16637;
	G28687<=G27434 or G16638;
	G28688<=G27435 or G16639;
	G28690<=G27436 or G16641;
	G28691<=G27437 or G16642;
	G28698<=G27451 or G16666;
	G28699<=G27452 or G16667;
	G28700<=G27454 or G16668;
	G28701<=G27455 or G16669;
	G28702<=G27457 or G16670;
	G28704<=G27459 or G16671;
	G28705<=G27460 or G16672;
	G28707<=G27461 or G16673;
	G28708<=G27462 or G16674;
	G28715<=G27480 or G16700;
	G28716<=G27481 or G13887;
	G28717<=G27482 or G16701;
	G28718<=G27483 or G16702;
	G28719<=G27485 or G16703;
	G28720<=G27486 or G16704;
	G28721<=G27488 or G16705;
	G28723<=G27490 or G16706;
	G28724<=G27491 or G16707;
	G28727<=G27500 or G16729;
	G28728<=G27501 or G16730;
	G28729<=G27502 or G16732;
	G28730<=G27503 or G13912;
	G28731<=G27504 or G16733;
	G28732<=G27505 or G16734;
	G28733<=G27507 or G16735;
	G28734<=G27508 or G16736;
	G28735<=G27510 or G16737;
	G28743<=G27517 or G16758;
	G28744<=G27518 or G16759;
	G28745<=G27519 or G16760;
	G28746<=G27520 or G16762;
	G28747<=G27521 or G13942;
	G28748<=G27522 or G16763;
	G28749<=G27523 or G16764;
	G28750<=G27525 or G16765;
	G28751<=G27526 or G16766;
	G28772<=G27534 or G16802;
	G28773<=G27535 or G16803;
	G28774<=G27536 or G16804;
	G28775<=G27537 or G16806;
	G28776<=G27538 or G13974;
	G28777<=G27539 or G16807;
	G28778<=G27540 or G16808;
	G28814<=G27545 or G16841;
	G28815<=G27546 or G16842;
	G28816<=G27547 or G16843;
	G28817<=G27548 or G16845;
	G28818<=G27549 or G13998;
	G28850<=G27557 or G16869;
	G28851<=G27558 or G16870;
	G28852<=G27559 or G16871;
	G28884<=G27568 or G16885;
	G29068<=G27628 or G17119;
	G29078<=G27633 or G26572;
	G29105<=G27645 or G17134;
	G29114<=G27646 or G26602;
	G29143<=G27650 or G17146;
	G29148<=G27651 or G26606;
	G29166<=G27653 or G17153;
	G29168<=G27658 or G26613;
	G29176<=G27661 or G17177;
	G29197<=G27187 or G27163;
	G29222<=G28252 or G18105;
	G29223<=G28341 or G18131;
	G29224<=G28919 or G18156;
	G29225<=G28451 or G18158;
	G29226<=G28455 or G18159;
	G29227<=G28456 or G18169;
	G29228<=G28426 or G18173;
	G29229<=G28532 or G18191;
	G29230<=G28107 or G18202;
	G29231<=G28301 or G18229;
	G29232<=G28183 or G18231;
	G29233<=G28171 or G18234;
	G29234<=G28415 or G18239;
	G29235<=G28110 or G18260;
	G29236<=G28313 or G18287;
	G29237<=G28185 or G18289;
	G29238<=G28178 or G18292;
	G29239<=G28427 or G18297;
	G29240<=G28655 or G18328;
	G29241<=G28638 or G18332;
	G29242<=G28674 or G18354;
	G29243<=G28657 or G18358;
	G29244<=G28692 or G18380;
	G29245<=G28676 or G18384;
	G29246<=G28710 or G18406;
	G29247<=G28694 or G18410;
	G29248<=G28677 or G18434;
	G29249<=G28658 or G18438;
	G29250<=G28695 or G18460;
	G29251<=G28679 or G18464;
	G29252<=G28712 or G18486;
	G29253<=G28697 or G18490;
	G29254<=G28725 or G18512;
	G29255<=G28714 or G18516;
	G29256<=G28597 or G18533;
	G29257<=G28228 or G18600;
	G29258<=G28238 or G18601;
	G29259<=G28304 or G18603;
	G29260<=G28315 or G18604;
	G29261<=G28247 or G18605;
	G29262<=G28327 or G18608;
	G29263<=G28239 or G18617;
	G29264<=G28248 or G18618;
	G29265<=G28318 or G18620;
	G29266<=G28330 or G18621;
	G29267<=G28257 or G18622;
	G29268<=G28343 or G18625;
	G29269<=G28249 or G18634;
	G29270<=G28258 or G18635;
	G29271<=G28333 or G18637;
	G29272<=G28346 or G18638;
	G29273<=G28269 or G18639;
	G29274<=G28360 or G18642;
	G29275<=G28165 or G21868;
	G29276<=G28616 or G18709;
	G29277<=G28440 or G18710;
	G29278<=G28626 or G18740;
	G29279<=G28442 or G18741;
	G29280<=G28530 or G18742;
	G29281<=G28541 or G18743;
	G29282<=G28617 or G18745;
	G29283<=G28627 or G18746;
	G29284<=G28554 or G18747;
	G29285<=G28639 or G18750;
	G29286<=G28542 or G18759;
	G29287<=G28555 or G18760;
	G29288<=G28630 or G18762;
	G29289<=G28642 or G18763;
	G29290<=G28569 or G18764;
	G29291<=G28660 or G18767;
	G29292<=G28556 or G18776;
	G29293<=G28570 or G18777;
	G29294<=G28645 or G18779;
	G29295<=G28663 or G18780;
	G29296<=G28586 or G18781;
	G29297<=G28683 or G18784;
	G29298<=G28571 or G18793;
	G29299<=G28587 or G18794;
	G29300<=G28666 or G18796;
	G29301<=G28686 or G18797;
	G29302<=G28601 or G18798;
	G29303<=G28703 or G18801;
	G29304<=G28588 or G18810;
	G29305<=G28602 or G18811;
	G29306<=G28689 or G18813;
	G29307<=G28706 or G18814;
	G29308<=G28612 or G18815;
	G29309<=G28722 or G18818;
	G29313<=G28284 or G27270;
	G29319<=G28812 or G14453;
	G29325<=G28813 or G27820;
	G29366<=G13738 or G28439;
	G29373<=G13832 or G28453;
	G29476<=G28108 or G28112;
	G29478<=G28111 or G22160;
	G29479<=G28113 or G28116;
	G29480<=G28115 or G22172;
	G29481<=G28117 or G28125;
	G29482<=G28524 or G27588;
	G29483<=G25801 or G28130;
	G29484<=G28124 or G22191;
	G29485<=G28535 or G27594;
	G29486<=G28537 or G27595;
	G29487<=G25815 or G28133;
	G29488<=G28547 or G27600;
	G29489<=G28550 or G27601;
	G29490<=G25832 or G28136;
	G29495<=G28563 or G27614;
	G29496<=G28567 or G27615;
	G29501<=G28583 or G27634;
	G29502<=G28139 or G25871;
	G29504<=G28143 or G25875;
	G29506<=G28148 or G25880;
	G29508<=G28152 or G27041;
	G29520<=G28291 or G28281 or G28264 or G28254;
	G29529<=G28303 or G28293 or G28283 or G28267;
	G29539<=G2864 or G28220;
	G29583<=G28182 or G27099;
	G29643<=G28192 or G27145;
	G29692<=G28197 or G10873;
	G29706<=G28198 or G27208;
	G29716<=G28199 or G15856;
	G29717<=G28200 or G10883;
	G29730<=G28150 or G28141;
	G29734<=G28201 or G15872;
	G29735<=G28202 or G10898;
	G29741<=G28205 or G15883;
	G29748<=G28210 or G28214;
	G29753<=G28213 or G22720;
	G29754<=G28215 or G28218;
	G29756<=G22717 or G28223;
	G29763<=G28217 or G22762;
	G29764<=G28219 or G28226;
	G29768<=G22760 or G28229;
	G29775<=G25966 or G28232;
	G29776<=G28225 or G22846;
	G29777<=G28227 or G28234;
	G29786<=G22843 or G28240;
	G29790<=G25975 or G28242;
	G29791<=G28233 or G22859;
	G29792<=G28235 or G28244;
	G29793<=G28237 or G27247;
	G29801<=G25987 or G28251;
	G29802<=G28243 or G22871;
	G29813<=G26020 or G28261;
	G29848<=G28260 or G26077;
	G29849<=G26049 or G28273;
	G29864<=G28272 or G26086;
	G29879<=G28289 or G26096;
	G29892<=G28300 or G26120;
	G29904<=G28312 or G26146;
	G29914<=G22531 or G22585 or I28147;
	G30081<=G28454 or G11366;
	G30092<=G28466 or G16699;
	G30093<=G28467 or G11397;
	G30103<=G28477 or G16731;
	G30104<=G28478 or G11427;
	G30114<=G28488 or G16761;
	G30115<=G28489 or G11449;
	G30127<=G28494 or G16805;
	G30128<=G28495 or G11497;
	G30141<=G28499 or G16844;
	G30163<=G23381 or G28523;
	G30176<=G23392 or G28531;
	G30189<=G23401 or G28543;
	G30201<=G23412 or G28557;
	G30214<=G23424 or G28572;
	G30270<=G28624 or G27664;
	G30279<=G28637 or G27668;
	G30286<=G28191 or G28186;
	G30287<=G28653 or G27677;
	G30291<=G28672 or G27685;
	G30293<=G28236 or G27246;
	G30298<=G28245 or G27251;
	G30300<=G28246 or G27252;
	G30304<=G28255 or G27259;
	G30307<=G28256 or G27260;
	G30311<=G28265 or G27265;
	G30314<=G28268 or G27266;
	G30317<=G29208 or I28566 or I28567;
	G30333<=G29834 or G21699;
	G30334<=G29837 or G18143;
	G30335<=G29746 or G18174;
	G30336<=G29324 or G18203;
	G30337<=G29334 or G18220;
	G30338<=G29613 or G18240;
	G30339<=G29629 or G18244;
	G30340<=G29377 or G18245;
	G30341<=G29380 or G18246;
	G30342<=G29330 or G18261;
	G30343<=G29344 or G18278;
	G30344<=G29630 or G18298;
	G30345<=G29644 or G18302;
	G30346<=G29381 or G18303;
	G30347<=G29383 or G18304;
	G30348<=G30083 or G18329;
	G30349<=G30051 or G18333;
	G30350<=G30118 or G18334;
	G30351<=G30084 or G18339;
	G30352<=G30094 or G18340;
	G30353<=G30095 or G18355;
	G30354<=G30064 or G18359;
	G30355<=G30131 or G18360;
	G30356<=G30096 or G18365;
	G30357<=G30107 or G18366;
	G30358<=G30108 or G18381;
	G30359<=G30075 or G18385;
	G30360<=G30145 or G18386;
	G30361<=G30109 or G18391;
	G30362<=G30120 or G18392;
	G30363<=G30121 or G18407;
	G30364<=G30086 or G18411;
	G30365<=G30158 or G18412;
	G30366<=G30122 or G18417;
	G30367<=G30133 or G18418;
	G30368<=G30098 or G18435;
	G30369<=G30066 or G18439;
	G30370<=G30135 or G18440;
	G30371<=G30099 or G18445;
	G30372<=G30110 or G18446;
	G30373<=G30111 or G18461;
	G30374<=G30078 or G18465;
	G30375<=G30149 or G18466;
	G30376<=G30112 or G18471;
	G30377<=G30124 or G18472;
	G30378<=G30125 or G18487;
	G30379<=G30089 or G18491;
	G30380<=G30161 or G18492;
	G30381<=G30126 or G18497;
	G30382<=G30137 or G18498;
	G30383<=G30138 or G18513;
	G30384<=G30101 or G18517;
	G30385<=G30172 or G18518;
	G30386<=G30139 or G18523;
	G30387<=G30151 or G18524;
	G30388<=G30023 or G18534;
	G30389<=G29969 or G18554;
	G30390<=G29985 or G18555;
	G30391<=G30080 or G18557;
	G30392<=G30091 or G18558;
	G30393<=G29986 or G21748;
	G30394<=G29805 or G21753;
	G30395<=G29841 or G21754;
	G30396<=G29856 or G21755;
	G30397<=G29747 or G21756;
	G30398<=G29749 or G21757;
	G30399<=G29757 or G21758;
	G30400<=G29766 or G21759;
	G30401<=G29782 or G21760;
	G30402<=G29871 or G21761;
	G30403<=G29750 or G21762;
	G30404<=G29758 or G21763;
	G30405<=G29767 or G21764;
	G30406<=G29783 or G21765;
	G30407<=G29794 or G21766;
	G30408<=G29806 or G21767;
	G30409<=G29842 or G21768;
	G30410<=G29857 or G21769;
	G30411<=G29872 or G21770;
	G30412<=G29885 or G21771;
	G30413<=G30001 or G21772;
	G30414<=G30002 or G21794;
	G30415<=G29843 or G21799;
	G30416<=G29858 or G21800;
	G30417<=G29874 or G21801;
	G30418<=G29751 or G21802;
	G30419<=G29759 or G21803;
	G30420<=G29769 or G21804;
	G30421<=G29784 or G21805;
	G30422<=G29795 or G21806;
	G30423<=G29887 or G21807;
	G30424<=G29760 or G21808;
	G30425<=G29770 or G21809;
	G30426<=G29785 or G21810;
	G30427<=G29796 or G21811;
	G30428<=G29807 or G21812;
	G30429<=G29844 or G21813;
	G30430<=G29859 or G21814;
	G30431<=G29875 or G21815;
	G30432<=G29888 or G21816;
	G30433<=G29899 or G21817;
	G30434<=G30024 or G21818;
	G30435<=G30025 or G21840;
	G30436<=G29860 or G21845;
	G30437<=G29876 or G21846;
	G30438<=G29890 or G21847;
	G30439<=G29761 or G21848;
	G30440<=G29771 or G21849;
	G30441<=G29787 or G21850;
	G30442<=G29797 or G21851;
	G30443<=G29808 or G21852;
	G30444<=G29901 or G21853;
	G30445<=G29772 or G21854;
	G30446<=G29788 or G21855;
	G30447<=G29798 or G21856;
	G30448<=G29809 or G21857;
	G30449<=G29845 or G21858;
	G30450<=G29861 or G21859;
	G30451<=G29877 or G21860;
	G30452<=G29891 or G21861;
	G30453<=G29902 or G21862;
	G30454<=G29909 or G21863;
	G30455<=G30041 or G21864;
	G30456<=G29378 or G21869;
	G30457<=G29369 or G21885;
	G30458<=G30005 or G24330;
	G30459<=G29314 or G21926;
	G30460<=G30207 or G21931;
	G30461<=G30219 or G21932;
	G30462<=G30228 or G21933;
	G30463<=G30140 or G21934;
	G30464<=G30152 or G21935;
	G30465<=G30164 or G21936;
	G30466<=G30174 or G21937;
	G30467<=G30185 or G21938;
	G30468<=G30238 or G21939;
	G30469<=G30153 or G21940;
	G30470<=G30165 or G21941;
	G30471<=G30175 or G21942;
	G30472<=G30186 or G21943;
	G30473<=G30196 or G21944;
	G30474<=G30208 or G21945;
	G30475<=G30220 or G21946;
	G30476<=G30229 or G21947;
	G30477<=G30239 or G21948;
	G30478<=G30248 or G21949;
	G30479<=G29320 or G21950;
	G30480<=G29321 or G21972;
	G30481<=G30221 or G21977;
	G30482<=G30230 or G21978;
	G30483<=G30241 or G21979;
	G30484<=G30154 or G21980;
	G30485<=G30166 or G21981;
	G30486<=G30177 or G21982;
	G30487<=G30187 or G21983;
	G30488<=G30197 or G21984;
	G30489<=G30250 or G21985;
	G30490<=G30167 or G21986;
	G30491<=G30178 or G21987;
	G30492<=G30188 or G21988;
	G30493<=G30198 or G21989;
	G30494<=G30209 or G21990;
	G30495<=G30222 or G21991;
	G30496<=G30231 or G21992;
	G30497<=G30242 or G21993;
	G30498<=G30251 or G21994;
	G30499<=G30261 or G21995;
	G30500<=G29326 or G21996;
	G30501<=G29327 or G22018;
	G30502<=G30232 or G22023;
	G30503<=G30243 or G22024;
	G30504<=G30253 or G22025;
	G30505<=G30168 or G22026;
	G30506<=G30179 or G22027;
	G30507<=G30190 or G22028;
	G30508<=G30199 or G22029;
	G30509<=G30210 or G22030;
	G30510<=G30263 or G22031;
	G30511<=G30180 or G22032;
	G30512<=G30191 or G22033;
	G30513<=G30200 or G22034;
	G30514<=G30211 or G22035;
	G30515<=G30223 or G22036;
	G30516<=G30233 or G22037;
	G30517<=G30244 or G22038;
	G30518<=G30254 or G22039;
	G30519<=G30264 or G22040;
	G30520<=G30272 or G22041;
	G30521<=G29331 or G22042;
	G30522<=G29332 or G22064;
	G30523<=G30245 or G22069;
	G30524<=G30255 or G22070;
	G30525<=G30266 or G22071;
	G30526<=G30181 or G22072;
	G30527<=G30192 or G22073;
	G30528<=G30202 or G22074;
	G30529<=G30212 or G22075;
	G30530<=G30224 or G22076;
	G30531<=G30274 or G22077;
	G30532<=G30193 or G22078;
	G30533<=G30203 or G22079;
	G30534<=G30213 or G22080;
	G30535<=G30225 or G22081;
	G30536<=G30234 or G22082;
	G30537<=G30246 or G22083;
	G30538<=G30256 or G22084;
	G30539<=G30267 or G22085;
	G30540<=G30275 or G22086;
	G30541<=G30281 or G22087;
	G30542<=G29337 or G22088;
	G30543<=G29338 or G22110;
	G30544<=G30257 or G22115;
	G30545<=G30268 or G22116;
	G30546<=G30277 or G22117;
	G30547<=G30194 or G22118;
	G30548<=G30204 or G22119;
	G30549<=G30215 or G22120;
	G30550<=G30226 or G22121;
	G30551<=G30235 or G22122;
	G30552<=G30283 or G22123;
	G30553<=G30205 or G22124;
	G30554<=G30216 or G22125;
	G30555<=G30227 or G22126;
	G30556<=G30236 or G22127;
	G30557<=G30247 or G22128;
	G30558<=G30258 or G22129;
	G30559<=G30269 or G22130;
	G30560<=G30278 or G22131;
	G30561<=G30284 or G22132;
	G30562<=G30289 or G22133;
	G30563<=G29347 or G22134;
	G30579<=G30173 or G14571;
	G30597<=G13564 or G29693;
	G30605<=G29529 or G29520;
	G30608<=G13604 or G29736;
	G30609<=G13633 or G29742;
	G30611<=G13671 or G29743;
	G30672<=G13737 or G29752;
	G30732<=G13778 or G29762;
	G30733<=G13807 or G29773;
	G30734<=G13808 or G29774;
	G30824<=G13833 or G29789;
	G30916<=G13853 or G29799;
	G30984<=G29765 or G29755;
	G31001<=G29360 or G28151;
	G31002<=G29362 or G28154;
	G31007<=G29364 or G28159;
	G31014<=G29367 or G28160;
	G31020<=G29375 or G28164;
	G31144<=G29477 or G28193;
	G31221<=G29494 or G28204;
	G31241<=G25959 or G29510;
	G31244<=G25963 or G29515;
	G31245<=G25964 or G29516;
	G31246<=G25965 or G29518;
	G31247<=G29513 or G13324;
	G31248<=G25970 or G29522;
	G31249<=G25971 or G29523;
	G31250<=G25972 or G29526;
	G31251<=G25973 or G29527;
	G31253<=G25980 or G29533;
	G31254<=G25981 or G29534;
	G31255<=G25982 or G29536;
	G31256<=G25983 or G29537;
	G31257<=G29531 or G28253;
	G31258<=G25991 or G29550;
	G31259<=G25992 or G29554;
	G31260<=G25993 or G29555;
	G31267<=G29548 or G28263;
	G31268<=G29552 or G28266;
	G31269<=G26024 or G29569;
	G31274<=G29565 or G28280;
	G31276<=G29567 or G28282;
	G31277<=G29570 or G28285;
	G31279<=G29571 or G29579;
	G31284<=G29575 or G28290;
	G31287<=G29578 or G28292;
	G31288<=G2955 or G29914;
	G31289<=G29580 or G29591;
	G31291<=G29581 or G29593;
	G31293<=G29582 or G28299;
	G31295<=G26090 or G29598;
	G31302<=G29590 or G28302;
	G31303<=G29592 or G29606;
	G31304<=G29594 or G29608;
	G31306<=G29595 or G29610;
	G31307<=G29596 or G28311;
	G31308<=G26101 or G29614;
	G31311<=G26103 or G29618;
	G31315<=G29607 or G29623;
	G31316<=G29609 or G29624;
	G31317<=G29611 or G29626;
	G31319<=G29612 or G28324;
	G31320<=G26125 or G29632;
	G31322<=G26128 or G29635;
	G31325<=G29625 or G29639;
	G31326<=G29627 or G29640;
	G31375<=G29628 or G28339;
	G31465<=G26156 or G29647;
	G31466<=G26160 or G29650;
	G31468<=G29641 or G29656;
	G31472<=G29642 or G28352;
	G31473<=G26180 or G29666;
	G31474<=G29668 or G13583;
	G31591<=G29358 or G29353;
	G31668<=G29924 or G28558;
	G31670<=G29937 or G28573;
	G31745<=G29959 or G29973;
	G31749<=G29974 or G29988;
	G31751<=G29975 or G29990;
	G31754<=G29989 or G30006;
	G31755<=G29991 or G30008;
	G31757<=G29992 or G30010;
	G31760<=G30007 or G30027;
	G31761<=G30009 or G30028;
	G31762<=G30011 or G30030;
	G31764<=G30015 or G30032;
	G31766<=G30029 or G30042;
	G31767<=G30031 or G30043;
	G31768<=G30033 or G30045;
	G31770<=G30034 or G30047;
	G31772<=G30035 or G28654;
	G31773<=G30044 or G30056;
	G31774<=G30046 or G30057;
	G31775<=G30048 or G30059;
	G31779<=G30050 or G28673;
	G31781<=G30058 or G30069;
	G31782<=G30060 or G30070;
	G31783<=I29351 or I29352;
	G31785<=G30071 or G30082;
	G31793<=G28031 or G30317;
	G31864<=G31271 or G21703;
	G31865<=G31149 or G21709;
	G31866<=G31252 or G18142;
	G31867<=G31238 or G18175;
	G31868<=G30600 or G18204;
	G31869<=G30592 or G18221;
	G31870<=G30607 or G18262;
	G31871<=G30596 or G18279;
	G31872<=G31524 or G18535;
	G31873<=G31270 or G21728;
	G31874<=G31016 or G21729;
	G31875<=G31066 or G21730;
	G31876<=G31125 or G21731;
	G31877<=G31278 or G21732;
	G31878<=G31015 or G21733;
	G31879<=G31475 or G21745;
	G31880<=G31280 or G21774;
	G31881<=G31018 or G21775;
	G31882<=G31115 or G21776;
	G31883<=G31132 or G21777;
	G31884<=G31290 or G21778;
	G31885<=G31017 or G21779;
	G31886<=G31481 or G21791;
	G31887<=G31292 or G21820;
	G31888<=G31067 or G21821;
	G31889<=G31118 or G21822;
	G31890<=G31143 or G21823;
	G31891<=G31305 or G21824;
	G31892<=G31019 or G21825;
	G31893<=G31490 or G21837;
	G31894<=G30671 or G21870;
	G31895<=G31505 or G24296;
	G31896<=G31242 or G24305;
	G31897<=G31237 or G24322;
	G31898<=G31707 or G21906;
	G31899<=G31470 or G21907;
	G31900<=G31484 or G21908;
	G31901<=G31516 or G21909;
	G31902<=G31744 or G21910;
	G31903<=G31374 or G21911;
	G31904<=G31780 or G21923;
	G31905<=G31746 or G21952;
	G31906<=G31477 or G21953;
	G31907<=G31492 or G21954;
	G31908<=G31519 or G21955;
	G31909<=G31750 or G21956;
	G31910<=G31471 or G21957;
	G31911<=G31784 or G21969;
	G31912<=G31752 or G21998;
	G31913<=G31485 or G21999;
	G31914<=G31499 or G22000;
	G31915<=G31520 or G22001;
	G31916<=G31756 or G22002;
	G31917<=G31478 or G22003;
	G31918<=G31786 or G22015;
	G31919<=G31758 or G22044;
	G31920<=G31493 or G22045;
	G31921<=G31508 or G22046;
	G31922<=G31525 or G22047;
	G31923<=G31763 or G22048;
	G31924<=G31486 or G22049;
	G31925<=G31789 or G22061;
	G31926<=G31765 or G22090;
	G31927<=G31500 or G22091;
	G31928<=G31517 or G22092;
	G31929<=G31540 or G22093;
	G31930<=G31769 or G22094;
	G31931<=G31494 or G22095;
	G31932<=G31792 or G22107;
	G31964<=G31654 or G14544;
	G32037<=G30566 or G29329;
	G32094<=G30612 or G29363;
	G32117<=G24482 or G30914;
	G32123<=G30915 or G30919;
	G32124<=G24488 or G30920;
	G32125<=G30918 or G29376;
	G32130<=G30921 or G30925;
	G32131<=G24495 or G30926;
	G32132<=G31487 or G31479;
	G32144<=G30927 or G30930;
	G32155<=G30935 or G29475;
	G32202<=G31069 or G13410;
	G32208<=G31120 or G29584;
	G32209<=G31122 or G29599;
	G32210<=G31123 or G29600;
	G32211<=G31124 or G29603;
	G32216<=G31128 or G29615;
	G32217<=G31129 or G29616;
	G32218<=G31130 or G29619;
	G32219<=G31131 or G29620;
	G32220<=G31139 or G29633;
	G32221<=G31140 or G29634;
	G32222<=G31141 or G29636;
	G32223<=G31142 or G29637;
	G32225<=G30576 or G29336;
	G32226<=G31145 or G29645;
	G32227<=G31146 or G29648;
	G32228<=G31147 or G29651;
	G32229<=G31148 or G29652;
	G32230<=G30589 or G29345;
	G32231<=G30590 or G29346;
	G32233<=G31150 or G29661;
	G32235<=G31151 or G29662;
	G32236<=G31152 or G29664;
	G32237<=G31153 or G29667;
	G32238<=G30594 or G29349;
	G32239<=G30595 or G29350;
	G32240<=G24757 or G31182;
	G32243<=G31166 or G29683;
	G32245<=G31167 or G29684;
	G32247<=G31168 or G29686;
	G32249<=G31169 or G29687;
	G32250<=G30598 or G29351;
	G32251<=G30599 or G29352;
	G32252<=G31183 or G31206;
	G32253<=G24771 or G31207;
	G32257<=G31184 or G29708;
	G32259<=G31185 or G29709;
	G32262<=G31186 or G29710;
	G32264<=G31187 or G29711;
	G32266<=G30604 or G29354;
	G32267<=G31208 or G31218;
	G32268<=G24785 or G31219;
	G32271<=G31209 or G29731;
	G32275<=G31210 or G29732;
	G32277<=G31211 or G29733;
	G32279<=G31220 or G31224;
	G32280<=G24790 or G31225;
	G32285<=G31222 or G29740;
	G32288<=G31226 or G31229;
	G32289<=G24796 or G31230;
	G32294<=G31231 or G31232;
	G32344<=G29804 or G31266;
	G32346<=G29838 or G31272;
	G32347<=G29839 or G31273;
	G32349<=G29840 or G31275;
	G32351<=G29851 or G31281;
	G32352<=G29852 or G31282;
	G32353<=G29853 or G31283;
	G32354<=G29854 or G31285;
	G32355<=G29855 or G31286;
	G32357<=G29865 or G31296;
	G32358<=G29866 or G31297;
	G32359<=G29867 or G31298;
	G32360<=G29868 or G31299;
	G32361<=G29869 or G31300;
	G32362<=G29870 or G31301;
	G32367<=G29880 or G31309;
	G32368<=G29881 or G31310;
	G32370<=G29882 or G31312;
	G32371<=G29883 or G31313;
	G32372<=G29884 or G31314;
	G32373<=G29894 or G31321;
	G32374<=G29895 or G31323;
	G32375<=G29896 or G31324;
	G32380<=G29907 or G31467;
	G32385<=G31480 or G29938;
	G32386<=G31488 or G29949;
	G32387<=G31489 or G29952;
	G32388<=G31495 or G29962;
	G32389<=G31496 or G29966;
	G32390<=G31501 or G29979;
	G32391<=G31502 or G29982;
	G32392<=G31513 or G30000;
	G32395<=G31523 or G30049;
	G32398<=G31526 or G30061;
	G32399<=G31527 or G30062;
	G32408<=G31541 or G30073;
	G32426<=G26105 or G26131 or G30613;
	G32427<=G8928 or G30583;
	G32429<=G30318 or G31794;
	G32454<=G30322 or G31795;
	G32976<=G32207 or G21704;
	G32977<=G32169 or G21710;
	G32978<=G32197 or G18145;
	G32979<=G32181 or G18177;
	G32980<=G32254 or G18198;
	G32981<=G32425 or G18206;
	G32982<=G31948 or G18208;
	G32983<=G31990 or G18222;
	G32984<=G31934 or G18264;
	G32985<=G31963 or G18266;
	G32986<=G31996 or G18280;
	G32987<=G32311 or G18323;
	G32988<=G32232 or G18325;
	G32989<=G32241 or G18326;
	G32990<=G32281 or G18341;
	G32991<=G32322 or G18349;
	G32992<=G32242 or G18351;
	G32993<=G32255 or G18352;
	G32994<=G32290 or G18367;
	G32995<=G32330 or G18375;
	G32996<=G32256 or G18377;
	G32997<=G32269 or G18378;
	G32998<=G32300 or G18393;
	G32999<=G32337 or G18401;
	G33000<=G32270 or G18403;
	G33001<=G32282 or G18404;
	G33002<=G32304 or G18419;
	G33003<=G32323 or G18429;
	G33004<=G32246 or G18431;
	G33005<=G32260 or G18432;
	G33006<=G32291 or G18447;
	G33007<=G32331 or G18455;
	G33008<=G32261 or G18457;
	G33009<=G32273 or G18458;
	G33010<=G32301 or G18473;
	G33011<=G32338 or G18481;
	G33012<=G32274 or G18483;
	G33013<=G32283 or G18484;
	G33014<=G32305 or G18499;
	G33015<=G32343 or G18507;
	G33016<=G32284 or G18509;
	G33017<=G32292 or G18510;
	G33018<=G32312 or G18525;
	G33019<=G32339 or G18536;
	G33020<=G32160 or G21734;
	G33021<=G32302 or G21749;
	G33022<=G32306 or G21750;
	G33023<=G32313 or G21751;
	G33024<=G32324 or G21752;
	G33025<=G32162 or G21780;
	G33026<=G32307 or G21795;
	G33027<=G32314 or G21796;
	G33028<=G32325 or G21797;
	G33029<=G32332 or G21798;
	G33030<=G32166 or G21826;
	G33031<=G32315 or G21841;
	G33032<=G32326 or G21842;
	G33033<=G32333 or G21843;
	G33034<=G32340 or G21844;
	G33035<=G32019 or G21872;
	G33036<=G32168 or G24309;
	G33037<=G32177 or G24310;
	G33038<=G32184 or G24311;
	G33039<=G32187 or G24312;
	G33040<=G32164 or G24313;
	G33041<=G32189 or G24323;
	G33042<=G32193 or G24324;
	G33043<=G32195 or G24325;
	G33044<=G32199 or G24327;
	G33045<=G32206 or G24328;
	G33046<=G32308 or G21912;
	G33047<=G31944 or G21927;
	G33048<=G31960 or G21928;
	G33049<=G31966 or G21929;
	G33050<=G31974 or G21930;
	G33051<=G32316 or G21958;
	G33052<=G31961 or G21973;
	G33053<=G31967 or G21974;
	G33054<=G31975 or G21975;
	G33055<=G31986 or G21976;
	G33056<=G32327 or G22004;
	G33057<=G31968 or G22019;
	G33058<=G31976 or G22020;
	G33059<=G31987 or G22021;
	G33060<=G31992 or G22022;
	G33061<=G32334 or G22050;
	G33062<=G31977 or G22065;
	G33063<=G31988 or G22066;
	G33064<=G31993 or G22067;
	G33065<=G32008 or G22068;
	G33066<=G32341 or G22096;
	G33067<=G31989 or G22111;
	G33068<=G31994 or G22112;
	G33069<=G32009 or G22113;
	G33070<=G32010 or G22114;
	G33076<=G32336 or G32446;
	G33115<=G32397 or G32401;
	G33116<=G32403 or G32411;
	G33118<=G32413 or G32418;
	G33119<=G32420 or G32428;
	G33123<=G31962 or G30577;
	G33149<=G32204 or I30717 or I30718;
	G33159<=G32016 or G30730;
	G33164<=G32203 or I30727 or I30728;
	G33176<=G32198 or I30734 or I30735;
	G33187<=G32014 or I30740 or I30741;
	G33197<=G32342 or I30745 or I30746;
	G33204<=G32317 or I30750 or I30751;
	G33212<=G32328 or I30755 or I30756;
	G33219<=G32335 or I30760 or I30761;
	G33227<=G32029 or G32031;
	G33231<=G32032 or G32036;
	G33232<=G32034 or G30936;
	G33234<=G32039 or G32043;
	G33235<=G32040 or G30982;
	G33236<=G32044 or G32045;
	G33238<=G32048 or G32051;
	G33240<=G32052 or G32068;
	G33251<=G32096 or G29509;
	G33253<=G32103 or G29511;
	G33254<=G32104 or G29512;
	G33255<=G32106 or G29514;
	G33256<=G32107 or G29517;
	G33257<=G32108 or G29519;
	G33259<=G32109 or G29521;
	G33260<=G32110 or G29524;
	G33261<=G32111 or G29525;
	G33262<=G32112 or G29528;
	G33265<=G32113 or G29530;
	G33266<=G32114 or G29532;
	G33267<=G32115 or G29535;
	G33268<=G32116 or G29538;
	G33270<=G32119 or G29547;
	G33271<=G32120 or G29549;
	G33272<=G32121 or G29551;
	G33273<=G32122 or G29553;
	G33274<=G32126 or G29563;
	G33275<=G32127 or G29564;
	G33276<=G32128 or G29566;
	G33277<=G32129 or G29568;
	G33278<=G32139 or G29572;
	G33279<=G32140 or G29573;
	G33280<=G32141 or G29574;
	G33281<=G32142 or G29576;
	G33282<=G32143 or G29577;
	G33283<=G31995 or G30318;
	G33286<=G32145 or G29585;
	G33287<=G32146 or G29586;
	G33288<=G32147 or G29587;
	G33289<=G32148 or G29588;
	G33290<=G32149 or G29589;
	G33291<=G32154 or G13477;
	G33292<=G32150 or G29601;
	G33293<=G32151 or G29602;
	G33294<=G32152 or G29604;
	G33295<=G32153 or G29605;
	G33296<=G32156 or G29617;
	G33297<=G32157 or G29621;
	G33298<=G32158 or G29622;
	G33303<=G32159 or G29638;
	G33310<=G29631 or G32165;
	G33312<=G29646 or G32170;
	G33313<=G29649 or G32171;
	G33314<=G29663 or G32174;
	G33315<=G29665 or G32175;
	G33316<=G29685 or G32178;
	G33317<=G29688 or G32179;
	G33318<=G31969 or G32434;
	G33321<=G29712 or G32182;
	G33323<=G31936 or G32442;
	G33380<=G32234 or G29926;
	G33383<=G32244 or G29940;
	G33384<=G32248 or G29943;
	G33386<=G32258 or G29951;
	G33387<=G32263 or G29954;
	G33389<=G32272 or G29964;
	G33390<=G32276 or G29968;
	G33393<=G32286 or G29984;
	G33534<=G33186 or G21700;
	G33535<=G33233 or G21711;
	G33536<=G33241 or G21715;
	G33537<=G33244 or G21716;
	G33538<=G33252 or G18144;
	G33539<=G33245 or G18178;
	G33540<=G33099 or G18207;
	G33541<=G33101 or G18223;
	G33542<=G33102 or G18265;
	G33543<=G33106 or G18281;
	G33544<=G33392 or G18317;
	G33545<=G33399 or G18324;
	G33546<=G33402 or G18327;
	G33547<=G33349 or G18331;
	G33548<=G33327 or G18336;
	G33549<=G33328 or G18337;
	G33550<=G33342 or G18338;
	G33551<=G33446 or G18342;
	G33552<=G33400 or G18343;
	G33553<=G33403 or G18350;
	G33554<=G33407 or G18353;
	G33555<=G33355 or G18357;
	G33556<=G33329 or G18362;
	G33557<=G33331 or G18363;
	G33558<=G33350 or G18364;
	G33559<=G33073 or G18368;
	G33560<=G33404 or G18369;
	G33561<=G33408 or G18376;
	G33562<=G33414 or G18379;
	G33563<=G33361 or G18383;
	G33564<=G33332 or G18388;
	G33565<=G33338 or G18389;
	G33566<=G33356 or G18390;
	G33567<=G33081 or G18394;
	G33568<=G33409 or G18395;
	G33569<=G33415 or G18402;
	G33570<=G33420 or G18405;
	G33571<=G33367 or G18409;
	G33572<=G33339 or G18414;
	G33573<=G33343 or G18415;
	G33574<=G33362 or G18416;
	G33575<=G33086 or G18420;
	G33576<=G33401 or G18423;
	G33577<=G33405 or G18430;
	G33578<=G33410 or G18433;
	G33579<=G33357 or G18437;
	G33580<=G33330 or G18442;
	G33581<=G33333 or G18443;
	G33582<=G33351 or G18444;
	G33583<=G33074 or G18448;
	G33584<=G33406 or G18449;
	G33585<=G33411 or G18456;
	G33586<=G33416 or G18459;
	G33587<=G33363 or G18463;
	G33588<=G33334 or G18468;
	G33589<=G33340 or G18469;
	G33590<=G33358 or G18470;
	G33591<=G33082 or G18474;
	G33592<=G33412 or G18475;
	G33593<=G33417 or G18482;
	G33594<=G33421 or G18485;
	G33595<=G33368 or G18489;
	G33596<=G33341 or G18494;
	G33597<=G33344 or G18495;
	G33598<=G33364 or G18496;
	G33599<=G33087 or G18500;
	G33600<=G33418 or G18501;
	G33601<=G33422 or G18508;
	G33602<=G33425 or G18511;
	G33603<=G33372 or G18515;
	G33604<=G33345 or G18520;
	G33605<=G33352 or G18521;
	G33606<=G33369 or G18522;
	G33607<=G33091 or G18526;
	G33608<=G33322 or G18537;
	G33609<=G33239 or G18615;
	G33610<=G33242 or G18616;
	G33611<=G33243 or G18632;
	G33612<=G33247 or G18633;
	G33613<=G33248 or G18649;
	G33614<=G33249 or G18650;
	G33615<=G33113 or G21871;
	G33616<=G33237 or G24314;
	G33617<=G33263 or G24326;
	G33618<=G33353 or G18757;
	G33619<=G33359 or G18758;
	G33620<=G33360 or G18774;
	G33621<=G33365 or G18775;
	G33622<=G33366 or G18791;
	G33623<=G33370 or G18792;
	G33624<=G33371 or G18808;
	G33625<=G33373 or G18809;
	G33626<=G33374 or G18825;
	G33627<=G33376 or G18826;
	G33628<=G33071 or G32450;
	G33685<=G32396 or G33423;
	G33692<=G32400 or G33428;
	G33694<=G32402 or G33429;
	G33699<=G32409 or G33433;
	G33703<=G32410 or G33434;
	G33706<=G32412 or G33440;
	G33709<=G32414 or G33441;
	G33714<=G32419 or G33450;
	G33732<=G33104 or G32011;
	G33733<=G33105 or G32012;
	G33788<=G33122 or G32041;
	G33791<=G33379 or G32430;
	G33794<=G33126 or G32053;
	G33891<=G33264 or G33269;
	G33914<=G33305 or G33311;
	G33945<=G32430 or G33455;
	G33946<=G32434 or G33456;
	G33947<=G32438 or G33457;
	G33948<=G32442 or G33458;
	G33949<=G32446 or G33459;
	G33950<=G32450 or G33460;
	G33951<=G33469 or I31838 or I31839;
	G33952<=G33478 or I31843 or I31844;
	G33953<=G33487 or I31848 or I31849;
	G33954<=G33496 or I31853 or I31854;
	G33955<=G33505 or I31858 or I31859;
	G33956<=G33514 or I31863 or I31864;
	G33957<=G33523 or I31868 or I31869;
	G33958<=G33532 or I31873 or I31874;
	G33960<=G33759 or G21701;
	G33961<=G33789 or G21712;
	G33962<=G33822 or G18123;
	G33963<=G33830 or G18124;
	G33964<=G33817 or G18146;
	G33965<=G33805 or G18179;
	G33966<=G33837 or G18318;
	G33967<=G33842 or G18319;
	G33968<=G33855 or G18320;
	G33969<=G33864 or G18321;
	G33970<=G33868 or G18322;
	G33971<=G33890 or G18330;
	G33972<=G33941 or G18335;
	G33973<=G33840 or G18344;
	G33974<=G33846 or G18345;
	G33975<=G33860 or G18346;
	G33976<=G33869 or G18347;
	G33977<=G33876 or G18348;
	G33978<=G33892 or G18356;
	G33979<=G33942 or G18361;
	G33980<=G33843 or G18370;
	G33981<=G33856 or G18371;
	G33982<=G33865 or G18372;
	G33983<=G33877 or G18373;
	G33984<=G33881 or G18374;
	G33985<=G33896 or G18382;
	G33986<=G33639 or G18387;
	G33987<=G33847 or G18396;
	G33988<=G33861 or G18397;
	G33989<=G33870 or G18398;
	G33990<=G33882 or G18399;
	G33991<=G33885 or G18400;
	G33992<=G33900 or G18408;
	G33993<=G33646 or G18413;
	G33994<=G33841 or G18424;
	G33995<=G33848 or G18425;
	G33996<=G33862 or G18426;
	G33997<=G33871 or G18427;
	G33998<=G33878 or G18428;
	G33999<=G33893 or G18436;
	G34000<=G33943 or G18441;
	G34001<=G33844 or G18450;
	G34002<=G33857 or G18451;
	G34003<=G33866 or G18452;
	G34004<=G33879 or G18453;
	G34005<=G33883 or G18454;
	G34006<=G33897 or G18462;
	G34007<=G33640 or G18467;
	G34008<=G33849 or G18476;
	G34009<=G33863 or G18477;
	G34010<=G33872 or G18478;
	G34011<=G33884 or G18479;
	G34012<=G33886 or G18480;
	G34013<=G33901 or G18488;
	G34014<=G33647 or G18493;
	G34015<=G33858 or G18502;
	G34016<=G33867 or G18503;
	G34017<=G33880 or G18504;
	G34018<=G33887 or G18505;
	G34019<=G33889 or G18506;
	G34020<=G33904 or G18514;
	G34021<=G33652 or G18519;
	G34022<=G33873 or G18538;
	G34023<=G33796 or G24320;
	G34024<=G33807 or G24331;
	G34025<=G33927 or G18672;
	G34026<=G33715 or G18682;
	G34027<=G33718 or G18683;
	G34028<=G33720 or G18684;
	G34029<=G33798 or G18703;
	G34030<=G33727 or G18704;
	G34031<=G33735 or G18705;
	G34032<=G33816 or G18706;
	G34033<=G33821 or G18708;
	G34034<=G33719 or G18713;
	G34035<=G33721 or G18714;
	G34036<=G33722 or G18715;
	G34037<=G33803 or G18734;
	G34038<=G33731 or G18735;
	G34039<=G33743 or G18736;
	G34040<=G33818 or G18737;
	G34041<=G33829 or G18739;
	G34043<=G33903 or G33905;
	G34046<=G33906 or G33908;
	G34055<=G33909 or G33910;
	G34057<=G33911 or G33915;
	G34064<=G33919 or G33922;
	G34090<=G33676 or G33680;
	G34095<=G33681 or G33687;
	G34099<=G33684 or G33689;
	G34100<=G33690 or G33697;
	G34101<=G33693 or G33700;
	G34103<=G33701 or G33707;
	G34107<=G33710 or G33121;
	G34125<=G33724 or G33124;
	G34127<=G33657 or G32438;
	G34148<=G33758 or G19656;
	G34149<=G33760 or G19674;
	G34153<=G33899 or G33451;
	G34158<=G33784 or G19740;
	G34166<=G33785 or G19752;
	G34167<=G33786 or G19768;
	G34168<=G33787 or G19784;
	G34170<=G33790 or G19855;
	G34172<=G33795 or G19914;
	G34189<=G33801 or G33808;
	G34190<=G33802 or G33810;
	G34193<=G33809 or G33814;
	G34194<=G33811 or G33815;
	G34199<=G33820 or G33828;
	G34204<=G33832 or G33833;
	G34206<=G33834 or G33836;
	G34207<=G33835 or G33304;
	G34231<=G33898 or G33902;
	G34232<=G33451 or G33944;
	G34233<=G32455 or G33951;
	G34234<=G32520 or G33952;
	G34235<=G32585 or G33953;
	G34236<=G32650 or G33954;
	G34237<=G32715 or G33955;
	G34238<=G32780 or G33956;
	G34239<=G32845 or G33957;
	G34240<=G32910 or G33958;
	G34249<=G34110 or G21702;
	G34250<=G34111 or G21713;
	G34251<=G34157 or G18147;
	G34252<=G34146 or G18180;
	G34253<=G34171 or G24300;
	G34254<=G34116 or G24301;
	G34255<=G34120 or G24302;
	G34256<=G34173 or G24303;
	G34257<=G34226 or G18674;
	G34258<=G34211 or G18675;
	G34259<=G34066 or G18679;
	G34260<=G34113 or G18680;
	G34261<=G34074 or G18688;
	G34262<=G34075 or G18697;
	G34263<=G34078 or G18699;
	G34264<=G34081 or G18701;
	G34265<=G34117 or G18711;
	G34266<=G34076 or G18719;
	G34267<=G34079 or G18728;
	G34268<=G34082 or G18730;
	G34269<=G34083 or G18732;
	G34273<=G27765 or G34203;
	G34274<=G27822 or G34205;
	G34278<=G26829 or G34212;
	G34280<=G26833 or G34213;
	G34282<=G26838 or G34214;
	G34283<=G26839 or G34215;
	G34286<=G26842 or G34216;
	G34288<=G26846 or G34217;
	G34289<=G26847 or G34218;
	G34290<=G26848 or G34219;
	G34292<=G26853 or G34223;
	G34293<=G26854 or G34224;
	G34294<=G26855 or G34225;
	G34297<=G26858 or G34228;
	G34300<=G26864 or G34230;
	G34303<=G25768 or G34045;
	G34305<=G25775 or G34050;
	G34306<=G25782 or G34054;
	G34314<=G25831 or G34061;
	G34318<=G25850 or G34063;
	G34321<=G25866 or G34065;
	G34330<=G34069 or G33717;
	G34331<=G27121 or G34072;
	G34332<=G34071 or G33723;
	G34347<=G25986 or G34102;
	G34349<=G26019 or G34104;
	G34350<=G26048 or G34106;
	G34352<=G26079 or G34109;
	G34353<=G26088 or G34114;
	G34366<=G26257 or G34133;
	G34368<=G26274 or G34135;
	G34369<=G26279 or G34136;
	G34372<=G26287 or G34137;
	G34373<=G26292 or G34138;
	G34374<=G26294 or G34139;
	G34376<=G26301 or G34140;
	G34377<=G26304 or G34141;
	G34379<=G26312 or G34143;
	G34399<=G34178 or G25067;
	G34402<=G34179 or G25084;
	G34403<=G34180 or G25085;
	G34404<=G34182 or G25102;
	G34405<=G34183 or G25103;
	G34406<=G34184 or G25123;
	G34407<=G34185 or G25124;
	G34411<=G34186 or G25142;
	G34412<=G34187 or G25143;
	G34416<=G34191 or G25159;
	G34417<=G27678 or G34196;
	G34421<=G27686 or G34198;
	G34438<=G34348 or G18150;
	G34439<=G34344 or G18181;
	G34440<=G34364 or G24226;
	G34441<=G34381 or G18540;
	G34442<=G34380 or G18542;
	G34443<=G34385 or G18545;
	G34444<=G34389 or G18546;
	G34445<=G34382 or G18548;
	G34446<=G34390 or G18550;
	G34447<=G34363 or G18552;
	G34448<=G34365 or G18553;
	G34449<=G34279 or G18662;
	G34450<=G34281 or G18663;
	G34451<=G34393 or G18664;
	G34452<=G34401 or G18665;
	G34453<=G34410 or G18666;
	G34454<=G34414 or G18667;
	G34455<=G34284 or G18668;
	G34456<=G34395 or G18669;
	G34457<=G34394 or G18670;
	G34458<=G34396 or G18671;
	G34459<=G34415 or G18673;
	G34460<=G34301 or G18677;
	G34461<=G34291 or G18681;
	G34462<=G34334 or G18685;
	G34463<=G34338 or G18686;
	G34464<=G34340 or G18687;
	G34465<=G34295 or G18712;
	G34466<=G34337 or G18716;
	G34467<=G34341 or G18717;
	G34468<=G34342 or G18718;
	G34494<=G26849 or G34413;
	G34535<=G34309 or G34073;
	G34537<=G34324 or G34084;
	G34598<=G34541 or G18136;
	G34599<=G34542 or G18149;
	G34600<=G34538 or G18182;
	G34601<=G34488 or G18211;
	G34602<=G34489 or G18269;
	G34603<=G34561 or G15075;
	G34604<=G34563 or G15076;
	G34605<=G34566 or G15077;
	G34606<=G34564 or G15080;
	G34607<=G34567 or G15081;
	G34608<=G34568 or G15082;
	G34609<=G34503 or G18563;
	G34610<=G34507 or G18564;
	G34611<=G34508 or G18565;
	G34612<=G34514 or G18566;
	G34613<=G34515 or G18567;
	G34614<=G34518 or G18568;
	G34615<=G34516 or G18576;
	G34616<=G34519 or G18577;
	G34617<=G34526 or G18579;
	G34618<=G34527 or G18580;
	G34619<=G34528 or G18581;
	G34620<=G34529 or G18582;
	G34621<=G34517 or G18583;
	G34622<=G34520 or G18584;
	G34623<=G34525 or G18585;
	G34624<=G34509 or G18592;
	G34625<=G34532 or G18610;
	G34626<=G34533 or G18627;
	G34627<=G34534 or G18644;
	G34628<=G34493 or G18653;
	G34629<=G34495 or G18654;
	G34630<=G34560 or G15117;
	G34631<=G34562 or G15118;
	G34632<=G34565 or G15119;
	G34633<=G34481 or G18690;
	G34634<=G34483 or G18691;
	G34635<=G34485 or G18692;
	G34636<=G34476 or G18693;
	G34637<=G34478 or G18694;
	G34638<=G34484 or G18721;
	G34639<=G34486 or G18722;
	G34640<=G34487 or G18723;
	G34641<=G34479 or G18724;
	G34642<=G34482 or G18725;
	G34643<=G34554 or G18752;
	G34644<=G34555 or G18769;
	G34645<=G34556 or G18786;
	G34646<=G34557 or G18803;
	G34647<=G34558 or G18820;
	G34649<=G33111 or G34492;
	G34657<=G33114 or G34497;
	G34663<=G32028 or G34500;
	G34693<=G34513 or G34310;
	G34695<=G34523 or G34322;
	G34708<=G33381 or G34572;
	G34719<=G34701 or G18133;
	G34720<=G34694 or G18134;
	G34721<=G34696 or G18135;
	G34722<=G34707 or G18137;
	G34723<=G34710 or G18139;
	G34724<=G34702 or G18152;
	G34725<=G34700 or G18183;
	G34726<=G34665 or G18212;
	G34727<=G34655 or G18213;
	G34728<=G34661 or G18214;
	G34729<=G34666 or G18270;
	G34730<=G34658 or G18271;
	G34731<=G34662 or G18272;
	G34732<=G34686 or G18593;
	G34733<=G34678 or G18651;
	G34734<=G34681 or G18652;
	G34735<=G34709 or G15116;
	G34761<=G34679 or G34506;
	G34762<=G34687 or G34524;
	G34781<=G33431 or G34715;
	G34783<=G33110 or G34667;
	G34790<=G34774 or G18151;
	G34791<=G34771 or G18184;
	G34792<=G34750 or G18569;
	G34793<=G34744 or G18570;
	G34794<=G34746 or G18571;
	G34795<=G34753 or G18572;
	G34796<=G34745 or G18573;
	G34797<=G34747 or G18574;
	G34798<=G34754 or G18575;
	G34799<=G34751 or G18578;
	G34800<=G34752 or G18586;
	G34801<=G34756 or G18588;
	G34802<=G34757 or G18589;
	G34803<=G34758 or G18590;
	G34804<=G34740 or G18591;
	G34805<=G34748 or G18594;
	G34806<=G34763 or G18595;
	G34807<=G34764 or G18596;
	G34808<=G34765 or G18599;
	G34809<=G33677 or G34738;
	G34819<=G34741 or G34684;
	G34826<=G34742 or G34685;
	G34843<=G33924 or G34782;
	G34849<=G34842 or G18154;
	G34850<=G34841 or G18185;
	G34856<=G34811 or G34743;
	G34880<=G34867 or G18153;
	G34881<=G34866 or G18187;
	G34882<=G34876 or G18659;
	G34884<=G34858 or G21666;
	G34887<=G34865 or G21670;
	G34890<=G34863 or G21674;
	G34894<=G34862 or G21678;
	G34897<=G34861 or G21682;
	G34900<=G34860 or G21686;
	G34903<=G34859 or G21690;
	G34906<=G34857 or G21694;
	G34911<=G34909 or G18188;
	G34931<=G2984 or G34912;
	G34957<=G34948 or G21662;
	G34970<=G34868 or G34961;
	G34971<=G34869 or G34962;
	G34974<=G34870 or G34963;
	G34975<=G34871 or G34964;
	G34976<=G34872 or G34965;
	G34977<=G34873 or G34966;
	G34978<=G34874 or G34967;
	G34979<=G34875 or G34968;
	G34980<=G34969 or G18587;
	G35000<=G34953 or G34999;
	I12583<=G1157 or G1239 or G990;
	I12611<=G1500 or G1582 or G1333;
	I12782<=G4188 or G4194 or G4197 or G4200;
	I12783<=G4204 or G4207 or G4210 or G4180;
	I12902<=G4235 or G4232 or G4229 or G4226;
	I12903<=G4222 or G4219 or G4216 or G4213;
	I18385<=G14413 or G14391 or G14360;
	I18417<=G14444 or G14414 or G14392;
	I18421<=G14447 or G14417 or G14395;
	I18449<=G14512 or G14445 or G14415;
	I18452<=G14514 or G14448 or G14418;
	I18492<=G14538 or G14513 or G14446;
	I18495<=G14539 or G14515 or G14449;
	I18543<=G14568 or G14540 or G14516;
	I22267<=G20236 or G20133 or G20111;
	I22280<=G20271 or G20150 or G20134;
	I22298<=G20371 or G20161 or G20151;
	I22830<=G21429 or G21338 or G21307;
	I22852<=G21459 or G21350 or G21339;
	I22880<=G21509 or G21356 or G21351;
	I22912<=G21555 or G21364 or G21357;
	I22958<=G21603 or G21386 or G21365;
	I23162<=G19919 or G19968 or G20014 or G20841;
	I23163<=G20982 or G21127 or G21193 or G21256;
	I23755<=G22904 or G22927 or G22980 or G23444;
	I23756<=G23457 or G23480 or G23494 or G23511;
	I24117<=G23088 or G23154 or G23172;
	I25612<=G25567 or G25568 or G25569 or G25570;
	I25613<=G25571 or G25572 or G25573 or G25574;
	I25736<=G12 or G22150 or G20277;
	I26522<=G19890 or G19935 or G19984 or G26365;
	I26523<=G20720 or G20857 or G20998 or G21143;
	I26643<=G27073 or G27058 or G27045 or G27040;
	I26644<=G27057 or G27044 or G27039 or G27032;
	I26741<=G22881 or G22905 or G22928 or G27402;
	I26742<=G23430 or G23445 or G23458 or G23481;
	I28147<=G2946 or G24561 or G28220;
	I28566<=G29201 or G29202 or G29203 or G28035;
	I28567<=G29204 or G29205 or G29206 or G29207;
	I29351<=G29328 or G29323 or G29316 or G30316;
	I29352<=G29322 or G29315 or G30315 or G30308;
	I29985<=G29385 or G31376 or G30735 or G30825;
	I29986<=G31070 or G31194 or G30614 or G30673;
	I30054<=G29385 or G31376 or G30735 or G30825;
	I30055<=G31070 or G31170 or G30614 or G30673;
	I30123<=G29385 or G31376 or G30735 or G30825;
	I30124<=G31070 or G31154 or G30614 or G30673;
	I30192<=G29385 or G31376 or G30735 or G30825;
	I30193<=G31070 or G30614 or G30673 or G31528;
	I30261<=G29385 or G31376 or G30735 or G30825;
	I30262<=G31672 or G31710 or G31021 or G30937;
	I30330<=G29385 or G31376 or G30735 or G30825;
	I30331<=G31672 or G31710 or G31021 or G30937;
	I30399<=G29385 or G31376 or G30735 or G30825;
	I30400<=G31021 or G30937 or G31327 or G30614;
	I30468<=G29385 or G31376 or G30735 or G30825;
	I30469<=G31672 or G31710 or G31021 or G30937;
	I30717<=G31787 or G32200 or G31940 or G31949;
	I30718<=G32348 or G32356 or G32097 or G32020;
	I30727<=G31759 or G32196 or G31933 or G31941;
	I30728<=G32345 or G32350 or G32056 or G32018;
	I30734<=G31790 or G32191 or G32086 or G32095;
	I30735<=G32369 or G32376 or G32089 or G32035;
	I30740<=G31776 or G32188 or G32083 or G32087;
	I30741<=G32085 or G32030 or G32224 or G32013;
	I30745<=G31777 or G32321 or G32069 or G32084;
	I30746<=G32047 or G31985 or G31991 or G32309;
	I30750<=G31788 or G32310 or G32054 or G32070;
	I30751<=G32042 or G32161 or G31943 or G31959;
	I30755<=G30564 or G32303 or G32049 or G32055;
	I30756<=G32088 or G32163 or G32098 or G32105;
	I30760<=G31778 or G32295 or G32046 or G32050;
	I30761<=G32071 or G32167 or G32067 or G32082;
	I31838<=G33461 or G33462 or G33463 or G33464;
	I31839<=G33465 or G33466 or G33467 or G33468;
	I31843<=G33470 or G33471 or G33472 or G33473;
	I31844<=G33474 or G33475 or G33476 or G33477;
	I31848<=G33479 or G33480 or G33481 or G33482;
	I31849<=G33483 or G33484 or G33485 or G33486;
	I31853<=G33488 or G33489 or G33490 or G33491;
	I31854<=G33492 or G33493 or G33494 or G33495;
	I31858<=G33497 or G33498 or G33499 or G33500;
	I31859<=G33501 or G33502 or G33503 or G33504;
	I31863<=G33506 or G33507 or G33508 or G33509;
	I31864<=G33510 or G33511 or G33512 or G33513;
	I31868<=G33515 or G33516 or G33517 or G33518;
	I31869<=G33519 or G33520 or G33521 or G33522;
	I31873<=G33524 or G33525 or G33526 or G33527;
	I31874<=G33528 or G33529 or G33530 or G33531;
	G7139<= not (G5406 or G5366);
	G7142<= not (G6573 or G6565);
	G7158<= not (G5752 or G5712);
	G7175<= not (G6098 or G6058);
	G7192<= not (G6444 or G6404);
	G7304<= not (G1183 or G1171);
	G7352<= not (G1526 or G1514);
	G7499<= not (G333 or G355);
	G7567<= not (G979 or G990);
	G7601<= not (G1322 or G1333);
	G7661<= not (G1211 or G1216 or G1221 or G1205);
	G7675<= not (G1554 or G1559 or G1564 or G1548);
	G7781<= not (G4064 or G4057);
	G8086<= not (G168 or G174 or G182);
	G8131<= not (G4776 or G4801 or G4793);
	G8177<= not (G4966 or G4991 or G4983);
	G8182<= not (G405 or G392);
	G8720<= not (G358 or G365);
	G8864<= not (G3179 or G3171);
	G8906<= not (G3530 or G3522);
	G8933<= not (G4709 or G4785);
	G8958<= not (G3881 or G3873);
	G8984<= not (G4899 or G4975);
	G9015<= not (G3050 or G3010);
	G9061<= not (G3401 or G3361);
	G9100<= not (G3752 or G3712);
	G9586<= not (G1668 or G1592);
	G9602<= not (G4688 or G4681 or G4674 or G4646);
	G9640<= not (G1802 or G1728);
	G9649<= not (G2227 or G2153);
	G9664<= not (G4878 or G4871 or G4864 or G4836);
	G9694<= not (G1936 or G1862);
	G9700<= not (G2361 or G2287);
	G9755<= not (G2070 or G1996);
	G9762<= not (G2495 or G2421);
	G9835<= not (G2629 or G2555);
	G10123<= not (G4294 or G4297);
	G10179<= not (G2098 or G1964 or G1830 or G1696);
	G10205<= not (G2657 or G2523 or G2389 or G2255);
	G10266<= not (G5188 or G5180);
	G10281<= not (G5535 or G5527);
	G10312<= not (G5881 or G5873);
	G10318<= not (G25 or G22);
	G10338<= not (G5062 or G5022);
	G10341<= not (G6227 or G6219);
	G10421<= not (G6227 or G9518);
	G10488<= not (G4616 or G7133 or G10336);
	G10491<= not (G6573 or G9576);
	G10510<= not (G7183 or G4593 or G4584);
	G10555<= not (G7227 or G4601 or G4608);
	G10615<= not (G1636 or G7308);
	G10649<= not (G1183 or G8407);
	G10666<= not (G8462 or G1171);
	G10671<= not (G1526 or G8466);
	G10695<= not (G8462 or G8407);
	G10699<= not (G8526 or G1514);
	G10709<= not (G7499 or G351);
	G10715<= not (G8526 or G8466);
	G10760<= not (G1046 or G7479);
	G10793<= not (G1389 or G7503);
	G10799<= not (G347 or G7541);
	G10801<= not (G1041 or G7479);
	G10803<= not (G1384 or G7503);
	G10808<= not (G8509 or G7611);
	G10819<= not (G7479 or G1041);
	G10821<= not (G7503 or G1384);
	G10831<= not (G7690 or G7827);
	G10862<= not (G7701 or G7840);
	G10884<= not (G7650 or G8451);
	G10893<= not (G1189 or G7715 or G7749);
	G10899<= not (G4064 or G8451);
	G10918<= not (G1532 or G7751 or G7778);
	G10922<= not (G7650 or G4057);
	G11006<= not (G7686 or G7836);
	G11012<= not (G7693 or G7846);
	G11039<= not (G9056 or G9092);
	G11107<= not (G9095 or G9177);
	G11119<= not (G9180 or G9203);
	G11148<= not (G8052 or G9197 or G9174 or G9050);
	G11171<= not (G8088 or G9226 or G9200 or G9091);
	G11184<= not (G513 or G9040);
	G11185<= not (G8038 or G8183 or G6804);
	G11191<= not (G4776 or G4801 or G9030);
	G11194<= not (G3288 or G6875);
	G11201<= not (G4125 or G7765);
	G11203<= not (G4966 or G4991 or G9064);
	G11207<= not (G3639 or G6905);
	G11213<= not (G4776 or G7892 or G9030);
	G11216<= not (G7998 or G8037);
	G11217<= not (G8531 or G6875);
	G11225<= not (G3990 or G6928);
	G11231<= not (G7928 or G4801 or G4793);
	G11232<= not (G4966 or G7898 or G9064);
	G11238<= not (G8584 or G6905);
	G11248<= not (G7953 or G4991 or G4983);
	G11252<= not (G8620 or G3057);
	G11255<= not (G8623 or G6928);
	G11261<= not (G7928 or G4801 or G9030);
	G11270<= not (G8431 or G8434);
	G11273<= not (G3061 or G8620);
	G11276<= not (G8534 or G8691);
	G11280<= not (G8647 or G3408);
	G11283<= not (G7953 or G4991 or G9064);
	G11303<= not (G8497 or G8500);
	G11306<= not (G3412 or G8647);
	G11309<= not (G8587 or G8728);
	G11313<= not (G8669 or G3759);
	G11345<= not (G8477 or G8479);
	G11346<= not (G7980 or G7964);
	G11357<= not (G8558 or G8561);
	G11360<= not (G3763 or G8669);
	G11363<= not (G8626 or G8751);
	G11384<= not (G8538 or G8540);
	G11385<= not (G8021 or G7985);
	G11414<= not (G8591 or G8593);
	G11415<= not (G8080 or G8026);
	G11435<= not (G8107 or G3171);
	G11448<= not (G4191 or G8790);
	G11469<= not (G650 or G9903 or G645);
	G11473<= not (G8107 or G8059);
	G11483<= not (G8165 or G3522);
	G11493<= not (G8964 or G8967);
	G11514<= not (G10295 or G3161 or G3155);
	G11527<= not (G8165 or G8114);
	G11537<= not (G8229 or G3873);
	G11563<= not (G8059 or G8011);
	G11566<= not (G3161 or G7964);
	G11571<= not (G10323 or G3512 or G3506);
	G11584<= not (G8229 or G8172);
	G11607<= not (G8848 or G8993 or G376);
	G11610<= not (G7980 or G3155);
	G11618<= not (G8114 or G8070);
	G11621<= not (G3512 or G7985);
	G11626<= not (G7121 or G3863 or G3857);
	G11653<= not (G7980 or G7964);
	G11658<= not (G8021 or G3506);
	G11666<= not (G8172 or G8125);
	G11669<= not (G3863 or G8026);
	G11692<= not (G8021 or G7985);
	G11697<= not (G8080 or G3857);
	G11715<= not (G8080 or G8026);
	G11729<= not (G3179 or G8059);
	G11747<= not (G3530 or G8114);
	G11755<= not (G4709 or G8796);
	G11763<= not (G3881 or G8172);
	G11771<= not (G8921 or G4185);
	G11773<= not (G8883 or G4785);
	G11780<= not (G4899 or G8822);
	G11797<= not (G8883 or G8796);
	G11804<= not (G8938 or G4975);
	G11834<= not (G8938 or G8822);
	G11846<= not (G7635 or G7518 or G7548);
	G11862<= not (G7134 or G7150);
	G11869<= not (G7649 or G7534 or G7581);
	G11885<= not (G7153 or G7167);
	G11891<= not (G812 or G9166);
	G11907<= not (G7170 or G7184);
	G11913<= not (G7197 or G9166);
	G11924<= not (G7187 or G7209);
	G11932<= not (G843 or G9166);
	G11935<= not (G9485 or G7267);
	G11940<= not (G2712 or G10084);
	G11945<= not (G7212 or G7228);
	G11950<= not (G9220 or G9166);
	G11954<= not (G9538 or G7314);
	G11958<= not (G9543 or G7327);
	G11972<= not (G9591 or G7361);
	G11976<= not (G9595 or G7379);
	G11995<= not (G9645 or G7410);
	G11999<= not (G9654 or G7423);
	G12002<= not (G5297 or G7004);
	G12017<= not (G9969 or G9586);
	G12025<= not (G9705 or G7461);
	G12026<= not (G9417 or G9340);
	G12029<= not (G5644 or G7028);
	G12046<= not (G10036 or G9640);
	G12050<= not (G10038 or G9649);
	G12059<= not (G9853 or G7004);
	G12067<= not (G5990 or G7051);
	G12081<= not (G10079 or G9694);
	G12085<= not (G10082 or G9700);
	G12093<= not (G9924 or G7028);
	G12101<= not (G6336 or G7074);
	G12113<= not (G1648 or G8187);
	G12117<= not (G10113 or G9755);
	G12121<= not (G10117 or G9762);
	G12123<= not (G6856 or G2748);
	G12126<= not (G9989 or G5069);
	G12129<= not (G9992 or G7051);
	G12137<= not (G6682 or G7097);
	G12146<= not (G1783 or G8241);
	G12150<= not (G2208 or G8259);
	G12154<= not (G10155 or G9835);
	G12160<= not (G9721 or G9724);
	G12163<= not (G5073 or G9989);
	G12166<= not (G9856 or G10124);
	G12170<= not (G10047 or G5413);
	G12173<= not (G10050 or G7074);
	G12189<= not (G1917 or G8302);
	G12193<= not (G2342 or G8316);
	G12198<= not (G9797 or G9800);
	G12201<= not (G5417 or G10047);
	G12204<= not (G9927 or G10160);
	G12208<= not (G10096 or G5759);
	G12211<= not (G10099 or G7097);
	G12223<= not (G2051 or G8365);
	G12226<= not (G2476 or G8373);
	G12228<= not (G10222 or G10206 or G10184 or G10335);
	G12234<= not (G9776 or G9778);
	G12235<= not (G9234 or G9206);
	G12246<= not (G9880 or G9883);
	G12249<= not (G5763 or G10096);
	G12252<= not (G9995 or G10185);
	G12256<= not (G10136 or G6105);
	G12288<= not (G2610 or G8418);
	G12296<= not (G9860 or G9862);
	G12297<= not (G9269 or G9239);
	G12308<= not (G9951 or G9954);
	G12311<= not (G6109 or G10136);
	G12314<= not (G10053 or G10207);
	G12318<= not (G10172 or G6451);
	G12333<= not (G1624 or G8139);
	G12346<= not (G9931 or G9933);
	G12347<= not (G9321 or G9274);
	G12358<= not (G10019 or G10022);
	G12361<= not (G6455 or G10172);
	G12364<= not (G10102 or G10224);
	G12371<= not (G1760 or G8195);
	G12374<= not (G2185 or G8205);
	G12377<= not (G6856 or G2748 or G9708);
	G12405<= not (G9374 or G5180);
	G12418<= not (G9999 or G10001);
	G12419<= not (G9402 or G9326);
	G12432<= not (G1894 or G8249);
	G12435<= not (G9012 or G8956 or G8904 or G8863);
	G12437<= not (G2319 or G8267);
	G12443<= not (G9374 or G9300);
	G12453<= not (G9444 or G5527);
	G12466<= not (G10057 or G10059);
	G12467<= not (G9472 or G9407);
	G12479<= not (G2028 or G8310);
	G12483<= not (G2453 or G8324);
	G12486<= not (G9055 or G9013 or G8957 or G8905);
	G12492<= not (G7704 or G5170 or G5164);
	G12505<= not (G9444 or G9381);
	G12515<= not (G9511 or G5873);
	G12540<= not (G2587 or G8381);
	G12550<= not (G9300 or G9259);
	G12553<= not (G5170 or G9206);
	G12558<= not (G7738 or G5517 or G5511);
	G12571<= not (G9511 or G9451);
	G12581<= not (G9569 or G6219);
	G12591<= not (G504 or G9040);
	G12593<= not (G9234 or G5164);
	G12601<= not (G9381 or G9311);
	G12604<= not (G5517 or G9239);
	G12609<= not (G7766 or G5863 or G5857);
	G12622<= not (G9569 or G9518);
	G12632<= not (G9631 or G6565);
	G12645<= not (G4467 or G6961);
	G12646<= not (G9234 or G9206);
	G12651<= not (G9269 or G5511);
	G12659<= not (G9451 or G9392);
	G12662<= not (G5863 or G9274);
	G12667<= not (G7791 or G6209 or G6203);
	G12680<= not (G9631 or G9576);
	G12695<= not (G9269 or G9239);
	G12700<= not (G9321 or G5857);
	G12708<= not (G9518 or G9462);
	G12711<= not (G6209 or G9326);
	G12716<= not (G7812 or G6555 or G6549);
	G12729<= not (G1657 or G8139);
	G12739<= not (G9321 or G9274);
	G12744<= not (G9402 or G6203);
	G12752<= not (G9576 or G9529);
	G12755<= not (G6555 or G9407);
	G12772<= not (G5188 or G9300);
	G12780<= not (G9402 or G9326);
	G12785<= not (G9472 or G6549);
	G12798<= not (G5535 or G9381);
	G12806<= not (G9472 or G9407);
	G12821<= not (G7132 or G10223 or G7149 or G10261);
	G12824<= not (G5881 or G9451);
	G12846<= not (G6837 or G10430);
	G12847<= not (G6838 or G10430);
	G12848<= not (G6839 or G10430);
	G12849<= not (G6840 or G10430);
	G12850<= not (G10430 or G6845);
	G12851<= not (G6846 or G10430);
	G12852<= not (G6847 or G10430);
	G12853<= not (G6848 or G10430);
	G12854<= not (G6849 or G10430);
	G12855<= not (G10430 or G6854);
	G12856<= not (G10430 or G6855);
	G12858<= not (G10365 or G10430);
	G12970<= not (G10555 or G10510 or G10488);
	G12980<= not (G7909 or G10741);
	G13004<= not (G7933 or G10741);
	G13005<= not (G7939 or G10762);
	G13013<= not (G7957 or G10762);
	G13021<= not (G7544 or G10741);
	G13031<= not (G7301 or G10741);
	G13032<= not (G7577 or G10762);
	G13044<= not (G7349 or G10762);
	G13056<= not (G7400 or G10741);
	G13076<= not (G7443 or G10741);
	G13078<= not (G7446 or G10762);
	G13094<= not (G7487 or G10762);
	G13110<= not (G7841 or G10741);
	G13114<= not (G7528 or G10741);
	G13125<= not (G7863 or G10762);
	G13129<= not (G7553 or G10762);
	G13202<= not (G8347 or G10511);
	G13325<= not (G7841 or G10741);
	G13326<= not (G10929 or G10905);
	G13335<= not (G7851 or G10741);
	G13336<= not (G11330 or G11011);
	G13341<= not (G7863 or G10762);
	G13342<= not (G10961 or G10935);
	G13377<= not (G7873 or G10762);
	G13378<= not (G11374 or G11017);
	G13480<= not (G3017 or G11858);
	G13500<= not (G8480 or G12641);
	G13501<= not (G3368 or G11881);
	G13512<= not (G9077 or G12527);
	G13517<= not (G8541 or G12692);
	G13518<= not (G3719 or G11903);
	G13539<= not (G8594 or G12735);
	G13568<= not (G8046 or G12527);
	G13603<= not (G8009 or G10721);
	G13622<= not (G278 or G11166);
	G13631<= not (G8068 or G10733);
	G13661<= not (G528 or G11185);
	G13670<= not (G8123 or G10756);
	G13698<= not (G528 or G12527 or G11185);
	G13700<= not (G3288 or G11615);
	G13730<= not (G3639 or G11663);
	G13765<= not (G8531 or G11615);
	G13772<= not (G3990 or G11702);
	G13796<= not (G9158 or G12527);
	G13799<= not (G8584 or G11663);
	G13806<= not (G11245 or G4076);
	G13824<= not (G8623 or G11702);
	G13831<= not (G11245 or G7666);
	G13852<= not (G11320 or G8347);
	G13872<= not (G8745 or G11083);
	G13883<= not (G4709 or G4785 or G11155);
	G13908<= not (G4709 or G8796 or G11155);
	G13910<= not (G4899 or G4975 or G11173);
	G13913<= not (G8859 or G11083);
	G13919<= not (G3347 or G11276);
	G13937<= not (G8883 or G4785 or G11155);
	G13939<= not (G4899 or G8822 or G11173);
	G13944<= not (G10262 or G12259);
	G13946<= not (G8651 or G11083);
	G13947<= not (G8948 or G11083);
	G13954<= not (G8663 or G11276);
	G13959<= not (G3698 or G11309);
	G13970<= not (G8883 or G8796 or G11155);
	G13971<= not (G8938 or G4975 or G11173);
	G13989<= not (G8697 or G11309);
	G13994<= not (G4049 or G11363);
	G13996<= not (G8938 or G8822 or G11173);
	G14000<= not (G8766 or G12259);
	G14001<= not (G739 or G11083);
	G14002<= not (G8681 or G11083);
	G14003<= not (G9003 or G11083);
	G14027<= not (G8734 or G11363);
	G14033<= not (G8808 or G12259);
	G14036<= not (G8725 or G11083);
	G14037<= not (G8748 or G11083);
	G14064<= not (G9214 or G12259);
	G14090<= not (G8851 or G12259);
	G14091<= not (G8854 or G12259);
	G14092<= not (G8774 or G11083);
	G14093<= not (G8833 or G11083);
	G14094<= not (G8770 or G11083);
	G14121<= not (G8891 or G12259);
	G14122<= not (G8895 or G12259);
	G14124<= not (G8830 or G11083);
	G14145<= not (G8945 or G12259);
	G14163<= not (G8997 or G12259);
	G14164<= not (G9000 or G12259);
	G14165<= not (G8951 or G11083);
	G14176<= not (G9044 or G12259);
	G14178<= not (G8899 or G11083);
	G14181<= not (G9083 or G12259);
	G14188<= not (G9162 or G12259);
	G14194<= not (G5029 or G10515);
	G14211<= not (G9779 or G10823);
	G14212<= not (G5373 or G10537);
	G14227<= not (G9863 or G10838);
	G14228<= not (G5719 or G10561);
	G14247<= not (G9934 or G10869);
	G14248<= not (G6065 or G10578);
	G14253<= not (G10032 or G12259 or G9217);
	G14271<= not (G10002 or G10874);
	G14272<= not (G6411 or G10598);
	G14278<= not (G562 or G12259 or G9217);
	G14291<= not (G9839 or G12155);
	G14306<= not (G10060 or G10887);
	G14313<= not (G12016 or G9250);
	G14320<= not (G9257 or G11111);
	G14334<= not (G12044 or G9337);
	G14335<= not (G12045 or G9283);
	G14337<= not (G12049 or G9284);
	G14339<= not (G12289 or G2735);
	G14347<= not (G9309 or G11123);
	G14360<= not (G12078 or G9484);
	G14361<= not (G12079 or G9413);
	G14362<= not (G12080 or G9338);
	G14364<= not (G12083 or G9415);
	G14365<= not (G12084 or G9339);
	G14367<= not (G9547 or G12289);
	G14382<= not (G9390 or G11139);
	G14391<= not (G12112 or G9585);
	G14392<= not (G12114 or G9537);
	G14393<= not (G12115 or G9488);
	G14394<= not (G12116 or G9414);
	G14395<= not (G12118 or G9542);
	G14396<= not (G12119 or G9489);
	G14397<= not (G12120 or G9416);
	G14399<= not (G5297 or G12598);
	G14411<= not (G9460 or G11160);
	G14413<= not (G11914 or G9638);
	G14414<= not (G12145 or G9639);
	G14415<= not (G12147 or G9590);
	G14416<= not (G12148 or G9541);
	G14417<= not (G12149 or G9648);
	G14418<= not (G12151 or G9594);
	G14419<= not (G12152 or G9546);
	G14420<= not (G12153 or G9490);
	G14425<= not (G5644 or G12656);
	G14437<= not (G9527 or G11178);
	G14444<= not (G11936 or G9692);
	G14445<= not (G12188 or G9693);
	G14446<= not (G12190 or G9644);
	G14447<= not (G11938 or G9698);
	G14448<= not (G12192 or G9699);
	G14449<= not (G12194 or G9653);
	G14450<= not (G12195 or G9598);
	G14490<= not (G9853 or G12598);
	G14497<= not (G5990 or G12705);
	G14512<= not (G11955 or G9753);
	G14513<= not (G12222 or G9754);
	G14514<= not (G11959 or G9760);
	G14515<= not (G12225 or G9761);
	G14516<= not (G12227 or G9704);
	G14522<= not (G9924 or G12656);
	G14529<= not (G6336 or G12749);
	G14538<= not (G11973 or G9828);
	G14539<= not (G11977 or G9833);
	G14540<= not (G12287 or G9834);
	G14549<= not (G9992 or G12705);
	G14556<= not (G6682 or G12790);
	G14568<= not (G12000 or G9915);
	G14575<= not (G10050 or G12749);
	G14602<= not (G10099 or G12790);
	G14611<= not (G12333 or G9749);
	G14640<= not (G12371 or G9824);
	G14642<= not (G12374 or G9829);
	G14678<= not (G12432 or G9907);
	G14679<= not (G12437 or G9911);
	G14687<= not (G5352 or G12166);
	G14707<= not (G10143 or G12259);
	G14712<= not (G12479 or G9971);
	G14713<= not (G12483 or G9974);
	G14726<= not (G10090 or G12166);
	G14731<= not (G5698 or G12204);
	G14751<= not (G10622 or G10617 or G10609 or G10603);
	G14752<= not (G12540 or G10040);
	G14754<= not (G12821 or G2988);
	G14767<= not (G10130 or G12204);
	G14772<= not (G6044 or G12252);
	G14792<= not (G10653 or G10623 or G10618 or G10611);
	G14793<= not (G2988 or G12228);
	G14816<= not (G10166 or G12252);
	G14821<= not (G6390 or G12314);
	G14867<= not (G10191 or G12314);
	G14872<= not (G6736 or G12364);
	G14911<= not (G10213 or G12364);
	G14914<= not (G12822 or G12797);
	G14988<= not (G10816 or G10812 or G10805);
	G15049<= not (G13350 or G6799);
	G15050<= not (G12834 or G13350);
	G15051<= not (G6801 or G13350);
	G15052<= not (G12835 or G13350);
	G15053<= not (G12836 or G13350);
	G15054<= not (G12837 or G13350);
	G15055<= not (G6808 or G13350);
	G15056<= not (G6809 or G13350);
	G15057<= not (G6810 or G13350);
	G15058<= not (G12838 or G13350);
	G15059<= not (G12839 or G13350);
	G15060<= not (G13350 or G6814);
	G15061<= not (G6815 or G13394);
	G15062<= not (G6817 or G13394);
	G15063<= not (G6818 or G13394);
	G15064<= not (G6820 or G13394);
	G15065<= not (G13394 or G12840);
	G15066<= not (G12841 or G13394);
	G15067<= not (G12842 or G13394);
	G15068<= not (G6826 or G13416);
	G15069<= not (G6828 or G13416);
	G15070<= not (G6829 or G13416);
	G15071<= not (G6831 or G13416);
	G15072<= not (G13416 or G12843);
	G15073<= not (G12844 or G13416);
	G15074<= not (G12845 or G13416);
	G15086<= not (G13144 or G12859);
	G15087<= not (G12860 or G13144);
	G15088<= not (G13144 or G6874);
	G15089<= not (G13144 or G12861);
	G15090<= not (G13144 or G12862);
	G15091<= not (G13177 or G12863);
	G15092<= not (G12864 or G13177);
	G15093<= not (G13177 or G6904);
	G15094<= not (G13177 or G12865);
	G15095<= not (G13177 or G12866);
	G15096<= not (G13191 or G12867);
	G15097<= not (G12868 or G13191);
	G15098<= not (G13191 or G6927);
	G15099<= not (G13191 or G12869);
	G15100<= not (G13191 or G12870);
	G15101<= not (G12871 or G14591);
	G15102<= not (G14591 or G6954);
	G15106<= not (G12872 or G10430);
	G15120<= not (G12873 or G13605);
	G15121<= not (G12874 or G13605);
	G15122<= not (G6959 or G13605);
	G15123<= not (G6975 or G13605);
	G15126<= not (G12878 or G13605);
	G15127<= not (G12879 or G13605);
	G15128<= not (G13638 or G12880);
	G15129<= not (G6984 or G13638);
	G15130<= not (G13638 or G6985);
	G15131<= not (G12881 or G13638);
	G15132<= not (G12882 or G13638);
	G15133<= not (G12883 or G13638);
	G15134<= not (G13638 or G12884);
	G15135<= not (G6990 or G13638);
	G15136<= not (G13680 or G12885);
	G15137<= not (G6992 or G13680);
	G15138<= not (G13680 or G6993);
	G15139<= not (G12886 or G13680);
	G15140<= not (G12887 or G13680);
	G15141<= not (G12888 or G13680);
	G15142<= not (G13680 or G12889);
	G15143<= not (G6998 or G13680);
	G15144<= not (G13716 or G12890);
	G15145<= not (G12891 or G13716);
	G15146<= not (G13716 or G7003);
	G15147<= not (G13716 or G12892);
	G15148<= not (G13716 or G12893);
	G15149<= not (G13745 or G12894);
	G15150<= not (G12895 or G13745);
	G15151<= not (G13745 or G7027);
	G15152<= not (G13745 or G12896);
	G15153<= not (G13745 or G12897);
	G15154<= not (G13782 or G12898);
	G15155<= not (G12899 or G13782);
	G15156<= not (G13782 or G7050);
	G15157<= not (G13782 or G12900);
	G15158<= not (G13782 or G12901);
	G15159<= not (G13809 or G12902);
	G15160<= not (G12903 or G13809);
	G15161<= not (G13809 or G7073);
	G15162<= not (G13809 or G12904);
	G15163<= not (G13809 or G12905);
	G15164<= not (G13835 or G12906);
	G15165<= not (G12907 or G13835);
	G15166<= not (G13835 or G7096);
	G15167<= not (G13835 or G12908);
	G15168<= not (G13835 or G12909);
	G15170<= not (G7118 or G14279);
	G15372<= not (G817 or G14279);
	G15508<= not (G10320 or G14279);
	G15570<= not (G822 or G14279);
	G15578<= not (G7216 or G14279);
	G15585<= not (G11862 or G14194);
	G15594<= not (G10614 or G13026 or G7285);
	G15608<= not (G11885 or G14212);
	G15628<= not (G11907 or G14228);
	G15647<= not (G11924 or G14248);
	G15669<= not (G11945 or G14272);
	G15718<= not (G13858 or G11330);
	G15724<= not (G13858 or G11374);
	G15754<= not (G341 or G7440 or G13385);
	G15825<= not (G7666 or G13217);
	G15992<= not (G10929 or G13846);
	G16024<= not (G14216 or G11890);
	G16027<= not (G10929 or G13260);
	G16044<= not (G10961 or G13861);
	G16066<= not (G10929 or G13307);
	G16072<= not (G10961 or G13273);
	G16090<= not (G10961 or G13315);
	G16183<= not (G9223 or G13545);
	G16198<= not (G9247 or G13574);
	G16201<= not (G13462 or G4704);
	G16209<= not (G13478 or G4749);
	G16210<= not (G13479 or G4894);
	G16215<= not (G1211 or G13545);
	G16219<= not (G13498 or G4760);
	G16220<= not (G13499 or G4939);
	G16226<= not (G8052 or G13545);
	G16227<= not (G1554 or G13574);
	G16231<= not (G13515 or G4771);
	G16232<= not (G13516 or G4950);
	G16237<= not (G8088 or G13574);
	G16242<= not (G13529 or G4961);
	G16246<= not (G13551 or G11169);
	G16268<= not (G7913 or G13121);
	G16272<= not (G13580 or G11189);
	G16287<= not (G13622 or G11144);
	G16288<= not (G13794 or G417);
	G16292<= not (G7943 or G13134);
	G16313<= not (G8005 or G13600);
	G16424<= not (G8064 or G13628);
	G16476<= not (G8119 or G13667);
	G16479<= not (G14719 or G12490);
	G16488<= not (G13697 or G13656);
	G16581<= not (G13756 or G8086);
	G16646<= not (G13437 or G11020 or G11372);
	G17148<= not (G827 or G14279);
	G17174<= not (G9194 or G14279);
	G17175<= not (G1216 or G13545);
	G17180<= not (G1559 or G13574);
	G17190<= not (G723 or G14279);
	G17194<= not (G11039 or G13480);
	G17198<= not (G9282 or G14279);
	G17213<= not (G11107 or G13501);
	G17239<= not (G11119 or G13518);
	G17284<= not (G9253 or G14317);
	G17309<= not (G9305 or G14344);
	G17393<= not (G9386 or G14379);
	G17420<= not (G9456 or G14408);
	G17482<= not (G9523 or G14434);
	G17515<= not (G13221 or G10828);
	G17619<= not (G10179 or G12955);
	G17625<= not (G14541 or G12123);
	G17657<= not (G14751 or G12955);
	G17663<= not (G10205 or G12983);
	G17694<= not (G12435 or G12955);
	G17700<= not (G14792 or G12983);
	G17727<= not (G12486 or G12983);
	G17954<= not (G832 or G14279);
	G19063<= not (G7909 or G15674);
	G19070<= not (G16957 or G11720);
	G19140<= not (G7939 or G15695);
	G19209<= not (G12971 or G15614 or G11320);
	G19268<= not (G15979 or G962);
	G19338<= not (G16031 or G1306);
	G19388<= not (G17181 or G14256);
	G19400<= not (G17139 or G14206);
	G19401<= not (G17193 or G14296);
	G19402<= not (G15979 or G13133);
	G19413<= not (G17151 or G14221);
	G19422<= not (G16031 or G13141);
	G19430<= not (G17150 or G14220);
	G19436<= not (G17176 or G14233);
	G19444<= not (G17192 or G14295);
	G19453<= not (G17199 or G14316);
	G19778<= not (G16268 or G1061);
	G19793<= not (G16292 or G1404);
	G19853<= not (G15746 or G1052);
	G19873<= not (G15755 or G1395);
	G19880<= not (G16201 or G13634);
	G19887<= not (G3025 or G16275);
	G19890<= not (G16987 or G8058);
	G19906<= not (G16209 or G13672);
	G19907<= not (G16210 or G13676);
	G19919<= not (G16987 or G11205);
	G19932<= not (G3376 or G16296);
	G19935<= not (G17062 or G8113);
	G19951<= not (G16219 or G13709);
	G19953<= not (G16220 or G13712);
	G19968<= not (G17062 or G11223);
	G19981<= not (G3727 or G16316);
	G19984<= not (G17096 or G8171);
	G19997<= not (G16231 or G13739);
	G19999<= not (G16232 or G13742);
	G20000<= not (G13661 or G16264);
	G20014<= not (G17096 or G11244);
	G20027<= not (G16242 or G13779);
	G20149<= not (G17091 or G14185);
	G20183<= not (G17152 or G14222);
	G20234<= not (G17140 or G14207);
	G20390<= not (G17182 or G14257);
	G20717<= not (G5037 or G17217);
	G20720<= not (G17847 or G9299);
	G20841<= not (G17847 or G12027);
	G20854<= not (G5381 or G17243);
	G20857<= not (G17929 or G9380);
	G20982<= not (G17929 or G12065);
	G20995<= not (G5727 or G17287);
	G20998<= not (G18065 or G9450);
	G21062<= not (G9547 or G17297);
	G21127<= not (G18065 or G12099);
	G21140<= not (G6073 or G17312);
	G21143<= not (G15348 or G9517);
	G21193<= not (G15348 or G12135);
	G21206<= not (G6419 or G17396);
	G21209<= not (G15483 or G9575);
	G21250<= not (G9417 or G9340 or G17494);
	G21256<= not (G15483 or G12179);
	G21277<= not (G9417 or G9340 or G17467);
	G21284<= not (G16646 or G9690);
	G21389<= not (G10143 or G17748 or G12259);
	G21652<= not (G17619 or G17663);
	G21655<= not (G17657 or G17700);
	G21658<= not (G17694 or G17727);
	G22190<= not (G2827 or G18949);
	G22357<= not (G1024 or G19699);
	G22399<= not (G1367 or G19720);
	G22400<= not (G19345 or G15718);
	G22405<= not (G18957 or G20136 or G20114);
	G22448<= not (G1018 or G19699);
	G22450<= not (G19345 or G15724);
	G22488<= not (G19699 or G1002);
	G22491<= not (G1361 or G19720);
	G22513<= not (G1002 or G19699);
	G22514<= not (G19699 or G1018);
	G22517<= not (G19720 or G1345);
	G22521<= not (G1036 or G19699);
	G22522<= not (G19699 or G1024);
	G22523<= not (G1345 or G19720);
	G22524<= not (G19720 or G1361);
	G22535<= not (G19699 or G1030);
	G22536<= not (G1379 or G19720);
	G22537<= not (G19720 or G1367);
	G22539<= not (G1030 or G19699);
	G22540<= not (G19720 or G1373);
	G22545<= not (G1373 or G19720);
	G22654<= not (G7733 or G19506);
	G22929<= not (G19773 or G12970);
	G22983<= not (G979 or G16268 or G19853);
	G22993<= not (G1322 or G16292 or G19873);
	G23024<= not (G7936 or G19407);
	G23042<= not (G16581 or G19462 or G10685);
	G23051<= not (G7960 or G19427);
	G23052<= not (G8334 or G19916);
	G23063<= not (G16313 or G19887);
	G23079<= not (G8390 or G19965);
	G23108<= not (G16424 or G19932);
	G23124<= not (G8443 or G20011);
	G23135<= not (G16476 or G19981);
	G23204<= not (G10685 or G19462 or G16488);
	G23208<= not (G20035 or G16324);
	G23560<= not (G9607 or G20838);
	G23586<= not (G17284 or G20717);
	G23602<= not (G9672 or G20979);
	G23626<= not (G17309 or G20854);
	G23642<= not (G9733 or G21124);
	G23662<= not (G17393 or G20995);
	G23678<= not (G9809 or G21190);
	G23686<= not (G2767 or G21066);
	G23695<= not (G17420 or G21140);
	G23711<= not (G9892 or G21253);
	G23729<= not (G17482 or G21206);
	G23763<= not (G2795 or G21276);
	G23835<= not (G2791 or G21303);
	G23871<= not (G2811 or G21348);
	G23883<= not (G2779 or G21067);
	G23918<= not (G2799 or G21382);
	G23955<= not (G2823 or G18890);
	G23956<= not (G18957 or G18918 or G20136 or G20114);
	G24018<= not (I23162 or I23163);
	G24145<= not (G19402 or G19422);
	G24148<= not (G19268 or G19338);
	G24383<= not (G22409 or G22360);
	G24391<= not (G22190 or G14645);
	G24439<= not (G7400 or G22312);
	G24453<= not (G7446 or G22325);
	G24494<= not (G23513 or G23532);
	G24497<= not (G23533 or G23553);
	G24508<= not (G23577 or G23618);
	G24514<= not (G23619 or G23657);
	G24575<= not (G23498 or G23514);
	G24619<= not (G23554 or G23581);
	G24631<= not (G20516 or G20436 or G20219 or G22957);
	G24701<= not (G979 or G23024 or G19778);
	G24720<= not (G1322 or G23051 or G19793);
	G24751<= not (G3034 or G23105);
	G24766<= not (G3385 or G23132);
	G24779<= not (G3736 or G23167);
	G24875<= not (G8725 or G23850 or G11083);
	G24953<= not (G10262 or G23978 or G12259);
	G24959<= not (G8858 or G23324);
	G24976<= not (G671 or G23324);
	G24990<= not (G8898 or G23324);
	G25004<= not (G676 or G23324);
	G25005<= not (G6811 or G23324);
	G25022<= not (G714 or G23324);
	G25141<= not (G22228 or G10334);
	G25144<= not (G5046 or G23623);
	G25160<= not (G5390 or G23659);
	G25175<= not (G5736 or G23692);
	G25189<= not (G6082 or G23726);
	G25203<= not (G6428 or G23756);
	G25247<= not (G23763 or G14645);
	G25317<= not (G9766 or G23782);
	G25321<= not (G23835 or G14645);
	G25407<= not (G23871 or G14645);
	G25446<= not (G23686 or G14645);
	G25447<= not (G23883 or G14645);
	G25501<= not (G23918 or G14645);
	G25504<= not (G22550 or G7222);
	G25521<= not (G23955 or G14645);
	G25540<= not (G22409 or G22360);
	G25769<= not (G25453 or G25414);
	G25770<= not (G25417 or G25377);
	G25776<= not (G7166 or G24380 or G24369);
	G25777<= not (G25482 or G25456);
	G25778<= not (G25459 or G25420);
	G25784<= not (G25507 or G25485);
	G25785<= not (G25488 or G25462);
	G25800<= not (G25518 or G25510);
	G25851<= not (G4311 or G24380 or G24369);
	G25887<= not (G24984 or G11706);
	G25932<= not (G7680 or G24528);
	G25944<= not (G7716 or G24591);
	G25947<= not (G1199 or G24591);
	G25948<= not (G7752 or G24609);
	G25950<= not (G1070 or G24591);
	G25952<= not (G1542 or G24609);
	G25954<= not (G7750 or G24591);
	G25956<= not (G1413 or G24609);
	G25958<= not (G7779 or G24609);
	G26098<= not (G9073 or G24732);
	G26162<= not (G23052 or G24751);
	G26183<= not (G23079 or G24766);
	G26209<= not (G23124 or G24779);
	G26212<= not (G23837 or G25408);
	G26247<= not (G7995 or G24732);
	G26256<= not (G23873 or G25479);
	G26267<= not (G8033 or G24732);
	G26268<= not (G283 or G24825);
	G26296<= not (G8287 or G24732);
	G26297<= not (G8519 or G24825);
	G26298<= not (G8297 or G24825);
	G26309<= not (G8575 or G24825);
	G26314<= not (G24808 or G24802);
	G26330<= not (G8631 or G24825);
	G26338<= not (G8458 or G24825);
	G26346<= not (G8522 or G24825);
	G26515<= not (G24843 or G24822);
	G26545<= not (G24881 or G24855);
	G26546<= not (G24858 or G24846);
	G26573<= not (G24897 or G24884);
	G26574<= not (G24887 or G24861);
	G26598<= not (G8990 or G13756 or G24732);
	G26603<= not (G24908 or G24900);
	G26609<= not (G146 or G24732);
	G26625<= not (G23560 or G25144);
	G26628<= not (G8990 or G24732);
	G26645<= not (G23602 or G25160);
	G26649<= not (G9037 or G24732);
	G26667<= not (G23642 or G25175);
	G26686<= not (G23678 or G25189);
	G26715<= not (G23711 or G25203);
	G26865<= not (G25328 or G25290);
	G26872<= not (G25411 or G25371);
	G26873<= not (G25374 or G25331);
	G26976<= not (G5016 or G25791);
	G26993<= not (G5360 or G25805);
	G27007<= not (G5706 or G25821);
	G27010<= not (G6052 or G25839);
	G27012<= not (G6398 or G25856);
	G27027<= not (G26398 or G26484);
	G27046<= not (G7544 or G25888);
	G27059<= not (G7577 or G25895);
	G27063<= not (G26485 or G26516);
	G27093<= not (G26712 or G26749);
	G27102<= not (G26750 or G26779);
	G27337<= not (G8334 or G26616);
	G27338<= not (G9291 or G26616);
	G27343<= not (G8005 or G26616);
	G27344<= not (G8390 or G26636);
	G27345<= not (G9360 or G26636);
	G27352<= not (G7975 or G26616);
	G27353<= not (G8097 or G26616);
	G27354<= not (G8064 or G26636);
	G27355<= not (G8443 or G26657);
	G27356<= not (G9429 or G26657);
	G27364<= not (G8426 or G26616);
	G27366<= not (G8016 or G26636);
	G27367<= not (G8155 or G26636);
	G27368<= not (G8119 or G26657);
	G27379<= not (G8492 or G26636);
	G27381<= not (G8075 or G26657);
	G27382<= not (G8219 or G26657);
	G27400<= not (G8553 or G26657);
	G27479<= not (G9056 or G26616);
	G27499<= not (G9095 or G26636);
	G27511<= not (G22137 or G26866 or G20277);
	G27516<= not (G9180 or G26657);
	G27528<= not (G8770 or G26352 or G11083);
	G27629<= not (G8891 or G26382 or G12259);
	G27647<= not (G3004 or G26616);
	G27652<= not (G3355 or G26636);
	G27659<= not (G3706 or G26657);
	G27703<= not (G9607 or G25791);
	G27704<= not (G7239 or G25791);
	G27717<= not (G9492 or G26745);
	G27720<= not (G9253 or G25791);
	G27721<= not (G9672 or G25805);
	G27722<= not (G7247 or G25805);
	G27731<= not (G9229 or G25791);
	G27732<= not (G9364 or G25791);
	G27733<= not (G9305 or G25805);
	G27734<= not (G9733 or G25821);
	G27735<= not (G7262 or G25821);
	G27766<= not (G9716 or G25791);
	G27768<= not (G9264 or G25805);
	G27769<= not (G9434 or G25805);
	G27770<= not (G9386 or G25821);
	G27771<= not (G9809 or G25839);
	G27772<= not (G7297 or G25839);
	G27823<= not (G9792 or G25805);
	G27825<= not (G9316 or G25821);
	G27826<= not (G9501 or G25821);
	G27827<= not (G9456 or G25839);
	G27828<= not (G9892 or G25856);
	G27829<= not (G7345 or G25856);
	G27875<= not (G9875 or G25821);
	G27877<= not (G9397 or G25839);
	G27878<= not (G9559 or G25839);
	G27879<= not (G9523 or G25856);
	G27924<= not (G9946 or G25839);
	G27926<= not (G9467 or G25856);
	G27927<= not (G9621 or G25856);
	G27954<= not (G10014 or G25856);
	G27960<= not (G7134 or G25791);
	G27966<= not (G7153 or G25805);
	G27969<= not (G7170 or G25821);
	G27973<= not (G7187 or G25839);
	G27982<= not (G7212 or G25856);
	G28031<= not (G21209 or I26522 or I26523);
	G28106<= not (G7812 or G26994);
	G28149<= not (G27598 or G27612);
	G28340<= not (G27439 or G26339);
	G28353<= not (G9073 or G27654 or G24732);
	G28414<= not (G27467 or G26347);
	G28425<= not (G27493 or G26351);
	G28444<= not (G8575 or G27463 or G24825);
	G28452<= not (G3161 or G27602);
	G28457<= not (G7980 or G27602);
	G28462<= not (G3512 or G27617);
	G28468<= not (G3155 or G10295 or G27602);
	G28469<= not (G3171 or G27602);
	G28470<= not (G8021 or G27617);
	G28475<= not (G3863 or G27635);
	G28476<= not (G27627 or G26547);
	G28480<= not (G8059 or G27602);
	G28481<= not (G3506 or G10323 or G27617);
	G28482<= not (G3522 or G27617);
	G28483<= not (G8080 or G27635);
	G28491<= not (G8114 or G27617);
	G28492<= not (G3857 or G7121 or G27635);
	G28493<= not (G3873 or G27635);
	G28496<= not (G3179 or G27602);
	G28498<= not (G8172 or G27635);
	G28509<= not (G8107 or G27602);
	G28510<= not (G3530 or G27617);
	G28514<= not (G8165 or G27617);
	G28515<= not (G3881 or G27635);
	G28519<= not (G8011 or G27602 or G10295);
	G28520<= not (G8229 or G27635);
	G28521<= not (G27649 or G26604);
	G28529<= not (G8070 or G27617 or G10323);
	G28540<= not (G8125 or G27635 or G7121);
	G28552<= not (G10295 or G27602);
	G28568<= not (G10323 or G27617);
	G28584<= not (G7121 or G27635);
	G28803<= not (G27730 or G22763);
	G28953<= not (G5170 or G27999);
	G28981<= not (G9234 or G27999);
	G28986<= not (G5517 or G28010);
	G29005<= not (G5164 or G7704 or G27999);
	G29006<= not (G5180 or G27999);
	G29007<= not (G9269 or G28010);
	G29012<= not (G5863 or G28020);
	G29032<= not (G9300 or G27999);
	G29033<= not (G5511 or G7738 or G28010);
	G29034<= not (G5527 or G28010);
	G29035<= not (G9321 or G28020);
	G29040<= not (G6209 or G26977);
	G29069<= not (G9381 or G28010);
	G29070<= not (G5857 or G7766 or G28020);
	G29071<= not (G5873 or G28020);
	G29072<= not (G9402 or G26977);
	G29077<= not (G6555 or G26994);
	G29104<= not (G5188 or G27999);
	G29106<= not (G9451 or G28020);
	G29107<= not (G6203 or G7791 or G26977);
	G29108<= not (G6219 or G26977);
	G29109<= not (G9472 or G26994);
	G29141<= not (G9374 or G27999);
	G29142<= not (G5535 or G28010);
	G29144<= not (G9518 or G26977);
	G29145<= not (G6549 or G7812 or G26994);
	G29146<= not (G6565 or G26994);
	G29164<= not (G9444 or G28010);
	G29165<= not (G5881 or G28020);
	G29167<= not (G9576 or G26994);
	G29173<= not (G9259 or G27999 or G7704);
	G29174<= not (G9511 or G28020);
	G29175<= not (G6227 or G26977);
	G29179<= not (G9311 or G28010 or G7738);
	G29180<= not (G9569 or G26977);
	G29181<= not (G6573 or G26994);
	G29183<= not (G9392 or G28020 or G7766);
	G29184<= not (G9631 or G26994);
	G29187<= not (G7704 or G27999);
	G29189<= not (G9462 or G26977 or G7791);
	G29191<= not (G7738 or G28010);
	G29193<= not (G9529 or G26994 or G7812);
	G29198<= not (G7766 or G28020);
	G29200<= not (G7791 or G26977);
	G29359<= not (G7528 or G28167);
	G29361<= not (G7553 or G28174);
	G29370<= not (G28585 or G28599);
	G29497<= not (G22763 or G28241);
	G29503<= not (G22763 or G28250);
	G29675<= not (G28380 or G8236 or G8354);
	G29705<= not (G28399 or G8284 or G8404);
	G29873<= not (G6875 or G28458);
	G29886<= not (G3288 or G28458);
	G29889<= not (G6905 or G28471);
	G29898<= not (G6895 or G28458);
	G29900<= not (G3639 or G28471);
	G29903<= not (G6928 or G28484);
	G29908<= not (G6918 or G28471);
	G29910<= not (G3990 or G28484);
	G29915<= not (G6941 or G28484);
	G29916<= not (G8681 or G28504 or G11083);
	G29933<= not (G8808 or G28500 or G12259);
	G30106<= not (G28739 or G7268);
	G30117<= not (G28739 or G7252);
	G30119<= not (G28761 or G7315);
	G30123<= not (G28768 or G7328);
	G30129<= not (G28739 or G14537);
	G30130<= not (G28761 or G7275);
	G30132<= not (G28789 or G7362);
	G30134<= not (G28768 or G7280);
	G30136<= not (G28799 or G7380);
	G30143<= not (G28761 or G14566);
	G30144<= not (G28789 or G7322);
	G30146<= not (G28833 or G7411);
	G30147<= not (G28768 or G14567);
	G30148<= not (G28799 or G7335);
	G30150<= not (G28846 or G7424);
	G30156<= not (G28789 or G14587);
	G30157<= not (G28833 or G7369);
	G30159<= not (G28799 or G14589);
	G30160<= not (G28846 or G7387);
	G30162<= not (G28880 or G7462);
	G30169<= not (G28833 or G14613);
	G30170<= not (G28846 or G14615);
	G30171<= not (G28880 or G7431);
	G30183<= not (G28880 or G14644);
	G30240<= not (G7004 or G28982);
	G30249<= not (G5297 or G28982);
	G30252<= not (G7028 or G29008);
	G30260<= not (G7018 or G28982);
	G30262<= not (G5644 or G29008);
	G30265<= not (G7051 or G29036);
	G30271<= not (G7041 or G29008);
	G30273<= not (G5990 or G29036);
	G30276<= not (G7074 or G29073);
	G30280<= not (G7064 or G29036);
	G30282<= not (G6336 or G29073);
	G30285<= not (G7097 or G29110);
	G30288<= not (G7087 or G29073);
	G30290<= not (G6682 or G29110);
	G30294<= not (G7110 or G29110);
	G30601<= not (G16279 or G29718);
	G30613<= not (G4507 or G29365);
	G30922<= not (G16662 or G29810);
	G30929<= not (G29803 or G29835);
	G30934<= not (G29836 or G29850);
	G31008<= not (G30004 or G30026);
	G31068<= not (G4801 or G29540);
	G31116<= not (G7892 or G29540);
	G31117<= not (G4991 or G29556);
	G31119<= not (G7898 or G29556);
	G31121<= not (G4776 or G29540);
	G31126<= not (G7928 or G29540);
	G31127<= not (G4966 or G29556);
	G31133<= not (G7953 or G29556);
	G31134<= not (G8033 or G29679 or G24732);
	G31233<= not (G8522 or G29778 or G24825);
	G31294<= not (G11326 or G29660);
	G31318<= not (G4785 or G29697);
	G31372<= not (G8796 or G29697);
	G31373<= not (G4975 or G29725);
	G31469<= not (G8822 or G29725);
	G31476<= not (G4709 or G29697);
	G31482<= not (G8883 or G29697);
	G31483<= not (G4899 or G29725);
	G31491<= not (G8938 or G29725);
	G31498<= not (G9030 or G29540);
	G31506<= not (G4793 or G29540);
	G31507<= not (G9064 or G29556);
	G31515<= not (G4983 or G29556);
	G31935<= not (G30583 or G4349);
	G31942<= not (G8977 or G30583);
	G31965<= not (G30583 or G4358);
	G31970<= not (G9024 or G30583);
	G32017<= not (G31504 or G23475);
	G32212<= not (G8859 or G31262 or G11083);
	G32296<= not (G9044 or G31509 or G12259);
	G32424<= not (G8721 or G31294);
	G32455<= not (G31566 or I29985 or I29986);
	G32520<= not (G31554 or I30054 or I30055);
	G32585<= not (G31542 or I30123 or I30124);
	G32650<= not (G31579 or I30192 or I30193);
	G32715<= not (G31327 or I30261 or I30262);
	G32780<= not (G31327 or I30330 or I30331);
	G32845<= not (G30673 or I30399 or I30400);
	G32910<= not (G31327 or I30468 or I30469);
	G33075<= not (G31997 or G7163);
	G33084<= not (G31978 or G7655);
	G33085<= not (G31978 or G4311);
	G33088<= not (G31997 or G7224);
	G33089<= not (G31978 or G4322);
	G33090<= not (G31997 or G4593);
	G33092<= not (G31978 or G4332);
	G33093<= not (G31997 or G4601);
	G33094<= not (G31950 or G4639);
	G33095<= not (G31997 or G7236);
	G33096<= not (G31997 or G4608);
	G33097<= not (G31950 or G4628);
	G33098<= not (G31997 or G4616);
	G33100<= not (G32172 or G31188);
	G33103<= not (G32176 or G31212);
	G33107<= not (G32180 or G31223);
	G33108<= not (G32183 or G31228);
	G33109<= not (G31997 or G4584);
	G33112<= not (G31240 or G32194);
	G33117<= not (G31261 or G32205);
	G33125<= not (G8606 or G32057);
	G33128<= not (G4653 or G32057);
	G33129<= not (G8630 or G32072);
	G33130<= not (G32265 or G31497);
	G33131<= not (G4659 or G32057);
	G33132<= not (G4843 or G32072);
	G33133<= not (G32278 or G31503);
	G33134<= not (G7686 or G32057);
	G33135<= not (G32090 or G8350);
	G33137<= not (G4849 or G32072);
	G33138<= not (G32287 or G31514);
	G33139<= not (G8650 or G32057);
	G33140<= not (G7693 or G32072);
	G33141<= not (G32099 or G8400);
	G33143<= not (G32293 or G31518);
	G33144<= not (G4664 or G32057);
	G33145<= not (G8677 or G32072);
	G33146<= not (G4669 or G32057);
	G33147<= not (G32090 or G7788);
	G33148<= not (G4854 or G32072);
	G33160<= not (G8672 or G32057);
	G33161<= not (G32090 or G7806);
	G33162<= not (G4859 or G32072);
	G33163<= not (G32099 or G7809);
	G33174<= not (G8714 or G32072);
	G33175<= not (G32099 or G7828);
	G33419<= not (G31978 or G7627);
	G33427<= not (G10278 or G31950);
	G33432<= not (G31997 or G6978);
	G33437<= not (G31997 or G10275);
	G33438<= not (G31950 or G4621);
	G33439<= not (G31950 or G4633);
	G33447<= not (G31978 or G7643);
	G33448<= not (G7785 or G31950);
	G33449<= not (G10311 or G31950);
	G33823<= not (G8774 or G33306 or G11083);
	G33851<= not (G8854 or G33299 or G12259);
	G34067<= not (G33859 or G11772);
	G34354<= not (G9003 or G34162 or G11083);
	G34359<= not (G9162 or G34174 or G12259);
	G34496<= not (G34370 or G27648);
	G34703<= not (G8899 or G34545 or G11083);
	G34737<= not (G34706 or G30003);
	G34912<= not (G34883 or G20277 or G20242 or G21370);
end RTL;
