-- File created by Bench2VHDL
-- Name: s13207
-- File: bench/s13207.bench
-- Timestamp: 2019-05-21T22:08:28.876525
--
-- Original File
-- =============
--	# s13207.1
--	# 62 inputs
--	# 152 outputs
--	# 638 D-type flipflops
--	# 5378 inverters
--	# 2573 gates (1114 ANDs + 849 NANDs + 512 ORs + 98 NORs)
--	
--	INPUT(g43)
--	INPUT(g49)
--	INPUT(g633)
--	INPUT(g634)
--	INPUT(g635)
--	INPUT(g645)
--	INPUT(g647)
--	INPUT(g648)
--	INPUT(g690)
--	INPUT(g694)
--	INPUT(g698)
--	INPUT(g702)
--	INPUT(g722)
--	INPUT(g723)
--	INPUT(g751)
--	INPUT(g752)
--	INPUT(g753)
--	INPUT(g754)
--	INPUT(g755)
--	INPUT(g756)
--	INPUT(g757)
--	INPUT(g781)
--	INPUT(g941)
--	INPUT(g962)
--	INPUT(g1000)
--	INPUT(g1008)
--	INPUT(g1016)
--	INPUT(g1080)
--	INPUT(g1234)
--	INPUT(g1553)
--	INPUT(g1554)
--	INPUT(g786)
--	INPUT(g1206)
--	INPUT(g929)
--	INPUT(g955)
--	INPUT(g795)
--	INPUT(g1194)
--	INPUT(g1198)
--	INPUT(g1202)
--	INPUT(g24)
--	INPUT(g1203)
--	INPUT(g1196)
--	INPUT(g29)
--	INPUT(g22)
--	INPUT(g28)
--	INPUT(g10)
--	INPUT(g23)
--	INPUT(g37)
--	INPUT(g26)
--	INPUT(g1)
--	INPUT(g27)
--	INPUT(g42)
--	INPUT(g11)
--	INPUT(g32)
--	INPUT(g41)
--	INPUT(g31)
--	INPUT(g45)
--	INPUT(g9)
--	INPUT(g44)
--	INPUT(g21)
--	INPUT(g30)
--	INPUT(g25)
--	
--	OUTPUT(g206)
--	OUTPUT(g291)
--	OUTPUT(g372)
--	OUTPUT(g453)
--	OUTPUT(g534)
--	OUTPUT(g594)
--	OUTPUT(g785)
--	OUTPUT(g1006)
--	OUTPUT(g1015)
--	OUTPUT(g1017)
--	OUTPUT(g1246)
--	OUTPUT(g1724)
--	OUTPUT(g1783)
--	OUTPUT(g1798)
--	OUTPUT(g1804)
--	OUTPUT(g1810)
--	OUTPUT(g1817)
--	OUTPUT(g1824)
--	OUTPUT(g1829)
--	OUTPUT(g1870)
--	OUTPUT(g1871)
--	OUTPUT(g1894)
--	OUTPUT(g1911)
--	OUTPUT(g1944)
--	OUTPUT(g2662)
--	OUTPUT(g2844)
--	OUTPUT(g2888)
--	OUTPUT(g3077)
--	OUTPUT(g3096)
--	OUTPUT(g3130)
--	OUTPUT(g3159)
--	OUTPUT(g3191)
--	OUTPUT(g3829)
--	OUTPUT(g3859)
--	OUTPUT(g3860)
--	OUTPUT(g4267)
--	OUTPUT(g4316)
--	OUTPUT(g4370)
--	OUTPUT(g4371)
--	OUTPUT(g4372)
--	OUTPUT(g4373)
--	OUTPUT(g4655)
--	OUTPUT(g4657)
--	OUTPUT(g4660)
--	OUTPUT(g4661)
--	OUTPUT(g4663)
--	OUTPUT(g4664)
--	OUTPUT(g5143)
--	OUTPUT(g5164)
--	OUTPUT(g5571)
--	OUTPUT(g5669)
--	OUTPUT(g5678)
--	OUTPUT(g5682)
--	OUTPUT(g5684)
--	OUTPUT(g5687)
--	OUTPUT(g5729)
--	OUTPUT(g6207)
--	OUTPUT(g6212)
--	OUTPUT(g6223)
--	OUTPUT(g6236)
--	OUTPUT(g6269)
--	OUTPUT(g6425)
--	OUTPUT(g6648)
--	OUTPUT(g6653)
--	OUTPUT(g6675)
--	OUTPUT(g6849)
--	OUTPUT(g6850)
--	OUTPUT(g6895)
--	OUTPUT(g6909)
--	OUTPUT(g7048)
--	OUTPUT(g7063)
--	OUTPUT(g7103)
--	OUTPUT(g7283)
--	OUTPUT(g7284)
--	OUTPUT(g7285)
--	OUTPUT(g7286)
--	OUTPUT(g7287)
--	OUTPUT(g7288)
--	OUTPUT(g7289)
--	OUTPUT(g7290)
--	OUTPUT(g7291)
--	OUTPUT(g7292)
--	OUTPUT(g7293)
--	OUTPUT(g7294)
--	OUTPUT(g7295)
--	OUTPUT(g7298)
--	OUTPUT(g7423)
--	OUTPUT(g7424)
--	OUTPUT(g7425)
--	OUTPUT(g7474)
--	OUTPUT(g7504)
--	OUTPUT(g7505)
--	OUTPUT(g7506)
--	OUTPUT(g7507)
--	OUTPUT(g7508)
--	OUTPUT(g7514)
--	OUTPUT(g7729)
--	OUTPUT(g7730)
--	OUTPUT(g7731)
--	OUTPUT(g7732)
--	OUTPUT(g8216)
--	OUTPUT(g8217)
--	OUTPUT(g8218)
--	OUTPUT(g8219)
--	OUTPUT(g8234)
--	OUTPUT(g8661)
--	OUTPUT(g8663)
--	OUTPUT(g8872)
--	OUTPUT(g8958)
--	OUTPUT(g9128)
--	OUTPUT(g9132)
--	OUTPUT(g9204)
--	OUTPUT(g9280)
--	OUTPUT(g9297)
--	OUTPUT(g9299)
--	OUTPUT(g9305)
--	OUTPUT(g9308)
--	OUTPUT(g9310)
--	OUTPUT(g9312)
--	OUTPUT(g9314)
--	OUTPUT(g9378)
--	OUTPUT(g7763)
--	OUTPUT(g1205)
--	OUTPUT(g3856)
--	OUTPUT(g3857)
--	OUTPUT(g3854)
--	OUTPUT(g1193)
--	OUTPUT(g1197)
--	OUTPUT(g1201)
--	OUTPUT(g6294)
--	OUTPUT(g6376)
--	OUTPUT(g1195)
--	OUTPUT(g6300)
--	OUTPUT(g6292)
--	OUTPUT(g6298)
--	OUTPUT(g6291)
--	OUTPUT(g6293)
--	OUTPUT(g6304)
--	OUTPUT(g6296)
--	OUTPUT(g6289)
--	OUTPUT(g6297)
--	OUTPUT(g6306)
--	OUTPUT(g6290)
--	OUTPUT(g6303)
--	OUTPUT(g6305)
--	OUTPUT(g6302)
--	OUTPUT(g6308)
--	OUTPUT(g6288)
--	OUTPUT(g6307)
--	OUTPUT(g6299)
--	OUTPUT(g6301)
--	OUTPUT(g6295)
--	
--	g397 = DFF(g4635)
--	g1271 = DFF(g5176)
--	g312 = DFF(g4618)
--	g273 = DFF(g4611)
--	g452 = DFF(g449)
--	g948 = DFF(g8664)
--	g629 = DFF(g6827)
--	g207 = DFF(g5733)
--	g1541 = DFF(g7778)
--	g1153 = DFF(g6856)
--	g940 = DFF(g5735)
--	g976 = DFF(g8864)
--	g498 = DFF(g9111)
--	g314 = DFF(g4620)
--	g1092 = DFF(g7520)
--	g454 = DFF(g4639)
--	g196 = DFF(g5731)
--	g535 = DFF(g3844)
--	g292 = DFF(g4613)
--	g772 = DFF(g6846)
--	g1375 = DFF(g6869)
--	g689 = DFF(g6371)
--	g183 = DFF(g6309)
--	g359 = DFF(g6336)
--	g1384 = DFF(g6881)
--	g1339 = DFF(g6865)
--	g20 = DFF(g6386)
--	g1424 = DFF(g3862)
--	g767 = DFF(g6841)
--	g393 = DFF(g4631)
--	g1077 = DFF(g7767)
--	g1231 = DFF(g1236)
--	g294 = DFF(g4615)
--	g1477 = DFF(g9036)
--	g4 = DFF(g9372)
--	g608 = DFF(g6806)
--	g1205 = DFF(g1204)
--	g465 = DFF(g6352)
--	g774 = DFF(g6848)
--	g921 = DFF(g916)
--	g1304 = DFF(g1312)
--	g243 = DFF(g6318)
--	g1499 = DFF(g7772)
--	g80 = DFF(g6778)
--	g1444 = DFF(g5185)
--	g1269 = DFF(g5740)
--	g600 = DFF(g6807)
--	g423 = DFF(g9105)
--	g771 = DFF(g6845)
--	g803 = DFF(g7757)
--	g843 = DFF(g2647)
--	g315 = DFF(g4621)
--	g455 = DFF(g4640)
--	g906 = DFF(g901)
--	g622 = DFF(g6821)
--	g891 = DFF(g3855)
--	g1014 = DFF(g1012)
--	g984 = DFF(g9133)
--	g117 = DFF(g5153)
--	g137 = DFF(g5150)
--	g527 = DFF(g9110)
--	g1513 = DFF(g1524)
--	g278 = DFF(g6323)
--	g1378 = DFF(g6880)
--	g718 = DFF(g7753)
--	g598 = DFF(g6797)
--	g1182 = DFF(g1160)
--	g1288 = DFF(g7527)
--	g1382 = DFF(g6888)
--	g179 = DFF(g5159)
--	g624 = DFF(g6831)
--	g48 = DFF(g9362)
--	g362 = DFF(g9093)
--	g878 = DFF(g890)
--	g270 = DFF(g9092)
--	g763 = DFF(g6836)
--	g710 = DFF(g7751)
--	g730 = DFF(g7754)
--	g295 = DFF(g4616)
--	g1037 = DFF(g7519)
--	g1102 = DFF(g6855)
--	g483 = DFF(g6356)
--	g775 = DFF(g7759)
--	g621 = DFF(g6819)
--	g1364 = DFF(g6878)
--	g1454 = DFF(g5187)
--	g1296 = DFF(g7304)
--	g5 = DFF(g9373)
--	g1532 = DFF(g7781)
--	g587 = DFF(g3852)
--	g741 = DFF(g9386)
--	g13 = DFF(g7308)
--	g606 = DFF(g6804)
--	g1012 = DFF(g6851)
--	g52 = DFF(g6781)
--	g646 = DFF(g4652)
--	g1412 = DFF(g5745)
--	g327 = DFF(g6332)
--	g1189 = DFF(g6392)
--	g1389 = DFF(g4658)
--	g1029 = DFF(g2654)
--	g1371 = DFF(g6868)
--	g1429 = DFF(g2671)
--	g398 = DFF(g4636)
--	g985 = DFF(g7515)
--	g354 = DFF(g4624)
--	g619 = DFF(g6817)
--	g113 = DFF(g5148)
--	g133 = DFF(g5149)
--	g180 = DFF(g5158)
--	g1138 = DFF(g7524)
--	g1309 = DFF(g1308)
--	g889 = DFF(g7101)
--	g390 = DFF(g6341)
--	g625 = DFF(g6823)
--	g417 = DFF(g9103)
--	g681 = DFF(g7748)
--	g437 = DFF(g6348)
--	g351 = DFF(g9100)
--	g1201 = DFF(g1200)
--	g109 = DFF(g6785)
--	g1049 = DFF(g8673)
--	g1098 = DFF(g6854)
--	g200 = DFF(g199)
--	g240 = DFF(g6317)
--	g479 = DFF(g4649)
--	g126 = DFF(g6789)
--	g596 = DFF(g6795)
--	g1268 = DFF(g5175)
--	g222 = DFF(g6313)
--	g420 = DFF(g9104)
--	g3 = DFF(g9360)
--	g58 = DFF(g7734)
--	g172 = DFF(g1270)
--	g387 = DFF(g6340)
--	g840 = DFF(g2648)
--	g365 = DFF(g9094)
--	g1486 = DFF(g8226)
--	g1504 = DFF(g7773)
--	g1185 = DFF(g1155)
--	g1385 = DFF(g6883)
--	g583 = DFF(g3851)
--	g822 = DFF(g7512)
--	g1025 = DFF(g8871)
--	g969 = DFF(g966)
--	g768 = DFF(g6842)
--	g174 = DFF(g7737)
--	g685 = DFF(g7749)
--	g1087 = DFF(g6853)
--	g355 = DFF(g4625)
--	g911 = DFF(g906)
--	g1226 = DFF(g6859)
--	g99 = DFF(g6783)
--	g1045 = DFF(g8224)
--	g1173 = DFF(g7526)
--	g1373 = DFF(g6871)
--	g186 = DFF(g3830)
--	g760 = DFF(g6833)
--	g959 = DFF(g5169)
--	g1369 = DFF(g6875)
--	g1007 = DFF(g8867)
--	g1459 = DFF(g3863)
--	g758 = DFF(g6840)
--	g480 = DFF(g6355)
--	g396 = DFF(g4634)
--	g612 = DFF(g6811)
--	g38 = DFF(g5746)
--	g632 = DFF(g6830)
--	g1415 = DFF(g5180)
--	g1227 = DFF(g7108)
--	g246 = DFF(g6319)
--	g449 = DFF(g3840)
--	g517 = DFF(g4651)
--	g118 = DFF(g6787)
--	g138 = DFF(g6792)
--	g16 = DFF(g1404)
--	g284 = DFF(g9086)
--	g142 = DFF(g6793)
--	g219 = DFF(g6312)
--	g426 = DFF(g9106)
--	g1388 = DFF(g6882)
--	g806 = DFF(g7510)
--	g846 = DFF(g2646)
--	g1428 = DFF(g2672)
--	g579 = DFF(g3850)
--	g1030 = DFF(g7518)
--	g614 = DFF(g6812)
--	g1430 = DFF(g4666)
--	g1247 = DFF(g6380)
--	g669 = DFF(g7745)
--	g110 = DFF(g109)
--	g130 = DFF(g6790)
--	g225 = DFF(g6314)
--	g281 = DFF(g9085)
--	g819 = DFF(g7761)
--	g1308 = DFF(g6385)
--	g611 = DFF(g6810)
--	g631 = DFF(g6829)
--	g1217 = DFF(g6377)
--	g104 = DFF(g6784)
--	g1365 = DFF(g6867)
--	g825 = DFF(g7513)
--	g1333 = DFF(g6863)
--	g474 = DFF(g4644)
--	g1396 = DFF(g4662)
--	g141 = DFF(g5151)
--	g1509 = DFF(g7774)
--	g766 = DFF(g6839)
--	g1018 = DFF(g8869)
--	g588 = DFF(g9031)
--	g1467 = DFF(g8875)
--	g317 = DFF(g4623)
--	g457 = DFF(g4642)
--	g486 = DFF(g6357)
--	g471 = DFF(g6354)
--	g1381 = DFF(g6887)
--	g1197 = DFF(g1196)
--	g513 = DFF(g9116)
--	g1397 = DFF(g6389)
--	g533 = DFF(g530)
--	g1021 = DFF(g8870)
--	g1421 = DFF(g5179)
--	g952 = DFF(g8668)
--	g1263 = DFF(g5737)
--	g580 = DFF(g6368)
--	g615 = DFF(g6813)
--	g1257 = DFF(g5738)
--	g46 = DFF(g8955)
--	g402 = DFF(g6343)
--	g998 = DFF(g1005)
--	g1041 = DFF(g7765)
--	g297 = DFF(g6324)
--	g954 = DFF(g8670)
--	g105 = DFF(g104)
--	g145 = DFF(g5152)
--	g212 = DFF(g4601)
--	g1368 = DFF(g6874)
--	g232 = DFF(g4606)
--	g990 = DFF(g7516)
--	g475 = DFF(g4645)
--	g33 = DFF(g5184)
--	g951 = DFF(g8667)
--	g799 = DFF(g7756)
--	g812 = DFF(g7758)
--	g567 = DFF(g6367)
--	g313 = DFF(g4619)
--	g333 = DFF(g6334)
--	g168 = DFF(g7742)
--	g214 = DFF(g4603)
--	g234 = DFF(g4608)
--	g652 = DFF(g646)
--	g1126 = DFF(g8674)
--	g1400 = DFF(g6390)
--	g1326 = DFF(g7306)
--	g92 = DFF(g6794)
--	g309 = DFF(g6328)
--	g211 = DFF(g4600)
--	g834 = DFF(g2650)
--	g231 = DFF(g4605)
--	g557 = DFF(g6366)
--	g1383 = DFF(g6889)
--	g1220 = DFF(g6378)
--	g158 = DFF(g7740)
--	g627 = DFF(g6825)
--	g661 = DFF(g7743)
--	g77 = DFF(g6777)
--	g831 = DFF(g2651)
--	g1327 = DFF(g7307)
--	g293 = DFF(g4614)
--	g1146 = DFF(g1612)
--	g89 = DFF(g92)
--	g150 = DFF(g7738)
--	g773 = DFF(g6847)
--	g859 = DFF(g8221)
--	g1240 = DFF(g1235)
--	g518 = DFF(g6361)
--	g1472 = DFF(g8960)
--	g1443 = DFF(g4667)
--	g436 = DFF(g4638)
--	g405 = DFF(g6344)
--	g1034 = DFF(g8957)
--	g1147 = DFF(g1146)
--	g374 = DFF(g4627)
--	g98 = DFF(g5146)
--	g563 = DFF(g9029)
--	g510 = DFF(g9115)
--	g530 = DFF(g3842)
--	g215 = DFF(g4604)
--	g235 = DFF(g4609)
--	g1013 = DFF(g1014)
--	g6 = DFF(g9374)
--	g55 = DFF(g7733)
--	g1317 = DFF(g5743)
--	g504 = DFF(g9113)
--	g665 = DFF(g7744)
--	g544 = DFF(g6365)
--	g371 = DFF(g368)
--	g62 = DFF(g7509)
--	g792 = DFF(g5162)
--	g468 = DFF(g6353)
--	g815 = DFF(g7760)
--	g1460 = DFF(g4668)
--	g553 = DFF(g9028)
--	g623 = DFF(g6822)
--	g501 = DFF(g9112)
--	g1190 = DFF(g8677)
--	g1390 = DFF(g4659)
--	g74 = DFF(g6776)
--	g1156 = DFF(g1081)
--	g318 = DFF(g6329)
--	g458 = DFF(g4643)
--	g342 = DFF(g9097)
--	g1250 = DFF(g7111)
--	g1163 = DFF(g2655)
--	g1363 = DFF(g6877)
--	g1432 = DFF(g5183)
--	g1053 = DFF(g8873)
--	g252 = DFF(g6321)
--	g330 = DFF(g6333)
--	g264 = DFF(g9090)
--	g1157 = DFF(g1156)
--	g1357 = DFF(g8675)
--	g375 = DFF(g4628)
--	g68 = DFF(g6774)
--	g852 = DFF(g2644)
--	g261 = DFF(g9089)
--	g516 = DFF(g4650)
--	g536 = DFF(g6363)
--	g979 = DFF(g7104)
--	g778 = DFF(g7296)
--	g199 = DFF(g3832)
--	g1292 = DFF(g7302)
--	g290 = DFF(g287)
--	g1084 = DFF(g7106)
--	g1439 = DFF(g5182)
--	g770 = DFF(g6844)
--	g1276 = DFF(g6384)
--	g890 = DFF(g7102)
--	g1004 = DFF(g7105)
--	g1404 = DFF(g1403)
--	g93 = DFF(g5145)
--	g2 = DFF(g9361)
--	g287 = DFF(g3836)
--	g560 = DFF(g6370)
--	g1224 = DFF(g6857)
--	g1320 = DFF(g7114)
--	g617 = DFF(g6815)
--	g316 = DFF(g4622)
--	g336 = DFF(g9095)
--	g933 = DFF(g5166)
--	g456 = DFF(g4641)
--	g345 = DFF(g9098)
--	g628 = DFF(g6826)
--	g8 = DFF(g9376)
--	g887 = DFF(g7099)
--	g789 = DFF(g7297)
--	g173 = DFF(g7736)
--	g550 = DFF(g9027)
--	g255 = DFF(g9087)
--	g949 = DFF(g8665)
--	g1244 = DFF(g2659)
--	g620 = DFF(g6818)
--	g1435 = DFF(g5181)
--	g477 = DFF(g4647)
--	g926 = DFF(g878)
--	g368 = DFF(g3838)
--	g855 = DFF(g8220)
--	g1214 = DFF(g5736)
--	g1110 = DFF(g7299)
--	g1310 = DFF(g1309)
--	g296 = DFF(g4617)
--	g972 = DFF(g2653)
--	g1402 = DFF(g6391)
--	g1236 = DFF(g1240)
--	g896 = DFF(g891)
--	g613 = DFF(g6820)
--	g566 = DFF(g3848)
--	g1394 = DFF(g6388)
--	g1489 = DFF(g7770)
--	g883 = DFF(g921)
--	g47 = DFF(g9389)
--	g971 = DFF(g5171)
--	g609 = DFF(g6808)
--	g103 = DFF(g5157)
--	g1254 = DFF(g6381)
--	g556 = DFF(g3847)
--	g1409 = DFF(g5178)
--	g626 = DFF(g6824)
--	g1229 = DFF(g7110)
--	g782 = DFF(g5734)
--	g237 = DFF(g6316)
--	g942 = DFF(g2652)
--	g228 = DFF(g6315)
--	g706 = DFF(g7750)
--	g746 = DFF(g8956)
--	g1462 = DFF(g8678)
--	g963 = DFF(g7764)
--	g129 = DFF(g5156)
--	g837 = DFF(g2649)
--	g599 = DFF(g6798)
--	g1192 = DFF(g1191)
--	g828 = DFF(g7762)
--	g1392 = DFF(g6387)
--	g492 = DFF(g6359)
--	g95 = DFF(g94)
--	g944 = DFF(g6372)
--	g195 = DFF(g3831)
--	g1431 = DFF(g2673)
--	g1252 = DFF(g2661)
--	g356 = DFF(g6335)
--	g953 = DFF(g8669)
--	g1176 = DFF(g5172)
--	g1376 = DFF(g6890)
--	g1005 = DFF(g1004)
--	g1405 = DFF(g5744)
--	g901 = DFF(g896)
--	g1270 = DFF(g1271)
--	g1225 = DFF(g6858)
--	g1073 = DFF(g9145)
--	g1324 = DFF(g7118)
--	g1069 = DFF(g9134)
--	g443 = DFF(g9101)
--	g1377 = DFF(g6891)
--	g377 = DFF(g4630)
--	g618 = DFF(g6816)
--	g602 = DFF(g6800)
--	g213 = DFF(g4602)
--	g233 = DFF(g4607)
--	g1199 = DFF(g6375)
--	g1399 = DFF(g3861)
--	g83 = DFF(g6779)
--	g888 = DFF(g7100)
--	g573 = DFF(g9033)
--	g399 = DFF(g6342)
--	g1245 = DFF(g1244)
--	g507 = DFF(g9114)
--	g547 = DFF(g9026)
--	g108 = DFF(g5147)
--	g610 = DFF(g6809)
--	g630 = DFF(g6828)
--	g1207 = DFF(g5173)
--	g249 = DFF(g6320)
--	g65 = DFF(g4598)
--	g916 = DFF(g911)
--	g936 = DFF(g5168)
--	g478 = DFF(g4648)
--	g604 = DFF(g6802)
--	g945 = DFF(g5170)
--	g1114 = DFF(g7521)
--	g100 = DFF(g99)
--	g429 = DFF(g9107)
--	g809 = DFF(g7511)
--	g849 = DFF(g2645)
--	g1408 = DFF(g5177)
--	g1336 = DFF(g6864)
--	g601 = DFF(g6799)
--	g122 = DFF(g6788)
--	g1065 = DFF(g9117)
--	g1122 = DFF(g8225)
--	g1228 = DFF(g7109)
--	g495 = DFF(g6360)
--	g1322 = DFF(g7116)
--	g1230 = DFF(g7300)
--	g1033 = DFF(g9034)
--	g267 = DFF(g9091)
--	g1195 = DFF(g6374)
--	g1395 = DFF(g1393)
--	g373 = DFF(g4626)
--	g274 = DFF(g4612)
--	g1266 = DFF(g5739)
--	g714 = DFF(g7752)
--	g734 = DFF(g7755)
--	g1142 = DFF(g8874)
--	g1342 = DFF(g7119)
--	g769 = DFF(g6843)
--	g1081 = DFF(g6852)
--	g1481 = DFF(g7769)
--	g1097 = DFF(g1185)
--	g543 = DFF(g3846)
--	g1154 = DFF(g1153)
--	g1354 = DFF(g7768)
--	g489 = DFF(g6358)
--	g874 = DFF(g4654)
--	g121 = DFF(g5154)
--	g591 = DFF(g9032)
--	g616 = DFF(g6814)
--	g1267 = DFF(g4656)
--	g1312 = DFF(g1311)
--	g605 = DFF(g6803)
--	g182 = DFF(g5161)
--	g1401 = DFF(g1399)
--	g950 = DFF(g8666)
--	g1329 = DFF(g2663)
--	g408 = DFF(g6345)
--	g871 = DFF(g5167)
--	g759 = DFF(g6832)
--	g146 = DFF(g7735)
--	g202 = DFF(g5732)
--	g440 = DFF(g6349)
--	g476 = DFF(g4646)
--	g184 = DFF(g6310)
--	g1149 = DFF(g7525)
--	g1398 = DFF(g1396)
--	g210 = DFF(g3834)
--	g394 = DFF(g4632)
--	g86 = DFF(g6780)
--	g570 = DFF(g9030)
--	g275 = DFF(g6322)
--	g303 = DFF(g6326)
--	g125 = DFF(g5155)
--	g181 = DFF(g5160)
--	g1524 = DFF(g6393)
--	g595 = DFF(g576)
--	g1319 = DFF(g7113)
--	g863 = DFF(g8222)
--	g1211 = DFF(g5174)
--	g966 = DFF(g8223)
--	g1186 = DFF(g1182)
--	g1386 = DFF(g6884)
--	g875 = DFF(g5165)
--	g1170 = DFF(g1173)
--	g1370 = DFF(g6876)
--	g201 = DFF(g200)
--	g1325 = DFF(g7305)
--	g1280 = DFF(g7112)
--	g1106 = DFF(g7107)
--	g1061 = DFF(g9035)
--	g1387 = DFF(g6885)
--	g762 = DFF(g6835)
--	g1461 = DFF(g4669)
--	g378 = DFF(g6337)
--	g1200 = DFF(g1199)
--	g1514 = DFF(g7775)
--	g1403 = DFF(g1402)
--	g1345 = DFF(g7528)
--	g1191 = DFF(g6373)
--	g1391 = DFF(g1390)
--	g185 = DFF(g4599)
--	g1307 = DFF(g3858)
--	g1159 = DFF(g1157)
--	g1223 = DFF(g6379)
--	g446 = DFF(g9102)
--	g1416 = DFF(g4665)
--	g395 = DFF(g4633)
--	g764 = DFF(g6837)
--	g1251 = DFF(g6860)
--	g216 = DFF(g6311)
--	g236 = DFF(g4610)
--	g205 = DFF(g3835)
--	g540 = DFF(g6364)
--	g576 = DFF(g3849)
--	g1537 = DFF(g7777)
--	g727 = DFF(g8228)
--	g999 = DFF(g8865)
--	g761 = DFF(g6834)
--	g1272 = DFF(g6383)
--	g1243 = DFF(g2660)
--	g1328 = DFF(g7309)
--	g1130 = DFF(g7522)
--	g1330 = DFF(g6862)
--	g114 = DFF(g6786)
--	g134 = DFF(g6791)
--	g1166 = DFF(g1167)
--	g524 = DFF(g9109)
--	g1366 = DFF(g6866)
--	g348 = DFF(g9099)
--	g1148 = DFF(g1147)
--	g1348 = DFF(g7529)
--	g1155 = DFF(g1154)
--	g1260 = DFF(g6382)
--	g7 = DFF(g9375)
--	g258 = DFF(g9088)
--	g521 = DFF(g6362)
--	g300 = DFF(g6325)
--	g765 = DFF(g6838)
--	g1118 = DFF(g7766)
--	g1167 = DFF(g1170)
--	g1318 = DFF(g6861)
--	g1367 = DFF(g6873)
--	g677 = DFF(g7747)
--	g376 = DFF(g4629)
--	g1057 = DFF(g8959)
--	g973 = DFF(g8672)
--	g1193 = DFF(g1192)
--	g1393 = DFF(g2664)
--	g1549 = DFF(g7780)
--	g1321 = DFF(g7115)
--	g1253 = DFF(g5741)
--	g1519 = DFF(g8227)
--	g584 = DFF(g6369)
--	g539 = DFF(g3845)
--	g324 = DFF(g6331)
--	g432 = DFF(g9108)
--	g1158 = DFF(g1159)
--	g321 = DFF(g6330)
--	g1311 = DFF(g1310)
--	g414 = DFF(g6347)
--	g1374 = DFF(g6872)
--	g94 = DFF(g6782)
--	g1284 = DFF(g7301)
--	g1545 = DFF(g7779)
--	g1380 = DFF(g6886)
--	g673 = DFF(g7746)
--	g607 = DFF(g6805)
--	g306 = DFF(g6327)
--	g943 = DFF(g8671)
--	g162 = DFF(g7741)
--	g411 = DFF(g6346)
--	g866 = DFF(g5163)
--	g1204 = DFF(g1203)
--	g1300 = DFF(g7303)
--	g384 = DFF(g6339)
--	g339 = DFF(g9096)
--	g459 = DFF(g6350)
--	g1323 = DFF(g7117)
--	g381 = DFF(g6338)
--	g1528 = DFF(g7776)
--	g1351 = DFF(g7530)
--	g597 = DFF(g6796)
--	g1372 = DFF(g6870)
--	g154 = DFF(g7739)
--	g435 = DFF(g4637)
--	g970 = DFF(g963)
--	g1134 = DFF(g7523)
--	g995 = DFF(g7517)
--	g190 = DFF(g201)
--	g1313 = DFF(g5742)
--	g603 = DFF(g6801)
--	g1494 = DFF(g7771)
--	g462 = DFF(g6351)
--	g1160 = DFF(g1163)
--	g1360 = DFF(g8676)
--	g1450 = DFF(g5186)
--	g187 = DFF(g5730)
--	g1179 = DFF(g1186)
--	g1379 = DFF(g6879)
--	g12 = DFF(g8662)
--	g71 = DFF(g6775)
--	
--	g1658 = NOT(g1313)
--	g1777 = NOT(g611)
--	I9325 = NOT(g4242)
--	I7758 = NOT(g2605)
--	g5652 = NOT(I10135)
--	I13502 = NOT(g7135)
--	g6895 = NOT(I12558)
--	g3880 = NOT(g2965)
--	g6837 = NOT(I12382)
--	I15824 = NOT(g9157)
--	g5843 = NOT(g5367)
--	I6112 = NOT(g4)
--	g7189 = NOT(I13109)
--	g8970 = NOT(I15414)
--	I6267 = NOT(g100)
--	g6062 = NOT(I10675)
--	I16126 = NOT(g9354)
--	I10519 = NOT(g5242)
--	I15181 = NOT(g8734)
--	I11443 = NOT(g6038)
--	I12436 = NOT(g6635)
--	I10675 = NOT(g5662)
--	g2547 = NOT(I6371)
--	I7365 = NOT(g3061)
--	I10154 = NOT(g5109)
--	g1611 = NOT(g1073)
--	I11278 = NOT(g5780)
--	g7171 = NOT(g7071)
--	I14154 = NOT(g7558)
--	I12274 = NOT(g6672)
--	g8224 = NOT(I14451)
--	g5834 = NOT(I10525)
--	g5971 = NOT(I10587)
--	g3978 = NOT(g3160)
--	I6676 = NOT(g1603)
--	g3612 = NOT(I7082)
--	I8520 = NOT(g3652)
--	g2892 = NOT(g2266)
--	I13469 = NOT(g7123)
--	I12346 = NOT(g6737)
--	I9636 = NOT(g4802)
--	I14637 = NOT(g8012)
--	g6788 = NOT(I12235)
--	g1799 = NOT(I5657)
--	g3935 = NOT(I7602)
--	I5933 = NOT(g1158)
--	g9207 = NOT(g9197)
--	I13039 = NOT(g6961)
--	I15426 = NOT(g8895)
--	g5598 = NOT(g4938)
--	g1674 = NOT(g1514)
--	g7281 = NOT(I13277)
--	g3982 = NOT(g3192)
--	g4666 = NOT(I8913)
--	I15190 = NOT(g8685)
--	g2945 = NOT(g2364)
--	g5121 = NOT(I9515)
--	g3128 = NOT(I6839)
--	g3629 = NOT(g2424)
--	g7297 = NOT(I13323)
--	g5670 = NOT(I10157)
--	I11815 = NOT(g6169)
--	g6842 = NOT(I12397)
--	g3130 = NOT(I6849)
--	g9088 = NOT(I15654)
--	g8789 = NOT(g8564)
--	g3542 = NOT(g1777)
--	I12292 = NOT(g6657)
--	g6298 = NOT(I11221)
--	g2709 = NOT(g1747)
--	I11677 = NOT(g6076)
--	g6392 = NOT(I11503)
--	g4648 = NOT(I8859)
--	I8829 = NOT(g4029)
--	I15546 = NOT(g9007)
--	g1680 = NOT(I5515)
--	I15211 = NOT(g8808)
--	g2340 = NOT(g1327)
--	I12409 = NOT(g6398)
--	g4655 = NOT(I8880)
--	g7745 = NOT(I14106)
--	g7138 = NOT(I12996)
--	I6703 = NOT(g1983)
--	g5938 = NOT(g5412)
--	g8771 = NOT(g8564)
--	g2478 = NOT(g31)
--	g5813 = NOT(I10472)
--	g7338 = NOT(I13432)
--	g2907 = NOT(g2289)
--	g1744 = NOT(g600)
--	g9215 = NOT(I15921)
--	g7109 = NOT(I12915)
--	g6854 = NOT(I12433)
--	I12635 = NOT(g6509)
--	g7309 = NOT(I13359)
--	g1802 = NOT(g628)
--	I10439 = NOT(g5214)
--	g2959 = NOT(g1926)
--	I14728 = NOT(g8152)
--	I8733 = NOT(g3996)
--	I14439 = NOT(g8063)
--	g2517 = NOT(I6348)
--	g4010 = NOT(g3097)
--	I7662 = NOT(g3642)
--	I9446 = NOT(g3926)
--	I8974 = NOT(g3871)
--	g5740 = NOT(I10277)
--	g5519 = NOT(I9929)
--	g9114 = NOT(I15732)
--	g1558 = NOT(I5435)
--	I7290 = NOT(g2936)
--	g2876 = NOT(g2231)
--	g9314 = NOT(I16058)
--	I11884 = NOT(g6091)
--	I9145 = NOT(g4264)
--	I6468 = NOT(g1917)
--	g5606 = NOT(g4748)
--	I8796 = NOT(g3934)
--	g7759 = NOT(I14148)
--	I14349 = NOT(g7588)
--	I11410 = NOT(g5845)
--	I12164 = NOT(g5847)
--	g695 = NOT(I5392)
--	g6708 = NOT(g6250)
--	I13410 = NOT(g7274)
--	I15625 = NOT(g9000)
--	g6520 = NOT(I11704)
--	g1901 = NOT(I5781)
--	g6219 = NOT(I10998)
--	g6640 = NOT(I11908)
--	I8980 = NOT(g4535)
--	g3902 = NOT(I7495)
--	I12891 = NOT(g6950)
--	I11479 = NOT(g6201)
--	I11666 = NOT(g5772)
--	g5687 = NOT(I10190)
--	g2915 = NOT(I6643)
--	I13666 = NOT(g7238)
--	g6252 = NOT(g5418)
--	g6812 = NOT(I12307)
--	g4372 = NOT(I8357)
--	g7049 = NOT(I12813)
--	g3512 = NOT(g1616)
--	I13478 = NOT(g7126)
--	g5586 = NOT(g4938)
--	g6958 = NOT(I12675)
--	I15943 = NOT(g9214)
--	g4618 = NOT(I8769)
--	I6716 = NOT(g1721)
--	g6376 = NOT(I11455)
--	g4667 = NOT(I8916)
--	I5981 = NOT(g459)
--	I8177 = NOT(g2810)
--	I7847 = NOT(g3798)
--	I16055 = NOT(g9291)
--	g9336 = NOT(I16084)
--	g2310 = NOT(I6087)
--	g7715 = NOT(I14022)
--	g1600 = NOT(g976)
--	g1574 = NOT(g681)
--	g1864 = NOT(g162)
--	g4566 = NOT(g2902)
--	I11556 = NOT(g6065)
--	g7098 = NOT(g6525)
--	I5997 = NOT(g114)
--	g6829 = NOT(I12358)
--	g7498 = NOT(I13672)
--	g2663 = NOT(I6460)
--	I12108 = NOT(g5939)
--	g6765 = NOT(I12164)
--	g3529 = NOT(g2323)
--	g8959 = NOT(I15391)
--	I6198 = NOT(g483)
--	g4693 = NOT(I8974)
--	I13580 = NOT(g7208)
--	g4134 = NOT(g3676)
--	g3649 = NOT(g2424)
--	I14139 = NOT(g7548)
--	I9416 = NOT(g4273)
--	I12283 = NOT(g6692)
--	g8482 = NOT(g8094)
--	g5525 = NOT(g4934)
--	g3851 = NOT(I7356)
--	g5645 = NOT(g4748)
--	I5353 = NOT(g3833)
--	g2402 = NOT(g29)
--	I7950 = NOT(g2774)
--	g2824 = NOT(g1688)
--	g1580 = NOT(g706)
--	g2236 = NOT(I5969)
--	g7584 = NOT(I13897)
--	g4555 = NOT(g2894)
--	g9065 = NOT(I15589)
--	I9642 = NOT(g4788)
--	g7539 = NOT(I13797)
--	I15411 = NOT(g8897)
--	I15527 = NOT(g9020)
--	I10415 = NOT(g5397)
--	I13084 = NOT(g7071)
--	g9322 = NOT(g9313)
--	g3964 = NOT(g3160)
--	g4792 = NOT(I9111)
--	g9230 = NOT(I15950)
--	g6225 = NOT(I11014)
--	I8781 = NOT(g3932)
--	I8898 = NOT(g4089)
--	g6073 = NOT(g5384)
--	g2877 = NOT(g2232)
--	g6796 = NOT(I12259)
--	g1736 = NOT(I5577)
--	I12091 = NOT(g5988)
--	g4621 = NOT(I8778)
--	g5607 = NOT(g4938)
--	g9033 = NOT(I15513)
--	g7162 = NOT(I13060)
--	g7268 = NOT(I13244)
--	g7019 = NOT(I12771)
--	I11740 = NOT(g6136)
--	g7362 = NOT(I13502)
--	g5158 = NOT(I9600)
--	I13740 = NOT(g7364)
--	I9654 = NOT(g4792)
--	I15894 = NOT(g9195)
--	g6324 = NOT(I11299)
--	I7723 = NOT(g3052)
--	g4113 = NOT(I7950)
--	g6069 = NOT(I10690)
--	g2556 = NOT(g1190)
--	g1889 = NOT(g1018)
--	I7101 = NOT(g2478)
--	I5901 = NOT(g52)
--	g2222 = NOT(I5939)
--	I13676 = NOT(g7256)
--	g9096 = NOT(I15678)
--	I8291 = NOT(g878)
--	I13373 = NOT(g7270)
--	g2928 = NOT(g2326)
--	g4202 = NOT(g2810)
--	g8663 = NOT(I14783)
--	I7605 = NOT(g2752)
--	I15714 = NOT(g9077)
--	g5587 = NOT(g4938)
--	g2930 = NOT(g2328)
--	I15315 = NOT(g8738)
--	I11800 = NOT(g6164)
--	g1871 = NOT(I5754)
--	g4908 = NOT(g4088)
--	g6377 = NOT(I11458)
--	g6206 = NOT(g5639)
--	g5311 = NOT(g4938)
--	g2899 = NOT(g2272)
--	g9195 = NOT(I15871)
--	g4094 = NOT(I7905)
--	I11936 = NOT(g5918)
--	g3872 = NOT(g2954)
--	I15202 = NOT(g8797)
--	g3652 = NOT(I7132)
--	g4567 = NOT(g2903)
--	g7728 = NOT(I14055)
--	g7486 = NOT(I13646)
--	g3843 = NOT(I7332)
--	g3989 = NOT(g3131)
--	I6186 = NOT(g138)
--	g7730 = NOT(I14061)
--	I9612 = NOT(g4776)
--	I10608 = NOT(g5701)
--	g5174 = NOT(I9648)
--	g8762 = NOT(g8585)
--	g7504 = NOT(I13692)
--	I15978 = NOT(g9235)
--	I14115 = NOT(g7563)
--	g7185 = NOT(I13099)
--	g4776 = NOT(I9081)
--	I7041 = NOT(g2401)
--	g6849 = NOT(I12418)
--	I9935 = NOT(g4812)
--	g4593 = NOT(g2939)
--	I11964 = NOT(g5971)
--	g3549 = NOT(g2404)
--	g3834 = NOT(I7305)
--	g3971 = NOT(I7688)
--	g7070 = NOT(g6562)
--	g2295 = NOT(g995)
--	I14052 = NOT(g7494)
--	g2237 = NOT(I5972)
--	g7470 = NOT(g7253)
--	I15741 = NOT(g9083)
--	g8657 = NOT(I14763)
--	g6781 = NOT(I12214)
--	g7425 = NOT(I13550)
--	g5180 = NOT(I9666)
--	g2844 = NOT(I6574)
--	I8215 = NOT(g3577)
--	g6898 = NOT(I12567)
--	g1838 = NOT(g1450)
--	g5591 = NOT(g4841)
--	g6900 = NOT(I12571)
--	g8222 = NOT(I14445)
--	I8886 = NOT(g4308)
--	g5832 = NOT(I10519)
--	I14813 = NOT(g8640)
--	g1795 = NOT(I5649)
--	g6797 = NOT(I12262)
--	g1737 = NOT(g597)
--	g2394 = NOT(I6270)
--	g9248 = NOT(I15978)
--	g1809 = NOT(g759)
--	I10973 = NOT(g5726)
--	I14798 = NOT(g8605)
--	g6245 = NOT(g5690)
--	g4360 = NOT(I8333)
--	I7368 = NOT(g3018)
--	g9255 = NOT(I15985)
--	g9081 = NOT(I15635)
--	I12948 = NOT(g6919)
--	I13909 = NOT(g7339)
--	I15735 = NOT(g9078)
--	g4521 = NOT(g2866)
--	I14184 = NOT(g7726)
--	g1672 = NOT(g1499)
--	I14674 = NOT(g7788)
--	g8464 = NOT(g8039)
--	g6291 = NOT(I11200)
--	I12702 = NOT(g6497)
--	g2557 = NOT(g940)
--	g4050 = NOT(g3080)
--	g4641 = NOT(I8838)
--	I11908 = NOT(g5918)
--	I12757 = NOT(g6577)
--	g9097 = NOT(I15681)
--	g2966 = NOT(g1856)
--	g5794 = NOT(I10421)
--	I5889 = NOT(g83)
--	g1643 = NOT(g1211)
--	I11569 = NOT(g6279)
--	g7131 = NOT(g6976)
--	g6344 = NOT(I11359)
--	g2471 = NOT(I6309)
--	g7006 = NOT(I12748)
--	g7331 = NOT(I13413)
--	I15196 = NOT(g8778)
--	I6636 = NOT(g1704)
--	I14732 = NOT(g8155)
--	g2242 = NOT(g985)
--	g6207 = NOT(I10962)
--	g3909 = NOT(I7520)
--	I11747 = NOT(g6123)
--	I12564 = NOT(g6720)
--	g8563 = NOT(I14662)
--	g2948 = NOT(g2366)
--	I11242 = NOT(g6183)
--	g7766 = NOT(I14169)
--	g6819 = NOT(I12328)
--	g7105 = NOT(I12903)
--	g3519 = NOT(g2185)
--	I10761 = NOT(g5302)
--	g7305 = NOT(I13347)
--	I7856 = NOT(g3805)
--	I7734 = NOT(g2595)
--	g2955 = NOT(I6703)
--	g7487 = NOT(I13649)
--	g5628 = NOT(g4748)
--	g1742 = NOT(g1486)
--	g6088 = NOT(I10708)
--	g6852 = NOT(I12427)
--	g5515 = NOT(g4923)
--	I12397 = NOT(g6764)
--	g6488 = NOT(I11652)
--	g4658 = NOT(I8889)
--	g7748 = NOT(I14115)
--	g4777 = NOT(I9084)
--	I10400 = NOT(g5201)
--	g5100 = NOT(I9484)
--	I9512 = NOT(g3985)
--	I13807 = NOT(g7320)
--	I11974 = NOT(g5956)
--	I12062 = NOT(g5988)
--	I14400 = NOT(g7677)
--	g2350 = NOT(I6166)
--	g9112 = NOT(I15726)
--	g7755 = NOT(I14136)
--	g9218 = NOT(I15930)
--	g1926 = NOT(g874)
--	I9823 = NOT(g5138)
--	g9312 = NOT(I16052)
--	g2038 = NOT(g809)
--	g4882 = NOT(g4069)
--	I14214 = NOT(g7576)
--	I12933 = NOT(g7018)
--	I9366 = NOT(g4350)
--	g7226 = NOT(g6937)
--	I11230 = NOT(g6140)
--	I11293 = NOT(g5824)
--	I10207 = NOT(g5075)
--	I13293 = NOT(g7159)
--	I12508 = NOT(g6593)
--	I11638 = NOT(g5847)
--	g6886 = NOT(I12529)
--	I6446 = NOT(g1812)
--	g4611 = NOT(I8748)
--	g291 = NOT(I5356)
--	I14005 = NOT(g7434)
--	g7045 = NOT(g6490)
--	I11416 = NOT(g5829)
--	I10538 = NOT(g5255)
--	I6003 = NOT(g228)
--	I9148 = NOT(g4354)
--	I13416 = NOT(g7165)
--	I5795 = NOT(g1236)
--	g9129 = NOT(I15765)
--	g2769 = NOT(g2424)
--	g7173 = NOT(g6980)
--	g9329 = NOT(g9317)
--	g6314 = NOT(I11269)
--	g7091 = NOT(g6525)
--	g7491 = NOT(I13653)
--	g6870 = NOT(I12481)
--	g3860 = NOT(I7383)
--	g2918 = NOT(g2310)
--	g3341 = NOT(I6936)
--	g1983 = NOT(I5839)
--	g6825 = NOT(I12346)
--	g6650 = NOT(g6213)
--	g7169 = NOT(I13075)
--	g7283 = NOT(I13281)
--	g1572 = NOT(g673)
--	g8955 = NOT(I15379)
--	I6695 = NOT(g2246)
--	g4541 = NOT(g2883)
--	g7059 = NOT(g6538)
--	g7920 = NOT(I14282)
--	g7578 = NOT(I13879)
--	g6008 = NOT(g5367)
--	I11835 = NOT(g6181)
--	g3691 = NOT(I7195)
--	I11014 = NOT(g5621)
--	g7459 = NOT(I13617)
--	g9221 = NOT(I15937)
--	I12205 = NOT(g6488)
--	I9463 = NOT(g3942)
--	g7718 = NOT(I14031)
--	g7767 = NOT(I14172)
--	g4153 = NOT(I8024)
--	g4680 = NOT(I8945)
--	I7688 = NOT(g3650)
--	g6136 = NOT(I10773)
--	g4353 = NOT(g3665)
--	I11586 = NOT(g6256)
--	I12912 = NOT(g7006)
--	g6336 = NOT(I11335)
--	I14100 = NOT(g7580)
--	I6223 = NOT(g330)
--	g8038 = NOT(g7694)
--	g6768 = NOT(I12173)
--	I8913 = NOT(g4306)
--	g7582 = NOT(I13891)
--	g6594 = NOT(I11796)
--	g1961 = NOT(g1345)
--	g3879 = NOT(g2963)
--	g4802 = NOT(I9129)
--	g7261 = NOT(I13225)
--	I14683 = NOT(g7825)
--	g3962 = NOT(g3131)
--	g5151 = NOT(I9579)
--	g7793 = NOT(I14234)
--	g3158 = NOT(I6853)
--	g3659 = NOT(g2293)
--	g6806 = NOT(I12289)
--	g5648 = NOT(g4748)
--	I6416 = NOT(g1794)
--	g3506 = NOT(g1781)
--	g7015 = NOT(I12763)
--	I12592 = NOT(g1008)
--	g4558 = NOT(g2897)
--	g9068 = NOT(I15598)
--	I7126 = NOT(g2494)
--	I5926 = NOT(g297)
--	I7400 = NOT(g3075)
--	I8859 = NOT(g3968)
--	I7326 = NOT(g2940)
--	I6115 = NOT(g134)
--	I6251 = NOT(g489)
--	g2921 = NOT(g2312)
--	g6065 = NOT(I10684)
--	g6887 = NOT(I12532)
--	g6122 = NOT(I10752)
--	I10882 = NOT(g5600)
--	g6228 = NOT(I11021)
--	I5754 = NOT(g966)
--	g3587 = NOT(g1964)
--	g6322 = NOT(I11293)
--	I11275 = NOT(g5768)
--	I9457 = NOT(g3940)
--	g8918 = NOT(I15340)
--	I16180 = NOT(g9387)
--	g6230 = NOT(I11025)
--	g7246 = NOT(I13196)
--	g8967 = NOT(I15405)
--	I13746 = NOT(g7311)
--	I13493 = NOT(g7132)
--	I9393 = NOT(g4266)
--	g4511 = NOT(g2841)
--	I15660 = NOT(g9062)
--	g2895 = NOT(g2268)
--	g6033 = NOT(g5384)
--	g2837 = NOT(g1780)
--	g7721 = NOT(g7344)
--	g5839 = NOT(I10532)
--	I9834 = NOT(g4782)
--	g4092 = NOT(I7899)
--	I13035 = NOT(g6964)
--	g3985 = NOT(I7712)
--	I12731 = NOT(g6579)
--	I11806 = NOT(g6275)
--	g4600 = NOT(I8715)
--	I7383 = NOT(g3465)
--	g4574 = NOT(g3466)
--	g6096 = NOT(g5317)
--	g6496 = NOT(I11662)
--	g1679 = NOT(I5512)
--	I8097 = NOT(g3237)
--	g5172 = NOT(I9642)
--	g5278 = NOT(I9794)
--	g6845 = NOT(I12406)
--	g7502 = NOT(I13682)
--	I15550 = NOT(g9008)
--	g9198 = NOT(g9187)
--	g3545 = NOT(g2344)
--	I8354 = NOT(g1163)
--	g738 = NOT(I5404)
--	g6195 = NOT(I10940)
--	g5618 = NOT(g5015)
--	g6137 = NOT(I10776)
--	g6891 = NOT(I12544)
--	g5143 = NOT(I9555)
--	g1831 = NOT(g689)
--	g6337 = NOT(I11338)
--	g3591 = NOT(g1789)
--	g3832 = NOT(I7299)
--	g4580 = NOT(g2919)
--	g9241 = NOT(I15971)
--	I7588 = NOT(g2584)
--	g3853 = NOT(I7362)
--	I14725 = NOT(g8145)
--	g7188 = NOT(I13106)
--	g5988 = NOT(I10592)
--	g2842 = NOT(g2209)
--	I9938 = NOT(g4878)
--	I10758 = NOT(g5662)
--	g1805 = NOT(I5667)
--	g6807 = NOT(I12292)
--	g1916 = NOT(g775)
--	g5693 = NOT(I10204)
--	g7216 = NOT(I13152)
--	g1749 = NOT(g371)
--	g2298 = NOT(I6072)
--	I14082 = NOT(g7539)
--	g6859 = NOT(I12448)
--	g2392 = NOT(g11)
--	I13193 = NOT(g7007)
--	g2485 = NOT(g62)
--	I11362 = NOT(g5821)
--	g7028 = NOT(g6525)
--	I13362 = NOT(g7265)
--	g3931 = NOT(I7592)
--	I8218 = NOT(g3002)
--	I15773 = NOT(g9126)
--	I6629 = NOT(g2052)
--	g4623 = NOT(I8784)
--	g7247 = NOT(I13199)
--	g1798 = NOT(I5654)
--	I6130 = NOT(g560)
--	g4076 = NOT(I7859)
--	g9319 = NOT(g9309)
--	I10940 = NOT(g5489)
--	g2941 = NOT(g2349)
--	I9606 = NOT(g4687)
--	g6342 = NOT(I11353)
--	g3905 = NOT(g3192)
--	I13475 = NOT(g7125)
--	g5621 = NOT(g4748)
--	I14848 = NOT(g8625)
--	g6255 = NOT(I11066)
--	g6815 = NOT(I12316)
--	I10804 = NOT(g5526)
--	I6800 = NOT(g2016)
--	I9687 = NOT(g4822)
--	g3630 = NOT(I7095)
--	g6481 = NOT(I11641)
--	I14804 = NOT(g8563)
--	g7741 = NOT(I14094)
--	g4651 = NOT(I8868)
--	g5113 = NOT(I9499)
--	g6692 = NOT(I12008)
--	g6097 = NOT(g5345)
--	I11437 = NOT(g5801)
--	I15839 = NOT(g9168)
--	g2520 = NOT(g41)
--	I15930 = NOT(g9209)
--	g2640 = NOT(g1584)
--	g9211 = NOT(I15909)
--	g6354 = NOT(I11389)
--	g4285 = NOT(I8233)
--	I8727 = NOT(g3944)
--	g9186 = NOT(I15836)
--	I5679 = NOT(g911)
--	g4500 = NOT(g2832)
--	g9386 = NOT(I16176)
--	g6960 = NOT(I12681)
--	I15965 = NOT(g9219)
--	I7944 = NOT(g3774)
--	g1579 = NOT(g703)
--	g1869 = NOT(g74)
--	g7108 = NOT(I12912)
--	I10135 = NOT(g4960)
--	g7308 = NOT(I13356)
--	I11347 = NOT(g5761)
--	g2958 = NOT(g2377)
--	I13347 = NOT(g7224)
--	g9026 = NOT(I15492)
--	I5831 = NOT(g1194)
--	g2376 = NOT(I6226)
--	g5494 = NOT(I9918)
--	g3750 = NOT(g2177)
--	I9570 = NOT(g4696)
--	I10406 = NOT(g5203)
--	I9341 = NOT(g4251)
--	I10962 = NOT(g5719)
--	g1752 = NOT(g603)
--	I14406 = NOT(g7681)
--	g3973 = NOT(g3097)
--	I9525 = NOT(g4413)
--	I11781 = NOT(g6284)
--	I12768 = NOT(g6718)
--	I15619 = NOT(g8998)
--	g9370 = NOT(I16138)
--	g1917 = NOT(I5795)
--	I9645 = NOT(g4900)
--	I15557 = NOT(g9010)
--	g2829 = NOT(g1785)
--	g9125 = NOT(I15753)
--	g4024 = NOT(g3160)
--	I11236 = NOT(g6148)
--	g2286 = NOT(I6042)
--	g6783 = NOT(I12220)
--	g7758 = NOT(I14145)
--	g7066 = NOT(I12839)
--	I10500 = NOT(g5234)
--	I16168 = NOT(g9381)
--	g7589 = NOT(I13912)
--	I6090 = NOT(g390)
--	g2911 = NOT(g2292)
--	g4795 = NOT(I9116)
--	I8932 = NOT(g4096)
--	I5422 = NOT(g1234)
--	g7466 = NOT(I13622)
--	g4809 = NOT(I9148)
--	g6267 = NOT(I11086)
--	g6312 = NOT(I11263)
--	g3969 = NOT(g3192)
--	I6166 = NOT(g480)
--	I14049 = NOT(g7493)
--	g9280 = NOT(I16006)
--	I11821 = NOT(g6170)
--	I12881 = NOT(g6478)
--	g1786 = NOT(g623)
--	g7365 = NOT(I13509)
--	g7048 = NOT(I12810)
--	I7347 = NOT(g2985)
--	g9083 = NOT(I15641)
--	g2270 = NOT(I6015)
--	g4477 = NOT(I8517)
--	g7448 = NOT(I13605)
--	I13063 = NOT(g6973)
--	g7711 = NOT(I14012)
--	g4523 = NOT(g2868)
--	g6676 = NOT(I11984)
--	I11790 = NOT(g6282)
--	g6293 = NOT(I11206)
--	I13264 = NOT(g7061)
--	I6148 = NOT(g5)
--	g7055 = NOT(g6517)
--	g8219 = NOT(I14436)
--	g4643 = NOT(I8844)
--	g3666 = NOT(g2134)
--	I9158 = NOT(g4256)
--	I13137 = NOT(g7027)
--	I6348 = NOT(g1354)
--	g2225 = NOT(I5948)
--	g6129 = NOT(I10758)
--	g8640 = NOT(I14728)
--	g7455 = NOT(I13613)
--	g6329 = NOT(I11314)
--	g6761 = NOT(I12154)
--	g2073 = NOT(g1254)
--	g5160 = NOT(I9606)
--	g7133 = NOT(I12983)
--	I7697 = NOT(g3052)
--	g9106 = NOT(I15708)
--	g7333 = NOT(I13419)
--	I13873 = NOT(g7342)
--	g9306 = NOT(I16036)
--	g6828 = NOT(I12355)
--	g1770 = NOT(g606)
--	g7774 = NOT(I14193)
--	g5521 = NOT(g4929)
--	g8958 = NOT(I15388)
--	g6830 = NOT(I12361)
--	g4634 = NOT(I8817)
--	g3648 = NOT(g2424)
--	g3875 = NOT(g2958)
--	g2324 = NOT(I6115)
--	g3530 = NOT(g2185)
--	I9111 = NOT(g4232)
--	g7196 = NOT(I13122)
--	g4742 = NOT(I9064)
--	g9061 = NOT(I15577)
--	I15601 = NOT(g8992)
--	g9187 = NOT(I15839)
--	g4104 = NOT(I7925)
--	I10605 = NOT(g5440)
--	I11422 = NOT(g5842)
--	g6592 = NOT(I11790)
--	g3655 = NOT(g1844)
--	I15187 = NOT(g8682)
--	I14273 = NOT(g7631)
--	I11209 = NOT(g6139)
--	I13422 = NOT(g7131)
--	I14106 = NOT(g7586)
--	I13209 = NOT(g6912)
--	g2540 = NOT(g1339)
--	I9615 = NOT(g4739)
--	g6221 = NOT(I11004)
--	I12003 = NOT(g6202)
--	g8765 = NOT(g8524)
--	g7538 = NOT(I13794)
--	I13834 = NOT(g7466)
--	I6463 = NOT(g1769)
--	I10463 = NOT(g5220)
--	I16084 = NOT(g9324)
--	g2177 = NOT(g1322)
--	g7780 = NOT(I14211)
--	g9027 = NOT(I15495)
--	g5724 = NOT(g4969)
--	g2377 = NOT(I6229)
--	I14463 = NOT(g8072)
--	I12779 = NOT(g6740)
--	g5179 = NOT(I9663)
--	g6703 = NOT(I12041)
--	g7509 = NOT(I13707)
--	g4926 = NOT(g4202)
--	I15937 = NOT(g9212)
--	g9200 = NOT(g9189)
--	I11021 = NOT(g5627)
--	I14234 = NOT(g7614)
--	g3884 = NOT(I7417)
--	g3839 = NOT(I7320)
--	g2287 = NOT(I6045)
--	g7018 = NOT(I12768)
--	g4273 = NOT(I8215)
--	g7067 = NOT(g6658)
--	g8974 = NOT(I15426)
--	I7317 = NOT(g2893)
--	g5658 = NOT(g4748)
--	I15791 = NOT(g9140)
--	g7418 = NOT(I13533)
--	g6624 = NOT(I11864)
--	g7467 = NOT(g7236)
--	g6953 = NOT(g6745)
--	I6118 = NOT(g243)
--	I14795 = NOT(g8604)
--	g8225 = NOT(I14454)
--	g5835 = NOT(I10528)
--	g7290 = NOT(I13302)
--	g4613 = NOT(I8754)
--	g6068 = NOT(I10687)
--	g1888 = NOT(g781)
--	I6872 = NOT(g2185)
--	g9145 = NOT(I15791)
--	g4044 = NOT(g2595)
--	g6468 = NOT(I11622)
--	I12945 = NOT(g7066)
--	I9591 = NOT(g4710)
--	g4444 = NOT(I8452)
--	g1787 = NOT(g625)
--	I6652 = NOT(g2016)
--	I11607 = NOT(g5767)
--	I6057 = NOT(g518)
--	I12826 = NOT(g6441)
--	I12999 = NOT(g7029)
--	I11320 = NOT(g5797)
--	I15666 = NOT(g9070)
--	I13320 = NOT(g7139)
--	I6457 = NOT(g1886)
--	g7493 = NOT(I13659)
--	g1675 = NOT(g1519)
--	g6677 = NOT(I11987)
--	g7256 = NOT(g7058)
--	I13274 = NOT(g6917)
--	I7775 = NOT(g3705)
--	g5611 = NOT(g4969)
--	g8324 = NOT(I14573)
--	g4572 = NOT(g2909)
--	I7922 = NOT(g3462)
--	g2898 = NOT(g2271)
--	I15478 = NOT(g8910)
--	g2900 = NOT(g2273)
--	g6866 = NOT(I12469)
--	I12672 = NOT(g6473)
--	I7581 = NOT(g3612)
--	I13122 = NOT(g7070)
--	g9107 = NOT(I15711)
--	g4543 = NOT(g2885)
--	I10421 = NOT(g5208)
--	I11464 = NOT(g6088)
--	g5799 = NOT(I10436)
--	I13565 = NOT(g7181)
--	I9794 = NOT(g4778)
--	I6834 = NOT(g287)
--	g9307 = NOT(g9300)
--	g2510 = NOT(g58)
--	g639 = NOT(I5374)
--	g2245 = NOT(g999)
--	g6149 = NOT(I10810)
--	g3988 = NOT(g3097)
--	I6686 = NOT(g2246)
--	g6349 = NOT(I11374)
--	g5674 = NOT(g5042)
--	g8177 = NOT(I14410)
--	g3693 = NOT(g2424)
--	I11034 = NOT(g5644)
--	g9223 = NOT(I15943)
--	I14163 = NOT(g7533)
--	g2291 = NOT(I6057)
--	I14012 = NOT(g7438)
--	I11641 = NOT(g5918)
--	g6848 = NOT(I12415)
--	I15580 = NOT(g8985)
--	I13797 = NOT(g7502)
--	I12331 = NOT(g6704)
--	g5541 = NOT(g4814)
--	g3548 = NOT(g2185)
--	g1684 = NOT(g1)
--	g1745 = NOT(g746)
--	g6198 = NOT(g5335)
--	g1639 = NOT(g1207)
--	g2344 = NOT(I6148)
--	g6855 = NOT(I12436)
--	g6398 = NOT(I11515)
--	I10541 = NOT(g5256)
--	I6121 = NOT(g321)
--	g7263 = NOT(I13231)
--	g2207 = NOT(I5920)
--	g5153 = NOT(I9585)
--	g5680 = NOT(g5101)
--	I12897 = NOT(g6962)
--	I12448 = NOT(g6569)
--	I12961 = NOT(g6921)
--	I9515 = NOT(g4301)
--	I9630 = NOT(g4867)
--	I14789 = NOT(g8544)
--	g2259 = NOT(g1325)
--	g9115 = NOT(I15735)
--	g4014 = NOT(I7769)
--	I7079 = NOT(g2532)
--	I12505 = NOT(g6612)
--	g9315 = NOT(I16061)
--	g1808 = NOT(g629)
--	g4885 = NOT(g4070)
--	I13635 = NOT(g7243)
--	g5744 = NOT(I10289)
--	g8199 = NOT(I14424)
--	g9047 = NOT(I15543)
--	g5802 = NOT(I10445)
--	g4660 = NOT(I8895)
--	g2923 = NOT(I6657)
--	I12717 = NOT(g6543)
--	g1707 = NOT(g955)
--	I14325 = NOT(g7713)
--	I10829 = NOT(g5224)
--	g8781 = NOT(g8585)
--	I10535 = NOT(g5254)
--	I5389 = NOT(g690)
--	I5706 = NOT(g901)
--	g8898 = NOT(I15308)
--	g4903 = NOT(g4084)
--	g7562 = NOT(I13858)
--	I15178 = NOT(g8753)
--	I10946 = NOT(g5563)
--	g8797 = NOT(I15003)
--	g6524 = NOT(I11710)
--	I14828 = NOT(g8639)
--	g6644 = NOT(g6208)
--	g8510 = NOT(I14643)
--	I13164 = NOT(g7086)
--	I5371 = NOT(g633)
--	g7723 = NOT(I14042)
--	I14121 = NOT(g7587)
--	g2215 = NOT(g1416)
--	I15953 = NOT(g9215)
--	g6319 = NOT(I11284)
--	g7101 = NOT(I12891)
--	g2886 = NOT(g2240)
--	g3908 = NOT(I7517)
--	g7301 = NOT(I13335)
--	I7356 = NOT(g2843)
--	I13891 = NOT(g7336)
--	I15654 = NOT(g9057)
--	g4036 = NOT(g3192)
--	g6152 = NOT(I10815)
--	g6258 = NOT(g5427)
--	g6352 = NOT(I11383)
--	g6818 = NOT(I12325)
--	g1575 = NOT(g685)
--	g1865 = NOT(g1013)
--	I8483 = NOT(g3641)
--	g6867 = NOT(I12472)
--	g3567 = NOT(g2407)
--	I15417 = NOT(g8893)
--	g1715 = NOT(I5559)
--	g2314 = NOT(I6099)
--	I9440 = NOT(g4285)
--	I14291 = NOT(g7680)
--	I12433 = NOT(g6632)
--	g4335 = NOT(g3659)
--	I9123 = NOT(g4455)
--	I15334 = NOT(g8800)
--	g7751 = NOT(I14124)
--	g2870 = NOT(g2225)
--	g5492 = NOT(g4919)
--	I12148 = NOT(g5988)
--	I13109 = NOT(g7059)
--	g4382 = NOT(I8373)
--	g1833 = NOT(g770)
--	g5600 = NOT(g5128)
--	I13537 = NOT(g7152)
--	g5574 = NOT(g4969)
--	I8790 = NOT(g4020)
--	g6211 = NOT(g5645)
--	g2825 = NOT(I6553)
--	g2650 = NOT(I6434)
--	g6186 = NOT(I10919)
--	g6386 = NOT(I11485)
--	I12646 = NOT(g6493)
--	g7585 = NOT(I13900)
--	g9017 = NOT(I15475)
--	I9666 = NOT(g4931)
--	I15762 = NOT(g9039)
--	I12343 = NOT(g6731)
--	g4805 = NOT(I9136)
--	g6975 = NOT(I12712)
--	g4916 = NOT(g4202)
--	g4022 = NOT(I7785)
--	g3965 = NOT(I7676)
--	I5963 = NOT(g225)
--	g1584 = NOT(g738)
--	g6599 = NOT(I11809)
--	g1896 = NOT(g86)
--	g7441 = NOT(I13580)
--	I15423 = NOT(g8894)
--	g6026 = NOT(g5384)
--	I9528 = NOT(g4006)
--	g6426 = NOT(I11559)
--	I6860 = NOT(g2185)
--	g3264 = NOT(I6900)
--	I7053 = NOT(g2452)
--	I6341 = NOT(g1351)
--	I10506 = NOT(g5236)
--	g5580 = NOT(g4938)
--	I9648 = NOT(g4795)
--	g9234 = NOT(I15956)
--	I10028 = NOT(g4825)
--	g9128 = NOT(I15762)
--	g6614 = NOT(I11838)
--	g6370 = NOT(I11437)
--	I14028 = NOT(g7501)
--	g3933 = NOT(g3131)
--	I8904 = NOT(g4126)
--	g9330 = NOT(g9319)
--	g6325 = NOT(I11302)
--	g6821 = NOT(I12334)
--	g3521 = NOT(g2185)
--	g4560 = NOT(g2899)
--	I8446 = NOT(g3014)
--	g3050 = NOT(I6788)
--	g3641 = NOT(I7115)
--	I15909 = NOT(g9201)
--	I15543 = NOT(g9006)
--	g5736 = NOT(I10265)
--	g2943 = NOT(g2362)
--	g6984 = NOT(I12725)
--	g7168 = NOT(I13072)
--	g6939 = NOT(g6543)
--	g3996 = NOT(I7731)
--	I11796 = NOT(g6287)
--	I12412 = NOT(g6404)
--	I8841 = NOT(g3979)
--	g5623 = NOT(g4969)
--	g7772 = NOT(I14187)
--	g6083 = NOT(I10702)
--	g7058 = NOT(g6649)
--	I5957 = NOT(g110)
--	g2887 = NOT(g2241)
--	g4873 = NOT(I9217)
--	g4632 = NOT(I8811)
--	g7531 = NOT(I13773)
--	g4095 = NOT(I7908)
--	g5076 = NOT(I9446)
--	g8870 = NOT(I15196)
--	I8763 = NOT(g3947)
--	g4037 = NOT(g2845)
--	g6483 = NOT(I11645)
--	I12229 = NOT(g6659)
--	I9884 = NOT(g4868)
--	g2934 = NOT(I6676)
--	g5476 = NOT(g4907)
--	g7743 = NOT(I14100)
--	g4653 = NOT(I8874)
--	I6358 = NOT(g13)
--	g4102 = NOT(I7919)
--	g6636 = NOT(I11900)
--	I15568 = NOT(g8981)
--	I15747 = NOT(g9042)
--	I5865 = NOT(g1206)
--	g9213 = NOT(I15915)
--	g6106 = NOT(g5345)
--	g5175 = NOT(I9651)
--	g4579 = NOT(g2918)
--	I10649 = NOT(g5657)
--	I12011 = NOT(g5939)
--	g6306 = NOT(I11245)
--	I5715 = NOT(g896)
--	g7505 = NOT(I13695)
--	g5871 = NOT(I10558)
--	g3878 = NOT(g2962)
--	g8008 = NOT(g7559)
--	g4719 = NOT(I9021)
--	g6790 = NOT(I12241)
--	g7734 = NOT(I14073)
--	I6587 = NOT(g1708)
--	g3777 = NOT(g2170)
--	g7411 = NOT(g7202)
--	I9372 = NOT(g3902)
--	I10491 = NOT(g5231)
--	I15814 = NOT(g9154)
--	g3835 = NOT(I7308)
--	I16116 = NOT(g9350)
--	g6387 = NOT(I11488)
--	I11522 = NOT(g5847)
--	g2096 = NOT(g1226)
--	I9618 = NOT(g4742)
--	I12582 = NOT(g6745)
--	g5285 = NOT(g4841)
--	g6461 = NOT(I11607)
--	g8768 = NOT(g8585)
--	I13663 = NOT(g7235)
--	g3882 = NOT(g2970)
--	g2496 = NOT(g942)
--	I7626 = NOT(g3632)
--	g4917 = NOT(g4102)
--	I15974 = NOT(g9234)
--	I6615 = NOT(g1983)
--	g6756 = NOT(I12141)
--	g8972 = NOT(I15420)
--	I10770 = NOT(g5441)
--	I12310 = NOT(g6723)
--	g1897 = NOT(g789)
--	g9090 = NOT(I15660)
--	g6622 = NOT(I11858)
--	g7474 = NOT(I13628)
--	I8757 = NOT(g3921)
--	g6027 = NOT(g5384)
--	g7992 = NOT(g7557)
--	g4265 = NOT(g3591)
--	g3611 = NOT(I7079)
--	g6427 = NOT(I11562)
--	g2137 = NOT(I5889)
--	g2891 = NOT(g2265)
--	g5184 = NOT(I9678)
--	I15638 = NOT(g8978)
--	g9366 = NOT(I16126)
--	g2913 = NOT(g2307)
--	I12379 = NOT(g6768)
--	g5139 = NOT(I9543)
--	g5384 = NOT(I9837)
--	g6904 = NOT(g6426)
--	I12958 = NOT(g6920)
--	g9056 = NOT(I15562)
--	g8065 = NOT(I14338)
--	I8315 = NOT(g3691)
--	I8811 = NOT(g4022)
--	g6446 = NOT(I11591)
--	g8228 = NOT(I14463)
--	g3981 = NOT(I7706)
--	g5024 = NOT(I9360)
--	g6514 = NOT(I11696)
--	I6239 = NOT(g8)
--	g3674 = NOT(I7164)
--	g2807 = NOT(g1782)
--	I5362 = NOT(g3841)
--	I11326 = NOT(g5819)
--	I9555 = NOT(g4892)
--	g5795 = NOT(I10424)
--	g5737 = NOT(I10268)
--	I15391 = NOT(g8917)
--	g6403 = NOT(I11522)
--	I13326 = NOT(g7176)
--	g5809 = NOT(I10460)
--	I5419 = NOT(g1603)
--	I9804 = NOT(g5113)
--	I10262 = NOT(g5551)
--	I7683 = NOT(g2573)
--	g3997 = NOT(I7734)
--	I12742 = NOT(g6590)
--	g6345 = NOT(I11362)
--	g6841 = NOT(I12394)
--	I15510 = NOT(g8969)
--	I11040 = NOT(g5299)
--	I11948 = NOT(g5897)
--	I8874 = NOT(g3884)
--	g2266 = NOT(I6003)
--	g6763 = NOT(I12158)
--	I7778 = NOT(g3019)
--	I16142 = NOT(g9366)
--	g6391 = NOT(I11500)
--	g1006 = NOT(I5410)
--	g4296 = NOT(g3790)
--	I6853 = NOT(g2185)
--	g3238 = NOT(I6894)
--	I9621 = NOT(g4732)
--	g5477 = NOT(g4908)
--	g9260 = NOT(I15990)
--	g5523 = NOT(I9935)
--	I12681 = NOT(g6469)
--	I10719 = NOT(g5559)
--	g6637 = NOT(I11903)
--	g5643 = NOT(I10128)
--	I15014 = NOT(g8607)
--	g1801 = NOT(g618)
--	g4553 = NOT(g2891)
--	g9063 = NOT(I15583)
--	g6307 = NOT(I11248)
--	I15586 = NOT(g8987)
--	I15007 = NOT(g8627)
--	I8880 = NOT(g4303)
--	I14718 = NOT(g8068)
--	g3802 = NOT(g1832)
--	g7688 = NOT(g7406)
--	g6359 = NOT(I11404)
--	g6223 = NOT(I11008)
--	g2481 = NOT(I6317)
--	g8913 = NOT(I15329)
--	g1748 = NOT(g601)
--	g2692 = NOT(g1671)
--	g4012 = NOT(I7765)
--	g6858 = NOT(I12445)
--	g5742 = NOT(I10283)
--	g5551 = NOT(I9974)
--	g5099 = NOT(g4477)
--	g2497 = NOT(g945)
--	I12690 = NOT(g6467)
--	g2354 = NOT(I6178)
--	I16165 = NOT(g9377)
--	g2960 = NOT(g2381)
--	g4706 = NOT(I9005)
--	I9567 = NOT(g4693)
--	I7526 = NOT(g2752)
--	I5897 = NOT(g173)
--	I14573 = NOT(g8179)
--	I10247 = NOT(g5266)
--	g3901 = NOT(I7492)
--	g7000 = NOT(I12742)
--	I13509 = NOT(g7137)
--	I15720 = NOT(g9053)
--	g9318 = NOT(g9304)
--	g9367 = NOT(I16129)
--	I11933 = NOT(g5847)
--	g7126 = NOT(I12968)
--	I8935 = NOT(g4005)
--	I5425 = NOT(g1245)
--	g4029 = NOT(I7800)
--	g6251 = NOT(I11060)
--	g6315 = NOT(I11272)
--	g6811 = NOT(I12304)
--	g6642 = NOT(I11912)
--	g4371 = NOT(I8354)
--	I11851 = NOT(g6277)
--	g3511 = NOT(g1616)
--	g5754 = NOT(g5403)
--	g9057 = NOT(I15565)
--	I16006 = NOT(g9261)
--	g7760 = NOT(I14151)
--	I14388 = NOT(g7605)
--	I7850 = NOT(g2795)
--	g9193 = NOT(g9181)
--	g3092 = NOT(I6826)
--	I14777 = NOT(g8511)
--	g3492 = NOT(I6970)
--	g4281 = NOT(g2562)
--	g6874 = NOT(I12493)
--	g5613 = NOT(g4748)
--	I14251 = NOT(g7541)
--	g3574 = NOT(g1771)
--	g3864 = NOT(g2943)
--	g8342 = NOT(g8008)
--	I15340 = NOT(g8856)
--	g2267 = NOT(I6006)
--	g2312 = NOT(I6093)
--	g6654 = NOT(I11942)
--	g5444 = NOT(g5074)
--	g5269 = NOT(I9791)
--	I7702 = NOT(g3062)
--	I15684 = NOT(g9067)
--	g8481 = NOT(I14637)
--	I12128 = NOT(g5897)
--	g1578 = NOT(g699)
--	g1868 = NOT(I5747)
--	I9360 = NOT(g4257)
--	g2401 = NOT(g22)
--	I7919 = NOT(g3761)
--	I10032 = NOT(g1236)
--	g1718 = NOT(I5562)
--	g7779 = NOT(I14208)
--	g2293 = NOT(g888)
--	g6880 = NOT(I12511)
--	g4684 = NOT(I8949)
--	I9050 = NOT(g3881)
--	I11452 = NOT(g6071)
--	g6595 = NOT(g6083)
--	g4639 = NOT(I8832)
--	I5682 = NOT(g168)
--	I5766 = NOT(g1254)
--	I11047 = NOT(g5653)
--	I13574 = NOT(g7205)
--	g2329 = NOT(I6130)
--	I6440 = NOT(g1806)
--	g7023 = NOT(I12779)
--	g9121 = NOT(I15747)
--	g4963 = NOT(g4328)
--	g2761 = NOT(g1820)
--	I5801 = NOT(g1424)
--	g9321 = NOT(g9311)
--	g8960 = NOT(I15394)
--	g7423 = NOT(I13544)
--	g1582 = NOT(g714)
--	I11912 = NOT(g5897)
--	I11311 = NOT(g5760)
--	I13912 = NOT(g7359)
--	I13311 = NOT(g7162)
--	g2828 = NOT(g1980)
--	I12298 = NOT(g6697)
--	I6323 = NOT(g1342)
--	I14061 = NOT(g7546)
--	g1793 = NOT(g626)
--	I7561 = NOT(g2562)
--	g7588 = NOT(I13909)
--	I10766 = NOT(g5674)
--	g2727 = NOT(g2424)
--	g4808 = NOT(I9145)
--	g6978 = NOT(I12717)
--	g6612 = NOT(I11832)
--	g7161 = NOT(I13057)
--	g1015 = NOT(I5416)
--	g5729 = NOT(g5144)
--	g3968 = NOT(I7683)
--	g6243 = NOT(I11050)
--	g7361 = NOT(I13499)
--	I15193 = NOT(g8774)
--	I13051 = NOT(g6967)
--	I13072 = NOT(g6969)
--	g2746 = NOT(g2259)
--	I12737 = NOT(g6460)
--	g2221 = NOT(I5936)
--	g3076 = NOT(g1831)
--	g7127 = NOT(g6974)
--	g8783 = NOT(g8524)
--	g7327 = NOT(I13403)
--	I12232 = NOT(g6662)
--	g1664 = NOT(g1462)
--	I6151 = NOT(g12)
--	g1246 = NOT(I5425)
--	g2703 = NOT(g1809)
--	g8218 = NOT(I14433)
--	I8823 = NOT(g3965)
--	g5014 = NOT(I9344)
--	g206 = NOT(I5353)
--	g6328 = NOT(I11311)
--	g6130 = NOT(I10761)
--	g7146 = NOT(g6998)
--	g6542 = NOT(I11718)
--	g6330 = NOT(I11317)
--	g7346 = NOT(I13454)
--	g7633 = NOT(I13962)
--	g1721 = NOT(I5565)
--	I11350 = NOT(g5763)
--	g3871 = NOT(g2953)
--	I7970 = NOT(g3557)
--	I13350 = NOT(g7223)
--	I15475 = NOT(g8901)
--	g2932 = NOT(g2329)
--	g7103 = NOT(I12897)
--	I9271 = NOT(g4263)
--	g3651 = NOT(I7129)
--	g7303 = NOT(I13341)
--	I7925 = NOT(g2761)
--	g8676 = NOT(I14822)
--	g2624 = NOT(g1569)
--	g2953 = NOT(g2373)
--	I15222 = NOT(g8834)
--	g6800 = NOT(I12271)
--	g3285 = NOT(g1689)
--	I13152 = NOT(g6966)
--	g8761 = NOT(g8564)
--	g4604 = NOT(I8727)
--	I10451 = NOT(g5216)
--	I10472 = NOT(g5223)
--	I13846 = NOT(g7487)
--	g3500 = NOT(g1616)
--	I14451 = NOT(g8172)
--	g7732 = NOT(I14067)
--	I5407 = NOT(g4653)
--	I13731 = NOT(g7441)
--	I5920 = NOT(g219)
--	I6839 = NOT(g2185)
--	I5868 = NOT(g74)
--	I7320 = NOT(g2927)
--	g2677 = NOT(g1664)
--	g7753 = NOT(I14130)
--	g5178 = NOT(I9660)
--	g5679 = NOT(I10172)
--	I11413 = NOT(g5871)
--	I5718 = NOT(g896)
--	g7508 = NOT(I13704)
--	I13413 = NOT(g7127)
--	g6213 = NOT(I10976)
--	I5535 = NOT(g48)
--	g2866 = NOT(g2221)
--	g4584 = NOT(g3466)
--	I12445 = NOT(g6568)
--	g4539 = NOT(g2881)
--	g8746 = NOT(g8524)
--	g8221 = NOT(I14442)
--	g5335 = NOT(g4677)
--	g5831 = NOT(I10516)
--	g3838 = NOT(I7317)
--	g1689 = NOT(g855)
--	g2149 = NOT(I5894)
--	g2349 = NOT(I6163)
--	I12499 = NOT(g6597)
--	g7043 = NOT(g6543)
--	g9141 = NOT(g9129)
--	g5182 = NOT(I9672)
--	I10776 = NOT(g5576)
--	I12316 = NOT(g6736)
--	I9132 = NOT(g4284)
--	I6143 = NOT(g1217)
--	I9209 = NOT(g4349)
--	g7116 = NOT(I12936)
--	g1671 = NOT(g1494)
--	I7987 = NOT(g3528)
--	g5805 = NOT(I10448)
--	g5916 = NOT(g5384)
--	g5022 = NOT(g4438)
--	g2699 = NOT(g1674)
--	g4019 = NOT(I7778)
--	g6090 = NOT(g5529)
--	g4362 = NOT(g2810)
--	I11929 = NOT(g6190)
--	I12989 = NOT(g6932)
--	g3077 = NOT(I6805)
--	g7034 = NOT(g6525)
--	g5749 = NOT(g5207)
--	g6490 = NOT(I11656)
--	g6823 = NOT(I12340)
--	g7434 = NOT(I13565)
--	I14825 = NOT(g8651)
--	g3523 = NOT(g2407)
--	I14370 = NOT(g7603)
--	g6366 = NOT(I11425)
--	I12722 = NOT(g6611)
--	g7565 = NOT(I13865)
--	I7299 = NOT(g2961)
--	I5664 = NOT(g916)
--	g3643 = NOT(g2453)
--	I12924 = NOT(g6983)
--	I13583 = NOT(g7252)
--	g2241 = NOT(I5984)
--	g1564 = NOT(g642)
--	g7147 = NOT(g6904)
--	I16122 = NOT(g9353)
--	I10151 = NOT(g5007)
--	I10172 = NOT(g4873)
--	g7347 = NOT(I13457)
--	I15516 = NOT(g8977)
--	I9558 = NOT(g4597)
--	g5798 = NOT(I10433)
--	I14151 = NOT(g7555)
--	g1826 = NOT(g632)
--	I12271 = NOT(g6663)
--	I14172 = NOT(g7545)
--	g6148 = NOT(I10807)
--	g6649 = NOT(I11929)
--	I14996 = NOT(g8510)
--	g6348 = NOT(I11371)
--	I8989 = NOT(g4537)
--	g8677 = NOT(I14825)
--	g7533 = NOT(I13779)
--	g3634 = NOT(I7107)
--	I8193 = NOT(g3547)
--	g6155 = NOT(I10826)
--	I14844 = NOT(g8641)
--	g6851 = NOT(I12424)
--	g6355 = NOT(I11392)
--	I11787 = NOT(g6273)
--	I14394 = NOT(g7536)
--	I12753 = NOT(g6445)
--	g8866 = NOT(I15184)
--	g7210 = NOT(I13144)
--	g2644 = NOT(I6416)
--	g3499 = NOT(g2185)
--	I8971 = NOT(g4464)
--	I12145 = NOT(g5971)
--	g1638 = NOT(g1092)
--	I11302 = NOT(g5796)
--	I7738 = NOT(g3038)
--	g5873 = NOT(g5367)
--	I13302 = NOT(g7164)
--	g5037 = NOT(g4438)
--	g9111 = NOT(I15723)
--	I12199 = NOT(g6475)
--	g7013 = NOT(I12757)
--	g9311 = NOT(I16049)
--	g5437 = NOT(g5041)
--	I11827 = NOT(g6231)
--	g5653 = NOT(g4748)
--	g7413 = NOT(I13524)
--	I13743 = NOT(g7454)
--	g3926 = NOT(I7581)
--	g5302 = NOT(g5028)
--	I14420 = NOT(g7554)
--	I15208 = NOT(g8810)
--	g2818 = NOT(g1792)
--	g6063 = NOT(I10678)
--	g4070 = NOT(I7847)
--	I12529 = NOT(g6628)
--	g2867 = NOT(g2222)
--	g3754 = NOT(g2543)
--	I9600 = NOT(g4698)
--	g8198 = NOT(g7721)
--	g8747 = NOT(g8545)
--	g4025 = NOT(I7792)
--	I14318 = NOT(g7657)
--	g5719 = NOT(I10236)
--	I12696 = NOT(g6503)
--	g9374 = NOT(I16148)
--	I14227 = NOT(g7552)
--	I5689 = NOT(g906)
--	I7959 = NOT(g2793)
--	g1758 = NOT(g1084)
--	g1589 = NOT(g746)
--	I14025 = NOT(g7500)
--	I7517 = NOT(g3578)
--	I11803 = NOT(g6280)
--	I7082 = NOT(g2470)
--	g2893 = NOT(I6615)
--	I15726 = NOT(g9069)
--	g7117 = NOT(I12939)
--	g6279 = NOT(I11132)
--	g5917 = NOT(g5412)
--	g7317 = NOT(I13383)
--	I14058 = NOT(g7544)
--	g6720 = NOT(g6254)
--	I5428 = NOT(g49)
--	g6118 = NOT(g5549)
--	g6167 = NOT(I10862)
--	g6318 = NOT(I11281)
--	g1571 = NOT(g669)
--	g3983 = NOT(g2845)
--	g6367 = NOT(I11428)
--	g9180 = NOT(I15824)
--	g6872 = NOT(I12487)
--	g7601 = NOT(g7450)
--	I15607 = NOT(g8994)
--	g9380 = NOT(g9379)
--	g3862 = NOT(I7389)
--	g5042 = NOT(I9396)
--	g1711 = NOT(I5555)
--	g2274 = NOT(g782)
--	g6652 = NOT(I11936)
--	I12161 = NOT(g5971)
--	g4678 = NOT(I8935)
--	g3712 = NOT(g1952)
--	g8524 = NOT(g7855)
--	g6843 = NOT(I12400)
--	I15530 = NOT(g8972)
--	g5786 = NOT(I10403)
--	g4006 = NOT(I7749)
--	g2170 = NOT(g1229)
--	g1827 = NOT(g762)
--	g2614 = NOT(g1562)
--	g9020 = NOT(I15484)
--	g7775 = NOT(I14196)
--	g5164 = NOT(I9618)
--	g6393 = NOT(I11506)
--	g4635 = NOT(I8820)
--	g5364 = NOT(g5124)
--	I15565 = NOT(g8980)
--	g2325 = NOT(I6118)
--	g2821 = NOT(g1786)
--	I12259 = NOT(g6652)
--	I10377 = NOT(g5188)
--	g1774 = NOT(I5616)
--	I12708 = NOT(g6482)
--	g7581 = NOT(I13888)
--	I11662 = NOT(g5956)
--	I10739 = NOT(g5572)
--	g4087 = NOT(I7882)
--	g4105 = NOT(I7928)
--	g8152 = NOT(I14388)
--	I9076 = NOT(g4353)
--	g5054 = NOT(g4457)
--	g6834 = NOT(I12373)
--	g4801 = NOT(I9126)
--	g8867 = NOT(I15187)
--	I9889 = NOT(g4819)
--	I14739 = NOT(g8173)
--	g2939 = NOT(g2348)
--	g3961 = NOT(g3131)
--	g7060 = NOT(g6654)
--	I11890 = NOT(g6135)
--	g1803 = NOT(g758)
--	g7460 = NOT(g7172)
--	I15641 = NOT(g9017)
--	I6160 = NOT(g324)
--	g5725 = NOT(g4841)
--	g4748 = NOT(g4465)
--	I11482 = NOT(g6117)
--	g6598 = NOT(I11806)
--	g3927 = NOT(I7584)
--	I5609 = NOT(g16)
--	I11248 = NOT(g6149)
--	g1780 = NOT(g614)
--	I12244 = NOT(g6642)
--	I11710 = NOT(g6098)
--	I13710 = NOT(g7340)
--	g2636 = NOT(g1580)
--	g7739 = NOT(I14088)
--	g3014 = NOT(I6767)
--	I9651 = NOT(g4805)
--	g6321 = NOT(I11290)
--	g4226 = NOT(g3591)
--	g8386 = NOT(g8014)
--	I5883 = NOT(g80)
--	g2106 = NOT(I5883)
--	g8975 = NOT(I15429)
--	g3946 = NOT(g3097)
--	g2306 = NOT(I6075)
--	I13779 = NOT(g7406)
--	g9204 = NOT(I15894)
--	I15408 = NOT(g8896)
--	I15635 = NOT(g8976)
--	g6625 = NOT(I11867)
--	g1662 = NOT(g1412)
--	g2790 = NOT(g1793)
--	g7937 = NOT(I14285)
--	I7762 = NOT(g3029)
--	I12810 = NOT(g6607)
--	g6232 = NOT(I11031)
--	I11778 = NOT(g6180)
--	g3903 = NOT(I7498)
--	g9100 = NOT(I15690)
--	I12068 = NOT(g5847)
--	I10427 = NOT(g5210)
--	g7479 = NOT(I13635)
--	g9300 = NOT(I16026)
--	g5412 = NOT(I9850)
--	I10366 = NOT(g5715)
--	g6253 = NOT(g5403)
--	g6938 = NOT(I12635)
--	I14427 = NOT(g7835)
--	I5466 = NOT(g926)
--	g6813 = NOT(I12310)
--	g7294 = NOT(I13314)
--	g4373 = NOT(I8360)
--	g3513 = NOT(g2407)
--	I9139 = NOT(g4364)
--	g6909 = NOT(I12592)
--	g7190 = NOT(I13112)
--	g2622 = NOT(g1568)
--	I11945 = NOT(g5874)
--	I12337 = NOT(g6724)
--	I5365 = NOT(g3843)
--	I5861 = NOT(g1313)
--	I11356 = NOT(g5799)
--	I13356 = NOT(g7221)
--	g1816 = NOT(g767)
--	g5171 = NOT(I9639)
--	g4602 = NOT(I8721)
--	g7501 = NOT(I13679)
--	I11380 = NOT(g5822)
--	I10403 = NOT(g5202)
--	g5787 = NOT(I10406)
--	g4007 = NOT(I7752)
--	g2904 = NOT(g2287)
--	I14403 = NOT(g7679)
--	g7156 = NOT(I13042)
--	g5956 = NOT(I10582)
--	g6552 = NOT(I11722)
--	g7356 = NOT(I13484)
--	g4920 = NOT(g4105)
--	g6606 = NOT(I11824)
--	g4578 = NOT(g2917)
--	I11090 = NOT(g1000)
--	I7928 = NOT(g2873)
--	I11998 = NOT(g5918)
--	g8544 = NOT(I14657)
--	g3831 = NOT(I7296)
--	I11233 = NOT(g6147)
--	g2514 = NOT(g1330)
--	g4718 = NOT(I9018)
--	g8483 = NOT(g8038)
--	I8962 = NOT(g4553)
--	I7064 = NOT(g2458)
--	I11672 = NOT(g5971)
--	g1847 = NOT(g765)
--	I9672 = NOT(g4803)
--	I15711 = NOT(g9075)
--	I13672 = NOT(g7242)
--	I7899 = NOT(g3743)
--	g4535 = NOT(g2876)
--	g2403 = NOT(g1176)
--	g8636 = NOT(I14718)
--	g1685 = NOT(I5528)
--	g2145 = NOT(g1296)
--	g6687 = NOT(I12003)
--	g2345 = NOT(I6151)
--	g2841 = NOT(g2208)
--	I7785 = NOT(g3029)
--	g7704 = NOT(I14001)
--	g4582 = NOT(g2922)
--	g3805 = NOT(g1752)
--	g3916 = NOT(I7545)
--	g9323 = NOT(g9315)
--	g6586 = NOT(I11778)
--	g8790 = NOT(g8585)
--	g2695 = NOT(g1672)
--	g4015 = NOT(g3160)
--	g2637 = NOT(g1581)
--	I11449 = NOT(g6068)
--	I12918 = NOT(g7013)
--	g5684 = NOT(I10183)
--	g8061 = NOT(I14330)
--	g5745 = NOT(I10292)
--	I15492 = NOT(g8971)
--	g5639 = NOT(g4748)
--	I14127 = NOT(g7594)
--	g7163 = NOT(I13063)
--	g3947 = NOT(I7640)
--	I11897 = NOT(g6141)
--	g2307 = NOT(I6078)
--	I11961 = NOT(g5988)
--	g7032 = NOT(g6525)
--	g2536 = NOT(g1354)
--	g5109 = NOT(I9493)
--	I13897 = NOT(g7354)
--	g8756 = NOT(g8564)
--	g3798 = NOT(g1757)
--	g5309 = NOT(g4969)
--	g7432 = NOT(I13559)
--	g6141 = NOT(I10786)
--	g6860 = NOT(I12451)
--	g2359 = NOT(g1397)
--	g4664 = NOT(I8907)
--	I9499 = NOT(g4382)
--	g6341 = NOT(I11350)
--	I11404 = NOT(g5834)
--	g3560 = NOT(g2361)
--	g9351 = NOT(I16103)
--	g2223 = NOT(I5942)
--	I7844 = NOT(g3784)
--	I15982 = NOT(g9236)
--	g5808 = NOT(I10457)
--	g1562 = NOT(g636)
--	I6680 = NOT(g1558)
--	g6645 = NOT(I11917)
--	I16040 = NOT(g9285)
--	g4721 = NOT(I9025)
--	I14103 = NOT(g7584)
--	I11212 = NOT(g6146)
--	g2016 = NOT(I5852)
--	I7731 = NOT(g3029)
--	g5759 = NOT(I10350)
--	g8514 = NOT(g8040)
--	g3873 = NOT(g2956)
--	g3632 = NOT(I7101)
--	g3095 = NOT(I6831)
--	g1817 = NOT(I5689)
--	g3495 = NOT(g1616)
--	g3653 = NOT(g2459)
--	I8180 = NOT(g3529)
--	I12322 = NOT(g6751)
--	g8145 = NOT(I14381)
--	g2522 = NOT(g1342)
--	I14181 = NOT(g7725)
--	g7157 = NOT(I13045)
--	g2642 = NOT(g1588)
--	I8832 = NOT(g3936)
--	g6879 = NOT(I12508)
--	g7357 = NOT(I13487)
--	g6607 = NOT(I11827)
--	I12532 = NOT(g6594)
--	g3579 = NOT(g1929)
--	g3869 = NOT(I7400)
--	g6962 = NOT(I12687)
--	I8853 = NOT(g4034)
--	g6659 = NOT(I11955)
--	I12158 = NOT(g5956)
--	g6358 = NOT(I11401)
--	g6506 = NOT(I11680)
--	g1751 = NOT(g452)
--	I5847 = NOT(g1360)
--	I12561 = NOT(g6449)
--	I16183 = NOT(g9388)
--	g5604 = NOT(g4969)
--	I12295 = NOT(g6693)
--	g3917 = NOT(I7548)
--	g2654 = NOT(I6446)
--	I10190 = NOT(g4670)
--	g1585 = NOT(g724)
--	g4689 = NOT(I8966)
--	g6587 = NOT(I11781)
--	g9372 = NOT(I16142)
--	I15522 = NOT(g9018)
--	I15663 = NOT(g9066)
--	I14190 = NOT(g7531)
--	I9543 = NOT(g4279)
--	g6111 = NOT(g5453)
--	g8223 = NOT(I14448)
--	g6311 = NOT(I11260)
--	g5833 = NOT(I10522)
--	I7814 = NOT(g2605)
--	I13646 = NOT(g7245)
--	g9235 = NOT(I15959)
--	g4028 = NOT(I7797)
--	g2880 = NOT(g2234)
--	I7350 = NOT(g2971)
--	I6574 = NOT(g576)
--	g2595 = NOT(g1643)
--	I6864 = NOT(g2528)
--	I11971 = NOT(g6179)
--	g4030 = NOT(g3160)
--	g8016 = NOT(I14311)
--	g8757 = NOT(g8585)
--	g5584 = NOT(g4841)
--	g1673 = NOT(g1504)
--	g6374 = NOT(I11449)
--	I14211 = NOT(g7712)
--	g9134 = NOT(I15776)
--	I15553 = NOT(g9009)
--	I13369 = NOT(g7268)
--	g2272 = NOT(I6021)
--	I14088 = NOT(g7585)
--	g4564 = NOT(I8665)
--	I11368 = NOT(g5833)
--	g8642 = NOT(I14732)
--	I5562 = NOT(g1300)
--	I12364 = NOT(g6714)
--	I7769 = NOT(g3038)
--	g5162 = NOT(I9612)
--	g3770 = NOT(g2551)
--	g5268 = NOT(I9788)
--	I9014 = NOT(g3864)
--	g5362 = NOT(I9823)
--	I10497 = NOT(g5233)
--	I15536 = NOT(g9004)
--	g1772 = NOT(g607)
--	g6380 = NOT(I11467)
--	I9660 = NOT(g4806)
--	g6591 = NOT(I11787)
--	I15702 = NOT(g9064)
--	I13850 = NOT(g7328)
--	g6832 = NOT(I12367)
--	I5817 = NOT(g1081)
--	g2982 = NOT(g1848)
--	g8874 = NOT(I15208)
--	g3532 = NOT(g2407)
--	I7967 = NOT(g2787)
--	g7778 = NOT(I14205)
--	g1743 = NOT(g598)
--	g2234 = NOT(I5963)
--	g6853 = NOT(I12430)
--	g2128 = NOT(g1284)
--	g4638 = NOT(I8829)
--	g2629 = NOT(g1574)
--	g6020 = NOT(g5367)
--	g2328 = NOT(I6127)
--	I10987 = NOT(g5609)
--	I12289 = NOT(g6702)
--	I5605 = NOT(g58)
--	I10250 = NOT(g5268)
--	g7735 = NOT(I14076)
--	g4609 = NOT(I8742)
--	g6507 = NOT(I11683)
--	g4308 = NOT(I8277)
--	g1011 = NOT(I5413)
--	I13228 = NOT(g6892)
--	g9113 = NOT(I15729)
--	g6794 = NOT(I12253)
--	g1856 = NOT(g774)
--	I12571 = NOT(g6729)
--	g9313 = NOT(I16055)
--	I11011 = NOT(g5693)
--	I5751 = NOT(g963)
--	g5086 = NOT(I9460)
--	g8880 = NOT(I15218)
--	g3189 = NOT(I6864)
--	I13716 = NOT(g7331)
--	g5730 = NOT(I10247)
--	g7475 = NOT(I13631)
--	I16072 = NOT(g9303)
--	g3990 = NOT(g3160)
--	g2554 = NOT(I6376)
--	I14338 = NOT(g7581)
--	g5185 = NOT(I9681)
--	g4589 = NOT(g2930)
--	I10969 = NOT(g5606)
--	g9094 = NOT(I15672)
--	g7627 = NOT(I13956)
--	g3888 = NOT(g3097)
--	I15062 = NOT(g8632)
--	g6905 = NOT(I12586)
--	g3029 = NOT(g1929)
--	g7292 = NOT(I13308)
--	g3787 = NOT(g1842)
--	g8017 = NOT(g7692)
--	g6628 = NOT(I11880)
--	I15933 = NOT(g9210)
--	g7526 = NOT(I13758)
--	g5470 = NOT(g4899)
--	g5897 = NOT(I10569)
--	g3956 = NOT(g2845)
--	g5025 = NOT(I9363)
--	g6515 = NOT(g6125)
--	I11627 = NOT(g5874)
--	g6630 = NOT(I11884)
--	g4571 = NOT(g2908)
--	I12687 = NOT(g6745)
--	g3675 = NOT(I7167)
--	I12976 = NOT(g6928)
--	g1573 = NOT(g677)
--	g1863 = NOT(g68)
--	g6300 = NOT(I11227)
--	I13112 = NOT(g7021)
--	g7603 = NOT(I13940)
--	I11050 = NOT(g5335)
--	I11958 = NOT(g5874)
--	g7039 = NOT(g6543)
--	I9422 = NOT(g4360)
--	I8351 = NOT(g1160)
--	g8234 = NOT(I14489)
--	g4455 = NOT(g3811)
--	g2902 = NOT(g2285)
--	g7439 = NOT(I13574)
--	I12643 = NOT(g6501)
--	I5368 = NOT(g3853)
--	I11386 = NOT(g5764)
--	g1569 = NOT(g661)
--	g453 = NOT(I5362)
--	I5772 = NOT(g1240)
--	g2490 = NOT(I6326)
--	I6024 = NOT(g544)
--	I5531 = NOT(g866)
--	g2366 = NOT(I6198)
--	I12669 = NOT(g6477)
--	g7583 = NOT(I13894)
--	g7702 = NOT(I13997)
--	g4196 = NOT(I8097)
--	g5678 = NOT(I10169)
--	I6795 = NOT(g1683)
--	I10503 = NOT(g5235)
--	g3684 = NOT(g2180)
--	g3639 = NOT(g2424)
--	g4803 = NOT(I9132)
--	g6973 = NOT(I12708)
--	g5006 = NOT(I9333)
--	g3338 = NOT(g1901)
--	g8800 = NOT(I15010)
--	g3963 = NOT(I7672)
--	g9360 = NOT(I16116)
--	I15574 = NOT(g8983)
--	g4538 = NOT(g2880)
--	g1688 = NOT(I5535)
--	g2148 = NOT(g1304)
--	I15205 = NOT(g8809)
--	g2649 = NOT(I6431)
--	g4780 = NOT(I9089)
--	g1857 = NOT(g889)
--	g2348 = NOT(I6160)
--	I7788 = NOT(g2595)
--	g9050 = NOT(I15550)
--	g5682 = NOT(I10177)
--	g5766 = NOT(I10373)
--	g5087 = NOT(I9463)
--	g1976 = NOT(g1269)
--	g6969 = NOT(I12702)
--	I15912 = NOT(g9193)
--	I9095 = NOT(g4283)
--	g5801 = NOT(I10442)
--	g3808 = NOT(g1827)
--	g7276 = NOT(I13264)
--	g5487 = NOT(I9907)
--	I14315 = NOT(g7676)
--	I6643 = NOT(g1970)
--	I11793 = NOT(g6188)
--	I11428 = NOT(g5813)
--	I12424 = NOT(g6446)
--	I13428 = NOT(g7167)
--	g3707 = NOT(g2226)
--	g6323 = NOT(I11296)
--	I14819 = NOT(g8647)
--	g4662 = NOT(I8901)
--	g2698 = NOT(g1673)
--	g4018 = NOT(I7775)
--	I12558 = NOT(g6449)
--	I14202 = NOT(g7708)
--	I8172 = NOT(g3524)
--	I14257 = NOT(g7716)
--	I9579 = NOT(g4713)
--	g2964 = NOT(I6716)
--	I14055 = NOT(g7495)
--	I16020 = NOT(g9264)
--	g9379 = NOT(I16161)
--	I7392 = NOT(g3230)
--	g5755 = NOT(g5494)
--	I15592 = NOT(g8989)
--	I15756 = NOT(g9081)
--	g7527 = NOT(I13761)
--	I14070 = NOT(g7714)
--	g3957 = NOT(I7662)
--	I12544 = NOT(g6617)
--	I6099 = NOT(g584)
--	I9752 = NOT(g4705)
--	g4093 = NOT(I7902)
--	g8512 = NOT(g8094)
--	I8282 = NOT(g3515)
--	I16046 = NOT(g9288)
--	g1760 = NOT(I5605)
--	g4493 = NOT(I8543)
--	g7764 = NOT(I14163)
--	g6351 = NOT(I11380)
--	g6648 = NOT(I11926)
--	g6875 = NOT(I12496)
--	g7546 = NOT(I13822)
--	g3865 = NOT(g2944)
--	I10384 = NOT(g5193)
--	g6655 = NOT(I11945)
--	g5445 = NOT(g5059)
--	g5173 = NOT(I9645)
--	I11317 = NOT(g5787)
--	g3604 = NOT(g2407)
--	I13317 = NOT(g7211)
--	g5491 = NOT(g4918)
--	g3498 = NOT(g1616)
--	I14067 = NOT(g7550)
--	I14094 = NOT(g7593)
--	g4381 = NOT(g3466)
--	g8649 = NOT(I14743)
--	g6010 = NOT(I10608)
--	g3833 = NOT(I7302)
--	I11129 = NOT(g5418)
--	g2872 = NOT(I6590)
--	g1924 = NOT(g174)
--	g5169 = NOT(I9633)
--	g4685 = NOT(I8952)
--	g4197 = NOT(g3591)
--	I10801 = NOT(g5463)
--	g6410 = NOT(I11533)
--	g7224 = NOT(I13164)
--	I7520 = NOT(g2734)
--	g4021 = NOT(g3131)
--	g5007 = NOT(I9336)
--	I13057 = NOT(g6968)
--	I14801 = NOT(g8608)
--	g2652 = NOT(I6440)
--	g1779 = NOT(g612)
--	g2057 = NOT(I5868)
--	I7640 = NOT(g3062)
--	I12124 = NOT(g5847)
--	I12678 = NOT(g6516)
--	g6884 = NOT(I12523)
--	g2843 = NOT(I6571)
--	g7120 = NOT(I12948)
--	g5059 = NOT(I9419)
--	g6839 = NOT(I12388)
--	g2457 = NOT(g24)
--	g5578 = NOT(g4841)
--	g5868 = NOT(I10555)
--	g7320 = NOT(I13388)
--	g2989 = NOT(g1843)
--	g3539 = NOT(g2424)
--	g3896 = NOT(I7473)
--	I11245 = NOT(g6143)
--	g5459 = NOT(g4882)
--	I14019 = NOT(g7480)
--	g2393 = NOT(I6267)
--	g5718 = NOT(g4841)
--	I12460 = NOT(g6674)
--	I12939 = NOT(g7022)
--	I11323 = NOT(g5808)
--	g1977 = NOT(g1357)
--	I11299 = NOT(g5786)
--	I13323 = NOT(g7145)
--	I14196 = NOT(g7534)
--	I13299 = NOT(g7163)
--	I14695 = NOT(g8016)
--	g7277 = NOT(I13267)
--	g1588 = NOT(g741)
--	I11533 = NOT(g5847)
--	g2834 = NOT(I6564)
--	g2971 = NOT(I6723)
--	I13533 = NOT(g7220)
--	g8063 = NOT(I14334)
--	g5582 = NOT(g4969)
--	I15405 = NOT(g8902)
--	g6278 = NOT(I11129)
--	g8463 = NOT(g8094)
--	g2686 = NOT(g1667)
--	g6372 = NOT(I11443)
--	g7789 = NOT(I14224)
--	g5261 = NOT(g4748)
--	g3019 = NOT(g2007)
--	g9132 = NOT(I15770)
--	g5793 = NOT(I10418)
--	I12065 = NOT(g5897)
--	I8202 = NOT(g3560)
--	g9332 = NOT(g9322)
--	g6618 = NOT(g6003)
--	g1665 = NOT(g1467)
--	g6143 = NOT(I10796)
--	g7516 = NOT(I13728)
--	I7765 = NOT(g2595)
--	g6343 = NOT(I11356)
--	g4562 = NOT(g3466)
--	g6235 = NOT(I11034)
--	g5015 = NOT(I9347)
--	g3052 = NOT(g2096)
--	g9209 = NOT(g9199)
--	g9353 = NOT(I16107)
--	I7911 = NOT(g2767)
--	I10457 = NOT(g5218)
--	I8094 = NOT(g2976)
--	g7771 = NOT(I14184)
--	I14457 = NOT(g8093)
--	g6566 = NOT(I11740)
--	g4631 = NOT(I8808)
--	I13737 = NOT(g7446)
--	g372 = NOT(I5359)
--	I15583 = NOT(g8986)
--	g7299 = NOT(I13329)
--	g4257 = NOT(I8190)
--	g6693 = NOT(I12011)
--	g6134 = NOT(g5428)
--	g8619 = NOT(I14695)
--	g7547 = NOT(I13825)
--	g6334 = NOT(I11329)
--	g4301 = NOT(I8264)
--	g5246 = NOT(I9760)
--	g2625 = NOT(g1570)
--	g8872 = NOT(I15202)
--	g2232 = NOT(I5957)
--	g4605 = NOT(I8730)
--	g3086 = NOT(g1852)
--	g2253 = NOT(g1323)
--	g2938 = NOT(g2347)
--	g3728 = NOT(g2202)
--	I14001 = NOT(g7433)
--	I13261 = NOT(g7041)
--	I11880 = NOT(g5748)
--	g6555 = NOT(I11729)
--	g6804 = NOT(I12283)
--	I7473 = NOT(g3546)
--	g2909 = NOT(g2291)
--	I6946 = NOT(g1887)
--	I10256 = NOT(g5401)
--	g6792 = NOT(I12247)
--	I11512 = NOT(g5874)
--	g1732 = NOT(g1439)
--	I9675 = NOT(g4807)
--	I13512 = NOT(g7138)
--	g3881 = NOT(g2969)
--	I5383 = NOT(g647)
--	I10280 = NOT(g5488)
--	g8971 = NOT(I15417)
--	g7738 = NOT(I14085)
--	g4585 = NOT(g2925)
--	I8264 = NOT(g3653)
--	g6621 = NOT(I11855)
--	g1944 = NOT(I5817)
--	g3897 = NOT(g3131)
--	g4041 = NOT(g2605)
--	I12915 = NOT(g7000)
--	g9092 = NOT(I15666)
--	I8360 = NOT(g1186)
--	g6313 = NOT(I11266)
--	g7078 = NOT(g6683)
--	g7340 = NOT(I13438)
--	I7377 = NOT(g3189)
--	I10157 = NOT(g5109)
--	I13831 = NOT(g7322)
--	I6036 = NOT(g130)
--	I14157 = NOT(g7547)
--	I12277 = NOT(g6681)
--	I6178 = NOT(g1220)
--	g4673 = NOT(I8928)
--	g6202 = NOT(I10949)
--	g8670 = NOT(I14804)
--	I9684 = NOT(g4813)
--	g7035 = NOT(g6543)
--	I13499 = NOT(g7134)
--	I15803 = NOT(g9148)
--	I9639 = NOT(g4685)
--	g7517 = NOT(I13731)
--	I7287 = NOT(g2561)
--	g6094 = NOT(I10716)
--	I14231 = NOT(g7566)
--	I9791 = NOT(g4779)
--	I6831 = NOT(g2185)
--	g5028 = NOT(I9372)
--	g4669 = NOT(I8922)
--	g1565 = NOT(g649)
--	I8724 = NOT(g3927)
--	g5671 = NOT(I10160)
--	I11722 = NOT(g5772)
--	I12782 = NOT(g6463)
--	I13722 = NOT(g7442)
--	I16090 = NOT(g9336)
--	I6805 = NOT(g1603)
--	g3635 = NOT(g1949)
--	I13924 = NOT(g7365)
--	I5633 = NOT(g891)
--	g1681 = NOT(g929)
--	g6776 = NOT(I12199)
--	I7781 = NOT(g2605)
--	I6422 = NOT(g1805)
--	g6593 = NOT(I11793)
--	g4890 = NOT(g4075)
--	I12352 = NOT(g6752)
--	I13432 = NOT(g7280)
--	g2525 = NOT(I6354)
--	g3801 = NOT(I7262)
--	I14763 = NOT(g7834)
--	I13271 = NOT(g7067)
--	g2645 = NOT(I6419)
--	I8835 = NOT(g3954)
--	g5826 = NOT(I10503)
--	I12418 = NOT(g6572)
--	I7797 = NOT(g3019)
--	g8606 = NOT(I14683)
--	I12170 = NOT(g5956)
--	g4011 = NOT(I7762)
--	I11461 = NOT(g6094)
--	g9076 = NOT(I15622)
--	g5741 = NOT(I10280)
--	g7110 = NOT(I12918)
--	I5732 = NOT(g859)
--	g6264 = NOT(g5403)
--	g7310 = NOT(I13362)
--	I11031 = NOT(g5335)
--	I13031 = NOT(g6984)
--	g5638 = NOT(g4748)
--	g6360 = NOT(I11407)
--	g2879 = NOT(I6597)
--	I13199 = NOT(g7025)
--	I11736 = NOT(g6076)
--	I11887 = NOT(g5918)
--	g9375 = NOT(I16151)
--	I7344 = NOT(g2964)
--	g2962 = NOT(g2382)
--	g5609 = NOT(g4748)
--	I15003 = NOT(g8633)
--	I8799 = NOT(g3951)
--	g2659 = NOT(g1655)
--	g6050 = NOT(g5246)
--	I12167 = NOT(g5939)
--	g2506 = NOT(I6341)
--	g1820 = NOT(g621)
--	I6437 = NOT(g1784)
--	I11696 = NOT(g5971)
--	g7236 = NOT(g6944)
--	I6302 = NOT(g1313)
--	g3091 = NOT(g1603)
--	I13843 = NOT(g7326)
--	I16026 = NOT(g9267)
--	g7762 = NOT(I14157)
--	g3491 = NOT(g1800)
--	g4080 = NOT(I7867)
--	I14076 = NOT(g7577)
--	I14085 = NOT(g7583)
--	g4573 = NOT(g2911)
--	I11764 = NOT(g6056)
--	g5758 = NOT(I10347)
--	I13764 = NOT(g7479)
--	g6724 = NOT(I12088)
--	I11365 = NOT(g5826)
--	g2275 = NOT(g990)
--	g2311 = NOT(I6090)
--	I9539 = NOT(g4018)
--	g6179 = NOT(I10896)
--	I13365 = NOT(g7267)
--	g5466 = NOT(g4890)
--	g4713 = NOT(I9014)
--	I10243 = NOT(g5026)
--	g6379 = NOT(I11464)
--	I11132 = NOT(g5624)
--	g7590 = NOT(I13915)
--	g9184 = NOT(I15830)
--	I13869 = NOT(g7338)
--	I5565 = NOT(g1296)
--	g2615 = NOT(g1563)
--	g6878 = NOT(I12505)
--	g5165 = NOT(I9621)
--	g4569 = NOT(g2906)
--	g5571 = NOT(I10032)
--	g3920 = NOT(g3097)
--	I12022 = NOT(g5874)
--	g3578 = NOT(I7053)
--	g3868 = NOT(g2948)
--	g2174 = NOT(g1319)
--	g6289 = NOT(I11194)
--	g6777 = NOT(I12202)
--	I8802 = NOT(g3963)
--	g6658 = NOT(g6224)
--	g2374 = NOT(I6220)
--	g5448 = NOT(g5137)
--	g1922 = NOT(g1251)
--	I9162 = NOT(g4272)
--	g7556 = NOT(I13846)
--	I13161 = NOT(g7080)
--	I10773 = NOT(g5708)
--	g5055 = NOT(g4477)
--	I12313 = NOT(g6730)
--	g6835 = NOT(I12376)
--	g2985 = NOT(I6733)
--	I9419 = NOT(g3916)
--	I10268 = NOT(g5471)
--	g1581 = NOT(g710)
--	g5827 = NOT(I10506)
--	I12748 = NOT(g6585)
--	g6882 = NOT(I12517)
--	I6042 = NOT(g237)
--	I15651 = NOT(g9056)
--	I15672 = NOT(g9047)
--	g3582 = NOT(g2407)
--	g2284 = NOT(I6036)
--	I5914 = NOT(g1097)
--	I13225 = NOT(g7095)
--	g7064 = NOT(I12829)
--	g2239 = NOT(I5978)
--	I7314 = NOT(g2916)
--	I10180 = NOT(g4721)
--	I16148 = NOT(g9368)
--	g1597 = NOT(g973)
--	g9077 = NOT(I15625)
--	g2180 = NOT(g1318)
--	g5846 = NOT(g5367)
--	g2380 = NOT(I6242)
--	I13258 = NOT(g6907)
--	I12900 = NOT(g6947)
--	I7870 = NOT(g2827)
--	I8901 = NOT(g4122)
--	g2832 = NOT(g2184)
--	I12466 = NOT(g6687)
--	g5396 = NOT(g4692)
--	I5413 = NOT(g1016)
--	g1784 = NOT(I5636)
--	g6799 = NOT(I12268)
--	I6054 = NOT(g465)
--	g2020 = NOT(I5855)
--	I10930 = NOT(g5600)
--	I15513 = NOT(g8970)
--	I11043 = NOT(g5648)
--	I6454 = NOT(g1868)
--	I12101 = NOT(g5971)
--	I6770 = NOT(g1590)
--	g6674 = NOT(I11978)
--	I13244 = NOT(g7033)
--	g7563 = NOT(I13861)
--	g8111 = NOT(I14374)
--	g5780 = NOT(I10387)
--	g4000 = NOT(g3131)
--	I10694 = NOT(g5445)
--	g4126 = NOT(I7981)
--	I10965 = NOT(g5719)
--	g6997 = NOT(I12737)
--	g7295 = NOT(I13317)
--	g2794 = NOT(g2185)
--	I11069 = NOT(g5671)
--	g9104 = NOT(I15702)
--	I5936 = NOT(g222)
--	g9099 = NOT(I15687)
--	I6532 = NOT(g1694)
--	g9304 = NOT(g9298)
--	g2931 = NOT(I6669)
--	g3721 = NOT(I7211)
--	g6238 = NOT(I11043)
--	I6553 = NOT(g2246)
--	g5662 = NOT(g5027)
--	I13810 = NOT(g7312)
--	g8174 = NOT(I14403)
--	g6332 = NOT(I11323)
--	I15717 = NOT(g9051)
--	I11955 = NOT(g5988)
--	g5418 = NOT(g5100)
--	g5467 = NOT(g4891)
--	I9025 = NOT(g4462)
--	g6353 = NOT(I11386)
--	g7194 = NOT(I13118)
--	I13879 = NOT(g7332)
--	I9425 = NOT(g3917)
--	g655 = NOT(I5383)
--	g2905 = NOT(I6629)
--	I6012 = NOT(g384)
--	g6744 = NOT(I12124)
--	g7731 = NOT(I14064)
--	g6802 = NOT(I12277)
--	g8284 = NOT(I14531)
--	g2628 = NOT(g1573)
--	g3502 = NOT(g1616)
--	g8545 = NOT(g7905)
--	I6189 = NOT(g249)
--	g2630 = NOT(g1575)
--	g5493 = NOT(g4920)
--	g8180 = NOT(g7719)
--	I14279 = NOT(g7700)
--	g4608 = NOT(I8739)
--	g4924 = NOT(g4113)
--	I5775 = NOT(g1240)
--	g7966 = NOT(I14291)
--	g2100 = NOT(g1227)
--	g3940 = NOT(I7623)
--	I10469 = NOT(g5222)
--	I11967 = NOT(g5971)
--	I11994 = NOT(g6195)
--	g7471 = NOT(g7233)
--	I15723 = NOT(g9065)
--	g9044 = NOT(I15536)
--	g1942 = NOT(g828)
--	I6029 = NOT(g1207)
--	g4023 = NOT(I7788)
--	I8736 = NOT(g4008)
--	I10286 = NOT(g5519)
--	I6371 = NOT(g33)
--	g1704 = NOT(I5548)
--	g5181 = NOT(I9669)
--	I12008 = NOT(g5897)
--	I9678 = NOT(g4808)
--	I15433 = NOT(g8911)
--	g5847 = NOT(I10552)
--	I6956 = NOT(g1907)
--	g6901 = NOT(g6525)
--	I14039 = NOT(g7449)
--	g4588 = NOT(g2929)
--	I11425 = NOT(g5872)
--	g5685 = NOT(I10186)
--	g5197 = NOT(g4938)
--	I13425 = NOT(g7166)
--	g5397 = NOT(g5076)
--	I8889 = NOT(g4311)
--	g6511 = NOT(I11693)
--	g703 = NOT(I5398)
--	I11458 = NOT(g6063)
--	I15811 = NOT(g9151)
--	I10815 = NOT(g5418)
--	I12454 = NOT(g6581)
--	g2973 = NOT(g1854)
--	g1810 = NOT(I5676)
--	g3430 = NOT(I6956)
--	g4665 = NOT(I8910)
--	I12712 = NOT(g6543)
--	g4051 = NOT(g3093)
--	g6092 = NOT(g5317)
--	I13918 = NOT(g7361)
--	I15971 = NOT(g9233)
--	I8871 = NOT(g3869)
--	I14187 = NOT(g7728)
--	g7150 = NOT(g6952)
--	I14677 = NOT(g7791)
--	g7350 = NOT(I13466)
--	g6864 = NOT(I12463)
--	I7195 = NOT(g1795)
--	g2969 = NOT(g2393)
--	I13444 = NOT(g7282)
--	g6714 = NOT(I12068)
--	g7773 = NOT(I14190)
--	g4146 = NOT(I8011)
--	g7009 = NOT(I12753)
--	g4633 = NOT(I8814)
--	g2323 = NOT(I6112)
--	I10937 = NOT(g5560)
--	I6963 = NOT(g1558)
--	g1568 = NOT(g658)
--	I6109 = NOT(g1214)
--	I6791 = NOT(g1967)
--	g4103 = NOT(I7922)
--	I12567 = NOT(g6721)
--	I6309 = NOT(g1336)
--	g4303 = NOT(I8268)
--	I11086 = NOT(g5397)
--	I7807 = NOT(g2595)
--	g3910 = NOT(I7523)
--	I12238 = NOT(g6637)
--	g7769 = NOT(I14178)
--	I10169 = NOT(g4873)
--	I7859 = NOT(g2804)
--	g4696 = NOT(I8983)
--	g1912 = NOT(g1524)
--	g5631 = NOT(g4938)
--	g7836 = NOT(I14260)
--	I14169 = NOT(g7715)
--	g5723 = NOT(g4938)
--	g4732 = NOT(I9034)
--	g5101 = NOT(g4259)
--	I12382 = NOT(g6772)
--	I5356 = NOT(g3837)
--	g2528 = NOT(g1260)
--	I14410 = NOT(g7697)
--	g2351 = NOT(g792)
--	g2648 = NOT(I6428)
--	I8838 = NOT(g3967)
--	I12176 = NOT(g5939)
--	I8024 = NOT(g3076)
--	I12675 = NOT(g6510)
--	g6736 = NOT(I12108)
--	g8750 = NOT(g8524)
--	I10479 = NOT(g5227)
--	g6968 = NOT(I12699)
--	g2655 = NOT(g1611)
--	g8973 = NOT(I15423)
--	g1929 = NOT(g1224)
--	I12154 = NOT(g5874)
--	I5942 = NOT(g300)
--	I9369 = NOT(g3901)
--	g7229 = NOT(g6938)
--	g6623 = NOT(I11861)
--	g7993 = NOT(I14298)
--	I7255 = NOT(g1955)
--	g6076 = NOT(g5287)
--	I14015 = NOT(g7440)
--	I9407 = NOT(g4232)
--	g6889 = NOT(I12538)
--	I11656 = NOT(g5772)
--	I13656 = NOT(g7228)
--	g3589 = NOT(I7061)
--	g8040 = NOT(g7699)
--	I11353 = NOT(g5788)
--	g9036 = NOT(I15522)
--	g4443 = NOT(I8449)
--	I13353 = NOT(g7231)
--	I11680 = NOT(g5939)
--	g8969 = NOT(I15411)
--	I8477 = NOT(g3014)
--	g9178 = NOT(I15814)
--	g9378 = NOT(I16158)
--	I13144 = NOT(g7031)
--	g4116 = NOT(I7959)
--	g6375 = NOT(I11452)
--	g6871 = NOT(I12484)
--	g4316 = NOT(I8291)
--	I5954 = NOT(g89)
--	g2884 = NOT(g2238)
--	g3861 = NOT(I7386)
--	g5041 = NOT(I9393)
--	g3048 = NOT(I6784)
--	g4034 = NOT(I7811)
--	I9582 = NOT(g4694)
--	I8205 = NOT(g2655)
--	g6651 = NOT(I11933)
--	g9182 = NOT(g9178)
--	I5432 = NOT(g1176)
--	g4565 = NOT(g2901)
--	g8666 = NOT(I14792)
--	g9382 = NOT(I16168)
--	I15959 = NOT(g9217)
--	I15379 = NOT(g8882)
--	I8742 = NOT(g3919)
--	g2372 = NOT(I6214)
--	g3774 = NOT(g1770)
--	I13631 = NOT(g7248)
--	I5568 = NOT(g1409)
--	g8875 = NOT(I15211)
--	g3846 = NOT(I7341)
--	g2618 = NOT(g1566)
--	g1683 = NOT(g795)
--	I16129 = NOT(g9355)
--	g6384 = NOT(I11479)
--	g2235 = NOT(I5966)
--	g2343 = NOT(g1392)
--	g6139 = NOT(I10780)
--	g5168 = NOT(I9630)
--	I12439 = NOT(g6566)
--	g5669 = NOT(I10154)
--	g4697 = NOT(I8986)
--	g6339 = NOT(I11344)
--	g4914 = NOT(g4093)
--	I14531 = NOT(g8178)
--	g2282 = NOT(g1400)
--	I7112 = NOT(g2546)
--	g1778 = NOT(g613)
--	g1894 = NOT(I5772)
--	g5058 = NOT(I9416)
--	g6838 = NOT(I12385)
--	g4596 = NOT(g3466)
--	I8754 = NOT(g3911)
--	g6024 = NOT(g5494)
--	I14178 = NOT(g7562)
--	g4013 = NOT(g3131)
--	g2134 = NOT(g1317)
--	g6795 = NOT(I12256)
--	g3780 = NOT(g1847)
--	I10186 = NOT(g5129)
--	g6737 = NOT(I12111)
--	g2334 = NOT(I6143)
--	I15681 = NOT(g9063)
--	g6809 = NOT(I12298)
--	I8273 = NOT(g2976)
--	I12349 = NOT(g6742)
--	g5743 = NOT(I10286)
--	I6419 = NOT(g1799)
--	I10373 = NOT(g5722)
--	g1782 = NOT(g624)
--	I7676 = NOT(g2584)
--	g2548 = NOT(g1351)
--	I7293 = NOT(g2955)
--	I12906 = NOT(g6918)
--	I15429 = NOT(g8899)
--	I7129 = NOT(g2495)
--	I13023 = NOT(g7040)
--	g1661 = NOT(g1405)
--	I7329 = NOT(g2920)
--	I11224 = NOT(g6255)
--	g6672 = NOT(I11974)
--	g2555 = NOT(g936)
--	g6231 = NOT(I11028)
--	g3018 = NOT(I6770)
--	I11308 = NOT(g5759)
--	g2804 = NOT(g1796)
--	I12304 = NOT(g6711)
--	g9095 = NOT(I15675)
--	I13308 = NOT(g7169)
--	g5734 = NOT(I10259)
--	g1949 = NOT(g1292)
--	g6523 = NOT(I11707)
--	I9502 = NOT(g3972)
--	g3994 = NOT(g3192)
--	I8983 = NOT(g4536)
--	g9102 = NOT(I15696)
--	g9208 = NOT(g9198)
--	I15765 = NOT(g9039)
--	g9302 = NOT(g9281)
--	I8862 = NOT(g3981)
--	g6205 = NOT(g5628)
--	I14334 = NOT(g7578)
--	g8172 = NOT(I14397)
--	I15690 = NOT(g9074)
--	g2621 = NOT(g1567)
--	I8712 = NOT(g4007)
--	I7592 = NOT(g2712)
--	g5074 = NOT(I9440)
--	g3093 = NOT(g1686)
--	I6728 = NOT(g1959)
--	I8543 = NOT(g2810)
--	g5474 = NOT(g4904)
--	g1646 = NOT(g1214)
--	g7298 = NOT(I13326)
--	g4601 = NOT(I8718)
--	I7746 = NOT(g3591)
--	g6634 = NOT(I11894)
--	g8667 = NOT(I14795)
--	I13816 = NOT(g7455)
--	g8235 = NOT(I14492)
--	g2313 = NOT(I6096)
--	g6742 = NOT(I12120)
--	g1603 = NOT(I5471)
--	g6104 = NOT(g5345)
--	I14964 = NOT(g8406)
--	g6304 = NOT(I11239)
--	I15504 = NOT(g8967)
--	g2202 = NOT(g1321)
--	I12138 = NOT(g5874)
--	g4922 = NOT(g4111)
--	I10587 = NOT(g5439)
--	I13752 = NOT(g7315)
--	I11374 = NOT(g5844)
--	g3847 = NOT(I7344)
--	g2908 = NOT(g2290)
--	g5480 = NOT(g4913)
--	I6425 = NOT(g1811)
--	g5713 = NOT(g4841)
--	g4581 = NOT(g2921)
--	I12415 = NOT(g6410)
--	g3700 = NOT(g2514)
--	g9042 = NOT(I15530)
--	g2494 = NOT(g9)
--	I7953 = NOT(g3542)
--	g6754 = NOT(I12135)
--	g1583 = NOT(g718)
--	g5569 = NOT(I10028)
--	g4597 = NOT(I8706)
--	I9564 = NOT(g4703)
--	I5894 = NOT(g86)
--	I11669 = NOT(g5918)
--	g7708 = NOT(I14005)
--	I13669 = NOT(g7240)
--	g9233 = NOT(I15953)
--	g7520 = NOT(I13740)
--	g8792 = NOT(I14996)
--	I11260 = NOT(g5779)
--	g6613 = NOT(I11835)
--	g3950 = NOT(g3131)
--	g4784 = NOT(I9095)
--	I10569 = NOT(g5417)
--	g4739 = NOT(I9053)
--	I11392 = NOT(g5800)
--	g1952 = NOT(g1333)
--	I9910 = NOT(g4681)
--	g6269 = NOT(I11090)
--	g5688 = NOT(I10193)
--	I6006 = NOT(g306)
--	I15533 = NOT(g9002)
--	g2965 = NOT(g2384)
--	g6983 = NOT(I12722)
--	g1616 = NOT(I5478)
--	I14747 = NOT(g8175)
--	g7176 = NOT(I13084)
--	I5475 = NOT(g1084)
--	I7716 = NOT(g3038)
--	g6572 = NOT(I11764)
--	g6862 = NOT(I12457)
--	I11559 = NOT(g6065)
--	g4079 = NOT(I7864)
--	I11525 = NOT(g5874)
--	I11488 = NOT(g6034)
--	I13559 = NOT(g7177)
--	g3562 = NOT(I7044)
--	I12484 = NOT(g6621)
--	I9609 = NOT(g4780)
--	g2264 = NOT(I5997)
--	g6712 = NOT(I12062)
--	g7405 = NOT(I13518)
--	g4668 = NOT(I8919)
--	I6087 = NOT(g318)
--	I6305 = NOT(g1333)
--	g3631 = NOT(I7098)
--	g7829 = NOT(I14251)
--	g2360 = NOT(g1435)
--	g2933 = NOT(I6673)
--	g3723 = NOT(g2096)
--	I12609 = NOT(g6571)
--	g7286 = NOT(I13290)
--	g7765 = NOT(I14166)
--	I7198 = NOT(g2509)
--	I10807 = NOT(g5294)
--	g5000 = NOT(I9325)
--	I5646 = NOT(g883)
--	g8094 = NOT(g7705)
--	I14807 = NOT(g8603)
--	g2641 = NOT(g1587)
--	I14974 = NOT(g8442)
--	I9217 = NOT(g4443)
--	I10639 = NOT(g5224)
--	g4501 = NOT(g2801)
--	g6729 = NOT(g6263)
--	g6961 = NOT(I12684)
--	I13544 = NOT(g1167)
--	g3605 = NOT(g1938)
--	I13865 = NOT(g7333)
--	g2996 = NOT(g1828)
--	I9466 = NOT(g3943)
--	g5760 = NOT(I10353)
--	g9189 = NOT(I15845)
--	g7733 = NOT(I14070)
--	I12921 = NOT(g6993)
--	I13713 = NOT(g7341)
--	g9389 = NOT(I16183)
--	g1970 = NOT(I5831)
--	I6226 = NOT(g408)
--	g7270 = NOT(I13250)
--	I8805 = NOT(g3976)
--	I10265 = NOT(g5468)
--	I8916 = NOT(g4195)
--	g1925 = NOT(g825)
--	g8776 = NOT(g8585)
--	g2724 = NOT(g1814)
--	g7225 = NOT(g6936)
--	g7610 = NOT(g7450)
--	g9029 = NOT(I15501)
--	g6014 = NOT(I10614)
--	I14416 = NOT(g7727)
--	g2379 = NOT(I6239)
--	I13610 = NOT(g7227)
--	I12813 = NOT(g6607)
--	I16145 = NOT(g9367)
--	g6885 = NOT(I12526)
--	I6045 = NOT(g309)
--	g4704 = NOT(I9001)
--	I13042 = NOT(g6963)
--	g6660 = NOT(I11958)
--	g6946 = NOT(I12649)
--	I13255 = NOT(g7057)
--	g2878 = NOT(g2233)
--	I13189 = NOT(g7002)
--	I7644 = NOT(g2584)
--	g5183 = NOT(I9675)
--	I13679 = NOT(g7259)
--	g7124 = NOT(g6896)
--	I12973 = NOT(g6927)
--	g5608 = NOT(g4969)
--	I9333 = NOT(g4245)
--	g2289 = NOT(I6051)
--	g6903 = NOT(I12582)
--	g2777 = NOT(g1797)
--	g9281 = NOT(I16009)
--	g5779 = NOT(I10384)
--	I10579 = NOT(g5433)
--	I9774 = NOT(g4678)
--	g4250 = NOT(I8177)
--	g2882 = NOT(g2236)
--	I11686 = NOT(g6076)
--	I11939 = NOT(g6015)
--	I7867 = NOT(g2818)
--	g9297 = NOT(I16017)
--	I13460 = NOT(g7263)
--	g4032 = NOT(I7807)
--	I11383 = NOT(g5827)
--	g2271 = NOT(I6018)
--	I9396 = NOT(g3908)
--	I13383 = NOT(g7275)
--	g1789 = NOT(g1034)
--	g7206 = NOT(I13134)
--	I6578 = NOT(g1603)
--	I6868 = NOT(g530)
--	I5616 = NOT(g979)
--	g6036 = NOT(I10643)
--	I13267 = NOT(g6913)
--	g6378 = NOT(I11461)
--	I6767 = NOT(g1933)
--	g5161 = NOT(I9609)
--	I16132 = NOT(g9356)
--	I10442 = NOT(g5215)
--	I15498 = NOT(g8974)
--	g1987 = NOT(I5842)
--	g1771 = NOT(g609)
--	I7211 = NOT(g1742)
--	g7287 = NOT(I13293)
--	I14442 = NOT(g8065)
--	g6135 = NOT(I10770)
--	I5404 = NOT(g722)
--	g4568 = NOT(g2904)
--	I7386 = NOT(g3013)
--	g5665 = NOT(g4748)
--	g9109 = NOT(I15717)
--	g5051 = NOT(I9407)
--	g6335 = NOT(I11332)
--	g6831 = NOT(I12364)
--	g9309 = NOT(I16043)
--	g3531 = NOT(g1616)
--	g5127 = NOT(I9525)
--	g2674 = NOT(g1675)
--	g6288 = NOT(I11191)
--	g6382 = NOT(I11473)
--	I16161 = NOT(g9363)
--	g8179 = NOT(I14416)
--	I9018 = NOT(g3872)
--	g3743 = NOT(g1776)
--	I7599 = NOT(g2734)
--	I15924 = NOT(g9207)
--	I6015 = NOT(g437)
--	I12400 = NOT(g6767)
--	g4357 = NOT(g3679)
--	g5146 = NOT(I9564)
--	g6805 = NOT(I12286)
--	g5633 = NOT(g4895)
--	I11218 = NOT(g6161)
--	I12214 = NOT(g6507)
--	g7781 = NOT(I14214)
--	g2238 = NOT(I5975)
--	g2332 = NOT(g926)
--	I10430 = NOT(g5211)
--	I13837 = NOT(g7324)
--	g3856 = NOT(I7371)
--	g2680 = NOT(g1665)
--	I14430 = NOT(g7836)
--	g2209 = NOT(I5926)
--	g2353 = NOT(g871)
--	I9493 = NOT(g4426)
--	g4929 = NOT(g4120)
--	g9201 = NOT(g9183)
--	I12328 = NOT(g6760)
--	I15753 = NOT(g9080)
--	g5696 = NOT(I10207)
--	g8882 = NOT(I15222)
--	g1945 = NOT(g1081)
--	g6947 = NOT(I12652)
--	g7510 = NOT(I13710)
--	g7245 = NOT(I13193)
--	g6798 = NOT(I12265)
--	I12538 = NOT(g6606)
--	g1738 = NOT(g741)
--	g3074 = NOT(I6800)
--	I16043 = NOT(g9285)
--	g5732 = NOT(I10253)
--	g7291 = NOT(I13305)
--	g3992 = NOT(I7723)
--	I14035 = NOT(g7310)
--	I15199 = NOT(g8792)
--	I10684 = NOT(g5258)
--	I11455 = NOT(g6087)
--	g4626 = NOT(I8793)
--	I8233 = NOT(g3588)
--	I11470 = NOT(g6095)
--	g5240 = NOT(I9752)
--	g7344 = NOT(g7150)
--	I13617 = NOT(g7276)
--	g5072 = NOT(g4457)
--	g9098 = NOT(I15684)
--	I13915 = NOT(g7360)
--	g8799 = NOT(I15007)
--	I12241 = NOT(g6640)
--	I14142 = NOT(g7551)
--	g1907 = NOT(g52)
--	g5472 = NOT(I9892)
--	I9021 = NOT(g4489)
--	g6873 = NOT(I12490)
--	g7207 = NOT(I13137)
--	g6632 = NOT(I11890)
--	g6095 = NOT(I10719)
--	g3080 = NOT(g1679)
--	g8674 = NOT(I14816)
--	g6037 = NOT(I10646)
--	g3573 = NOT(g2424)
--	I15696 = NOT(g9050)
--	g3863 = NOT(I7392)
--	I5789 = NOT(g1524)
--	g1959 = NOT(g1252)
--	g2901 = NOT(g2284)
--	g7259 = NOT(g7060)
--	g6653 = NOT(I11939)
--	I13277 = NOT(g7078)
--	g6102 = NOT(g5345)
--	g6208 = NOT(I10965)
--	g6302 = NOT(I11233)
--	g8541 = NOT(g8094)
--	I13075 = NOT(g6958)
--	g2511 = NOT(g1328)
--	I7061 = NOT(g2457)
--	g6869 = NOT(I12478)
--	g1876 = NOT(g77)
--	I12771 = NOT(g6735)
--	I11467 = NOT(g6064)
--	I11494 = NOT(g6037)
--	I13595 = NOT(g7216)
--	g7488 = NOT(g7225)
--	I12235 = NOT(g6634)
--	g2092 = NOT(g1225)
--	g5434 = NOT(g5112)
--	I10193 = NOT(g4670)
--	I11037 = NOT(g5299)
--	I14130 = NOT(g7592)
--	I14193 = NOT(g7532)
--	g6752 = NOT(I12131)
--	g5147 = NOT(I9567)
--	I13782 = NOT(g7498)
--	I11984 = NOT(g6246)
--	g8802 = NOT(I15014)
--	I11419 = NOT(g5835)
--	I6428 = NOT(g1818)
--	g9019 = NOT(I15481)
--	g9362 = NOT(I16122)
--	I13419 = NOT(g7277)
--	g3857 = NOT(I7374)
--	g7951 = NOT(I14288)
--	I8706 = NOT(g3828)
--	g3976 = NOT(I7697)
--	I15225 = NOT(g8689)
--	I15708 = NOT(g9072)
--	I13822 = NOT(g7459)
--	I10475 = NOT(g5529)
--	I9301 = NOT(g4295)
--	g7114 = NOT(I12930)
--	I11266 = NOT(g5794)
--	g4661 = NOT(I8898)
--	g6786 = NOT(I12229)
--	I7145 = NOT(g2501)
--	I6564 = NOT(g2073)
--	g4075 = NOT(I7856)
--	I5945 = NOT(g333)
--	I8787 = NOT(g4012)
--	g4475 = NOT(g3818)
--	g5596 = NOT(g4841)
--	g1663 = NOT(g1416)
--	I6826 = NOT(g2185)
--	g6364 = NOT(I11419)
--	g7870 = NOT(I14270)
--	g5013 = NOT(I9341)
--	g4627 = NOT(I8796)
--	I5709 = NOT(g901)
--	g8511 = NOT(I14646)
--	g9086 = NOT(I15648)
--	g1824 = NOT(I5706)
--	I5478 = NOT(g1148)
--	g6296 = NOT(I11215)
--	I11194 = NOT(g6243)
--	g4646 = NOT(I8853)
--	I7107 = NOT(g2480)
--	g2623 = NOT(g1585)
--	g6725 = NOT(I12091)
--	I9585 = NOT(g4697)
--	I10347 = NOT(g5706)
--	I10253 = NOT(g5240)
--	g5820 = NOT(I10485)
--	I7359 = NOT(g2871)
--	g9185 = NOT(I15833)
--	g4084 = NOT(I7875)
--	g4603 = NOT(I8724)
--	I5435 = NOT(g1461)
--	g7336 = NOT(I13428)
--	I13524 = NOT(g7151)
--	I15657 = NOT(g9059)
--	g9385 = NOT(I16173)
--	g8864 = NOT(I15178)
--	I15068 = NOT(g8638)
--	g7768 = NOT(I14175)
--	g1590 = NOT(I5466)
--	g1877 = NOT(g595)
--	I11401 = NOT(g5828)
--	g6553 = NOT(I11725)
--	g9070 = NOT(I15604)
--	g7594 = NOT(I13927)
--	I8745 = NOT(g3929)
--	I10236 = NOT(g5014)
--	g2375 = NOT(I6223)
--	g2871 = NOT(I6587)
--	I12725 = NOT(g6565)
--	g3220 = NOT(g1889)
--	I15337 = NOT(g8802)
--	g2651 = NOT(I6437)
--	I6217 = NOT(g105)
--	g6012 = NOT(g5367)
--	g1556 = NOT(g65)
--	I13118 = NOT(g7068)
--	g3779 = NOT(g2511)
--	g4583 = NOT(g2924)
--	I11864 = NOT(g5753)
--	I14175 = NOT(g7718)
--	g2285 = NOT(I6039)
--	I7115 = NOT(g2547)
--	g6189 = NOT(I10930)
--	I8808 = NOT(g4014)
--	g6389 = NOT(I11494)
--	I7811 = NOT(g3019)
--	I16158 = NOT(g9363)
--	I9669 = NOT(g4909)
--	I13749 = NOT(g7313)
--	g7887 = NOT(I14273)
--	g7122 = NOT(I12958)
--	g4919 = NOT(g4104)
--	g3977 = NOT(g3160)
--	I6571 = NOT(g1711)
--	g6888 = NOT(I12535)
--	I6048 = NOT(g387)
--	I10516 = NOT(g5241)
--	g5581 = NOT(g4969)
--	I14264 = NOT(g7698)
--	g3588 = NOT(g2379)
--	I9531 = NOT(g4463)
--	g2184 = NOT(I5911)
--	I6711 = NOT(g1726)
--	g6371 = NOT(I11440)
--	g1785 = NOT(g615)
--	g6787 = NOT(I12232)
--	g8968 = NOT(I15408)
--	g2384 = NOT(I6254)
--	I11704 = NOT(g6076)
--	g5060 = NOT(I9422)
--	I13704 = NOT(g7352)
--	I11305 = NOT(g5807)
--	g9331 = NOT(g9321)
--	g6956 = NOT(I12669)
--	I13305 = NOT(g7168)
--	g5460 = NOT(g4684)
--	g5597 = NOT(g4969)
--	I11254 = NOT(g5793)
--	g7433 = NOT(I13562)
--	g6675 = NOT(I11981)
--	g4616 = NOT(I8763)
--	I11809 = NOT(g6285)
--	I11900 = NOT(g5847)
--	g4561 = NOT(g2900)
--	g3051 = NOT(I6791)
--	I13900 = NOT(g7356)
--	I6333 = NOT(g1345)
--	I13466 = NOT(g7122)
--	I9505 = NOT(g4300)
--	g1563 = NOT(g639)
--	g2424 = NOT(g1329)
--	I12141 = NOT(g5897)
--	g2795 = NOT(g1801)
--	I8449 = NOT(g3630)
--	I12652 = NOT(g6664)
--	g9087 = NOT(I15651)
--	g9105 = NOT(I15705)
--	g5784 = NOT(I10397)
--	g4004 = NOT(g2845)
--	I15010 = NOT(g8584)
--	I15918 = NOT(g9211)
--	g9305 = NOT(I16033)
--	g5739 = NOT(I10274)
--	I8865 = NOT(g4032)
--	g7496 = NOT(I13666)
--	g4527 = NOT(g3466)
--	g7550 = NOT(I13834)
--	g6297 = NOT(I11218)
--	g3999 = NOT(I7738)
--	g4647 = NOT(I8856)
--	g8175 = NOT(I14406)
--	I8715 = NOT(g3903)
--	I7595 = NOT(g2573)
--	g8871 = NOT(I15199)
--	g3633 = NOT(I7104)
--	g2672 = NOT(I6471)
--	g2231 = NOT(I5954)
--	g7137 = NOT(I12993)
--	I14208 = NOT(g7711)
--	g8651 = NOT(I14747)
--	g2477 = NOT(g25)
--	I16017 = NOT(g9264)
--	g2643 = NOT(g1589)
--	g6684 = NOT(I11998)
--	I12135 = NOT(g5988)
--	g6639 = NOT(g6198)
--	g5668 = NOT(I10151)
--	g6338 = NOT(I11341)
--	I15598 = NOT(g8991)
--	I6509 = NOT(g1684)
--	g5294 = NOT(g5087)
--	g4503 = NOT(I8565)
--	g5840 = NOT(I10535)
--	g6963 = NOT(I12690)
--	I7978 = NOT(g3574)
--	g6791 = NOT(I12244)
--	g2205 = NOT(g13)
--	I12406 = NOT(g6773)
--	g6309 = NOT(I11254)
--	g5190 = NOT(g4938)
--	g4925 = NOT(g4114)
--	I5657 = NOT(g921)
--	I12361 = NOT(g6765)
--	I7417 = NOT(g3659)
--	g3732 = NOT(g2533)
--	I6018 = NOT(g462)
--	g1557 = NOT(I5432)
--	g2634 = NOT(g1578)
--	g3753 = NOT(g2540)
--	I10614 = NOT(g5302)
--	g6808 = NOT(I12295)
--	I9573 = NOT(g4701)
--	g9045 = NOT(I15539)
--	I10436 = NOT(g5213)
--	g724 = NOT(I5401)
--	I14614 = NOT(g7832)
--	g7266 = NOT(I13238)
--	g2551 = NOT(g1360)
--	I14436 = NOT(g7904)
--	g2104 = NOT(I5879)
--	g3944 = NOT(I7635)
--	I11693 = NOT(g6076)
--	g5156 = NOT(I9594)
--	g9373 = NOT(I16145)
--	g9091 = NOT(I15663)
--	g4120 = NOT(I7967)
--	I16023 = NOT(g9267)
--	I7629 = NOT(g3633)
--	g6759 = NOT(I12148)
--	I10274 = NOT(g5524)
--	I14073 = NOT(g7627)
--	I6093 = NOT(g468)
--	I8268 = NOT(g2801)
--	I13009 = NOT(g6935)
--	g1948 = NOT(g1250)
--	g8809 = NOT(I15065)
--	g7142 = NOT(I13012)
--	g6201 = NOT(I10946)
--	g2926 = NOT(g2325)
--	g7342 = NOT(I13444)
--	I11008 = NOT(g5693)
--	g9369 = NOT(I16135)
--	I10565 = NOT(g5402)
--	g6957 = NOT(I12672)
--	g7255 = NOT(I13209)
--	g4617 = NOT(I8766)
--	I8452 = NOT(g2816)
--	g649 = NOT(I5380)
--	g8672 = NOT(I14810)
--	g3316 = NOT(I6930)
--	g9059 = NOT(I15571)
--	I11476 = NOT(g6194)
--	I11485 = NOT(g6137)
--	I7800 = NOT(g2605)
--	g6449 = NOT(I11596)
--	g2273 = NOT(I6024)
--	g1814 = NOT(g630)
--	g6865 = NOT(I12466)
--	I7554 = NOT(g2573)
--	g7097 = NOT(I12881)
--	g7726 = NOT(I14049)
--	I13454 = NOT(g7147)
--	g7497 = NOT(I13669)
--	I10292 = NOT(g5577)
--	g2044 = NOT(I5861)
--	g7354 = NOT(I13478)
--	g5163 = NOT(I9615)
--	g6604 = NOT(I11818)
--	g5810 = NOT(I10463)
--	I13570 = NOT(g7198)
--	I6021 = NOT(g495)
--	g6498 = NOT(I11666)
--	g2269 = NOT(I6012)
--	g1773 = NOT(g610)
--	I8486 = NOT(g2824)
--	I10409 = NOT(g5204)
--	g4547 = NOT(g3466)
--	g5053 = NOT(g4438)
--	g6833 = NOT(I12370)
--	I8730 = NOT(g3987)
--	g3533 = NOT(g2397)
--	g5453 = NOT(g4680)
--	g2862 = NOT(I6578)
--	I15631 = NOT(g9003)
--	I12463 = NOT(g6682)
--	g4892 = NOT(I9250)
--	I11239 = NOT(g6173)
--	g2712 = NOT(g2039)
--	I14136 = NOT(g7633)
--	g9227 = NOT(I15947)
--	g1769 = NOT(I5609)
--	I9126 = NOT(g3870)
--	I7902 = NOT(g2709)
--	g2543 = NOT(g1348)
--	g6896 = NOT(I12561)
--	I13238 = NOT(g6900)
--	I9760 = NOT(g4838)
--	g3013 = NOT(I6764)
--	g1918 = NOT(g822)
--	g1967 = NOT(g1432)
--	g7112 = NOT(I12924)
--	g7267 = NOT(I13241)
--	I5966 = NOT(g278)
--	g5157 = NOT(I9597)
--	g2961 = NOT(I6711)
--	g4738 = NOT(I9050)
--	g8754 = NOT(g8524)
--	I5471 = NOT(g1029)
--	g6019 = NOT(g5367)
--	g6362 = NOT(I11413)
--	I13185 = NOT(g7020)
--	I6723 = NOT(g2052)
--	I13092 = NOT(g7047)
--	g7293 = NOT(I13311)
--	g2927 = NOT(I6663)
--	I12514 = NOT(g6605)
--	I5948 = NOT(g378)
--	g3936 = NOT(I7605)
--	I13518 = NOT(g7141)
--	g7129 = NOT(I12973)
--	I15571 = NOT(g8982)
--	I15308 = NOT(g8799)
--	g1822 = NOT(g761)
--	g7329 = NOT(I13407)
--	g7761 = NOT(I14154)
--	g4907 = NOT(g4087)
--	g2885 = NOT(g2239)
--	g4035 = NOT(I7814)
--	g2660 = NOT(I6451)
--	g2946 = NOT(g2365)
--	I12421 = NOT(g6486)
--	I14109 = NOT(g7590)
--	g7727 = NOT(I14052)
--	I15495 = NOT(g8973)
--	g4482 = NOT(I8520)
--	I7964 = NOT(g3488)
--	g2903 = NOT(g2286)
--	g5626 = NOT(g4748)
--	g7592 = NOT(I13921)
--	I8766 = NOT(g3960)
--	I9588 = NOT(g4704)
--	g6486 = NOT(I11648)
--	I8105 = NOT(g3339)
--	I10283 = NOT(g5643)
--	g4656 = NOT(I8883)
--	g7746 = NOT(I14109)
--	g6730 = NOT(I12098)
--	g9188 = NOT(I15842)
--	g7221 = NOT(I13157)
--	I15687 = NOT(g9071)
--	g9388 = NOT(I16180)
--	g3922 = NOT(I7561)
--	I15985 = NOT(g9237)
--	I14492 = NOT(g7829)
--	g9216 = NOT(I15924)
--	g6385 = NOT(I11482)
--	g6881 = NOT(I12514)
--	I12541 = NOT(g6614)
--	I8748 = NOT(g3997)
--	g4915 = NOT(g4094)
--	I11215 = NOT(g6156)
--	g9028 = NOT(I15498)
--	g6070 = NOT(g5317)
--	I11729 = NOT(g5772)
--	g1895 = NOT(I5775)
--	g6897 = NOT(I12564)
--	g1837 = NOT(g1007)
--	I13577 = NOT(g7186)
--	g9030 = NOT(I15504)
--	g6025 = NOT(g5367)
--	I6673 = NOT(g2246)
--	g6425 = NOT(I11556)
--	I14381 = NOT(g7596)
--	I13728 = NOT(g7439)
--	g5683 = NOT(I10180)
--	I12325 = NOT(g6755)
--	I9633 = NOT(g4800)
--	g2288 = NOT(I6048)
--	I7118 = NOT(g2484)
--	I7167 = NOT(g2505)
--	I14091 = NOT(g7589)
--	g2382 = NOT(I6248)
--	g7068 = NOT(g6556)
--	I12829 = NOT(g6441)
--	I12535 = NOT(g6599)
--	I15669 = NOT(g9045)
--	g3784 = NOT(g1768)
--	I10796 = NOT(g5397)
--	g8014 = NOT(g7564)
--	I9103 = NOT(g4374)
--	I12358 = NOT(g6761)
--	I13438 = NOT(g7143)
--	g3739 = NOT(g2536)
--	I6669 = NOT(g1698)
--	g4663 = NOT(I8904)
--	I6368 = NOT(g20)
--	g2916 = NOT(I6646)
--	I15842 = NOT(g9171)
--	I8373 = NOT(g3783)
--	g5735 = NOT(I10262)
--	g1788 = NOT(g984)
--	g3995 = NOT(I7728)
--	g3937 = NOT(g2845)
--	g8903 = NOT(I15315)
--	g3079 = NOT(g1603)
--	g5782 = NOT(I10393)
--	g4002 = NOT(g3192)
--	I10390 = NOT(g5195)
--	I13906 = NOT(g7358)
--	I11284 = NOT(g5795)
--	I13284 = NOT(g7156)
--	g6131 = NOT(g5529)
--	g7576 = NOT(I13873)
--	g6331 = NOT(I11320)
--	g5075 = NOT(I9443)
--	g3840 = NOT(I7323)
--	g2947 = NOT(I6695)
--	g7716 = NOT(I14025)
--	g7149 = NOT(I13031)
--	g2798 = NOT(g1787)
--	I11622 = NOT(g5847)
--	g1842 = NOT(g764)
--	g7349 = NOT(I13463)
--	g6635 = NOT(I11897)
--	I13622 = NOT(g7279)
--	g9108 = NOT(I15714)
--	g3390 = NOT(I6949)
--	g9308 = NOT(I16040)
--	I8868 = NOT(g4035)
--	g5627 = NOT(g4673)
--	g6682 = NOT(I11994)
--	g6766 = NOT(I12167)
--	g6087 = NOT(I10705)
--	I12173 = NOT(g5918)
--	g8178 = NOT(I14413)
--	g6305 = NOT(I11242)
--	g6801 = NOT(I12274)
--	I6856 = NOT(g449)
--	g4590 = NOT(g2932)
--	I10522 = NOT(g5243)
--	I15830 = NOT(g9180)
--	I8718 = NOT(g3909)
--	g3501 = NOT(g2185)
--	I9443 = NOT(g4564)
--	g5526 = NOT(g5086)
--	g7198 = NOT(I13126)
--	g4657 = NOT(I8886)
--	g7747 = NOT(I14112)
--	g7855 = NOT(I14267)
--	g9217 = NOT(I15927)
--	g2873 = NOT(g1779)
--	g1854 = NOT(g773)
--	g2632 = NOT(g1576)
--	I9116 = NOT(g4297)
--	I8261 = NOT(g3643)
--	g4556 = NOT(g2895)
--	g9066 = NOT(I15592)
--	I13653 = NOT(g7246)
--	g5084 = NOT(g4477)
--	g5603 = NOT(g4938)
--	g1941 = NOT(I5812)
--	I6474 = NOT(g1941)
--	g2495 = NOT(g26)
--	I8793 = NOT(g3923)
--	I9034 = NOT(g4317)
--	g2653 = NOT(I6443)
--	g7241 = NOT(I13185)
--	g6755 = NOT(I12138)
--	g2208 = NOT(I5923)
--	g3942 = NOT(I7629)
--	I12760 = NOT(g6685)
--	g5439 = NOT(g5058)
--	g4928 = NOT(g4119)
--	I10862 = NOT(g5364)
--	g6226 = NOT(g5658)
--	g4930 = NOT(g4121)
--	g8916 = NOT(I15334)
--	g2869 = NOT(g2224)
--	I15610 = NOT(g8995)
--	I15705 = NOT(g9068)
--	I10949 = NOT(g5513)
--	g9048 = NOT(I15546)
--	g4899 = NOT(g4080)
--	g4464 = NOT(I8486)
--	I9347 = NOT(g3896)
--	g1708 = NOT(I5552)
--	I9681 = NOT(g4811)
--	g7524 = NOT(I13752)
--	g6173 = NOT(I10882)
--	g2752 = NOT(g2389)
--	g3954 = NOT(I7655)
--	g6373 = NOT(I11446)
--	I10702 = NOT(g5529)
--	I15678 = NOT(g9060)
--	g9133 = NOT(I15773)
--	g2917 = NOT(g2309)
--	g9333 = NOT(g9323)
--	g7119 = NOT(I12945)
--	g1812 = NOT(I5682)
--	g7319 = NOT(g7124)
--	I14904 = NOT(g8629)
--	I8721 = NOT(g3918)
--	g1958 = NOT(g786)
--	g2265 = NOT(I6000)
--	g6369 = NOT(I11434)
--	g7352 = NOT(I13472)
--	g7577 = NOT(I13876)
--	g6007 = NOT(g5494)
--	I12927 = NOT(g7014)
--	g9196 = NOT(g9185)
--	g7717 = NOT(I14028)
--	g6059 = NOT(g5317)
--	g6868 = NOT(I12475)
--	g5616 = NOT(g4938)
--	g3568 = NOT(g1935)
--	g8873 = NOT(I15205)
--	I13484 = NOT(g7128)
--	g1829 = NOT(I5715)
--	g8632 = NOT(I14712)
--	I5842 = NOT(g68)
--	I15065 = NOT(g8636)
--	g6767 = NOT(I12170)
--	g2364 = NOT(I6192)
--	I12649 = NOT(g6457)
--	g2233 = NOT(I5960)
--	I10183 = NOT(g5129)
--	g1911 = NOT(I5789)
--	I10397 = NOT(g5200)
--	g7211 = NOT(I13147)
--	I5392 = NOT(g694)
--	g3912 = NOT(g3192)
--	I14397 = NOT(g7686)
--	g4089 = NOT(I7888)
--	I12903 = NOT(g6905)
--	g2454 = NOT(I6294)
--	I11200 = NOT(g6251)
--	g8869 = NOT(I15193)
--	g4489 = NOT(g2826)
--	g2770 = NOT(g2210)
--	g6793 = NOT(I12250)
--	I10509 = NOT(g5237)
--	g9018 = NOT(I15478)
--	g4557 = NOT(g2896)
--	g5764 = NOT(I10369)
--	g7599 = NOT(g7450)
--	g9067 = NOT(I15595)
--	g1974 = NOT(g803)
--	I10933 = NOT(g5668)
--	g7274 = NOT(I13258)
--	I15218 = NOT(g8801)
--	g6015 = NOT(I10617)
--	g4071 = NOT(I7850)
--	I6000 = NOT(g202)
--	I7341 = NOT(g2931)
--	g2532 = NOT(I6358)
--	g8752 = NOT(g8564)
--	g6227 = NOT(I11018)
--	g3929 = NOT(I7588)
--	I13921 = NOT(g7362)
--	I6326 = NOT(g1443)
--	I14851 = NOT(g8630)
--	g8917 = NOT(I15337)
--	g1796 = NOT(g617)
--	g4242 = NOT(I8161)
--	g7125 = NOT(I12965)
--	g9093 = NOT(I15669)
--	I8428 = NOT(g3611)
--	g6246 = NOT(I11055)
--	I7691 = NOT(g3651)
--	I15160 = NOT(g8631)
--	I13813 = NOT(g7314)
--	g8042 = NOT(I14325)
--	g5224 = NOT(g5114)
--	g7280 = NOT(I13274)
--	g8442 = NOT(I14623)
--	g6721 = NOT(g6257)
--	g8786 = NOT(g8545)
--	g5120 = NOT(I9512)
--	I12262 = NOT(g6656)
--	g2389 = NOT(g1230)
--	g9181 = NOT(g9177)
--	g2706 = NOT(g1821)
--	g7544 = NOT(I13816)
--	I8826 = NOT(g4023)
--	g9381 = NOT(I16165)
--	I5812 = NOT(g1243)
--	g7483 = NOT(g7226)
--	I15915 = NOT(g9194)
--	I9460 = NOT(g3941)
--	I9597 = NOT(g4738)
--	I6183 = NOT(g6)
--	g4350 = NOT(I8315)
--	g2888 = NOT(I6608)
--	I6608 = NOT(g1612)
--	g9197 = NOT(g9186)
--	I6220 = NOT(g126)
--	I10574 = NOT(g5426)
--	g2371 = NOT(g944)
--	I8910 = NOT(g4200)
--	g2787 = NOT(g1807)
--	g4438 = NOT(I8446)
--	g7106 = NOT(I12906)
--	I11732 = NOT(g6076)
--	g5617 = NOT(g4969)
--	g8770 = NOT(g8545)
--	g6502 = NOT(I11672)
--	I14205 = NOT(g7710)
--	g7306 = NOT(I13350)
--	g5789 = NOT(I10412)
--	g4009 = NOT(I7758)
--	g2956 = NOT(g2375)
--	I16119 = NOT(g9351)
--	I14311 = NOT(g7566)
--	g7790 = NOT(I14227)
--	g5516 = NOT(g4924)
--	I15595 = NOT(g8990)
--	g6940 = NOT(I12639)
--	I5911 = NOT(g216)
--	I8308 = NOT(g3674)
--	g7061 = NOT(g6650)
--	g7187 = NOT(I13103)
--	I7311 = NOT(g2879)
--	g5987 = NOT(g5294)
--	g1849 = NOT(I5732)
--	g3778 = NOT(g2145)
--	I13692 = NOT(g7343)
--	I13761 = NOT(g7418)
--	g642 = NOT(I5377)
--	I8883 = NOT(g4198)
--	g7756 = NOT(I14139)
--	g6388 = NOT(I11491)
--	I10592 = NOT(g5444)
--	g5299 = NOT(I9804)
--	I9840 = NOT(g4702)
--	g3735 = NOT(g1961)
--	g4918 = NOT(g4103)
--	g6216 = NOT(I10987)
--	g1781 = NOT(g622)
--	I6051 = NOT(g440)
--	I7374 = NOT(g3084)
--	I10780 = NOT(g5445)
--	g8012 = NOT(I14305)
--	I6127 = NOT(g471)
--	I6451 = NOT(g1895)
--	g6028 = NOT(g5529)
--	I14780 = NOT(g8284)
--	I12247 = NOT(g6646)
--	g6671 = NOT(I11971)
--	g7904 = NOT(I14276)
--	g1797 = NOT(g627)
--	g2639 = NOT(g1583)
--	g7046 = NOT(I12806)
--	I11329 = NOT(g5825)
--	g3075 = NOT(g2216)
--	g2963 = NOT(g2383)
--	g4229 = NOT(I8140)
--	I10350 = NOT(g5707)
--	I13329 = NOT(g7247)
--	g7446 = NOT(I13595)
--	g7514 = NOT(I13722)
--	g3949 = NOT(I7644)
--	g2309 = NOT(I6084)
--	g9101 = NOT(I15693)
--	I7545 = NOT(g3589)
--	I12388 = NOT(g6403)
--	g9301 = NOT(g9260)
--	g4822 = NOT(I9177)
--	g7145 = NOT(I13023)
--	g8029 = NOT(I14318)
--	I7380 = NOT(g3461)
--	g7345 = NOT(I13451)
--	I12098 = NOT(g5956)
--	g8787 = NOT(g8564)
--	I16036 = NOT(g9282)
--	I7832 = NOT(g2768)
--	g5738 = NOT(I10271)
--	g6826 = NOT(I12349)
--	g7763 = NOT(I14160)
--	g3526 = NOT(g2185)
--	g8956 = NOT(I15382)
--	g3998 = NOT(g3097)
--	g8675 = NOT(I14819)
--	g5709 = NOT(g4841)
--	I8333 = NOT(g3721)
--	g6741 = NOT(I12117)
--	I15589 = NOT(g8988)
--	g3084 = NOT(I6820)
--	g3603 = NOT(g2092)
--	I5377 = NOT(g635)
--	g785 = NOT(I5407)
--	g5478 = NOT(g5025)
--	I13241 = NOT(g7030)
--	I14413 = NOT(g7723)
--	g1694 = NOT(g21)
--	g7107 = NOT(I12909)
--	g4921 = NOT(g4202)
--	g7307 = NOT(I13353)
--	g3850 = NOT(I7353)
--	I15836 = NOT(g9165)
--	g2957 = NOT(g2376)
--	I8196 = NOT(g3654)
--	g7159 = NOT(I13051)
--	I7931 = NOT(g2780)
--	g1852 = NOT(g887)
--	g1923 = NOT(I5801)
--	I6072 = NOT(g1211)
--	g6108 = NOT(g5345)
--	g7359 = NOT(I13493)
--	I9250 = NOT(g4134)
--	g5435 = NOT(g5121)
--	g6308 = NOT(I11251)
--	g5517 = NOT(g4925)
--	g5690 = NOT(g4748)
--	I9363 = NOT(g4258)
--	g7223 = NOT(I13161)
--	g5482 = NOT(g4915)
--	g1701 = NOT(I5545)
--	g6883 = NOT(I12520)
--	I9053 = NOT(g4327)
--	g8684 = NOT(I14848)
--	g3583 = NOT(g2128)
--	g4895 = NOT(g4078)
--	g8639 = NOT(I14725)
--	I6443 = NOT(g1774)
--	g7757 = NOT(I14142)
--	I7905 = NOT(g2863)
--	I11683 = NOT(g5988)
--	g4620 = NOT(I8775)
--	g8791 = NOT(g8585)
--	g4462 = NOT(I8480)
--	g2498 = NOT(I6333)
--	g6217 = NOT(g5649)
--	g3919 = NOT(I7554)
--	g6758 = NOT(I12145)
--	g6589 = NOT(g6083)
--	g1886 = NOT(I5766)
--	I7204 = NOT(g2520)
--	I16009 = NOT(g9261)
--	I15616 = NOT(g8997)
--	I5781 = NOT(g979)
--	g2833 = NOT(I6561)
--	g7522 = NOT(I13746)
--	g7115 = NOT(I12933)
--	g7251 = NOT(I13203)
--	g8808 = NOT(I15062)
--	I6434 = NOT(g1830)
--	g3952 = NOT(I7651)
--	g7315 = NOT(I13373)
--	g7811 = NOT(I14238)
--	g7047 = NOT(g6498)
--	g9368 = NOT(I16132)
--	I8994 = NOT(g4565)
--	I10046 = NOT(g4840)
--	g6861 = NOT(I12454)
--	g6365 = NOT(I11422)
--	g2584 = NOT(g1646)
--	I14046 = NOT(g7492)
--	g4788 = NOT(I9103)
--	g6048 = NOT(g5246)
--	I11515 = NOT(g5897)
--	I11991 = NOT(g5939)
--	g2539 = NOT(I6363)
--	g2896 = NOT(g2269)
--	g3561 = NOT(I7041)
--	g9058 = NOT(I15568)
--	I13515 = NOT(g7152)
--	g8759 = NOT(g8524)
--	I13882 = NOT(g7350)
--	g6711 = NOT(I12059)
--	g1870 = NOT(I5751)
--	I11407 = NOT(g5841)
--	I13407 = NOT(g7271)
--	g1825 = NOT(I5709)
--	g6827 = NOT(I12352)
--	g3527 = NOT(g1616)
--	g8957 = NOT(I15385)
--	g6133 = NOT(I10766)
--	g6333 = NOT(I11326)
--	I14282 = NOT(g7709)
--	g3647 = NOT(g2424)
--	I9929 = NOT(g5052)
--	g2162 = NOT(I5901)
--	I7973 = NOT(g3071)
--	g2268 = NOT(I6009)
--	g6774 = NOT(I12193)
--	g2362 = NOT(I6186)
--	I12629 = NOT(g6523)
--	g3764 = NOT(g2039)
--	g4085 = NOT(I7878)
--	I12451 = NOT(g6524)
--	g6846 = NOT(I12409)
--	I12472 = NOT(g6591)
--	I12220 = NOT(g6645)
--	g8865 = NOT(I15181)
--	g3546 = NOT(I7029)
--	g5002 = NOT(g4335)
--	I14743 = NOT(g8174)
--	I8847 = NOT(g4025)
--	g2052 = NOT(I5865)
--	g5402 = NOT(g5000)
--	g5824 = NOT(I10497)
--	g7595 = NOT(I13930)
--	g6803 = NOT(I12280)
--	g2452 = NOT(g23)
--	g8604 = NOT(I14677)
--	g3503 = NOT(g2407)
--	g3970 = NOT(g2845)
--	g1768 = NOT(g605)
--	g9074 = NOT(I15616)
--	g6538 = NOT(I11714)
--	I13441 = NOT(g7146)
--	I5852 = NOT(g1202)
--	I5923 = NOT(g252)
--	I11206 = NOT(g6133)
--	I7323 = NOT(g2905)
--	g6780 = NOT(I12211)
--	g6509 = NOT(I11689)
--	g1806 = NOT(I5670)
--	g1943 = NOT(g1025)
--	I6820 = NOT(g1707)
--	g7243 = NOT(I13189)
--	I6936 = NOT(g1878)
--	I11725 = NOT(g6036)
--	I12776 = NOT(g6739)
--	I13725 = NOT(g7437)
--	g2728 = NOT(g2256)
--	g2486 = NOT(g959)
--	g6662 = NOT(I11964)
--	g6018 = NOT(g5494)
--	I6317 = NOT(g1339)
--	g1887 = NOT(g83)
--	I16176 = NOT(g9385)
--	I13758 = NOT(g7414)
--	I15693 = NOT(g9048)
--	I12355 = NOT(g6756)
--	I13435 = NOT(g7170)
--	g1934 = NOT(g154)
--	g2185 = NOT(I5914)
--	g6290 = NOT(I11197)
--	g4640 = NOT(I8835)
--	g2881 = NOT(g2235)
--	I7648 = NOT(g2712)
--	I16154 = NOT(g9370)
--	I7875 = NOT(g3819)
--	I12370 = NOT(g6758)
--	g4031 = NOT(I7804)
--	g7130 = NOT(I12976)
--	I7655 = NOT(g2734)
--	g3617 = NOT(g1655)
--	g6093 = NOT(g5345)
--	I11744 = NOT(g6120)
--	g7542 = NOT(I13810)
--	g2470 = NOT(g42)
--	g7330 = NOT(I13410)
--	g2897 = NOT(g2270)
--	g6493 = NOT(I11659)
--	g6256 = NOT(I11069)
--	I12151 = NOT(g5847)
--	g6816 = NOT(I12319)
--	g5785 = NOT(I10400)
--	I12996 = NOT(g6934)
--	g4005 = NOT(I7746)
--	I13940 = NOT(g7355)
--	I8101 = NOT(g3259)
--	I8817 = NOT(g3935)
--	I14662 = NOT(g7783)
--	g3987 = NOT(I7716)
--	g3771 = NOT(g1853)
--	I11848 = NOT(g6159)
--	I9782 = NOT(g4720)
--	I11398 = NOT(g5823)
--	I12367 = NOT(g6754)
--	I12394 = NOT(g6759)
--	I6060 = NOT(g580)
--	g6381 = NOT(I11470)
--	g4286 = NOT(g3790)
--	I11652 = NOT(g5939)
--	g6847 = NOT(I12412)
--	I6460 = NOT(g2104)
--	I6597 = NOT(g1970)
--	I10482 = NOT(g5228)
--	g3547 = NOT(g2345)
--	g6700 = NOT(g6244)
--	g6397 = NOT(I11512)
--	I10552 = NOT(g5396)
--	I8751 = NOT(g4009)
--	g3892 = NOT(g3131)
--	I11263 = NOT(g5784)
--	I10204 = NOT(g5060)
--	I9627 = NOT(g4777)
--	g2131 = NOT(g1300)
--	I6784 = NOT(g2052)
--	g2006 = NOT(g806)
--	g2331 = NOT(g933)
--	I12319 = NOT(g6741)
--	g4733 = NOT(g4202)
--	I11332 = NOT(g5832)
--	g5844 = NOT(I10545)
--	I13332 = NOT(g7241)
--	g6263 = NOT(g5688)
--	g4270 = NOT(g2573)
--	I5972 = NOT(g356)
--	g2635 = NOT(g1579)
--	g1807 = NOT(g619)
--	g6950 = NOT(I12659)
--	g8881 = NOT(g8683)
--	g9126 = NOT(I15756)
--	g4610 = NOT(I8745)
--	g2105 = NOT(g1444)
--	I7667 = NOT(g3052)
--	g3945 = NOT(g3097)
--	I12059 = NOT(g5874)
--	I10786 = NOT(g5452)
--	I12025 = NOT(g5918)
--	g2487 = NOT(I6323)
--	I9084 = NOT(g4358)
--	g5731 = NOT(I10250)
--	I9603 = NOT(g4719)
--	I13962 = NOT(g7413)
--	I14786 = NOT(g8606)
--	g7512 = NOT(I13716)
--	I9484 = NOT(g3957)
--	g3991 = NOT(g3160)
--	g7090 = NOT(g6525)
--	I6294 = NOT(g1330)
--	I9850 = NOT(g4798)
--	g594 = NOT(I5368)
--	I10356 = NOT(g5711)
--	I15382 = NOT(g8883)
--	I11500 = NOT(g6219)
--	g6562 = NOT(I11736)
--	g7366 = NOT(I13512)
--	g4069 = NOT(I7844)
--	I15519 = NOT(g9019)
--	g5071 = NOT(g4438)
--	g3078 = NOT(g1603)
--	g3340 = NOT(g2474)
--	I10826 = NOT(g5434)
--	I15675 = NOT(g9058)
--	I10380 = NOT(g5448)
--	g5705 = NOT(g4841)
--	g5471 = NOT(I9889)
--	g7056 = NOT(g6520)
--	g6631 = NOT(I11887)
--	g4540 = NOT(g2882)
--	g2226 = NOT(g1320)
--	I7548 = NOT(g3590)
--	I10998 = NOT(g5672)
--	I12044 = NOT(g5847)
--	g6723 = NOT(I12085)
--	g7456 = NOT(g7174)
--	I13048 = NOT(g6956)
--	g7529 = NOT(I13767)
--	g6257 = NOT(g5685)
--	g3959 = NOT(g3097)
--	g1815 = NOT(g760)
--	g6101 = NOT(g5317)
--	g7148 = NOT(I13028)
--	g6817 = NOT(I12322)
--	g9183 = NOT(g9161)
--	g6301 = NOT(I11230)
--	g7348 = NOT(I13460)
--	g3517 = NOT(g2283)
--	I11004 = NOT(g5613)
--	g3082 = NOT(g1680)
--	g9383 = NOT(g9380)
--	I8772 = NOT(g4011)
--	I7804 = NOT(g3029)
--	g9220 = NOT(g9205)
--	I11221 = NOT(g6167)
--	g7155 = NOT(I13039)
--	g7355 = NOT(I13481)
--	g6605 = NOT(I11821)
--	I7792 = NOT(g3038)
--	I12301 = NOT(g6703)
--	g8678 = NOT(I14828)
--	g1726 = NOT(g158)
--	g3876 = NOT(g3466)
--	g8131 = NOT(I14378)
--	I12120 = NOT(g5939)
--	g2373 = NOT(I6217)
--	g2091 = NOT(g819)
--	g8406 = NOT(I14614)
--	I13613 = NOT(g7273)
--	g1960 = NOT(g1268)
--	g5814 = NOT(I10475)
--	g7260 = NOT(g7064)
--	g6751 = NOT(I12128)
--	g5150 = NOT(I9576)
--	I8011 = NOT(g3225)
--	I9561 = NOT(g4695)
--	g8682 = NOT(I14844)
--	g8766 = NOT(g8545)
--	g5038 = NOT(g4457)
--	I5395 = NOT(g698)
--	I8856 = NOT(g3955)
--	g2283 = NOT(I6033)
--	g7063 = NOT(I12826)
--	I12699 = NOT(g6504)
--	g9161 = NOT(I15803)
--	I16138 = NOT(g9358)
--	I13106 = NOT(g7056)
--	g9361 = NOT(I16119)
--	g2007 = NOT(g1223)
--	I13605 = NOT(g7197)
--	I10448 = NOT(g5335)
--	g7463 = NOT(g7239)
--	g5009 = NOT(g4344)
--	g2407 = NOT(I6286)
--	I6163 = NOT(g402)
--	I14448 = NOT(g7792)
--	g2920 = NOT(I6652)
--	g2868 = NOT(g2223)
--	I6363 = NOT(g16)
--	I15501 = NOT(g8975)
--	g9051 = NOT(I15553)
--	I15729 = NOT(g9073)
--	g2459 = NOT(I6299)
--	I15577 = NOT(g8984)
--	g4898 = NOT(g4079)
--	g6441 = NOT(I11586)
--	I13463 = NOT(g7264)
--	g9127 = NOT(I15759)
--	g2767 = NOT(I6509)
--	g4900 = NOT(I9258)
--	g1783 = NOT(I5633)
--	I7908 = NOT(g3516)
--	g5769 = NOT(I10380)
--	I11951 = NOT(g5847)
--	I11371 = NOT(g5840)
--	g8755 = NOT(g8545)
--	g636 = NOT(I5371)
--	g7279 = NOT(I13271)
--	g8226 = NOT(I14457)
--	g5836 = NOT(g5529)
--	g4510 = NOT(g2840)
--	I13234 = NOT(g6898)
--	g4245 = NOT(I8172)
--	I12427 = NOT(g6553)
--	g7720 = NOT(I14035)
--	g7118 = NOT(I12942)
--	g5918 = NOT(I10574)
--	g2793 = NOT(I6532)
--	g7367 = NOT(I13515)
--	I12632 = NOT(g6514)
--	g9103 = NOT(I15699)
--	g9303 = NOT(g9301)
--	g1676 = NOT(g727)
--	g2015 = NOT(g33)
--	I8480 = NOT(g3640)
--	g6368 = NOT(I11431)
--	g7057 = NOT(g6644)
--	g8173 = NOT(I14400)
--	g4344 = NOT(g3124)
--	g6772 = NOT(I12187)
--	I6157 = NOT(g246)
--	I12403 = NOT(g6769)
--	I12547 = NOT(g6708)
--	g1828 = NOT(g769)
--	g2664 = NOT(I6463)
--	g2246 = NOT(I5989)
--	g4259 = NOT(I8196)
--	g5822 = NOT(I10491)
--	g6890 = NOT(I12541)
--	g7549 = NOT(I13831)
--	g1830 = NOT(I5718)
--	g4694 = NOT(I8977)
--	I15622 = NOT(g8999)
--	g1727 = NOT(g596)
--	g3590 = NOT(I7064)
--	g3877 = NOT(g2960)
--	I10433 = NOT(g5212)
--	I5692 = NOT(g906)
--	g8602 = NOT(g8094)
--	I10387 = NOT(g5194)
--	I12226 = NOT(g6636)
--	I14433 = NOT(g8061)
--	g7686 = NOT(I13979)
--	g8407 = NOT(g8013)
--	g4088 = NOT(I7885)
--	I12481 = NOT(g6616)
--	g9072 = NOT(I15610)
--	g3657 = NOT(I7145)
--	g4923 = NOT(g4112)
--	g2721 = NOT(g1803)
--	g6505 = NOT(I11677)
--	g8868 = NOT(I15190)
--	I14148 = NOT(g7543)
--	g6011 = NOT(g5494)
--	I5960 = NOT(g187)
--	g1746 = NOT(g290)
--	I14097 = NOT(g7595)
--	g6856 = NOT(I12439)
--	g4701 = NOT(I8994)
--	I10646 = NOT(g5364)
--	g8767 = NOT(g8564)
--	g9043 = NOT(I15533)
--	g3556 = NOT(I7036)
--	I13012 = NOT(g7071)
--	I10343 = NOT(g5704)
--	I14646 = NOT(g7790)
--	g3928 = NOT(g3097)
--	I16052 = NOT(g9291)
--	g8582 = NOT(g8094)
--	g9116 = NOT(I15738)
--	g6074 = NOT(g5317)
--	g3930 = NOT(g3097)
--	g2502 = NOT(I6337)
--	g9316 = NOT(g9302)
--	I11473 = NOT(g6069)
--	I13541 = NOT(g7209)
--	g4886 = NOT(g4071)
--	I10369 = NOT(g5716)
--	g9034 = NOT(I15516)
--	I12490 = NOT(g6625)
--	g8015 = NOT(g7689)
--	g2940 = NOT(I6686)
--	g8227 = NOT(I14460)
--	g4114 = NOT(I7953)
--	g7253 = NOT(g7049)
--	I11359 = NOT(g5810)
--	I12376 = NOT(g6766)
--	I12385 = NOT(g6397)
--	I13359 = NOT(g7255)
--	I9892 = NOT(g4879)
--	g5462 = NOT(g4886)
--	g2689 = NOT(g1670)
--	g6573 = NOT(g5868)
--	g6863 = NOT(I12460)
--	I11920 = NOT(g5874)
--	I12980 = NOT(g6929)
--	I7878 = NOT(g2829)
--	g8664 = NOT(I14786)
--	I8760 = NOT(g3931)
--	I11434 = NOT(g5789)
--	g3563 = NOT(g2007)
--	I10412 = NOT(g5205)
--	g2216 = NOT(I5933)
--	g6713 = NOT(I12065)
--	g1677 = NOT(g1532)
--	g7519 = NOT(I13737)
--	g7740 = NOT(I14091)
--	g4650 = NOT(I8865)
--	I7658 = NOT(g2562)
--	I5401 = NOT(g723)
--	I12888 = NOT(g6948)
--	I13828 = NOT(g7321)
--	I5676 = NOT(g911)
--	I14133 = NOT(g7574)
--	g2671 = NOT(I6468)
--	g9210 = NOT(g9200)
--	g1576 = NOT(g691)
--	g6569 = NOT(I11747)
--	g1866 = NOT(g71)
--	I7882 = NOT(g2700)
--	g5788 = NOT(I10409)
--	g4008 = NOT(I7755)
--	I10896 = NOT(g5475)
--	I6894 = NOT(g1863)
--	I11344 = NOT(g5820)
--	g3844 = NOT(I7335)
--	I13344 = NOT(g7210)
--	I15484 = NOT(g8918)
--	g1848 = NOT(g772)
--	I10716 = NOT(g5537)
--	I13682 = NOT(g7251)
--	g4594 = NOT(g2941)
--	g5842 = NOT(I10541)
--	g2826 = NOT(g2183)
--	g1747 = NOT(g599)
--	g1855 = NOT(g866)
--	I6075 = NOT(g2)
--	g6857 = NOT(I12442)
--	g7586 = NOT(I13903)
--	I9907 = NOT(g4837)
--	I13173 = NOT(g7089)
--	g5192 = NOT(g4841)
--	I10582 = NOT(g5437)
--	g3557 = NOT(g1773)
--	g5085 = NOT(I9457)
--	g4806 = NOT(I9139)
--	I7981 = NOT(g3555)
--	I6949 = NOT(g2148)
--	I12190 = NOT(g5918)
--	g3966 = NOT(g3160)
--	I8977 = NOT(g3877)
--	g2910 = NOT(I6636)
--	g3071 = NOT(g1948)
--	g3705 = NOT(I7204)
--	g9117 = NOT(I15741)
--	I12520 = NOT(g6622)
--	g2638 = NOT(g1582)
--	g4065 = NOT(I7838)
--	g9317 = NOT(g9306)
--	I8161 = NOT(g3517)
--	g8689 = NOT(I14857)
--	g4122 = NOT(I7973)
--	I15921 = NOT(g9206)
--	g4465 = NOT(g3677)
--	g7141 = NOT(I13009)
--	I14925 = NOT(g8381)
--	g3948 = NOT(g3131)
--	g4934 = NOT(g4125)
--	g7341 = NOT(I13441)
--	g8216 = NOT(I14427)
--	I6646 = NOT(g2246)
--	g2308 = NOT(I6081)
--	I7132 = NOT(g2554)
--	I13134 = NOT(g7017)
--	I7332 = NOT(g2947)
--	I8665 = NOT(g3051)
--	I12211 = NOT(g6502)
--	I14112 = NOT(g7560)
--	g6326 = NOT(I11305)
--	g7525 = NOT(I13755)
--	g7710 = NOT(I14009)
--	g3955 = NOT(I7658)
--	I7680 = NOT(g2712)
--	I11506 = NOT(g6189)
--	I14378 = NOT(g7691)
--	g2883 = NOT(g2237)
--	I6084 = NOT(g240)
--	I7353 = NOT(g2833)
--	g8671 = NOT(I14807)
--	I11028 = NOT(g5642)
--	I13506 = NOT(g7148)
--	I12088 = NOT(g5874)
--	I6039 = NOT(g207)
--	g4033 = NOT(g3192)
--	I13028 = NOT(g7087)
--	g6760 = NOT(I12151)
--	I14603 = NOT(g7827)
--	g5520 = NOT(g4928)
--	I15184 = NOT(g8684)
--	g4096 = NOT(I7911)
--	g8564 = NOT(g7951)
--	g3038 = NOT(g2092)
--	g1818 = NOT(I5692)
--	g1577 = NOT(g695)
--	g1867 = NOT(g878)
--	g9060 = NOT(I15574)
--	I9310 = NOT(g4268)
--	I7558 = NOT(g2734)
--	I10681 = NOT(g5686)
--	g5812 = NOT(I10469)
--	g6183 = NOT(I10914)
--	g7158 = NOT(I13048)
--	g2365 = NOT(I6195)
--	I12659 = NOT(g6459)
--	g6383 = NOT(I11476)
--	g7358 = NOT(I13490)
--	g5176 = NOT(I9654)
--	g4195 = NOT(I8094)
--	I9663 = NOT(g4809)
--	g6220 = NOT(I11001)
--	g7506 = NOT(I13698)
--	I15732 = NOT(g9076)
--	g4891 = NOT(g4076)
--	I13927 = NOT(g7366)
--	g4913 = NOT(g4092)
--	I12250 = NOT(g6651)
--	g658 = NOT(I5386)
--	g8910 = NOT(I15324)
--	I16100 = NOT(g9338)
--	g6779 = NOT(I12208)
--	I14857 = NOT(g8657)
--	g3769 = NOT(g2548)
--	I6952 = NOT(g1896)
--	g8638 = NOT(I14722)
--	g3836 = NOT(I7311)
--	g5829 = NOT(I10512)
--	g7587 = NOT(I13906)
--	I13649 = NOT(g7281)
--	g5286 = NOT(g4714)
--	g1975 = NOT(g1253)
--	I5747 = NOT(g1260)
--	g4807 = NOT(I9142)
--	g6977 = NOT(g6664)
--	g7111 = NOT(I12921)
--	I5855 = NOT(g71)
--	I5398 = NOT(g702)
--	g3918 = NOT(I7551)
--	g2774 = NOT(g1813)
--	g7275 = NOT(I13261)
--	g7311 = NOT(I13365)
--	g3967 = NOT(I7680)
--	I6561 = NOT(g1715)
--	I11648 = NOT(g6028)
--	I10690 = NOT(g5538)
--	g6588 = NOT(g5836)
--	I11491 = NOT(g6010)
--	I11903 = NOT(g5939)
--	g9079 = NOT(I15631)
--	I13903 = NOT(g7357)
--	g8883 = NOT(I15225)
--	g6161 = NOT(I10842)
--	I7492 = NOT(g3561)
--	g6361 = NOT(I11410)
--	g4266 = NOT(I8202)
--	g2396 = NOT(g1033)
--	I7864 = NOT(g3812)
--	I10548 = NOT(g5260)
--	I13755 = NOT(g7317)
--	g5733 = NOT(I10256)
--	g7174 = NOT(g7097)
--	g6051 = NOT(g5246)
--	g3993 = NOT(g3192)
--	g8217 = NOT(I14430)
--	I13770 = NOT(g7491)
--	I11981 = NOT(g6246)
--	I9657 = NOT(g4784)
--	I12968 = NOT(g6925)
--	g1821 = NOT(g631)
--	I15329 = NOT(g8793)
--	g6327 = NOT(I11308)
--	g2780 = NOT(I6517)
--	I6764 = NOT(g1955)
--	g3822 = NOT(g1815)
--	g5610 = NOT(g4938)
--	g2509 = NOT(g37)
--	I15539 = NOT(g9005)
--	g5073 = NOT(g4477)
--	g5796 = NOT(I10427)
--	I8565 = NOT(g3071)
--	g5473 = NOT(g4903)
--	g7284 = NOT(I13284)
--	g6146 = NOT(I10801)
--	g4081 = NOT(I7870)
--	g7239 = NOT(g6945)
--	g6346 = NOT(I11365)
--	g7545 = NOT(I13819)
--	I6970 = NOT(g1872)
--	g2662 = NOT(I6457)
--	g5124 = NOT(I9520)
--	g7180 = NOT(I13092)
--	g6103 = NOT(g5317)
--	g4692 = NOT(I8971)
--	g7591 = NOT(I13918)
--	g6303 = NOT(I11236)
--	g2467 = NOT(I6305)
--	I9064 = NOT(g4302)
--	I13767 = NOT(g7486)
--	I13794 = NOT(g7346)
--	I11395 = NOT(g5812)
--	g5469 = NOT(g4898)
--	g2290 = NOT(I6054)
--	I7262 = NOT(g2514)
--	I10128 = NOT(g4688)
--	g6696 = NOT(I12022)
--	g3921 = NOT(I7558)
--	I9785 = NOT(g4747)
--	I5577 = NOT(g172)
--	g4960 = NOT(g4259)
--	g7420 = NOT(I13537)
--	I11633 = NOT(g5897)
--	g5177 = NOT(I9657)
--	I12894 = NOT(g7009)
--	g7507 = NOT(I13701)
--	g8774 = NOT(I14964)
--	g5206 = NOT(g4938)
--	I7623 = NOT(g3631)
--	g2256 = NOT(g1324)
--	I11191 = NOT(g6155)
--	g2816 = NOT(g1685)
--	I13719 = NOT(g7334)
--	g6508 = NOT(I11686)
--	g6944 = NOT(I12643)
--	g3837 = NOT(I7314)
--	g6072 = NOT(g5345)
--	I11718 = NOT(g6115)
--	g3062 = NOT(g2100)
--	I14298 = NOT(g7678)
--	g9032 = NOT(I15510)
--	I5386 = NOT(g648)
--	g3462 = NOT(g1743)
--	g1756 = NOT(g533)
--	g2381 = NOT(I6245)
--	I5975 = NOT(g381)
--	I11832 = NOT(g6274)
--	g8780 = NOT(g8524)
--	g9053 = NOT(I15557)
--	I12202 = NOT(g6481)
--	g4112 = NOT(I7947)
--	g7905 = NOT(I14279)
--	g4267 = NOT(I8205)
--	g2700 = NOT(g1744)
--	I7651 = NOT(g2573)
--	I16107 = NOT(g9337)
--	I8820 = NOT(g3952)
--	I11440 = NOT(g6009)
--	g2397 = NOT(g1272)
--	I12496 = NOT(g6592)
--	g5199 = NOT(g4841)
--	g1904 = NOT(g1021)
--	I12111 = NOT(g5956)
--	g6316 = NOT(I11275)
--	g7515 = NOT(I13725)
--	I11861 = NOT(g5747)
--	g8662 = NOT(I14780)
--	g5781 = NOT(I10390)
--	g4001 = NOT(g3160)
--	g6034 = NOT(I10639)
--	g8018 = NOT(I14315)
--	I13861 = NOT(g7330)
--	I9089 = NOT(g4566)
--	g8067 = NOT(I14342)
--	g2263 = NOT(g1394)
--	g7100 = NOT(I12888)
--	I13247 = NOT(g6906)
--	I6299 = NOT(g47)
--	g7300 = NOT(I13332)
--	I11389 = NOT(g5766)
--	I11926 = NOT(g6190)
--	I12986 = NOT(g6931)
--	g5797 = NOT(I10430)
--	I15414 = NOT(g8900)
--	I13045 = NOT(g6955)
--	g6147 = NOT(I10804)
--	I5984 = NOT(g540)
--	g9157 = NOT(g9141)
--	g6347 = NOT(I11368)
--	I5939 = NOT(g275)
--	I13099 = NOT(g7054)
--	g3842 = NOT(I7329)
--	I13388 = NOT(g7149)
--	g8093 = NOT(I14370)
--	g6681 = NOT(I11991)
--	I11701 = NOT(g5772)
--	g8493 = NOT(g8041)
--	I13701 = NOT(g7349)
--	I10512 = NOT(g5238)
--	g3085 = NOT(g1945)
--	I8775 = NOT(g4019)
--	I7838 = NOT(g2781)
--	I8922 = NOT(g4229)
--	I11251 = NOT(g6152)
--	I11272 = NOT(g5758)
--	g7750 = NOT(I14121)
--	g3485 = NOT(g1737)
--	g2562 = NOT(g1652)
--	g1695 = NOT(g778)
--	g6697 = NOT(I12025)
--	g1637 = NOT(g1087)
--	g5144 = NOT(I9558)
--	g4592 = NOT(g2938)
--	g5344 = NOT(I9819)
--	g6210 = NOT(I10969)
--	I5636 = NOT(g891)
--	g2631 = NOT(g1586)
--	g4746 = NOT(I9076)
--	I12877 = NOT(g6700)
--	g8181 = NOT(I14420)
--	g6596 = NOT(I11800)
--	g5207 = NOT(g4673)
--	g8381 = NOT(I14603)
--	g3854 = NOT(I7365)
--	g2817 = NOT(g1849)
--	g3941 = NOT(I7626)
--	I7672 = NOT(g3062)
--	I16135 = NOT(g9357)
--	g4703 = NOT(I8998)
--	g5819 = NOT(I10482)
--	g8685 = NOT(I14851)
--	g7440 = NOT(I13577)
--	I10445 = NOT(g5418)
--	I7523 = NOT(g2562)
--	I14445 = NOT(g8067)
--	I12196 = NOT(g6471)
--	I6078 = NOT(g95)
--	g2605 = NOT(g1639)
--	I13140 = NOT(g6954)
--	I9350 = NOT(g4503)
--	g7123 = NOT(I12961)
--	g8421 = NOT(g8017)
--	g5088 = NOT(I9466)
--	I8784 = NOT(g3949)
--	I13997 = NOT(g7432)
--	I8739 = NOT(g3910)
--	g1757 = NOT(g604)
--	g5488 = NOT(I9910)
--	g4932 = NOT(g4202)
--	I12526 = NOT(g6626)
--	I15759 = NOT(g9082)
--	g5701 = NOT(g5120)
--	g6820 = NOT(I12331)
--	g4624 = NOT(I8787)
--	I9009 = NOT(g4591)
--	I6959 = NOT(g1558)
--	g3520 = NOT(g1616)
--	g6936 = NOT(I12629)
--	g3219 = NOT(I6872)
--	I6517 = NOT(g1687)
--	g3640 = NOT(I7112)
--	I16049 = NOT(g9288)
--	g6117 = NOT(I10739)
--	g1811 = NOT(I5679)
--	g6317 = NOT(I11278)
--	I7551 = NOT(g2712)
--	I7104 = NOT(g2479)
--	g3812 = NOT(g1750)
--	I12457 = NOT(g6671)
--	g7528 = NOT(I13764)
--	I14722 = NOT(g8076)
--	g7151 = NOT(I13035)
--	g3958 = NOT(g3097)
--	g7351 = NOT(I13469)
--	g4677 = NOT(I8932)
--	g6601 = NOT(g6083)
--	g7530 = NOT(I13770)
--	I12866 = NOT(g6483)
--	I8190 = NOT(g3545)
--	g8562 = NOT(g8094)
--	I9918 = NOT(g4968)
--	I10271 = NOT(g5487)
--	g5114 = NOT(I9502)
--	g4576 = NOT(g2913)
--	I15940 = NOT(g9213)
--	I13447 = NOT(g7261)
--	g8631 = NOT(I14709)
--	g2673 = NOT(I6474)
--	g6775 = NOT(I12196)
--	g3829 = NOT(I7290)
--	g6922 = NOT(g6525)
--	I5763 = NOT(g1207)
--	g3911 = NOT(I7526)
--	I6214 = NOT(g7)
--	g6581 = NOT(I11773)
--	g5825 = NOT(I10500)
--	I14342 = NOT(g7582)
--	g8605 = NOT(I14680)
--	I14145 = NOT(g7542)
--	I12256 = NOT(g6647)
--	I14031 = NOT(g7448)
--	g4198 = NOT(I8101)
--	I7044 = NOT(g2402)
--	g6597 = NOT(I11803)
--	g9075 = NOT(I15619)
--	I13451 = NOT(g7262)
--	I13472 = NOT(g7266)
--	I14199 = NOT(g7704)
--	I12280 = NOT(g6684)
--	g3974 = NOT(g3131)
--	I6663 = NOT(g2246)
--	I13628 = NOT(g7248)
--	g8751 = NOT(g8545)
--	g2458 = NOT(g30)
--	I5359 = NOT(g3839)
--	g6784 = NOT(I12223)
--	g2743 = NOT(g1808)
--	g3610 = NOT(g2424)
--	g2890 = NOT(g2264)
--	g5768 = NOT(I10377)
--	I10528 = NOT(g5245)
--	I16033 = NOT(g9282)
--	g8585 = NOT(g7993)
--	g1612 = NOT(I5475)
--	I10393 = NOT(g5196)
--	g7172 = NOT(g7092)
--	g1017 = NOT(I5419)
--	I7712 = NOT(g3657)
--	I14330 = NOT(g7538)
--	g2505 = NOT(g28)
--	g8041 = NOT(g7701)
--	I15962 = NOT(g9218)
--	g2011 = NOT(I5847)
--	g3124 = NOT(g1857)
--	g5806 = NOT(I10451)
--	I5416 = NOT(g8868)
--	g1935 = NOT(g1280)
--	g3980 = NOT(g3192)
--	g6937 = NOT(I12632)
--	g7143 = NOT(g6996)
--	I11591 = NOT(g5814)
--	g2734 = NOT(g2170)
--	g7343 = NOT(I13447)
--	I13776 = NOT(g7497)
--	g9039 = NOT(I15527)
--	g4524 = NOT(g2869)
--	g6294 = NOT(I11209)
--	g6840 = NOT(I12391)
--	g4644 = NOT(I8847)
--	I6590 = NOT(g2467)
--	I13147 = NOT(g7024)
--	g8673 = NOT(I14813)
--	g3540 = NOT(g2424)
--	I15833 = NOT(g9162)
--	g4119 = NOT(I7964)
--	I9837 = NOT(g4781)
--	g6190 = NOT(I10933)
--	g2074 = NOT(I5872)
--	I6657 = NOT(g1701)
--	g6390 = NOT(I11497)
--	g7134 = NOT(I12986)
--	I12885 = NOT(g6946)
--	g7334 = NOT(I13422)
--	I13825 = NOT(g7318)
--	g2992 = NOT(g1833)
--	g4258 = NOT(I8193)
--	I11858 = NOT(g6165)
--	g4577 = NOT(g2914)
--	g6501 = NOT(I11669)
--	g7548 = NOT(I13828)
--	g8669 = NOT(I14801)
--	g4867 = NOT(I9209)
--	I13858 = NOT(g7329)
--	I14709 = NOT(g8198)
--	I10259 = NOT(g5362)
--	g6156 = NOT(I10829)
--	I12511 = NOT(g6598)
--	g6356 = NOT(I11395)
--	g5433 = NOT(g5024)
--	I10708 = NOT(g5545)
--	g7555 = NOT(I13843)
--	g1800 = NOT(g1477)
--	I12763 = NOT(g6686)
--	g3287 = NOT(I6911)
--	g8772 = NOT(g8585)
--	I7885 = NOT(g2837)
--	I5654 = NOT(g921)
--	I8357 = NOT(g1182)
--	I6930 = NOT(g1876)
--	g2573 = NOT(g1649)
--	g2863 = NOT(g1778)
--	g7792 = NOT(I14231)
--	g2480 = NOT(g44)
--	I15613 = NOT(g8996)
--	I9788 = NOT(g4711)
--	g8743 = NOT(g8524)
--	g3849 = NOT(I7350)
--	g6704 = NOT(I12044)
--	I15947 = NOT(g9221)
--	g5845 = NOT(I10548)
--	g4599 = NOT(I8712)
--	g5137 = NOT(I9539)
--	g5395 = NOT(I9840)
--	g8856 = NOT(I15160)
--	g7113 = NOT(I12927)
--	g3898 = NOT(g3160)
--	g8734 = NOT(I14904)
--	g4026 = NOT(g3192)
--	g7313 = NOT(I13369)
--	g4274 = NOT(I8218)
--	g4426 = NOT(I8428)
--	I7036 = NOT(g2454)
--	g6250 = NOT(g5679)
--	g6810 = NOT(I12301)
--	g4614 = NOT(I8757)
--	g6363 = NOT(I11416)
--	g4370 = NOT(I8351)
--	I5978 = NOT(g414)
--	g3510 = NOT(g2185)
--	I10810 = NOT(g5403)
--	g6032 = NOT(g5494)
--	I11446 = NOT(g6062)
--	g4125 = NOT(I7978)
--	I14810 = NOT(g8481)
--	I11227 = NOT(g6130)
--	g6432 = NOT(I11569)
--	g5807 = NOT(I10454)
--	I14657 = NOT(g7782)
--	g7094 = NOT(g6525)
--	I12307 = NOT(g6712)
--	I11025 = NOT(g5638)
--	I12085 = NOT(g5971)
--	g2976 = NOT(I6728)
--	I7335 = NOT(g2910)
--	g1823 = NOT(g768)
--	g7494 = NOT(g7260)
--	g7518 = NOT(I13734)
--	g5266 = NOT(I9782)
--	g6568 = NOT(I11744)
--	g4544 = NOT(g2886)
--	I11203 = NOT(g6129)
--	I5542 = NOT(g1272)
--	I13203 = NOT(g7088)
--	g7776 = NOT(I14199)
--	g1649 = NOT(g1217)
--	I7749 = NOT(g3692)
--	g7593 = NOT(I13924)
--	g3819 = NOT(g1748)
--	g4636 = NOT(I8823)
--	g3694 = NOT(g2174)
--	g2326 = NOT(I6121)
--	I14792 = NOT(g8583)
--	I9520 = NOT(g3995)
--	g6357 = NOT(I11398)
--	g4106 = NOT(I7931)
--	I15507 = NOT(g8968)
--	I12942 = NOT(g7023)
--	g3852 = NOT(I7359)
--	I6471 = NOT(g1923)
--	g3923 = NOT(I7564)
--	g4306 = NOT(I8273)
--	I8778 = NOT(g3922)
--	I11281 = NOT(g5785)
--	I12268 = NOT(g6661)
--	g9320 = NOT(g9307)
--	g5481 = NOT(g4914)
--	g3488 = NOT(g1727)
--	I7947 = NOT(g3485)
--	I13281 = NOT(g7155)
--	g1698 = NOT(I5542)
--	I6242 = NOT(g1554)
--	I16173 = NOT(g9382)
--	I12655 = NOT(g6458)
--	I11377 = NOT(g5811)
--	g7264 = NOT(I13234)
--	g5726 = NOT(I10243)
--	g5154 = NOT(I9588)
--	I10919 = NOT(g5479)
--	I9005 = NOT(g4585)
--	g7160 = NOT(I13054)
--	g7360 = NOT(I13496)
--	I11562 = NOT(g5939)
--	I11645 = NOT(g5874)
--	I13562 = NOT(g7179)
--	g7521 = NOT(I13743)
--	g4622 = NOT(I8781)
--	g4027 = NOT(g2845)
--	g2183 = NOT(I5908)
--	g3951 = NOT(I7648)
--	g7050 = NOT(g6618)
--	I6254 = NOT(g536)
--	g2383 = NOT(I6251)
--	g2924 = NOT(g2314)
--	I12839 = NOT(g6630)
--	I12930 = NOT(g7019)
--	I8949 = NOT(g4116)
--	I7632 = NOT(g3634)
--	I7095 = NOT(g2539)
--	I12993 = NOT(g6933)
--	I10545 = NOT(g5259)
--	g6626 = NOT(I11870)
--	I11290 = NOT(g5818)
--	I13290 = NOT(g7158)
--	I7495 = NOT(g3562)
--	I14079 = NOT(g7579)
--	g4904 = NOT(g4085)
--	g4200 = NOT(I8105)
--	I13698 = NOT(g7348)
--	I7302 = NOT(g2825)
--	I12965 = NOT(g6924)
--	I12131 = NOT(g5918)
--	g9299 = NOT(I16023)
--	I6009 = NOT(g359)
--	g3870 = NOT(g3466)
--	I8998 = NOT(g4576)
--	I5512 = NOT(g557)
--	g4003 = NOT(g3192)
--	I9974 = NOT(g4676)
--	g5112 = NOT(I9496)
--	g3825 = NOT(g1826)
--	g3650 = NOT(I7126)
--	g5267 = NOT(I9785)
--	I12487 = NOT(g6623)
--	g4841 = NOT(g4250)
--	g2161 = NOT(g1454)
--	I8084 = NOT(g3706)
--	g1652 = NOT(g1220)
--	g2361 = NOT(I6183)
--	I7752 = NOT(g3591)
--	I12502 = NOT(g6604)
--	g4191 = NOT(I8084)
--	g1843 = NOT(g771)
--	g8760 = NOT(g8545)
--	g3008 = NOT(g1816)
--	I8850 = NOT(g4031)
--	g2665 = NOT(g1661)
--	g7289 = NOT(I13299)
--	g7777 = NOT(I14202)
--	g6683 = NOT(g6237)
--	g5401 = NOT(I9845)
--	I10125 = NOT(g5127)
--	g4695 = NOT(I8980)
--	I10532 = NOT(g5253)
--	g4637 = NOT(I8826)
--	I5649 = NOT(g1389)
--	g7835 = NOT(I14257)
--	g2327 = NOT(I6124)
--	g5129 = NOT(I9531)
--	g6778 = NOT(I12205)
--	g5761 = NOT(I10356)
--	g3768 = NOT(g2253)
--	I10783 = NOT(g5542)
--	g6894 = NOT(g6525)
--	I13403 = NOT(g7269)
--	I13547 = NOT(g1170)
--	g4307 = NOT(g3700)
--	g4536 = NOT(g2877)
--	g2999 = NOT(g1823)
--	I14783 = NOT(g8324)
--	g3972 = NOT(I7691)
--	g1686 = NOT(I5531)
--	g5828 = NOT(I10509)
--	g2346 = NOT(I6154)
--	g2633 = NOT(g1577)
--	I12469 = NOT(g6586)
--	g9244 = NOT(I15974)
--	I10561 = NOT(g5265)
--	I6229 = NOT(g486)
--	g8608 = NOT(I14687)
--	g8220 = NOT(I14439)
--	I10353 = NOT(g5710)
--	I12286 = NOT(g6696)
--	g6782 = NOT(I12217)
--	I7164 = NOT(g2157)
--	I10295 = NOT(g5523)
--	I8919 = NOT(g4196)
--	g3943 = NOT(I7632)
--	g9140 = NOT(I15784)
--	I9177 = NOT(g4299)
--	g9078 = NOT(I15628)
--	g9340 = NOT(I16090)
--	I13481 = NOT(g7254)
--	g5592 = NOT(g4969)
--	I14680 = NOT(g7810)
--	g6661 = NOT(I11961)
--	g6075 = NOT(g5345)
--	g4016 = NOT(g3192)
--	I8952 = NOT(g4197)
--	g699 = NOT(I5395)
--	I12038 = NOT(g5847)
--	g5746 = NOT(I10295)
--	g6475 = NOT(I11633)
--	g9035 = NOT(I15519)
--	g1670 = NOT(g1489)
--	g3465 = NOT(I6963)
--	g8977 = NOT(I15433)
--	I7296 = NOT(g2915)
--	g3934 = NOT(I7599)
--	g9082 = NOT(I15638)
--	g3230 = NOT(I6887)
--	g4522 = NOT(g2867)
--	g4115 = NOT(I7956)
--	g4251 = NOT(I8180)
--	g6292 = NOT(I11203)
--	I12187 = NOT(g5897)
--	g4811 = NOT(I9158)
--	g4642 = NOT(I8841)
--	g7541 = NOT(I13807)
--	g2944 = NOT(g2363)
--	g2240 = NOT(I5981)
--	g1938 = NOT(g1288)
--	g1813 = NOT(g620)
--	g6646 = NOT(I11920)
--	g7132 = NOT(I12980)
--	I8986 = NOT(g4552)
--	g8665 = NOT(I14789)
--	g7332 = NOT(I13416)
--	I13490 = NOT(g7130)
--	g1909 = NOT(g998)
--	g7353 = NOT(I13475)
--	g6603 = NOT(I11815)
--	g3096 = NOT(I6834)
--	I5872 = NOT(g77)
--	I13956 = NOT(g7499)
--	g5468 = NOT(I9884)
--	g6850 = NOT(I12421)
--	g3496 = NOT(I6974)
--	g7744 = NOT(I14103)
--	g4654 = NOT(I8877)
--	I13103 = NOT(g7055)
--	g3845 = NOT(I7338)
--	g2316 = NOT(I6109)
--	g9214 = NOT(I15918)
--	I5989 = NOT(g1460)
--	I7389 = NOT(g3496)
--	I11824 = NOT(g6283)
--	g5677 = NOT(I10166)
--	I7706 = NOT(g2584)
--	I13888 = NOT(g7335)
--	g3891 = NOT(g3097)
--	I8925 = NOT(g4482)
--	g3913 = NOT(g2834)
--	I10289 = NOT(g5569)
--	g9110 = NOT(I15720)
--	g9310 = NOT(I16046)
--	g6702 = NOT(I12038)
--	g7558 = NOT(I13850)
--	I7888 = NOT(g3505)
--	g4595 = NOT(g2942)
--	g4537 = NOT(g2878)
--	I15927 = NOT(g9208)
--	I7029 = NOT(g2392)
--	g1687 = NOT(g10)
--	I7371 = NOT(g3050)
--	g2347 = NOT(I6157)
--	I12666 = NOT(g6476)
--	g5149 = NOT(I9573)
--	I14288 = NOT(g7705)
--	I14224 = NOT(g7722)
--	I9344 = NOT(g4341)
--	I12217 = NOT(g6631)
--	I7956 = NOT(g2810)
--	g1586 = NOT(g730)
--	I6788 = NOT(g1681)
--	I12478 = NOT(g6603)
--	g2533 = NOT(g1336)
--	g8753 = NOT(I14925)
--	g3859 = NOT(I7380)
--	g4612 = NOT(I8751)
--	g7511 = NOT(I13713)
--	g4017 = NOT(g2845)
--	I15648 = NOT(g9044)
--	g2914 = NOT(g2308)
--	I8277 = NOT(g3504)
--	g5198 = NOT(g4969)
--	I9819 = NOT(g4691)
--	g8072 = NOT(I14349)
--	g9236 = NOT(I15962)
--	g2210 = NOT(g1326)
--	g6616 = NOT(I11848)
--	g4935 = NOT(g4202)
--	g7092 = NOT(I12866)
--	I5670 = NOT(g941)
--	I15604 = NOT(g8993)
--	g7492 = NOT(I13656)
--	I14816 = NOT(g8642)
--	g1570 = NOT(g665)
--	g1860 = NOT(g162)
--	g8443 = NOT(g8015)
--	I6192 = NOT(g327)
--	g7574 = NOT(I13869)
--	g6004 = NOT(g5494)
--	I15770 = NOT(g9121)
--	I10687 = NOT(g5674)
--	g4629 = NOT(I8802)
--	I10976 = NOT(g5726)
--	g6404 = NOT(I11525)
--	I12223 = NOT(g6655)
--	g4328 = NOT(g3086)
--	I14687 = NOT(g7826)
--	g7714 = NOT(I14019)
--	g6647 = NOT(I11923)
--	g4130 = NOT(I7987)
--	g4542 = NOT(g2884)
--	I10752 = NOT(g5618)
--	g3815 = NOT(g1822)
--	I7338 = NOT(g2923)
--	g6764 = NOT(I12161)
--	I14374 = NOT(g7693)
--	I10643 = NOT(g5267)
--	g3692 = NOT(I7198)
--	I13088 = NOT(g7045)
--	g9222 = NOT(I15940)
--	I14643 = NOT(g7837)
--	g2936 = NOT(I6680)
--	g3497 = NOT(g2185)
--	g5524 = NOT(I9938)
--	g7580 = NOT(I13885)
--	g4800 = NOT(I9123)
--	g5644 = NOT(g4748)
--	I15845 = NOT(g9174)
--	g3960 = NOT(I7667)
--	I8892 = NOT(g4115)
--	g1879 = NOT(I5763)
--	g4554 = NOT(g2892)
--	I11497 = NOT(g6014)
--	g9064 = NOT(I15586)
--	I15990 = NOT(g9239)
--	I5552 = NOT(g1284)
--	g7262 = NOT(I13228)
--	g5152 = NOT(I9582)
--	g5258 = NOT(I9774)
--	I14260 = NOT(g7717)
--	g7736 = NOT(I14079)
--	g5818 = NOT(I10479)
--	I10842 = NOT(g5701)
--	g6224 = NOT(I11011)
--	g5577 = NOT(I10046)
--	I14668 = NOT(g7787)
--	I11659 = NOT(g5897)
--	g5717 = NOT(g4969)
--	I13126 = NOT(g6949)
--	I13659 = NOT(g7232)
--	I8945 = NOT(g4106)
--	I11987 = NOT(g6278)
--	g6320 = NOT(I11287)
--	I12373 = NOT(g6763)
--	I6431 = NOT(g1825)
--	I13250 = NOT(g7036)
--	I14489 = NOT(g7829)
--	g2922 = NOT(g2313)
--	g1587 = NOT(g734)
--	g3783 = NOT(I7255)
--	g8013 = NOT(g7561)
--	I10525 = NOT(g5244)
--	I10488 = NOT(g5230)
--	I16061 = NOT(g9294)
--	I10424 = NOT(g5209)
--	g7476 = NOT(g7229)
--	I8709 = NOT(g4191)
--	g3979 = NOT(I7702)
--	I14424 = NOT(g7652)
--	I6376 = NOT(g38)
--	g5186 = NOT(I9684)
--	I10558 = NOT(g5264)
--	I8140 = NOT(g3429)
--	I12936 = NOT(g7015)
--	g9237 = NOT(I15965)
--	I9136 = NOT(g4280)
--	I11296 = NOT(g5831)
--	I9336 = NOT(g4493)
--	g6617 = NOT(I11851)
--	g6789 = NOT(I12238)
--	I13296 = NOT(g7161)
--	g4512 = NOT(g2842)
--	g2460 = NOT(I6302)
--	I7098 = NOT(g2477)
--	I8907 = NOT(g4095)
--	I11338 = NOT(g5798)
--	g7722 = NOT(I14039)
--	I12334 = NOT(g6713)
--	I13338 = NOT(g7190)
--	I9594 = NOT(g4718)
--	I7498 = NOT(g2752)
--	g5026 = NOT(I9366)
--	I6286 = NOT(g1307)
--	g3676 = NOT(g2380)
--	g9194 = NOT(g9182)
--	g5426 = NOT(g5013)
--	I6911 = NOT(g1869)
--	I8517 = NOT(g3014)
--	g7285 = NOT(I13287)
--	g2784 = NOT(g2340)
--	g5170 = NOT(I9636)
--	g3761 = NOT(g1772)
--	g4056 = NOT(g3082)
--	g7500 = NOT(I13676)
--	I11060 = NOT(g5453)
--	g9089 = NOT(I15657)
--	I13060 = NOT(g6959)
--	g6299 = NOT(I11224)
--	g5821 = NOT(I10488)
--	I11197 = NOT(g6122)
--	g3828 = NOT(I7287)
--	g4649 = NOT(I8862)
--	I7584 = NOT(g3062)
--	I11855 = NOT(g5751)
--	I6733 = NOT(g1718)
--	g3830 = NOT(I7293)
--	I6974 = NOT(g2528)
--	I15388 = NOT(g8898)
--	I15324 = NOT(g8779)
--	I6270 = NOT(g492)
--	g2937 = NOT(g2346)
--	I11870 = NOT(g5752)
--	g7139 = NOT(I12999)
--	g9071 = NOT(I15607)
--	g5939 = NOT(I10579)
--	I10705 = NOT(g5463)
--	g6892 = NOT(I12547)
--	g1832 = NOT(g763)
--	g2479 = NOT(g32)
--	g7339 = NOT(I13435)
--	I13527 = NOT(g7217)
--	g2668 = NOT(g1662)
--	I14042 = NOT(g7470)
--	g1853 = NOT(g766)
--	g2840 = NOT(g2207)
--	g4698 = NOT(I8989)
--	g8775 = NOT(g8564)
--	g3746 = NOT(g2100)
--	g5083 = NOT(g4457)
--	g7838 = NOT(I14264)
--	I5879 = NOT(g1267)
--	g7024 = NOT(I12782)
--	g7424 = NOT(I13547)
--	I7362 = NOT(g2933)
--	I12909 = NOT(g7046)
--	I14270 = NOT(g7703)
--	g7737 = NOT(I14082)
--	I10678 = NOT(g5566)
--	I6124 = NOT(g399)
--	g8581 = NOT(g8094)
--	I14124 = NOT(g7591)
--	g6945 = NOT(I12646)
--	I12117 = NOT(g5918)
--	g1794 = NOT(I5646)
--	I11503 = NOT(g6220)
--	g2501 = NOT(g27)
--	I11867 = NOT(g6286)
--	I11894 = NOT(g5956)
--	I10460 = NOT(g5219)
--	I13894 = NOT(g7353)
--	g4463 = NOT(I8483)
--	I14460 = NOT(g7789)
--	g6244 = NOT(g5670)
--	g7077 = NOT(g6676)
--	I9496 = NOT(g3971)
--	g7231 = NOT(I13173)
--	g3932 = NOT(I7595)
--	g5790 = NOT(I10415)
--	g7523 = NOT(I13749)
--	I9845 = NOT(g4728)
--	g6140 = NOT(I10783)
--	g3953 = NOT(g3160)
--	g6340 = NOT(I11347)
--	I11714 = NOT(g5772)
--	g9350 = NOT(I16100)
--	g5187 = NOT(I9687)
--	g5061 = NOT(I9425)
--	I14267 = NOT(g7695)
--	I14294 = NOT(g7553)
--	g6478 = NOT(I11638)
--	g8784 = NOT(g8545)
--	g2942 = NOT(g2350)
--	g5461 = NOT(g4885)
--	g4279 = NOT(g3340)
--	I11707 = NOT(g5988)
--	g7205 = NOT(I13131)
--	I13707 = NOT(g7420)
--	I13819 = NOT(g7426)
--	g5756 = NOT(I10343)
--	g6035 = NOT(g5494)
--	g6959 = NOT(I12678)
--	I7728 = NOT(g3675)
--	I11257 = NOT(g5805)
--	g5622 = NOT(g4938)
--	g4619 = NOT(I8772)
--	g5027 = NOT(I9369)
--	g6517 = NOT(I11701)
--	I11818 = NOT(g6276)
--	g3677 = NOT(g2485)
--	g5427 = NOT(g5115)
--	I15871 = NOT(g9184)
--	I11055 = NOT(g5696)
--	I13979 = NOT(g7415)
--	I5374 = NOT(g634)
--	I13496 = NOT(g7133)
--	g7742 = NOT(I14097)
--	g4652 = NOT(I8871)
--	g7551 = NOT(I13837)
--	g7104 = NOT(I12900)
--	g6876 = NOT(I12499)
--	g7099 = NOT(I12885)
--	g4057 = NOT(I7832)
--	g7304 = NOT(I13344)
--	g8668 = NOT(I14798)
--	I11978 = NOT(g6186)
--	I6849 = NOT(g368)
--	g3866 = NOT(g2945)
--	g2954 = NOT(g2374)
--	g4457 = NOT(I8477)
--	g7499 = NOT(g7258)
--	I8877 = NOT(g4274)
--	g2810 = NOT(g1922)
--	g2363 = NOT(I6189)
--	g6656 = NOT(I11948)
--	g9212 = NOT(I15912)
--	I12639 = NOT(g6506)
--	I16151 = NOT(g9369)
--	g3716 = NOT(g2522)
--	g5514 = NOT(g4922)
--	I5545 = NOT(g1276)
--	g5403 = NOT(g5088)
--	g5145 = NOT(I9561)
--	g2453 = NOT(I6291)
--	I5380 = NOT(g645)
--	g5841 = NOT(I10538)
--	g3848 = NOT(I7347)
--	g1750 = NOT(g602)
--	I6900 = NOT(g1866)
--	I12265 = NOT(g6660)
--	g7754 = NOT(I14133)
--	I10160 = NOT(g5139)
--	g5763 = NOT(I10366)
--	I9142 = NOT(g4236)
--	g5191 = NOT(g4969)
--	g8156 = NOT(I14394)
--	g3855 = NOT(I7368)
--	I14160 = NOT(g7549)
--	g3398 = NOT(I6952)
--	I8928 = NOT(g4153)
--	g7273 = NOT(I13255)
--	I6245 = NOT(g142)
--	I9081 = NOT(g4357)
--	I12391 = NOT(g6744)
--	g4598 = NOT(I8709)
--	g6110 = NOT(g5335)
--	g6310 = NOT(I11257)
--	I6291 = NOT(g46)
--	g7044 = NOT(g6543)
--	I10617 = NOT(g5677)
--	I15628 = NOT(g9001)
--	g4121 = NOT(I7970)
--	I5559 = NOT(g1292)
--	g2157 = NOT(I5897)
--	g7269 = NOT(I13247)
--	g6663 = NOT(I11967)
--	g4670 = NOT(I8925)
--	g5159 = NOT(I9603)
--	g4625 = NOT(I8790)
--	g7983 = NOT(I14294)
--	I10277 = NOT(g5472)
--	I11018 = NOT(g5626)
--	I13196 = NOT(g7008)
--	I7635 = NOT(g3052)
--	I13695 = NOT(g7345)
--	g6824 = NOT(I12343)
--	g7712 = NOT(I14015)
--	g1666 = NOT(g1472)
--	g3524 = NOT(g2306)
--	g4253 = NOT(g2734)
--	g2929 = NOT(g2327)
--	g4938 = NOT(I9310)
--	g6236 = NOT(I11037)
--	g4813 = NOT(I9162)
--	I12586 = NOT(g6643)
--	g7543 = NOT(I13813)
--	g5016 = NOT(I9350)
--	g5757 = NOT(g5261)
--	g8810 = NOT(I15068)
--	g3644 = NOT(g2131)
--	I7305 = NOT(g3048)
--	g8363 = NOT(g7992)
--	I15776 = NOT(g9127)
--	I16058 = NOT(g9294)
--	I10494 = NOT(g5232)
--	g4909 = NOT(I9271)
--	I12442 = NOT(g6542)
--	I5515 = NOT(g567)
--	I14623 = NOT(g7833)
--	I8844 = NOT(g3992)
--	g5522 = NOT(g4930)
--	g5115 = NOT(I9505)
--	g6877 = NOT(I12502)
--	g5811 = NOT(I10466)
--	g5642 = NOT(I10125)
--	g2626 = NOT(g1571)
--	g3577 = NOT(g2372)
--	g7534 = NOT(I13782)
--	g7729 = NOT(I14058)
--	g3867 = NOT(g2946)
--	I15950 = NOT(g9222)
--	I13457 = NOT(g7120)
--	g1655 = NOT(g1231)
--	g6657 = NOT(I11951)
--	I7755 = NOT(g3019)
--	g4552 = NOT(g2890)
--	g9062 = NOT(I15580)
--	I11917 = NOT(g5897)
--	g4606 = NOT(I8733)
--	g6556 = NOT(I11732)
--	I10418 = NOT(g5453)
--	g6222 = NOT(g5654)
--	I12041 = NOT(g5897)
--	g5874 = NOT(I10565)
--	I9001 = NOT(g4577)
--	I14822 = NOT(g8649)
--	g7014 = NOT(I12760)
--	g4687 = NOT(I8962)
--	I8966 = NOT(g4444)
--	I12430 = NOT(g6432)
--	I11001 = NOT(g5698)
--	g5654 = NOT(g4748)
--	I12493 = NOT(g6587)
--	g7414 = NOT(I13527)
--	I9129 = NOT(g4475)
--	I15394 = NOT(g8916)
--	g3975 = NOT(g3131)
--	g6064 = NOT(I10681)
--	g4586 = NOT(g2926)
--	g6899 = NOT(g6525)
--	g2683 = NOT(g1666)
--	g6785 = NOT(I12226)
--	I11689 = NOT(g5956)
--	I11923 = NOT(g5939)
--	I12340 = NOT(g6725)
--	I12983 = NOT(g6930)
--	g7513 = NOT(I13719)
--	I5969 = NOT(g303)
--	I12806 = NOT(g6602)
--	I12684 = NOT(g6472)
--	I7602 = NOT(g2562)
--	g2894 = NOT(g2267)
--	I15420 = NOT(g8881)
--	g4570 = NOT(g2907)
--	g4341 = NOT(I8308)
--	g9298 = NOT(I16020)
--	g9085 = NOT(I15645)
--	I8814 = NOT(g4028)
--	g1667 = NOT(g1481)
--	g4525 = NOT(g2870)
--	g4710 = NOT(I9009)
--	g7178 = NOT(I13088)
--	g2782 = NOT(g1616)
--	g6295 = NOT(I11212)
--	g1235 = NOT(I5422)
--	g5612 = NOT(g4814)
--	I12517 = NOT(g6613)
--	g6237 = NOT(I11040)
--	g4645 = NOT(I8850)
--	I13157 = NOT(g6997)
--	g2661 = NOT(I6454)
--	g5417 = NOT(g5006)
--	g1566 = NOT(g652)
--	g7135 = NOT(I12989)
--	g6844 = NOT(I12403)
--	g7335 = NOT(I13425)
--	I11066 = NOT(g5460)
--	I13066 = NOT(g6957)
--	I13231 = NOT(g6897)
--	g7288 = NOT(I13296)
--	g6194 = NOT(I10937)
--	I5528 = NOT(g43)
--	g2627 = NOT(g1572)
--	I14118 = NOT(g7565)
--	g5128 = NOT(I9528)
--	I9624 = NOT(g4746)
--	g2292 = NOT(I6060)
--	I14022 = NOT(g7443)
--	g6089 = NOT(g5317)
--	I12193 = NOT(g6468)
--	g6731 = NOT(I12101)
--	g4607 = NOT(I8736)
--	I8769 = NOT(g3999)
--	I13876 = NOT(g7347)
--	I13885 = NOT(g7351)
--	g5542 = NOT(g5061)
--	g7022 = NOT(I12776)
--	g2646 = NOT(I6422)
--	g7422 = NOT(I13541)
--	g4659 = NOT(I8892)
--	g7749 = NOT(I14118)
--	g1555 = NOT(I5428)
--	I12523 = NOT(g6624)
--	g4358 = NOT(g3680)
--	g1804 = NOT(I5664)
--	I6887 = NOT(g2528)
--	g8683 = NOT(g8235)
--	I13854 = NOT(g7327)
--	g6071 = NOT(I10694)
--	g9219 = NOT(I15933)
--	g1792 = NOT(g616)
--	g2039 = NOT(g1228)
--	g3061 = NOT(I6795)
--	g3187 = NOT(I6860)
--	g6471 = NOT(I11627)
--	g8778 = NOT(I14974)
--	I14276 = NOT(g7720)
--	I14285 = NOT(g7625)
--	g2484 = NOT(g45)
--	g9031 = NOT(I15507)
--	g5800 = NOT(I10439)
--	I5410 = NOT(g8866)
--	g3461 = NOT(I6959)
--	g6242 = NOT(I11047)
--	I14305 = NOT(g7537)
--	g9252 = NOT(I15982)
--	g4587 = NOT(g2928)
--	I12475 = NOT(g6596)
--	I6033 = NOT(g3)
--	I9576 = NOT(g4706)
--	I10466 = NOT(g5221)
--	g6948 = NOT(I12655)
--	g4111 = NOT(I7944)
--	I5839 = NOT(g1198)
--	g7560 = NOT(I13854)
--	g4275 = NOT(g3790)
--	g4311 = NOT(I8282)
--	g9376 = NOT(I16154)
--	I15738 = NOT(g9079)
--	I15562 = NOT(g8979)
--	I15645 = NOT(g9043)
--	g6955 = NOT(I12666)
--	g4615 = NOT(I8760)
--	g3904 = NOT(g3160)
--	g8661 = NOT(I14777)
--	I10177 = NOT(g4721)
--	I15699 = NOT(g9061)
--	I6096 = NOT(g521)
--	g6254 = NOT(g5683)
--	g6814 = NOT(I12313)
--	g7095 = NOT(I12877)
--	g3514 = NOT(g2424)
--	g2919 = NOT(g2311)
--	g7037 = NOT(g6525)
--	g6150 = NOT(g5287)
--	g7495 = NOT(I13663)
--	g1908 = NOT(g812)
--	g7437 = NOT(I13570)
--	g6350 = NOT(I11377)
--	g7102 = NOT(I12894)
--	g7208 = NOT(I13140)
--	I6195 = NOT(g405)
--	g7302 = NOT(I13338)
--	I13550 = NOT(g1173)
--	g6038 = NOT(I10649)
--	I5667 = NOT(g916)
--	I11314 = NOT(g5781)
--	I6337 = NOT(g1348)
--	g3841 = NOT(I7326)
--	I13314 = NOT(g7160)
--	I11287 = NOT(g5806)
--	g2276 = NOT(I6029)
--	I12253 = NOT(g6427)
--	g6773 = NOT(I12190)
--	I13287 = NOT(g7157)
--	g1567 = NOT(g655)
--	I16103 = NOT(g9339)
--	g7579 = NOT(I13882)
--	I14064 = NOT(g7556)
--	g6009 = NOT(I10605)
--	g3191 = NOT(I6868)
--	g4545 = NOT(g2887)
--	g2616 = NOT(g1564)
--	g7719 = NOT(g7475)
--	g2561 = NOT(g1555)
--	g5490 = NOT(g4917)
--	g691 = NOT(I5389)
--	g5823 = NOT(I10494)
--	g534 = NOT(I5365)
--	g5166 = NOT(I9624)
--	I11596 = NOT(g6228)
--	g4591 = NOT(g2937)
--	g8603 = NOT(I14674)
--	I13054 = NOT(g6960)
--	g8039 = NOT(g7696)
--	g1776 = NOT(g608)
--	g6769 = NOT(I12176)
--	g7752 = NOT(I14127)
--	I11431 = NOT(g5782)
--	g9073 = NOT(I15613)
--	g6836 = NOT(I12379)
--	g4020 = NOT(I7781)
--	g6212 = NOT(I10973)
--	g2404 = NOT(g1276)
--	I5548 = NOT(g1280)
--	I8895 = NOT(g4130)
--	g2647 = NOT(I6425)
--	g5529 = NOT(g4689)
--	g3159 = NOT(I6856)
--	I10166 = NOT(g5016)
--	g5148 = NOT(I9570)
--	g3359 = NOT(I6946)
--	g5649 = NOT(g4748)
--	g6918 = NOT(I12609)
--	g6967 = NOT(I12696)
--	I5555 = NOT(g1288)
--	I11269 = NOT(g5756)
--	I14166 = NOT(g7702)
--	I14009 = NOT(g7436)
--	g2764 = NOT(g1802)
--	g7265 = NOT(g7077)
--	g9324 = NOT(I16072)
--	g7042 = NOT(g6543)
--	g2546 = NOT(I6368)
--	I11773 = NOT(g6262)
--	g5155 = NOT(I9591)
--	g4559 = NOT(g2898)
--	g9069 = NOT(I15601)
--	I11942 = NOT(g6015)
--	I11341 = NOT(g5809)
--	I13773 = NOT(g7496)
--	g3858 = NOT(I7377)
--	g7442 = NOT(I13583)
--	g8583 = NOT(I14668)
--	I13341 = NOT(g7207)
--	g4931 = NOT(I9301)
--	I6248 = NOT(g411)
--	I7564 = NOT(g2752)
--	I9258 = NOT(g4249)
--	g3757 = NOT(g1977)
--	g2970 = NOT(g2394)
--	g6229 = NOT(g5665)
--	I15481 = NOT(g8913)
--	I10485 = NOT(g5229)
--	g6993 = NOT(I12731)
--	g1933 = NOT(g1247)
--	g7164 = NOT(I13066)
--	g7364 = NOT(I13506)
--	I6081 = NOT(g118)
--	g2925 = NOT(g2324)
--	g9177 = NOT(I15811)
--	g7233 = NOT(g6940)
--	g9206 = NOT(g9196)
--	I10555 = NOT(g5529)
--	I10454 = NOT(g5217)
--	g6822 = NOT(I12337)
--	g3522 = NOT(g2407)
--	I14454 = NOT(g8177)
--	g7054 = NOT(g6511)
--	g2224 = NOT(I5945)
--	g3642 = NOT(I7118)
--	I13734 = NOT(g7422)
--	g3047 = NOT(g1736)
--	I10914 = NOT(g5448)
--	I11335 = NOT(g5839)
--	g7454 = NOT(I13610)
--	g4628 = NOT(I8799)
--	I14712 = NOT(g8059)
--	I13335 = NOT(g7206)
--	g7770 = NOT(I14181)
--	g5463 = NOT(g5085)
--	I6154 = NOT(g122)
--	g7296 = NOT(I13320)
--	I6354 = NOT(g1357)
--	g4630 = NOT(I8805)
--	I13930 = NOT(g7405)
--	g7725 = NOT(I14046)
--	I11838 = NOT(g6281)
--	I5908 = NOT(g196)
--	g4300 = NOT(I8261)
--	g7532 = NOT(I13776)
--	g1724 = NOT(I5568)
--	I7308 = NOT(g3074)
--	g3874 = NOT(g2957)
--	I12208 = NOT(g6496)
--	I13131 = NOT(g6951)
--	g3654 = NOT(g2521)
--	g9199 = NOT(g9188)
--	I15784 = NOT(g9125)
--	g8647 = NOT(I14739)
--	I15956 = NOT(g9216)
--	g2617 = NOT(g1565)
--	g2906 = NOT(g2288)
--	I15385 = NOT(g8880)
--	g1878 = NOT(g80)
--	g5167 = NOT(I9627)
--	I14238 = NOT(g7608)
--	g5367 = NOT(I9834)
--	g5872 = NOT(I10561)
--	I13487 = NOT(g7129)
--	
--	g7412 = AND(g7121, g4841)
--	g6462 = AND(g6215, g2424)
--	g8925 = AND(g4592, g8754)
--	g4969 = AND(g4362, g2216)
--	g7429 = AND(g1057, g7212)
--	g9144 = AND(g9123, g6096)
--	g9344 = AND(g9329, g6211)
--	g4123 = AND(g2627, g2617)
--	g8320 = AND(g4557, g7951)
--	I8431 = AND(g3430, g3398, g3359, g3341)
--	g9259 = AND(g9230, g5639)
--	g8277 = AND(g162, g8042)
--	I8005 = AND(g3430, g3398, g3359, g2106)
--	g4351 = AND(g309, g3131)
--	g8299 = AND(g591, g8181)
--	g6941 = AND(g1126, g6582)
--	g4410 = AND(g408, g3160)
--	g8892 = AND(g8681, g4969)
--	I7994 = AND(g3430, g3398, g3359, g3341)
--	g5552 = AND(g1114, g4832)
--	g8945 = AND(g4541, g8784)
--	g8738 = AND(g8619, g3338)
--	g6431 = AND(g5847, g5494)
--	g4172 = AND(I8057, I8058)
--	g7449 = AND(g7272, g6901)
--	g8709 = AND(g2818, g8386)
--	g6176 = AND(g1149, g5198)
--	g6005 = AND(g5557, g2407)
--	g4343 = AND(g306, g3131)
--	g8078 = AND(g7463, g7634)
--	g8340 = AND(g423, g7920)
--	g6405 = AND(g5956, g5494)
--	g4282 = AND(g3549, g3568)
--	g7604 = AND(g7456, g3466)
--	g1714 = AND(g1454, g1450)
--	g5570 = AND(g1759, g4841)
--	g8690 = AND(g3485, g8363)
--	g7833 = AND(g6461, g7601)
--	g4334 = AND(g225, g3097)
--	g8876 = AND(g8769, g6102)
--	g6733 = AND(g685, g5873)
--	g6974 = AND(g3613, g6505)
--	g4804 = AND(g952, g3876)
--	g8915 = AND(g8794, g8239)
--	g7419 = AND(g7230, g3530)
--	g8310 = AND(g573, g8181)
--	g4494 = AND(I8546, I8547)
--	g8824 = AND(g264, g8524)
--	g8877 = AND(g8773, g6104)
--	g6399 = AND(g5971, g5494)
--	I9330 = AND(g2784, g2770, g2746)
--	g9142 = AND(g9124, g6059)
--	g8928 = AND(g4595, g8757)
--	g5020 = AND(g579, g3937)
--	g4933 = AND(g2746, g2728, g4320, g2770)
--	g8930 = AND(g3866, g8760)
--	I8114 = AND(g2162, g2149, g2137, g2106)
--	g8064 = AND(g7483, g7634)
--	g7678 = AND(g7367, g4158)
--	g4724 = AND(g828, g4038)
--	g7087 = AND(g6440, g5311)
--	g4379 = AND(g399, g3160)
--	g8295 = AND(g4512, g7905)
--	g8237 = AND(g89, g8131)
--	g6923 = AND(g6570, g5612)
--	g4878 = AND(g2573, g2562, I9222)
--	g8844 = AND(g4056, g8602)
--	I8594 = AND(g3316, g2057, g2020, g1987)
--	I9166 = AND(g4041, g2595, g2584)
--	g8089 = AND(g840, g7658)
--	g8731 = AND(g2743, g8421)
--	g4271 = AND(g3666, g3684)
--	g6951 = AND(g5511, g6595)
--	g8071 = AND(g7540, g4969)
--	g8705 = AND(g2798, g8421)
--	g4799 = AND(g951, g4596)
--	I8033 = AND(g3430, g3398, g3359, g2106)
--	g8948 = AND(g4570, g8789)
--	g5969 = AND(g5564, g2424)
--	g7602 = AND(g7476, g3466)
--	g7007 = AND(g6627, g5072)
--	g5123 = AND(g516, g4033)
--	g4132 = AND(g2637, g2633)
--	I8496 = AND(g3316, g3287, g2020, g1987)
--	g4238 = AND(g2695, g2698, I8157)
--	g8814 = AND(g3880, g8463)
--	g6408 = AND(g669, g6019)
--	g8150 = AND(g846, g7658)
--	g4744 = AND(g3525, g4296)
--	g8438 = AND(g649, g7793)
--	g6972 = AND(g5661, g6498)
--	g7415 = AND(g7222, g5603)
--	g8836 = AND(g348, g8545)
--	g4901 = AND(g3723, g4288, I9261)
--	g6433 = AND(g778, g6134)
--	g8229 = AND(g8180, g5680)
--	g9349 = AND(g9340, g5690)
--	g8822 = AND(g417, g8564)
--	g6395 = AND(g2157, g6007)
--	g8921 = AND(g4579, g8747)
--	g7689 = AND(g7367, g4417)
--	g5334 = AND(g4887, g2424)
--	g5548 = AND(g1549, g4826)
--	g4968 = AND(g4403, g1760)
--	g6266 = AND(g1481, g5285)
--	g8837 = AND(g426, g8564)
--	g7030 = AND(g6705, g5723)
--	g8062 = AND(g7476, g7634)
--	g8620 = AND(g751, g8199)
--	g8462 = AND(g49, g8199)
--	g9119 = AND(g9049, g5345)
--	I8001 = AND(g2074, g3287, g2020, g1987)
--	g7564 = AND(g7367, g4172)
--	g9258 = AND(g9227, g5628)
--	I8401 = AND(g3316, g3287, g3264, g3238)
--	g4175 = AND(g1110, g3502)
--	g4375 = AND(g219, g3097)
--	g5313 = AND(g4820, g2407)
--	g6726 = AND(g5897, g5367)
--	g6154 = AND(g1499, g5713)
--	g8842 = AND(g429, g8564)
--	g7609 = AND(g7467, g3466)
--	g8298 = AND(g553, g8181)
--	g5094 = AND(g535, g4004)
--	g9274 = AND(g4748, g9255)
--	g4139 = AND(I8000, I8001)
--	g4384 = AND(g246, g3097)
--	g4838 = AND(g4517, g1760)
--	g8854 = AND(g443, g8564)
--	g7217 = AND(g1142, g6941)
--	g8941 = AND(g3882, g8776)
--	g4424 = AND(g489, g3192)
--	g6979 = AND(g5095, g6511)
--	g5593 = AND(g4110, g4969)
--	g6112 = AND(g5673, g4841, g5541)
--	g4077 = AND(g1284, g3582)
--	g6001 = AND(g5540, g2407)
--	g6401 = AND(g5971, g5367)
--	g8708 = AND(g3557, g8407)
--	g7827 = AND(g7575, g7173)
--	g5050 = AND(g587, g3970)
--	g1725 = AND(g1409, g1416)
--	g6727 = AND(g681, g5846)
--	g8405 = AND(g741, g8018)
--	g4099 = AND(g117, g3647)
--	g4304 = AND(g2784, g3779)
--	g8829 = AND(g267, g8524)
--	g8286 = AND(g180, g8156)
--	g8911 = AND(g8798, g7688)
--	g8733 = AND(g2996, g8493)
--	g8270 = AND(g110, g8131)
--	g8610 = AND(g665, g7887)
--	g9345 = AND(g9330, g6217)
--	g4269 = AND(g2354, g3563, I8209)
--	I8524 = AND(g3316, g2057, g3264, g1987)
--	g2781 = AND(g1600, g976)
--	g8069 = AND(g7456, g7634)
--	g4712 = AND(g1179, g4276)
--	g7181 = AND(g6124, g7039)
--	g9159 = AND(g9138, g6074)
--	g9359 = AND(g4748, g9340)
--	g8377 = AND(g507, g7966)
--	g7197 = AND(g7093, g5055)
--	g7700 = AND(g7367, g4494)
--	g7021 = AND(g3390, g6673)
--	g4729 = AND(g1504, g4059)
--	g4961 = AND(g377, g3904)
--	g9016 = AND(g8904, g8239)
--	g8287 = AND(g4500, g7855)
--	I8186 = AND(g3778, g3549, g3568, g3583)
--	g5132 = AND(I9534, I9535)
--	g8849 = AND(g513, g8585)
--	I7995 = AND(g2074, g3287, g2020, g3238)
--	g9251 = AND(g4748, g9230)
--	g4414 = AND(I8412, I8413)
--	g3313 = AND(g2334, g2316, g2298)
--	g7631 = AND(g7367, g4187)
--	g8291 = AND(g122, g8111)
--	g3094 = AND(g945, g1898)
--	g4436 = AND(g492, g3192)
--	g6577 = AND(g6142, g4160)
--	g7605 = AND(g7435, g5607)
--	g4378 = AND(g321, g3131)
--	g4135 = AND(I7994, I7995)
--	g5092 = AND(g456, g4002)
--	g4182 = AND(I8071, I8072)
--	g4288 = AND(g3563, g3579, g3603, I8240)
--	g9272 = AND(g4748, g9248)
--	g8259 = AND(g4538, g7855)
--	g5714 = AND(g1532, g4733)
--	g8088 = AND(g837, g7658)
--	g8852 = AND(g362, g8545)
--	g8923 = AND(g4587, g8751)
--	I8461 = AND(g3316, g3287, g2020, g3238)
--	g7041 = AND(g6734, g5206)
--	g4422 = AND(g411, g3160)
--	g8701 = AND(g2700, g8363)
--	g2768 = AND(g1597, g973)
--	g9328 = AND(g9324, g6465)
--	g4798 = AND(g4216, g1760)
--	g9130 = AND(g9054, g5345)
--	g6125 = AND(g5548, g4202)
--	g2972 = AND(g2397, g2407)
--	I8046 = AND(g2074, g2057, g3264, g1987)
--	g8951 = AND(g8785, g6072)
--	g8314 = AND(g443, g7920)
--	g4437 = AND(g540, g2845)
--	g8825 = AND(g342, g8545)
--	g8650 = AND(g591, g8094)
--	g4302 = AND(g3086, g3659, g3124)
--	g1728 = AND(g1432, g1439)
--	g8336 = AND(g420, g7920)
--	g6061 = AND(g5257, g1616)
--	g8943 = AND(g4560, g8781)
--	g6046 = AND(g1073, g5592)
--	I8115 = AND(g2074, g3287, g3264, g1987)
--	I8642 = AND(g3430, g3398, g3359, g2106)
--	g8322 = AND(g4559, g7993)
--	g6003 = AND(g3716, g5633, I10597)
--	g8934 = AND(g3873, g8766)
--	g9348 = AND(g9333, g6229)
--	g7713 = AND(g4403, g7367)
--	g6145 = AND(g1489, g5705)
--	g4054 = AND(g3767, g2424)
--	g4454 = AND(g544, g2845)
--	g5077 = AND(g236, g3988)
--	g4532 = AND(I8617, I8618)
--	g6107 = AND(g5478, g1849)
--	g8845 = AND(g432, g8564)
--	I9202 = AND(g2605, g4044, g2584)
--	g8337 = AND(g498, g7966)
--	g4412 = AND(g486, g3192)
--	g5104 = AND(g274, g4010)
--	g6757 = AND(g5874, g5412)
--	g9279 = AND(g9255, g5665)
--	g4389 = AND(g480, g3192)
--	I8612 = AND(g3430, g3398, g3359, g3341)
--	g6416 = AND(g710, g6026)
--	I8417 = AND(g3430, g3398, g3359, g2106)
--	g9118 = AND(g9046, g5345)
--	g4787 = AND(g953, g4547)
--	g6047 = AND(g1477, g5596)
--	g8266 = AND(g2157, g8042)
--	g6447 = AND(g734, g6073)
--	g4956 = AND(g295, g3892)
--	g2979 = AND(g1494, g1733)
--	g5044 = AND(g234, g3959)
--	g8081 = AND(g834, g7658)
--	g8815 = AND(g258, g8524)
--	g7183 = AND(g6132, g7042)
--	g7608 = AND(g7367, g4169)
--	g8692 = AND(g3462, g8363)
--	g8726 = AND(g2795, g8386)
--	g4138 = AND(g2638, g2634)
--	g4109 = AND(g990, g3790)
--	g4791 = AND(g949, g4562)
--	g4707 = AND(g812, g4062)
--	g6417 = AND(g718, g6027)
--	I8090 = AND(g3316, g2057, g2020, g3238)
--	I8490 = AND(g3430, g3398, g3359, g3341)
--	g4201 = AND(I8108, I8109)
--	g8267 = AND(g154, g8042)
--	g8312 = AND(g365, g7870)
--	g6629 = AND(g6023, g4841)
--	g4957 = AND(g2746, g2728, g4320)
--	g4049 = AND(g141, g3514)
--	I8456 = AND(g3316, g3287, g2020, g1987)
--	I8529 = AND(g3316, g2057, g3264, g3238)
--	g8293 = AND(g4510, g7855)
--	g8329 = AND(g527, g7966)
--	g7696 = AND(g7367, g4469)
--	g5513 = AND(g4889, g5071)
--	g4098 = AND(g985, g3790)
--	g6554 = AND(g5762, g1616)
--	g8828 = AND(g4573, g8541)
--	g8830 = AND(g345, g8545)
--	g8727 = AND(g2724, g8421)
--	g5436 = AND(g1541, g4926)
--	g7240 = AND(g6719, g6894)
--	I8063 = AND(g2162, g2149, g2137, g2106)
--	g8703 = AND(g3574, g8407)
--	g4268 = AND(g2216, g2655)
--	g8932 = AND(g3868, g8762)
--	g6166 = AND(g1509, g5725)
--	g8624 = AND(g754, g8199)
--	g8953 = AND(g8758, g6093)
--	g4052 = AND(g1276, g3522)
--	g8068 = AND(g7687, g5610)
--	g4452 = AND(g437, g3160)
--	g6056 = AND(g3760, g5286, g1695)
--	g6456 = AND(g6116, g2407)
--	I8057 = AND(g3430, g3398, g3359, g3341)
--	g7681 = AND(g7444, g5099)
--	g9158 = AND(g9137, g6070)
--	g5560 = AND(g3390, g5036)
--	g4086 = AND(g103, g3629)
--	g4728 = AND(g190, g4179)
--	g4486 = AND(I8528, I8529)
--	g8716 = AND(g3506, g8443)
--	g7596 = AND(g7428, g7028)
--	g4504 = AND(I8568, I8569)
--	g4185 = AND(g2636, g2632)
--	g9275 = AND(g9241, g5645)
--	g4385 = AND(g300, g3131)
--	g8848 = AND(g281, g8524)
--	g5579 = AND(g4090, g4841)
--	g4425 = AND(g536, g2845)
--	g2386 = AND(g1130, g1092)
--	g5442 = AND(g4679, g4202)
--	g6057 = AND(g1061, g5617)
--	g4131 = AND(g2630, g2622)
--	g8319 = AND(g255, g7838)
--	I8552 = AND(g3316, g2057, g3264, g1987)
--	g8258 = AND(g142, g8111)
--	g6971 = AND(g6424, g4969)
--	g8717 = AND(g2764, g8421)
--	g7597 = AND(g7316, g4841)
--	g7079 = AND(g4259, g6677)
--	g8274 = AND(g4580, g7951)
--	g4445 = AND(I8455, I8456)
--	g4091 = AND(g129, g3639)
--	g4491 = AND(g557, g2845)
--	g8325 = AND(g184, g8156)
--	g8821 = AND(g339, g8545)
--	g4169 = AND(I8052, I8053)
--	g5029 = AND(g212, g3945)
--	g4369 = AND(g580, g2845)
--	g8280 = AND(g114, g8111)
--	g8939 = AND(g3879, g8772)
--	g4407 = AND(g252, g3097)
--	g4059 = AND(g1499, g2979)
--	g4868 = AND(g4227, g4160)
--	g8306 = AND(g4525, g7951)
--	g4793 = AND(g3887, g4202)
--	g8461 = AND(g658, g7793)
--	g8622 = AND(g738, g7811)
--	g4246 = AND(g1106, g3226)
--	g8403 = AND(g639, g7793)
--	g8841 = AND(g351, g8545)
--	g5049 = AND(g474, g3969)
--	I8020 = AND(g2074, g3287, g2020, g1987)
--	g8695 = AND(g2709, g8363)
--	g8307 = AND(g432, g7920)
--	g9278 = AND(g9252, g5658)
--	g4388 = AND(g402, g3160)
--	g8359 = AND(g642, g7793)
--	g4216 = AND(I8114, I8115)
--	g9143 = AND(g9122, g6089)
--	g9343 = AND(g9328, g1738)
--	g7626 = AND(g7463, g3466)
--	g8858 = AND(g524, g8585)
--	g4430 = AND(I8436, I8437)
--	I9534 = AND(g3019, g3029, g3038, g3052)
--	g9334 = AND(g9318, g6205)
--	g8315 = AND(g4544, g7993)
--	g4826 = AND(g1545, g4239)
--	g6239 = AND(g1514, g5314)
--	g5019 = AND(g312, g3933)
--	g2935 = AND(g1612, g1077)
--	g7683 = AND(g1061, g7429)
--	g5452 = AND(g4876, g3499)
--	g8654 = AND(g570, g8094)
--	g6420 = AND(g5918, g5367)
--	g4108 = AND(g782, g3655)
--	g4883 = AND(g3746, g3723, g4288)
--	I8040 = AND(g3430, g3398, g3359, g3341)
--	g4066 = AND(g1280, g3532)
--	g8272 = AND(g158, g8042)
--	g4466 = AND(I8490, I8491)
--	g8978 = AND(g8909, g5587)
--	g8612 = AND(g673, g7887)
--	g3429 = AND(g1454, g1838, g1444)
--	g6204 = AND(g5542, g5294)
--	g4365 = AND(g237, g3097)
--	g4048 = AND(g1288, g3513)
--	g8935 = AND(g3874, g8767)
--	g5425 = AND(g1528, g4916)
--	g4448 = AND(I8460, I8461)
--	g4711 = AND(g190, g4072)
--	I8528 = AND(g3430, g3398, g3359, g2106)
--	g8328 = AND(g4571, g7993)
--	g4133 = AND(g2631, g2623)
--	g4333 = AND(g1087, g2782)
--	g8542 = AND(g661, g7887)
--	g8330 = AND(g261, g7838)
--	g4396 = AND(g459, g3192)
--	g9160 = AND(g9139, g6092)
--	g6040 = AND(g1462, g5578)
--	g5105 = AND(g354, g4013)
--	g7616 = AND(g7367, g4517)
--	g7561 = AND(g7367, g4163)
--	g4067 = AND(g133, g3539)
--	I8618 = AND(g2074, g3287, g3264, g3238)
--	I8143 = AND(g2674, g2677, g2680)
--	g3049 = AND(g2274, g1844)
--	g8090 = AND(g843, g7658)
--	g6151 = AND(g1494, g5709)
--	g8823 = AND(g4561, g8512)
--	g5045 = AND(g293, g3961)
--	g5091 = AND(g397, g4001)
--	g4181 = AND(g1142, g3512)
--	g8456 = AND(g703, g7811)
--	g9271 = AND(g4748, g9244)
--	g4397 = AND(g483, g3192)
--	g8851 = AND(g284, g8524)
--	g4421 = AND(g333, g3131)
--	g8698 = AND(g3774, g8342)
--	g8260 = AND(g138, g8111)
--	g5767 = AND(g5344, g3079)
--	g6172 = AND(g1514, g5192)
--	g9238 = AND(g4748, g9223)
--	g8720 = AND(g3825, g8421)
--	g4101 = AND(g108, g3649)
--	g8318 = AND(g183, g8156)
--	g8652 = AND(g563, g8094)
--	g8843 = AND(g507, g8585)
--	I8593 = AND(g3430, g3398, g3359, g2106)
--	g8457 = AND(g724, g7811)
--	I10597 = AND(g3769, g3754, g3735)
--	g1753 = AND(g819, g815)
--	g8686 = AND(g3819, g8342)
--	g7709 = AND(g7367, g4529)
--	g8321 = AND(g446, g7920)
--	g6908 = AND(g6478, g5246)
--	g4168 = AND(g1106, g3500)
--	g6567 = AND(g6265, g2424)
--	g4368 = AND(g318, g3131)
--	g8938 = AND(g3878, g8771)
--	g5428 = AND(g775, g4707)
--	g8813 = AND(g255, g8524)
--	g5030 = AND(g233, g3946)
--	g4058 = AND(g3656, g2407)
--	g4743 = AND(g3518, g4286)
--	g8740 = AND(g2966, g8493)
--	g6965 = AND(g55, g6489)
--	g4411 = AND(g462, g3192)
--	g8687 = AND(g3488, g8363)
--	g6160 = AND(g1504, g5718)
--	g3226 = AND(g1102, g1919)
--	g4074 = AND(g137, g3573)
--	g5108 = AND(g539, g4017)
--	g6641 = AND(g5939, g5494)
--	g7002 = AND(g6770, g5054)
--	g6996 = AND(g3678, g6552)
--	g5066 = AND(g395, g3978)
--	g8860 = AND(g527, g8585)
--	g8341 = AND(g501, g7966)
--	g8710 = AND(g2790, g8421)
--	g9384 = AND(g9383, g6245)
--	g8645 = AND(g550, g8094)
--	I8209 = AND(g2298, g2316, g2334)
--	g7657 = AND(g7367, g4201)
--	g8691 = AND(g3805, g8342)
--	g5048 = AND(g394, g3966)
--	g9024 = AND(g8884, g5317)
--	g8879 = AND(g8782, g6108)
--	g8607 = AND(g8154, g5616)
--	g8962 = AND(g8890, g5317)
--	g6611 = AND(g3390, g6249)
--	g1739 = AND(g803, g799)
--	g8275 = AND(g4581, g7993)
--	g8311 = AND(g4540, g7905)
--	g4400 = AND(g1138, g3614)
--	g6541 = AND(g6144, g3510)
--	I8574 = AND(g3316, g2057, g2020, g3238)
--	g5018 = AND(g232, g3930)
--	g5067 = AND(g454, g3980)
--	g5093 = AND(g477, g4003)
--	g9273 = AND(g4748, g9252)
--	g7557 = AND(g7367, g4147)
--	g4383 = AND(g222, g3097)
--	g4220 = AND(g3533, g3549, g3568, g3583)
--	g8380 = AND(g681, g7887)
--	g8832 = AND(g501, g8585)
--	g7071 = AND(g6639, g1872)
--	g4779 = AND(g4176, g1760)
--	g7705 = AND(g7367, g4514)
--	g8853 = AND(g365, g8545)
--	g7242 = AND(g7081, g6899)
--	g4423 = AND(g465, g3192)
--	g3188 = AND(g2298, g2316)
--	g5700 = AND(g1638, g4969)
--	g4361 = AND(g471, g3192)
--	g8931 = AND(g3867, g8761)
--	g4127 = AND(g2628, g2618)
--	g4451 = AND(g359, g3131)
--	g4327 = AND(g2959, g1867)
--	g6574 = AND(g1045, g5984)
--	g7038 = AND(g6466, g4841)
--	g8628 = AND(g753, g8199)
--	g8300 = AND(g126, g8111)
--	g9014 = AND(g8906, g8239)
--	g7212 = AND(g1053, g7010)
--	g5817 = AND(g5395, g3091)
--	g4472 = AND(g440, g3160)
--	g3466 = AND(g936, g2557)
--	g8440 = AND(g714, g7937)
--	I8523 = AND(g3430, g3398, g3359, g3341)
--	g5585 = AND(g4741, g4841)
--	I8643 = AND(g2074, g3287, g3264, g1987)
--	I9535 = AND(g3062, g2712, g4253, g2752)
--	g6175 = AND(g4332, g5614)
--	g8323 = AND(g524, g7966)
--	g9335 = AND(g9320, g6206)
--	g5441 = AND(g4870, g3497)
--	g4434 = AND(g356, g3131)
--	I9261 = AND(g3777, g3764, g3746)
--	g4147 = AND(I8014, I8015)
--	I8551 = AND(g3430, g3398, g3359, g2106)
--	g9022 = AND(g8887, g5317)
--	g4681 = AND(g4255, g3533)
--	g8151 = AND(g849, g7658)
--	g8648 = AND(g588, g8094)
--	g7837 = AND(g6470, g7610)
--	g5458 = AND(g4686, g1616)
--	g3509 = AND(g1637, g1616)
--	I8613 = AND(g2074, g3287, g3264, g1987)
--	g8839 = AND(g4050, g8581)
--	g9037 = AND(g8965, g5345)
--	g6643 = AND(g1860, g5868)
--	g4936 = AND(g214, g3888)
--	g4117 = AND(g2626, g2616)
--	g4317 = AND(g878, g3086, g1857, g3659)
--	g8278 = AND(g4589, g7993)
--	g7192 = AND(g7026, g3526)
--	g8282 = AND(g179, g8156)
--	g5080 = AND(g396, g3991)
--	g5573 = AND(g3011, g4841)
--	g8693 = AND(g3798, g8342)
--	g8334 = AND(g264, g7838)
--	I8014 = AND(g3430, g3398, g3359, g3341)
--	g1919 = AND(g1098, g1087)
--	g6044 = AND(g1467, g5584)
--	g7031 = AND(g3390, g6717)
--	g6444 = AND(g1676, g6125)
--	g7252 = AND(g3591, g6977)
--	g8621 = AND(g734, g7937)
--	g4937 = AND(g3086, g4309)
--	g8313 = AND(g4542, g7951)
--	g4840 = AND(g4235, g1980)
--	I8436 = AND(g3430, g3398, g3359, g2106)
--	g4190 = AND(g1122, g3527)
--	g4390 = AND(g560, g2845)
--	g5126 = AND(g556, g4037)
--	g9012 = AND(g8908, g8239)
--	I8288 = AND(g3666, g3684, g3694)
--	g4356 = AND(g468, g3192)
--	g9371 = AND(g9352, g5917)
--	g6414 = AND(g673, g6025)
--	g8264 = AND(g105, g8131)
--	g4163 = AND(I8040, I8041)
--	g8933 = AND(g4511, g8765)
--	g7177 = AND(g7016, g5586)
--	g4053 = AND(g1292, g3523)
--	g5588 = AND(g3028, g4969)
--	g4453 = AND(g495, g3192)
--	I8495 = AND(g3430, g3398, g3359, g2106)
--	I8437 = AND(g3316, g3287, g3264, g1987)
--	g6182 = AND(g1519, g5199)
--	g8724 = AND(g3822, g8464)
--	g8379 = AND(g691, g7793)
--	g7199 = AND(g1467, g7003)
--	g6916 = AND(g727, g6515)
--	g6022 = AND(g5595, g2424)
--	g8878 = AND(g8777, g6106)
--	g6422 = AND(g714, g6033)
--	g8289 = AND(g348, g7870)
--	g8835 = AND(g270, g8524)
--	g8271 = AND(g130, g8111)
--	g8611 = AND(g669, g7887)
--	g5043 = AND(g213, g3958)
--	I8296 = AND(g3666, g3684, g3707)
--	g6437 = AND(g859, g6050)
--	g5443 = AND(g1549, g4935)
--	g7694 = AND(g7367, g4448)
--	g5116 = AND(g355, g4021)
--	g8238 = AND(g100, g8131)
--	g5034 = AND(g583, g3956)
--	g8332 = AND(g417, g7920)
--	g7701 = AND(g7367, g4497)
--	g8153 = AND(g852, g7658)
--	g4778 = AND(g4169, g1760)
--	g8744 = AND(g3802, g8464)
--	g7215 = AND(g6111, g6984)
--	I8412 = AND(g3430, g3398, g3359, g3341)
--	g4782 = AND(g4187, g1760)
--	g6042 = AND(g1041, g5581)
--	I8029 = AND(g2074, g2057, g3264, g1987)
--	g8901 = AND(g8804, g5631)
--	g6054 = AND(g1057, g5611)
--	g4526 = AND(g2642, g741)
--	g7008 = AND(g6615, g5083)
--	g2889 = AND(g1612, g1077)
--	g7136 = AND(g4057, g6953)
--	g5117 = AND(g435, g4024)
--	g8714 = AND(g2873, g8407)
--	g9025 = AND(g8889, g5317)
--	I8109 = AND(g2074, g3287, g3264, g3238)
--	g4702 = AND(g4243, g1690)
--	g6412 = AND(g158, g6024)
--	g7228 = AND(g6688, g7090)
--	g6990 = AND(g799, g6517)
--	g8262 = AND(g4554, g7855)
--	g6171 = AND(g5363, g4841)
--	g8736 = AND(g3771, g8464)
--	g4276 = AND(g2216, g2618)
--	g6429 = AND(g168, g6035)
--	g7033 = AND(g6716, g5190)
--	g9131 = AND(g9055, g5345)
--	g8623 = AND(g755, g8199)
--	g8076 = AND(g7690, g3521)
--	g7096 = AND(g6677, g5101)
--	g8722 = AND(g2787, g8386)
--	g7195 = AND(g6984, g4226)
--	g1844 = AND(g792, g795)
--	g5937 = AND(g5562, g2407)
--	g5079 = AND(g375, g3990)
--	g4546 = AND(g2643, g746)
--	g5479 = AND(g5141, g5037)
--	g6745 = AND(g1872, g6198)
--	g8285 = AND(g118, g8111)
--	g9226 = AND(g9220, g5403)
--	g6109 = AND(g5453, g5335)
--	g4224 = AND(g2680, g2683, I8127)
--	g8384 = AND(g636, g7793)
--	g8339 = AND(g345, g7870)
--	g4320 = AND(g3728, g3750, g3768, I8299)
--	g8838 = AND(g504, g8585)
--	I8019 = AND(g3430, g3398, g3359, g2106)
--	g8737 = AND(g2992, g8493)
--	I8052 = AND(g2162, g2149, g2137, g2106)
--	g4906 = AND(g4320, g2728)
--	g4789 = AND(g2751, g4202)
--	g6049 = AND(g1045, g5597)
--	g8077 = AND(g859, g7616)
--	g7692 = AND(g7367, g4430)
--	g8643 = AND(g547, g8094)
--	g6715 = AND(g677, g5843)
--	g6098 = AND(g5681, g1247)
--	g5032 = AND(g313, g3950)
--	g5432 = AND(g1537, g4921)
--	g4299 = AND(g3233, g3358)
--	g9015 = AND(g8905, g8239)
--	g8742 = AND(g2973, g8493)
--	g8304 = AND(g4523, g7905)
--	g8926 = AND(g4593, g8755)
--	g6162 = AND(g1134, g5724)
--	g6268 = AND(g1092, g5309)
--	g7001 = AND(g3722, g6562)
--	g8273 = AND(g185, g8156)
--	g6419 = AND(g162, g6032)
--	g7676 = AND(g7367, g4216)
--	g6052 = AND(g1049, g5604)
--	g4078 = AND(g3753, g3732, g3712, g3700)
--	g8269 = AND(g4569, g7951)
--	g4959 = AND(g376, g3898)
--	I8006 = AND(g2074, g3287, g2020, g3238)
--	g4435 = AND(g414, g3160)
--	g4517 = AND(I8593, I8594)
--	g4690 = AND(g4081, g3078)
--	g4082 = AND(g1296, g3604)
--	g8712 = AND(g2804, g8386)
--	g8543 = AND(g706, g7887)
--	g7703 = AND(g7367, g4504)
--	g8729 = AND(g2999, g8493)
--	g8961 = AND(g8885, g5317)
--	g9247 = AND(g4748, g9227)
--	g8927 = AND(g4594, g8756)
--	I8045 = AND(g3430, g3398, g3359, g2106)
--	g5894 = AND(g1118, g5552)
--	g8660 = AND(g1069, g8147)
--	g8946 = AND(g4556, g8786)
--	g7677 = AND(g7503, g5073)
--	I8491 = AND(g3316, g2057, g3264, g3238)
--	g6006 = AND(g5575, g2424)
--	g4236 = AND(g3260, g3221)
--	g8513 = AND(g718, g7937)
--	g6406 = AND(g154, g6018)
--	g5475 = AND(g3801, g5022)
--	g3190 = AND(g1658, g2424)
--	g6105 = AND(g5618, g2817)
--	g4877 = AND(g3746, g3723, g4288, g3764)
--	g8378 = AND(g677, g7887)
--	g6487 = AND(g5750, g4969)
--	g7699 = AND(g7367, g4486)
--	g8335 = AND(g342, g7870)
--	g8831 = AND(g423, g8564)
--	g8288 = AND(g270, g7838)
--	g8382 = AND(g685, g7887)
--	g5484 = AND(g1037, g5096)
--	I8015 = AND(g2074, g2057, g3264, g3238)
--	g8749 = AND(g2989, g8493)
--	g4785 = AND(g1678, g4202)
--	g6045 = AND(g1472, g5591)
--	g5583 = AND(g1775, g4969)
--	g6091 = AND(g5712, g5038)
--	g8947 = AND(g4558, g8787)
--	g6407 = AND(g5956, g5367)
--	g6578 = AND(g6218, g3913)
--	g4194 = AND(I8089, I8090)
--	g8653 = AND(g573, g8094)
--	g4394 = AND(g381, g3160)
--	g8302 = AND(g4521, g7855)
--	g7186 = AND(g6600, g7044)
--	g6582 = AND(g1122, g5894)
--	g1733 = AND(g1489, g1481)
--	g8719 = AND(g2821, g8443)
--	g4705 = AND(g190, g3986)
--	g6415 = AND(g5988, g5367)
--	g7614 = AND(g7367, g4176)
--	g5970 = AND(g5605, g2424)
--	I8028 = AND(g3430, g3398, g3359, g3341)
--	g8265 = AND(g134, g8111)
--	g4955 = AND(g215, g3891)
--	g4254 = AND(g3583, g3568, g3549)
--	g4814 = AND(g150, g4265)
--	g4150 = AND(I8019, I8020)
--	g4038 = AND(g825, g2949)
--	g9021 = AND(g8886, g5317)
--	g8296 = AND(g351, g7870)
--	g4409 = AND(g384, g3160)
--	g8725 = AND(g3008, g8493)
--	I8108 = AND(g2162, g2149, g2137, g2106)
--	g6689 = AND(g1519, g6239)
--	g7027 = AND(g3390, g6698)
--	g5547 = AND(g4814, g1819)
--	g7427 = AND(g1472, g7199)
--	g1898 = AND(g959, g955)
--	I8589 = AND(g2074, g3287, g3264, g3238)
--	g6428 = AND(g5874, g5494)
--	g6430 = AND(g5874, g5384)
--	g7003 = AND(g1462, g6689)
--	I8455 = AND(g3430, g3398, g3359, g3341)
--	g7695 = AND(g7367, g4466)
--	g8281 = AND(g168, g8042)
--	g5078 = AND(g316, g3989)
--	g6638 = AND(g174, g5755)
--	g7536 = AND(g4414, g7367)
--	g8297 = AND(g429, g7920)
--	g5082 = AND(g476, g3994)
--	g8745 = AND(g2982, g8493)
--	g4837 = AND(g2573, g2562, I9202)
--	g8338 = AND(g570, g8181)
--	g8963 = AND(g8891, g5317)
--	g4062 = AND(g809, g2986)
--	g7416 = AND(g7140, g4969)
--	g8309 = AND(g550, g8181)
--	I8418 = AND(g3316, g3287, g3264, g3238)
--	g6448 = AND(g5918, g5384)
--	g6055 = AND(g5239, g4202)
--	g7654 = AND(g7367, g4142)
--	g4192 = AND(g1126, g3531)
--	g4392 = AND(g303, g3131)
--	g6196 = AND(g4927, g5615)
--	g6396 = AND(g661, g6008)
--	g8715 = AND(g2761, g8386)
--	g7537 = AND(g7363, g7411)
--	g8833 = AND(g4583, g8562)
--	g7017 = AND(g3390, g6706)
--	g7417 = AND(g7144, g1616)
--	g8584 = AND(g8146, g7034)
--	g9080 = AND(g9011, g5598)
--	g6418 = AND(g5897, g5494)
--	g6994 = AND(g3658, g6538)
--	g7128 = AND(g6926, g3047)
--	g8268 = AND(g4568, g7905)
--	g5064 = AND(g315, g3975)
--	g8362 = AND(g504, g7966)
--	g4958 = AND(g296, g3897)
--	g4176 = AND(I8063, I8064)
--	g4376 = AND(g243, g3097)
--	g7554 = AND(g7367, g4139)
--	g5563 = AND(g3390, g5070)
--	g1913 = AND(g1528, g1532)
--	g6021 = AND(g5594, g2424)
--	g6421 = AND(g5847, g5384)
--	g8728 = AND(g3815, g8464)
--	g8730 = AND(g2863, g8407)
--	g4225 = AND(g2686, g2689, g2692, g2695)
--	g8385 = AND(g695, g7811)
--	I8041 = AND(g2074, g2057, g2020, g3238)
--	g4073 = AND(g1300, g3567)
--	g4796 = AND(g950, g4584)
--	g8070 = AND(g863, g7616)
--	g5089 = AND(g273, g3998)
--	g4473 = AND(g518, g3192)
--	g5489 = AND(g4912, g5053)
--	g4124 = AND(g2641, g2640)
--	g4469 = AND(I8495, I8496)
--	g4377 = AND(g297, g3131)
--	I8058 = AND(g2074, g2057, g2020, g1987)
--	g8331 = AND(g339, g7870)
--	g9023 = AND(g8888, g5317)
--	g4287 = AND(g3563, g2334, g3579, I8237)
--	g7698 = AND(g7367, g4483)
--	g8087 = AND(g7471, g7634)
--	g8305 = AND(g362, g7870)
--	g4199 = AND(g93, g2769)
--	g5438 = AND(g1545, g4932)
--	g4781 = AND(g4182, g1760)
--	g6041 = AND(g5189, g4969)
--	g8748 = AND(g2721, g8483)
--	g9327 = AND(g9316, g5757)
--	g4797 = AND(g3893, g1616)
--	g9146 = AND(g9135, g6101)
--	g9346 = AND(g9331, g6222)
--	g3002 = AND(g871, g1834)
--	I8573 = AND(g3430, g3398, g3359, g2106)
--	g6168 = AND(g1138, g5191)
--	g7652 = AND(g7367, g4194)
--	g6058 = AND(g5561, g3501)
--	g7193 = AND(g6911, g1616)
--	I8569 = AND(g3316, g2057, g2020, g1987)
--	g6743 = AND(g730, g5916)
--	g4819 = AND(g2573, g2562, I9166)
--	g8283 = AND(g267, g7838)
--	g9240 = AND(g9223, g5261)
--	g8059 = AND(g7682, g7032)
--	g8920 = AND(g4578, g8746)
--	g8459 = AND(g655, g7793)
--	g6411 = AND(g5918, g5494)
--	g8718 = AND(g2774, g8386)
--	g7598 = AND(g7483, g3466)
--	g3222 = AND(g1537, g1913)
--	g8261 = AND(g174, g8042)
--	g6474 = AND(g6203, g2424)
--	g7625 = AND(g7367, g4182)
--	g8793 = AND(g8637, g5622)
--	g6992 = AND(g6610, g3519)
--	g7232 = AND(g6694, g7091)
--	I8000 = AND(g3430, g3398, g3359, g3341)
--	g4314 = AND(g3694, g3684, g3666)
--	I8400 = AND(g3430, g3398, g3359, g3341)
--	g9147 = AND(g9136, g6103)
--	g5062 = AND(g235, g3973)
--	g9347 = AND(g9332, g6226)
--	g4825 = AND(g4228, g1964)
--	g8721 = AND(g2703, g8464)
--	g7552 = AND(g7319, g5749)
--	g7606 = AND(g7471, g3466)
--	g4408 = AND(g330, g3131)
--	g9013 = AND(g8907, g8239)
--	g5298 = AND(g1912, g4814)
--	g6976 = AND(g4399, g6508)
--	g8940 = AND(g4543, g8775)
--	I8588 = AND(g3430, g3398, g3359, g3341)
--	g4230 = AND(g2683, g3491, I8143)
--	g6400 = AND(g150, g6011)
--	I8127 = AND(g2699, g2674, g2677)
--	g4433 = AND(g278, g3097)
--	g7691 = AND(g7367, g4427)
--	g5031 = AND(g292, g3948)
--	g7607 = AND(g7325, g4969)
--	g8826 = AND(g420, g8564)
--	g4395 = AND(g405, g3160)
--	g8741 = AND(g3787, g8464)
--	g5005 = AND(g2728, g4320, I9330)
--	g2827 = AND(g1889, g1690)
--	g6423 = AND(g5897, g5384)
--	g5765 = AND(g1695, g5428)
--	I8240 = AND(g2298, g2316, g2334, g2354)
--	I8072 = AND(g3316, g3287, g2020, g3238)
--	g8609 = AND(g7828, g4969)
--	g8308 = AND(g510, g7966)
--	g7615 = AND(g7488, g3466)
--	g3229 = AND(g1728, g2015)
--	g8066 = AND(g7488, g7634)
--	I8034 = AND(g2074, g2057, g3264, g3238)
--	g4142 = AND(I8005, I8006)
--	g4342 = AND(g228, g3097)
--	I9222 = AND(g4041, g4044, g2584)
--	g6999 = AND(g815, g6556)
--	g4255 = AND(g3605, g3644, g3635, I8186)
--	g6633 = AND(g5526, g5987)
--	g8711 = AND(g3542, g8407)
--	g5069 = AND(g566, g3983)
--	g4097 = AND(g2624, g2614)
--	g7832 = AND(g5343, g7599)
--	g4497 = AND(I8551, I8552)
--	g8455 = AND(g652, g7793)
--	g4154 = AND(g1098, g3495)
--	g8827 = AND(g498, g8585)
--	g8333 = AND(g563, g8181)
--	g6732 = AND(g5874, g5367)
--	g8846 = AND(g510, g8585)
--	g6753 = AND(g5939, g5384)
--	g7559 = AND(g7367, g4155)
--	I8413 = AND(g3316, g3287, g3264, g1987)
--	g5287 = AND(g786, g4724)
--	g4783 = AND(g948, g4527)
--	g6043 = AND(g1069, g5582)
--	g4312 = AND(g3666, g3684, g3694, g3707)
--	g7628 = AND(g7367, g4532)
--	g6434 = AND(g855, g6048)
--	g8290 = AND(g588, g8181)
--	g4129 = AND(g2629, g2621)
--	g8256 = AND(g95, g8131)
--	g4830 = AND(g4288, g3723)
--	g8816 = AND(g336, g8545)
--	g6914 = AND(g6483, g5246)
--	I8460 = AND(g3430, g3398, g3359, g2106)
--	g6013 = AND(g5589, g2424)
--	g6413 = AND(g5939, g5367)
--	g8700 = AND(g3784, g8342)
--	g7323 = AND(g4065, g7171)
--	g8263 = AND(g4555, g7905)
--	g8950 = AND(g4582, g8791)
--	g4068 = AND(g121, g3540)
--	I8079 = AND(g3316, g3287, g2020, g1987)
--	g5314 = AND(g1509, g4729)
--	g8723 = AND(g2706, g8421)
--	g8257 = AND(g146, g8042)
--	g8817 = AND(g4545, g8482)
--	g8301 = AND(g182, g8156)
--	g7010 = AND(g1049, g6574)
--	g6060 = AND(g1065, g5623)
--	g4699 = AND(g1557, g4276)
--	g6460 = AND(g6178, g2424)
--	g4398 = AND(g567, g2845)
--	g5008 = AND(g231, g3920)
--	g7278 = AND(g6965, g1745)
--	g6995 = AND(g6435, g1616)
--	g8441 = AND(g746, g8018)
--	g7235 = AND(g6699, g7094)
--	I8432 = AND(g3316, g3287, g2020, g3238)
--	g9084 = AND(g8964, g5345)
--	I8053 = AND(g3316, g3287, g3264, g3238)
--	g7282 = AND(g5830, g6939)
--	g5065 = AND(g374, g3977)
--	g5122 = AND(g436, g4030)
--	g4319 = AND(g3728, g3694, g3750, I8296)
--	g7693 = AND(g7367, g4445)
--	I8568 = AND(g3430, g3398, g3359, g3341)
--	g4352 = AND(g387, g3160)
--	g5033 = AND(g393, g3953)
--	I8157 = AND(g2686, g2689, g2692)
--	g8458 = AND(g756, g8199)
--	g5096 = AND(g1149, g4400)
--	g4186 = AND(g1118, g3520)
--	g9276 = AND(g9244, g5649)
--	g4386 = AND(g324, g3131)
--	g6954 = AND(g5518, g6601)
--	g8074 = AND(g855, g7616)
--	g6053 = AND(g1053, g5608)
--	g4083 = AND(g125, g3610)
--	g8080 = AND(g7467, g7634)
--	g4483 = AND(I8523, I8524)
--	g3259 = AND(g1976, g1960)
--	g8713 = AND(g2777, g8421)
--	g5142 = AND(g1677, g4202)
--	g6157 = AND(g1130, g5717)
--	g5081 = AND(g455, g3993)
--	g9120 = AND(g9052, g5345)
--	g4187 = AND(I8078, I8079)
--	g9277 = AND(g9248, g5654)
--	g4387 = AND(g378, g3160)
--	g8688 = AND(g3812, g8342)
--	g8857 = AND(g446, g8564)
--	g8976 = AND(g8903, g6588)
--	g4427 = AND(I8431, I8432)
--	g4514 = AND(I8588, I8589)
--	g5783 = AND(g1897, g5287)
--	g7724 = AND(g7337, g5938)
--	g7179 = AND(g6121, g7035)
--	g4403 = AND(I8400, I8401)
--	g8326 = AND(g258, g7838)
--	g4145 = AND(g2639, g2635)
--	g4391 = AND(g249, g3097)
--	g5001 = AND(g458, g3912)
--	g7658 = AND(g7367, g4150)
--	g4107 = AND(g2625, g2615)
--	g1834 = AND(g933, g929)
--	g7271 = AND(g6436, g6922)
--	g4159 = AND(g1102, g3498)
--	g8383 = AND(g730, g7937)
--	g8924 = AND(g4588, g8752)
--	g7611 = AND(g7367, g4507)
--	g8779 = AND(g8634, g7037)
--	g6949 = AND(g5483, g6589)
--	g4315 = AND(g3707, g3728, I8288)
--	g4047 = AND(g1272, g3503)
--	g8361 = AND(g426, g7920)
--	g6998 = AND(g4474, g6555)
--	g7238 = AND(g6707, g7098)
--	g5624 = AND(g5140, g2794)
--	g7680 = AND(g7367, g4166)
--	g8327 = AND(g336, g7870)
--	g6039 = AND(g1037, g5574)
--	g5068 = AND(g475, g3982)
--	g6439 = AND(g789, g6150)
--	I8546 = AND(g3430, g3398, g3359, g3341)
--	g8303 = AND(g284, g7838)
--	g8696 = AND(g3743, g8342)
--	g8732 = AND(g3808, g8464)
--	g4272 = AND(g3233, g3286)
--	g8944 = AND(g4539, g8783)
--	g5699 = AND(g1667, g4841)
--	g4417 = AND(I8417, I8418)
--	I8617 = AND(g3430, g3398, g3359, g2106)
--	g7600 = AND(g7460, g3466)
--	g4128 = AND(g98, g3693)
--	g3081 = AND(g1682, g1616)
--	g8316 = AND(g513, g7966)
--	I8299 = AND(g3666, g3684, g3694, g3707)
--	I8547 = AND(g3316, g2057, g2020, g3238)
--	g6970 = AND(g5035, g6490)
--	g8147 = AND(g1065, g7683)
--	g5119 = AND(g543, g4027)
--	g8697 = AND(g3761, g8342)
--	g8914 = AND(g8795, g8239)
--	g4902 = AND(g4304, g2770, g2746, g2728)
--	I8078 = AND(g2162, g2149, g2137, g2106)
--	g7175 = AND(g6893, g4841)
--	g5599 = AND(g4745, g4969)
--	g4490 = AND(g521, g3192)
--	g4823 = AND(g4238, g4230, g174)
--	g4166 = AND(I8045, I8046)
--	g8820 = AND(g261, g8524)
--	g4366 = AND(g216, g3097)
--	g8936 = AND(g3875, g8768)
--	g6771 = AND(g146, g6004)
--	g8317 = AND(g547, g8181)
--	g4529 = AND(I8612, I8613)
--	g5125 = AND(g517, g4036)
--	g7184 = AND(g6138, g7043)
--	g4155 = AND(I8028, I8029)
--	g5984 = AND(g1041, g5484)
--	g4355 = AND(g390, g3160)
--	g8922 = AND(g4586, g8750)
--	g6738 = AND(g5847, g5367)
--	g8060 = AND(g7535, g4841)
--	g5106 = AND(g398, g4015)
--	g6991 = AND(g5689, g6520)
--	g8460 = AND(g757, g8199)
--	g9038 = AND(g8966, g5345)
--	g8739 = AND(g3780, g8464)
--	g4720 = AND(g190, g4055)
--	g4118 = AND(g995, g3790)
--	g4167 = AND(g2783, g1616)
--	g4367 = AND(g240, g3097)
--	g4872 = AND(g1924, g4225, g4224)
--	g7634 = AND(g7367, g4549)
--	g8937 = AND(g4524, g8770)
--	g8079 = AND(g831, g7658)
--	g8294 = AND(g281, g7838)
--	g5046 = AND(g314, g3962)
--	g8840 = AND(g4590, g8582)
--	g4193 = AND(g145, g2727)
--	g4393 = AND(g327, g3131)
--	g4549 = AND(I8642, I8643)
--	g6915 = AND(g6493, g5246)
--	I8064 = AND(g3316, g3287, g3264, g1987)
--	g8942 = AND(g4522, g8780)
--	g2912 = AND(g1080, g1945)
--	g5107 = AND(g478, g4016)
--	g8704 = AND(g2829, g8386)
--	g6002 = AND(g5539, g2407)
--	g6402 = AND(g665, g6012)
--	g8954 = AND(g8763, g6097)
--	I8237 = AND(g2298, g2316, g2354)
--	g6762 = AND(g5847, g5412)
--	g4740 = AND(g2242, g4275)
--	g3258 = AND(g2298, g2316, g2334, g2354)
--	g5047 = AND(g373, g3964)
--	I8089 = AND(g2162, g2149, g2137, g2106)
--	g8912 = AND(g8796, g8239)
--	I8071 = AND(g2162, g2149, g2137, g2106)
--	g6464 = AND(g6177, g2424)
--	g8929 = AND(g3865, g8759)
--	g3614 = AND(g1134, g2386)
--	g7036 = AND(g6728, g5197)
--	g7679 = AND(g7447, g5084)
--	g8626 = AND(g752, g8199)
--	g3984 = AND(g2403, g3085)
--	g5017 = AND(g211, g3928)
--	g4691 = AND(g4219, g1690)
--	g2949 = AND(g822, g1753)
--	g7182 = AND(g6902, g4969)
--	g6394 = AND(g5988, g5494)
--	g4962 = AND(g457, g3905)
--	g4158 = AND(I8033, I8034)
--	g6966 = AND(g6580, g5580)
--	g8735 = AND(g2807, g8443)
--	g8075 = AND(g7460, g7634)
--	g8949 = AND(g4572, g8790)
--	g7632 = AND(g7445, g3548)
--	g7653 = AND(g7480, g5754)
--	g8292 = AND(g181, g8156)
--	g2952 = AND(g2474, g2215)
--	g6438 = AND(g4829, g6051)
--	g4284 = AND(g3260, g3314)
--	g4239 = AND(g1541, g3222)
--	g5090 = AND(g317, g4000)
--	g8646 = AND(g553, g8094)
--	g6409 = AND(g706, g6020)
--	g4180 = AND(g1114, g3511)
--	g9270 = AND(g4748, g9241)
--	g4380 = AND(g584, g2845)
--	g4832 = AND(g1110, g4246)
--	g8439 = AND(g699, g7811)
--	g2986 = AND(g806, g1739)
--	g4420 = AND(g275, g3097)
--	g4507 = AND(I8573, I8574)
--	g4794 = AND(g954, g4574)
--	g8702 = AND(g2837, g8386)
--	g8919 = AND(g4567, g8743)
--	g8952 = AND(g8788, g6075)
--	g8276 = AND(g150, g8042)
--	g5063 = AND(g294, g3974)
--	g4100 = AND(g113, g3648)
--	g7553 = AND(g7367, g4135)
--	g8404 = AND(g710, g7937)
--	g5118 = AND(g479, g4026)
--	g8764 = AND(g8231, g4969)
--	
--	g5057 = OR(g3939, g3925, g3915, g3907)
--	I14941 = OR(g8275, g8323, g8459, g8380)
--	g5193 = OR(g5017, g4366)
--	g9291 = OR(g9273, g6216)
--	g5549 = OR(g2935, g4712)
--	g7029 = OR(g6433, g5765)
--	g7787 = OR(g4791, g7602)
--	g6249 = OR(g4066, g5313)
--	g8906 = OR(g8088, g8062, g8699)
--	g5232 = OR(g5082, g4412)
--	g8987 = OR(g8927, g8826)
--	g5253 = OR(g5116, g4451)
--	g7791 = OR(g4796, g7606)
--	I8225 = OR(g3062, g2712, g2734, g2752)
--	I15250 = OR(g8238, g8265, g8272, g8292)
--	g8991 = OR(g8931, g8831)
--	I9107 = OR(g4133, g4145, g4138, g4132)
--	g9008 = OR(g8948, g8857)
--	g2214 = OR(g1376, g1377, g1378, g1379)
--	g7575 = OR(g7323, g7142)
--	g9136 = OR(g8952, g9131)
--	g8907 = OR(g8081, g8064, g8707)
--	g8082 = OR(g7654, g7628, g7611)
--	g5710 = OR(g4958, g4351)
--	I9047 = OR(g4155, g4147, g4139)
--	g9122 = OR(g8953, g9084)
--	g6270 = OR(g1000, g5335, g1909)
--	g6610 = OR(g4180, g6061)
--	g6124 = OR(g5432, g4789)
--	g6980 = OR(g6745, g6028)
--	I14484 = OR(g7993, g7966, g7793, g7811)
--	g9137 = OR(g8877, g9118)
--	g9337 = OR(g9240, g9327)
--	g7086 = OR(g4101, g6464)
--	I15055 = OR(I15051, I15052, I15053, I15054)
--	I15111 = OR(g7951, g7920, g7983, g8181)
--	g5545 = OR(g3617, g4824)
--	g7025 = OR(g6541, g3095)
--	g4264 = OR(g2490, g3315)
--	g8899 = OR(g8839, g8652)
--	g8785 = OR(g8623, g8656, I14985)
--	I15019 = OR(g7951, g7920, g7983, g8181)
--	g6144 = OR(g4175, g5458)
--	g9154 = OR(g9142, g9021)
--	g9354 = OR(g9275, g9344)
--	I15018 = OR(g7855, g7838, g7905, g7870)
--	g4179 = OR(g207, g3083)
--	g7682 = OR(g6044, g7412)
--	g6694 = OR(g6151, g5573)
--	g5204 = OR(g5033, g4379)
--	g9267 = OR(g9251, g6225)
--	g9001 = OR(g8941, g8846)
--	g8966 = OR(g8741, g8745, g8912, g8850)
--	g7445 = OR(g4192, g7193)
--	g5040 = OR(g3900, g3895, g3890, g4363)
--	g5440 = OR(g4790, g4786)
--	I15102 = OR(I15098, I15099, I15100, I15101)
--	g2229 = OR(g1371, g1372, g1373, g1374)
--	I14771 = OR(g7993, g7966, g7793, g7811)
--	I15231 = OR(g8701, g8715, g8730, g8720)
--	g8773 = OR(I14959, I14960)
--	g8009 = OR(g3591, g7406, g7566, I14302)
--	g8769 = OR(I14951, I14952)
--	g7227 = OR(g6992, g3128)
--	g6934 = OR(g6422, g6430)
--	g8993 = OR(g8933, g8835)
--	g6913 = OR(g6733, g6738)
--	g5235 = OR(g5091, g4422)
--	g5343 = OR(g4690, g2862)
--	I15085 = OR(g8363, g8342, g8407, g8386)
--	g5566 = OR(g3617, g4810)
--	I14759 = OR(g7937, g7887, g8029, g8018)
--	I15054 = OR(g8363, g8342, g8407, g8386)
--	I15243 = OR(I15239, I15240, I15241, I15242)
--	I14758 = OR(g7993, g7966, g7793, g7811)
--	g4736 = OR(g4532, g4517, I9044)
--	g8895 = OR(g8823, g8646)
--	g7428 = OR(g6040, g7175)
--	g9352 = OR(g9343, g4526)
--	g7826 = OR(g4804, g7626)
--	g8788 = OR(g8620, g8658, I14990)
--	g5202 = OR(g5031, g4377)
--	g5518 = OR(g4744, g4118)
--	g4737 = OR(g4135, g4529, g4514, I9047)
--	g7165 = OR(g6434, g6908)
--	g5264 = OR(g5125, g4490)
--	g8176 = OR(g7566, g1030, g6664, g6452)
--	g9387 = OR(g9349, g9384)
--	g2206 = OR(g1363, g1364, g1365, g1366)
--	I14951 = OR(g8328, g8316, g8455, g8378)
--	g9046 = OR(g8744, g8749, g9016, g8862)
--	g6932 = OR(g6417, g6423)
--	I15169 = OR(g8483, g8464, g8514)
--	g9003 = OR(g8943, g8849)
--	g8796 = OR(g8150, g8078, g8070, g8360)
--	g8980 = OR(g8920, g8815)
--	g6716 = OR(g6162, g5588)
--	g7421 = OR(g6745, g7202)
--	g6699 = OR(g6154, g5579)
--	g5238 = OR(g5094, g4425)
--	g4927 = OR(g4318, g1590)
--	g5209 = OR(g5044, g4384)
--	I15084 = OR(g7951, g7920, g7983, g8181)
--	I15110 = OR(g7855, g7838, g7905, g7870)
--	g8900 = OR(g8840, g8653)
--	g5511 = OR(g4743, g4109)
--	g6717 = OR(g4082, g6005)
--	g3160 = OR(g1751, g449)
--	g8886 = OR(g8727, g8812, I15254)
--	g2230 = OR(g1380, g1381, g1382, g1383)
--	I15242 = OR(g8697, g8714, g8718, g8719)
--	g5722 = OR(g5001, g4361)
--	g2845 = OR(g1877, g576)
--	I15230 = OR(g8274, g8321, g8298, g8696)
--	I15265 = OR(I15261, I15262, I15263, I15264)
--	g4786 = OR(g4107, g4097, g4124, I9099)
--	I13553 = OR(g1166, g1167, g1170)
--	g8887 = OR(I15265, g8819)
--	g7080 = OR(g4086, g6462)
--	g4364 = OR(g2952, g1725)
--	g9148 = OR(g9143, g9024)
--	I14767 = OR(g7937, g7887, g8029, g8018)
--	g9355 = OR(g9276, g9345)
--	g3541 = OR(g1663, g1421)
--	I14990 = OR(g8337, g8379, g8543)
--	g5231 = OR(g5081, g4411)
--	g5205 = OR(g5034, g4380)
--	g8891 = OR(g8705, g8811, I15297, I15298)
--	I15041 = OR(g7855, g7838, g7905, g7870)
--	g6115 = OR(g3617, g5558)
--	I15275 = OR(g8693, g8703, g8712, g8717)
--	g4297 = OR(g3617, g3602)
--	g7220 = OR(g1304, g7062)
--	g5572 = OR(g5051, g1236)
--	g8154 = OR(g6054, g7607)
--	I14766 = OR(g7993, g7966, g7793, g7811)
--	g6935 = OR(g6429, g6431)
--	I15165 = OR(g8483, g8464, g8514)
--	g8979 = OR(g8919, g8813)
--	g5036 = OR(g4047, g2972)
--	g3339 = OR(g1424, g2014)
--	I15253 = OR(g8698, g8711, g8722, g8716)
--	g7443 = OR(g7192, g3158)
--	I14754 = OR(g7937, g7887, g8029, g8018)
--	I15175 = OR(g8483, g8464, g8514)
--	I15264 = OR(g8700, g8708, g8726, g8731)
--	g9358 = OR(g9279, g9348)
--	g7697 = OR(g7419, g3187)
--	g6698 = OR(g4073, g6001)
--	g6964 = OR(g6447, g6448)
--	g5208 = OR(g5043, g4383)
--	g9174 = OR(g9147, g8963)
--	I15021 = OR(I15017, I15018, I15019, I15020)
--	g9239 = OR(g7653, g9226)
--	g5265 = OR(g5126, g4491)
--	I15073 = OR(g7951, g7920, g7983, g8181)
--	I15274 = OR(g8306, g8361, g8299, g8687)
--	g6457 = OR(g6196, g6209, g4937)
--	g5233 = OR(g5089, g4420)
--	g6686 = OR(g4068, g5970)
--	I15292 = OR(g8704, g8710, g8805)
--	g8893 = OR(g8814, g8643)
--	g7784 = OR(g7406, g6664, g3492, I14219)
--	g6121 = OR(g5425, g4785)
--	I14366 = OR(g7566, g1030, g6664)
--	g5706 = OR(g4955, g4342)
--	g6740 = OR(g4100, g6022)
--	g4283 = OR(g3587, g2665)
--	g8984 = OR(g8924, g8822)
--	I15109 = OR(g8131, g8111, g8042, g8156)
--	g9123 = OR(g8954, g9037)
--	I15283 = OR(g8291, g8276, g8325, g8330)
--	g5138 = OR(g4108, g3049)
--	g7810 = OR(g4799, g7609)
--	g7363 = OR(g7136, g6903)
--	I9099 = OR(g4127, g4123, g4117)
--	g9151 = OR(g9144, g8961)
--	g6525 = OR(g6112, g5547)
--	g6710 = OR(g55, g6264)
--	I6209 = OR(g911, g916, g921, g883)
--	g8904 = OR(g8090, g8080, g8706)
--	g5707 = OR(g4956, g4343)
--	I14980 = OR(g8362, g8403, g8610)
--	g9010 = OR(g8950, g8860)
--	g5201 = OR(g5030, g4376)
--	g8763 = OR(g8232, I14941, I14942)
--	I9044 = OR(g4150, g4142, g4549)
--	g8637 = OR(g6057, g8071)
--	g5715 = OR(g4961, g4355)
--	g9282 = OR(g9270, g6238)
--	I15040 = OR(g8131, g8111, g8042, g8156)
--	g5052 = OR(g4049, g4054)
--	I15252 = OR(g8320, g8307, g8317, g8692)
--	g7782 = OR(g4783, g7598)
--	g6931 = OR(g6416, g6421)
--	I14969 = OR(g8315, g8377, g8359, g8611)
--	g5070 = OR(g4052, g4058)
--	g2213 = OR(g1367, g1368, g1369, g1370)
--	g8982 = OR(g8922, g8820)
--	g4055 = OR(g187, g3012)
--	g8128 = OR(g7566, g6910, g6452)
--	I11603 = OR(g6193, g6197, g6175)
--	g9264 = OR(g9247, g6242)
--	g6440 = OR(g6268, g5700)
--	g6123 = OR(g3617, g5556)
--	I15051 = OR(g8131, g8111, g8042, g8156)
--	I15072 = OR(g7855, g7838, g7905, g7870)
--	I14496 = OR(g7937, g7887, g8029, g8018)
--	g8902 = OR(g8844, g8654)
--	I15152 = OR(g8483, g8464, g8514)
--	g8155 = OR(g7632, g3219)
--	g8964 = OR(g8915, g8863, I15400)
--	g5227 = OR(g5077, g4407)
--	I15020 = OR(g8363, g8342, g8407, g8386)
--	g5203 = OR(g5032, g4378)
--	I9029 = OR(g4504, g4494, g4430)
--	g8989 = OR(g8929, g8829)
--	I15113 = OR(I15109, I15110, I15111, I15112)
--	g8834 = OR(g7096, g8229)
--	g5188 = OR(g5008, g4365)
--	g7435 = OR(g6052, g7182)
--	g7690 = OR(g4181, g7417)
--	g5216 = OR(g5062, g4391)
--	g3131 = OR(g1749, g368)
--	g8909 = OR(g6043, g8764)
--	g4734 = OR(g4469, g4448, I9038)
--	g6933 = OR(g6419, g6428)
--	I14480 = OR(g7937, g7887, g8029, g8018)
--	g9285 = OR(g9271, g6221)
--	I6208 = OR(g891, g896, g901, g906)
--	g5217 = OR(g5063, g4392)
--	g9139 = OR(g8879, g9120)
--	g9339 = OR(g9259, g9335)
--	g5711 = OR(g4959, g4352)
--	g7222 = OR(g6049, g6971)
--	I14942 = OR(g8439, g8440, g8405, g8460)
--	g4688 = OR(g4193, g3190)
--	g5196 = OR(g5020, g4369)
--	g6132 = OR(g5436, g4793)
--	g8985 = OR(g8925, g8824)
--	g7089 = OR(g4128, g6474)
--	g5256 = OR(g5119, g4454)
--	I14468 = OR(g7937, g7887, g8029, g8018)
--	g8794 = OR(g8153, g8074, g8069, g8523)
--	g5021 = OR(g943, g4501)
--	g7254 = OR(g6923, g5298)
--	g6600 = OR(g5443, g6055)
--	g8905 = OR(g8089, g8087, g8694)
--	g7438 = OR(g7184, g6978)
--	g6580 = OR(g6039, g6041)
--	g6262 = OR(g4074, g5334)
--	I15229 = OR(g8262, g8303, g8268, g8312)
--	I14479 = OR(g7993, g7966, g7793, g7811)
--	I15228 = OR(g8270, g8258, g8281, g8273)
--	g4072 = OR(g196, g2995)
--	g9135 = OR(g8951, g9130)
--	g9288 = OR(g9272, g6235)
--	I15112 = OR(g8363, g8342, g8407, g8386)
--	g5673 = OR(g4823, g4872)
--	g7062 = OR(g4048, g6456)
--	g4413 = OR(g2371, g3285)
--	g8884 = OR(g8735, g8818, I15232)
--	g7788 = OR(g4794, g7604)
--	g8988 = OR(g8928, g8827)
--	g6926 = OR(g6406, g6411)
--	g8804 = OR(g6060, g8609)
--	g9054 = OR(g8724, g8729, g9013, g8680)
--	I15298 = OR(g8332, g8333, g8686, g8702)
--	g6543 = OR(g6125, g1553)
--	g8908 = OR(g8079, g8066, g8855)
--	I14772 = OR(g7937, g7887, g8029, g8018)
--	I15232 = OR(I15228, I15229, I15230, I15231)
--	I15261 = OR(g8256, g8271, g8267, g8286)
--	g6927 = OR(g6408, g6413)
--	g9171 = OR(g9146, g8962)
--	g8965 = OR(g8739, g8742, g8914, g8847)
--	g5220 = OR(g5066, g4395)
--	g6436 = OR(g6266, g5699)
--	g8996 = OR(g8936, g8838)
--	g9138 = OR(g8878, g9119)
--	g9338 = OR(g9258, g9334)
--	g8777 = OR(I14969, I14970)
--	g9049 = OR(g8732, g8737, g9015, g8861)
--	I15031 = OR(g7951, g7920, g7983, g8181)
--	g8981 = OR(g8921, g8816)
--	g1690 = OR(g1021, g1025, g1018)
--	g8997 = OR(g8937, g8841)
--	g6579 = OR(g6098, g1975)
--	g7088 = OR(g6638, g6641)
--	g6719 = OR(g6166, g6171)
--	g6917 = OR(g6743, g6753)
--	g9162 = OR(g9158, g9022)
--	g4735 = OR(g4427, g4414, g4403, I9041)
--	g9052 = OR(g8728, g8733, g9014, g8679)
--	g5210 = OR(g5045, g4385)
--	g2262 = OR(g1384, g1385, g1386, g1387)
--	I15043 = OR(g8363, g8342, g8407, g8386)
--	g7825 = OR(g4801, g7615)
--	g3760 = OR(I7232, I7233)
--	I9041 = OR(g4483, g4466, g4445)
--	g5317 = OR(g4727, g4737, g4735)
--	I14952 = OR(g8456, g8513, g8458, g8236)
--	g6706 = OR(g4077, g6002)
--	g7230 = OR(g4190, g6995)
--	g9006 = OR(g8946, g8853)
--	g8889 = OR(I15283, I15284, I15285)
--	I14834 = OR(g8483, g8464, g8514)
--	g7337 = OR(g7278, g4546)
--	g6138 = OR(g5438, g5442)
--	I15086 = OR(I15082, I15083, I15084, I15085)
--	g6707 = OR(g6160, g5585)
--	g8795 = OR(g8151, g8077, g8075, g8279)
--	g7248 = OR(g7079, g5652)
--	g1955 = OR(g1189, g16)
--	g5704 = OR(g4936, g4334)
--	g9007 = OR(g8947, g8854)
--	g7081 = OR(g6172, g6629)
--	g9261 = OR(g9238, g6227)
--	g8634 = OR(g6047, g8060)
--	I15017 = OR(g8131, g8111, g8042, g8156)
--	g7783 = OR(g4787, g7600)
--	g8613 = OR(g8082, g7616)
--	g8983 = OR(g8923, g8821)
--	g4876 = OR(g4159, g4167)
--	g6728 = OR(g6168, g5593)
--	g6470 = OR(g5817, g2934)
--	g8885 = OR(g8723, g8806, I15243)
--	I7232 = OR(g2367, g2352, g2378, g2330)
--	g9165 = OR(g9159, g9023)
--	I15042 = OR(g7951, g7920, g7983, g8181)
--	g9055 = OR(g8721, g8725, g9012, g8859)
--	g6445 = OR(g6105, g6107)
--	g7258 = OR(g7083, g5403, I13220)
--	g6602 = OR(g6058, g3092)
--	g4295 = OR(g2828, g2668)
--	I15030 = OR(g7855, g7838, g7905, g7870)
--	g6920 = OR(g6395, g6399)
--	g5561 = OR(g4168, g4797)
--	g6459 = OR(g6259, g6185, I11603)
--	g6718 = OR(g4083, g6006)
--	g7026 = OR(g4186, g6554)
--	I14933 = OR(g8385, g8404, g8441, g8462)
--	g7426 = OR(g1173, g7217, I13553)
--	g7170 = OR(g6916, g6444)
--	g7083 = OR(g5448, g6267, g6710)
--	I15075 = OR(I15071, I15072, I15073, I15074)
--	g8990 = OR(g8930, g8830)
--	g8888 = OR(I15276, g8807)
--	g7191 = OR(g7071, g6980)
--	g5244 = OR(g5107, g4436)
--	g5140 = OR(g4333, g3509)
--	g7016 = OR(g6042, g6487)
--	g9168 = OR(g9160, g9025)
--	I15276 = OR(I15272, I15273, I15274, I15275)
--	I15285 = OR(g8709, g8713, g8803)
--	g5214 = OR(g5049, g4389)
--	I15053 = OR(g7951, g7920, g7983, g8181)
--	I15254 = OR(I15250, I15251, I15252, I15253)
--	g4249 = OR(g3617, g1639)
--	g3986 = OR(g202, g3129)
--	I14302 = OR(g6664, g3492, g979)
--	g9011 = OR(g6046, g8892)
--	I15101 = OR(g8363, g8342, g8407, g8386)
--	g5236 = OR(g5092, g4423)
--	g7272 = OR(g6182, g7038)
--	g8896 = OR(g8828, g8648)
--	g5222 = OR(g5068, g4397)
--	g4812 = OR(g2490, g4237)
--	g4829 = OR(g863, g4051)
--	g6685 = OR(g4067, g5969)
--	g5237 = OR(g5093, g4424)
--	I15074 = OR(g8363, g8342, g8407, g8386)
--	I15239 = OR(g8264, g8260, g8277, g8301)
--	g5194 = OR(g5018, g4367)
--	g9000 = OR(g8940, g8845)
--	g8897 = OR(g8833, g8650)
--	g7166 = OR(g6437, g6914)
--	g5242 = OR(g5105, g4434)
--	g5254 = OR(g5117, g4452)
--	I14932 = OR(g8278, g8329, g8461, g8382)
--	g6585 = OR(g3617, g6119)
--	g6673 = OR(g4053, g5937)
--	g5212 = OR(g5047, g4387)
--	g7167 = OR(g6438, g6915)
--	g8091 = OR(g7215, g6452, I14366)
--	I15083 = OR(g7855, g7838, g7905, g7870)
--	g5229 = OR(g5079, g4409)
--	I15284 = OR(g8335, g8340, g8290, g8691)
--	g6458 = OR(g6184, g6259, g6174, g6214)
--	g7834 = OR(g7724, g6762)
--	g6734 = OR(g6176, g5599)
--	g4870 = OR(g4154, g3081)
--	g7687 = OR(g6053, g7416)
--	g6688 = OR(g6145, g5570)
--	I15052 = OR(g7855, g7838, g7905, g7870)
--	I14959 = OR(g8322, g8308, g8438, g8612)
--	g5708 = OR(g2889, g4699)
--	g5219 = OR(g5065, g4394)
--	g6924 = OR(g6400, g6405)
--	I15400 = OR(g8736, g8748, g8740)
--	g9294 = OR(g9274, g6230)
--	g8758 = OR(g8655, I14932, I14933)
--	g9356 = OR(g9277, g9346)
--	g7020 = OR(g3617, g6578)
--	I15241 = OR(g8269, g8314, g8309, g8695)
--	I15100 = OR(g7951, g7920, g7983, g8181)
--	g9363 = OR(g9359, g6210)
--	g6116 = OR(g5546, g4681)
--	g6565 = OR(g2396, g6131, g1603)
--	g8994 = OR(g8934, g8836)
--	g5245 = OR(g5108, g4437)
--	g9357 = OR(g9278, g9347)
--	g3192 = OR(g1756, g530)
--	g4727 = OR(g4417, g4172, g4163, I9029)
--	g7040 = OR(g6439, g5783)
--	g5259 = OR(g5122, g4472)
--	I14831 = OR(g8483, g8464, g8514)
--	I9038 = OR(g4507, g4497, g4486)
--	I15082 = OR(g8131, g8111, g8042, g8156)
--	g5215 = OR(g5050, g4390)
--	I14753 = OR(g7993, g7966, g7793, g7811)
--	g2368 = OR(I6208, I6209)
--	g4747 = OR(g3984, g2912)
--	I13220 = OR(g58, g6258, g5418)
--	I15263 = OR(g8313, g8297, g8310, g8690)
--	g6739 = OR(g4099, g6021)
--	I5757 = OR(g969, g970, g966, g963)
--	I8363 = OR(g2655, g1163, g1160)
--	I14960 = OR(g8621, g8622, g8628, g8230)
--	g5228 = OR(g5078, g4408)
--	g5230 = OR(g5080, g4410)
--	g8890 = OR(I15290, I15291, I15292)
--	I15273 = OR(g8287, g8334, g8295, g8339)
--	g5195 = OR(g5019, g4368)
--	g9004 = OR(g8944, g8851)
--	g7202 = OR(g6028, g7071)
--	I15033 = OR(I15029, I15030, I15031, I15032)
--	g8992 = OR(g8932, g8832)
--	I14970 = OR(g8457, g8383, g8626, g8233)
--	g4280 = OR(I8224, I8225)
--	g6912 = OR(g4199, g6567)
--	g5255 = OR(g5118, g4453)
--	g4790 = OR(g4185, g4131, g4129, I9107)
--	g6929 = OR(g6412, g6418)
--	g7450 = OR(g6090, g7195)
--	g1872 = OR(g971, g962, g972, I5757)
--	g5218 = OR(g5064, g4393)
--	g6735 = OR(g4091, g6013)
--	g5830 = OR(g5714, g5142)
--	I15291 = OR(g8331, g8336, g8338, g8688)
--	I7233 = OR(g2315, g2385, g2294, g2395)
--	g5221 = OR(g5067, g4396)
--	I15029 = OR(g8131, g8111, g8042, g8156)
--	g2043 = OR(g1263, g1257)
--	g8999 = OR(g8939, g8843)
--	g8146 = OR(g6045, g7597)
--	I8224 = OR(g3019, g3029, g3038, g3052)
--	g5716 = OR(g4962, g4356)
--	g6919 = OR(g6771, g6394)
--	g9002 = OR(g8942, g8848)
--	g6952 = OR(g6633, g6204)
--	I15240 = OR(g8259, g8294, g8263, g8305)
--	I14495 = OR(g7993, g7966, g7793, g7811)
--	g5241 = OR(g5104, g4433)
--	I14985 = OR(g8341, g8384, g8542)
--	g3097 = OR(g1746, g287)
--	I15262 = OR(g8293, g8283, g8304, g8289)
--	g6925 = OR(g6402, g6407)
--	g6120 = OR(g3617, g5555)
--	g5211 = OR(g5046, g4386)
--	g6906 = OR(g6715, g6726)
--	I15099 = OR(g7855, g7838, g7905, g7870)
--	I15098 = OR(g8131, g8111, g8042, g8156)
--	I15251 = OR(g8302, g8288, g8311, g8296)
--	I15272 = OR(g8237, g8300, g8261, g8282)
--	g5483 = OR(g4740, g4098)
--	I15032 = OR(g8363, g8342, g8407, g8386)
--	g6907 = OR(g6727, g6732)
--	g9009 = OR(g8949, g8858)
--	g8995 = OR(g8935, g8837)
--	I14219 = OR(g979, g7566, g1865)
--	g5200 = OR(g5029, g4375)
--	g5345 = OR(g4736, g4734)
--	g5223 = OR(g5069, g4398)
--	I15071 = OR(g8131, g8111, g8042, g8156)
--	I14467 = OR(g7993, g7966, g7793, g7811)
--	I15147 = OR(g8483, g8464, g8514)
--	g6590 = OR(g3617, g6153)
--	I15172 = OR(g8483, g8464, g8514)
--	g6928 = OR(g6409, g6415)
--	g6930 = OR(g6414, g6420)
--	g5537 = OR(g3617, g4835)
--	g7436 = OR(g7183, g6975)
--	g5243 = OR(g5106, g4435)
--	g5234 = OR(g5090, g4421)
--	I15044 = OR(I15040, I15041, I15042, I15043)
--	g6705 = OR(g6157, g5583)
--	g8894 = OR(g8817, g8645)
--	g8782 = OR(g8624, g8659, I14980)
--	g9005 = OR(g8945, g8852)
--	g5213 = OR(g5048, g4388)
--	I15290 = OR(g8285, g8266, g8318, g8326)
--	g4374 = OR(g1182, g1186, g1179, I8363)
--	g8998 = OR(g8938, g8842)
--	g9124 = OR(g8876, g9038)
--	g5698 = OR(g5057, g5040)
--	I14485 = OR(g7937, g7887, g8029, g8018)
--	g5260 = OR(g5123, g4473)
--	g9377 = OR(g9371, g6757)
--	g6921 = OR(g6396, g6401)
--	g8986 = OR(g8926, g8825)
--	I15297 = OR(g8280, g8257, g8319, g8327)
--	
--	I15888 = NAND(g9192, I15887)
--	I7466 = NAND(g2982, g1704)
--	I10092 = NAND(g4881, g2177)
--	g5686 = NAND(g5132, g1263)
--	I5521 = NAND(g1098, I5519)
--	g4528 = NAND(I8606, I8607)
--	g5625 = NAND(g2044, g4957)
--	I7538 = NAND(g2996, g1715)
--	I11143 = NAND(g5493, I11142)
--	I7467 = NAND(g2982, I7466)
--	g4839 = NAND(g1879, g4269)
--	I10906 = NAND(g5492, g2605)
--	I12575 = NAND(g6574, g1049)
--	I7181 = NAND(g795, I7179)
--	g4235 = NAND(g1415, g2668)
--	g6286 = NAND(I11178, I11179)
--	I7421 = NAND(g2525, g2703)
--	g5141 = NAND(I9548, I9549)
--	g6911 = NAND(I12597, I12598)
--	g4548 = NAND(I8636, I8637)
--	I15855 = NAND(g9168, g9165)
--	I11110 = NAND(g2734, I11108)
--	I11179 = NAND(g3019, I11177)
--	g6473 = NAND(g5269, g5988)
--	I6524 = NAND(g1102, I6522)
--	I11178 = NAND(g5466, I11177)
--	I8510 = NAND(g2517, g2807)
--	I8245 = NAND(g3506, I8243)
--	g4313 = NAND(g3712, g3700)
--	I11186 = NAND(g3029, I11184)
--	g6469 = NAND(g5918, g5278)
--	I13685 = NAND(g1977, g7237)
--	I6258 = NAND(g837, I6257)
--	g6177 = NAND(I10889, I10890)
--	I13800 = NAND(g7429, g1061)
--	I15819 = NAND(g9148, I15817)
--	I15818 = NAND(g9151, I15817)
--	I5600 = NAND(g1489, I5598)
--	g6287 = NAND(I11185, I11186)
--	I9978 = NAND(g4880, g2092)
--	I9243 = NAND(g4305, I9241)
--	I6274 = NAND(g840, I6273)
--	g5284 = NAND(g4344, g4335, g4963)
--	I10745 = NAND(g2100, I10743)
--	g5239 = NAND(I9746, I9747)
--	I9234 = NAND(g4310, I9233)
--	I6170 = NAND(g843, g911)
--	I13587 = NAND(g2556, g7234)
--	g6510 = NAND(g5278, g5874)
--	I6939 = NAND(g2161, g2051)
--	I11117 = NAND(g3062, I11115)
--	g5559 = NAND(g5132, g1257)
--	g3232 = NAND(g2298, g2276)
--	I7531 = NAND(g2487, g3787)
--	g3938 = NAND(I7610, I7611)
--	I7505 = NAND(g3802, I7503)
--	I7011 = NAND(g2333, I7009)
--	I11123 = NAND(g5517, I11122)
--	I11751 = NAND(g6112, I11750)
--	g6701 = NAND(I12032, I12033)
--	g4835 = NAND(I9195, I9196)
--	I13639 = NAND(g7257, I13638)
--	I10329 = NAND(g2562, I10327)
--	g6215 = NAND(I10981, I10982)
--	I6904 = NAND(g2105, g1838)
--	I13638 = NAND(g7257, g7069)
--	I10328 = NAND(g5467, I10327)
--	g5750 = NAND(I10314, I10315)
--	I7480 = NAND(g3808, I7478)
--	I11841 = NAND(g2548, g6158)
--	I7569 = NAND(g3780, I7567)
--	I9964 = NAND(g1938, I9963)
--	g3525 = NAND(I7010, I7011)
--	g4332 = NAND(g3681, g2368)
--	g7535 = NAND(I13786, I13787)
--	I6757 = NAND(g186, g1983)
--	I12051 = NAND(g5956, g5939)
--	g3358 = NAND(I6940, I6941)
--	I11116 = NAND(g5481, I11115)
--	I11615 = NAND(g6239, I11614)
--	I6522 = NAND(g1919, g1102)
--	I9057 = NAND(g4059, g1504)
--	I10991 = NAND(g5632, g2389)
--	I9549 = NAND(g4307, I9547)
--	I8255 = NAND(g3825, I8253)
--	g4492 = NAND(I8537, I8538)
--	g4714 = NAND(g4344, g4335, g4328)
--	I11142 = NAND(g5493, g3062)
--	I7423 = NAND(g2703, I7421)
--	I11165 = NAND(g3029, I11163)
--	I6234 = NAND(g896, I6232)
--	I10744 = NAND(g5550, I10743)
--	g5555 = NAND(I9979, I9980)
--	I10849 = NAND(g2595, I10847)
--	g4889 = NAND(I9242, I9243)
--	g4476 = NAND(I8511, I8512)
--	g6142 = NAND(I10790, I10791)
--	I10848 = NAND(g5490, I10847)
--	g4871 = NAND(g3635, g3605, g4220, g3644)
--	g6497 = NAND(g5278, g5847)
--	I7240 = NAND(g1658, I7239)
--	g5567 = NAND(g1879, g4883)
--	I10361 = NAND(g1118, I10359)
--	I7443 = NAND(g2973, g1701)
--	I13600 = NAND(g7244, I13598)
--	I9691 = NAND(g5096, g1037)
--	g6218 = NAND(I10992, I10993)
--	g4231 = NAND(g2276, g3258)
--	I11137 = NAND(g3052, I11135)
--	I7533 = NAND(g3787, I7531)
--	I11873 = NAND(g2543, g6187)
--	I12552 = NAND(g1462, I12550)
--	I9985 = NAND(g4836, g2096)
--	I11614 = NAND(g6239, g1519)
--	g7093 = NAND(I12870, I12871)
--	g9191 = NAND(I15856, I15857)
--	I6843 = NAND(g205, I6842)
--	I8119 = NAND(g1904, g3220)
--	I11122 = NAND(g5517, g2712)
--	I8152 = NAND(g38, I8150)
--	I7460 = NAND(g2506, I7459)
--	I14473 = NAND(g8147, I14472)
--	I10789 = NAND(g5512, g2170)
--	I7937 = NAND(g3614, g1138)
--	I11136 = NAND(g5476, I11135)
--	I6232 = NAND(g834, g896)
--	I7479 = NAND(g2502, I7478)
--	I10359 = NAND(g5552, g1118)
--	I6813 = NAND(g210, g2052)
--	g1759 = NAND(I5599, I5600)
--	g5558 = NAND(I10000, I10001)
--	I6740 = NAND(g195, I6739)
--	g4513 = NAND(I8582, I8583)
--	I11164 = NAND(g5469, I11163)
--	I8939 = NAND(g4239, I8938)
--	g6119 = NAND(I10744, I10745)
--	g7257 = NAND(I13214, I13215)
--	I7156 = NAND(g2331, g929)
--	g4679 = NAND(I8939, I8940)
--	I11575 = NAND(g5894, I11574)
--	g3518 = NAND(I6997, I6998)
--	I8636 = NAND(g2481, I8635)
--	g4831 = NAND(g3635, g3605, g4220)
--	I11109 = NAND(g5522, I11108)
--	g6893 = NAND(I12551, I12552)
--	I11108 = NAND(g5522, g2734)
--	g6274 = NAND(I11102, I11103)
--	I9151 = NAND(g3883, g1649)
--	I7453 = NAND(g3226, I7452)
--	g6170 = NAND(I10874, I10875)
--	I11750 = NAND(g6112, g1486)
--	I7568 = NAND(g2481, I7567)
--	g6280 = NAND(I11136, I11137)
--	I7157 = NAND(g2331, I7156)
--	I8637 = NAND(g2743, I8635)
--	g4869 = NAND(g4254, g3533)
--	I8536 = NAND(g2506, g2798)
--	I9278 = NAND(g4313, I9276)
--	g3658 = NAND(I7149, I7150)
--	g6187 = NAND(g5633, g3735, g3716)
--	I6275 = NAND(g906, I6273)
--	I9235 = NAND(g2180, I9233)
--	I10981 = NAND(g5625, I10980)
--	g2395 = NAND(I6274, I6275)
--	I9693 = NAND(g1037, I9691)
--	I9548 = NAND(g1952, I9547)
--	g7480 = NAND(I13639, I13640)
--	I10899 = NAND(g5520, g2752)
--	g1678 = NAND(I5506, I5507)
--	I11757 = NAND(g1758, g6118)
--	g5672 = NAND(g5056, g5039, g5023)
--	g6695 = NAND(I12016, I12017)
--	g3680 = NAND(I7187, I7188)
--	g1682 = NAND(I5520, I5521)
--	g6159 = NAND(I10835, I10836)
--	I8537 = NAND(g2506, I8536)
--	I13397 = NAND(g1057, I13395)
--	I6905 = NAND(g2105, I6904)
--	I8243 = NAND(g2011, g3506)
--	I8328 = NAND(g2721, I8326)
--	g2783 = NAND(I6523, I6524)
--	I9965 = NAND(g4869, I9963)
--	I6750 = NAND(g1733, g1494)
--	I13213 = NAND(g7065, g7082)
--	g5712 = NAND(I10224, I10225)
--	g4745 = NAND(I9070, I9071)
--	I11574 = NAND(g5894, g1122)
--	g4309 = NAND(g3002, g3124, g3659)
--	I10061 = NAND(g4910, I10060)
--	I7616 = NAND(g3008, g1721)
--	I8512 = NAND(g2807, I8510)
--	g3889 = NAND(I7437, I7438)
--	I10360 = NAND(g5552, I10359)
--	I8166 = NAND(g3231, I8164)
--	I7503 = NAND(g2498, g3802)
--	g3722 = NAND(I7215, I7216)
--	g4575 = NAND(I8679, I8680)
--	I15863 = NAND(g9174, I15862)
--	I13396 = NAND(g7212, I13395)
--	I14472 = NAND(g8147, g1069)
--	I14246 = NAND(g1065, I14244)
--	I7277 = NAND(g2497, g1898)
--	I10071 = NAND(g4954, g2253)
--	I6172 = NAND(g911, I6170)
--	I7617 = NAND(g3008, I7616)
--	g6902 = NAND(I12576, I12577)
--	I9153 = NAND(g1649, I9151)
--	g7316 = NAND(I13377, I13378)
--	g3231 = NAND(g1889, g1904)
--	I6134 = NAND(g846, I6133)
--	I12080 = NAND(g5971, I12078)
--	I7892 = NAND(g2979, I7891)
--	I8393 = NAND(g2949, I8392)
--	g1910 = NAND(g1435, g1439)
--	I13787 = NAND(g1477, I13785)
--	I12031 = NAND(g5918, g5897)
--	g5632 = NAND(g2276, g4901)
--	g5095 = NAND(I9476, I9477)
--	g4881 = NAND(g2460, g4315)
--	g2352 = NAND(I6171, I6172)
--	I7140 = NAND(g2397, I7138)
--	g6463 = NAND(g5918, g5278)
--	I7478 = NAND(g2502, g3808)
--	I8121 = NAND(g3220, I8119)
--	I6202 = NAND(g831, I6201)
--	I13640 = NAND(g7069, I13638)
--	g3613 = NAND(I7086, I7087)
--	g5752 = NAND(I10328, I10329)
--	I12869 = NAND(g2536, g6618)
--	I8253 = NAND(g2454, g3825)
--	I8938 = NAND(g4239, g1545)
--	I6776 = NAND(g1134, I6774)
--	I8606 = NAND(g2487, I8605)
--	I7214 = NAND(g815, g2091)
--	g4305 = NAND(g3712, g3700, g3732)
--	I9476 = NAND(g4038, I9475)
--	I13003 = NAND(g7010, I13002)
--	I6996 = NAND(g2275, g2242)
--	g5189 = NAND(I9692, I9693)
--	I13786 = NAND(g7427, I13785)
--	I6878 = NAND(g1910, I6876)
--	g3679 = NAND(I7180, I7181)
--	I8607 = NAND(g2764, I8605)
--	I8659 = NAND(g2471, I8658)
--	I9477 = NAND(g1942, I9475)
--	g4227 = NAND(I8133, I8134)
--	I6997 = NAND(g2275, I6996)
--	I12079 = NAND(g5988, I12078)
--	g6570 = NAND(I11751, I11752)
--	I12078 = NAND(g5988, g5971)
--	I12598 = NAND(g1126, I12596)
--	I10889 = NAND(g5590, I10888)
--	I10980 = NAND(g5625, g2210)
--	I10888 = NAND(g5590, g2259)
--	g2315 = NAND(I6103, I6104)
--	g4502 = NAND(I8559, I8560)
--	g6158 = NAND(g3735, g3716, g5633, g3754)
--	g5575 = NAND(I10039, I10040)
--	I11149 = NAND(g5473, g3038)
--	I8559 = NAND(g2502, I8558)
--	g6275 = NAND(I11109, I11110)
--	g6615 = NAND(I11842, I11843)
--	I7150 = NAND(g1974, I7148)
--	g5539 = NAND(I9947, I9948)
--	I7438 = NAND(g3822, I7436)
--	I7009 = NAND(g2295, g2333)
--	I15862 = NAND(g9174, g9171)
--	I12017 = NAND(g5847, I12015)
--	g6284 = NAND(I11164, I11165)
--	g6180 = NAND(I10900, I10901)
--	g4741 = NAND(I9058, I9059)
--	I9946 = NAND(g2128, g4905)
--	g4910 = NAND(g2460, g4314)
--	I10625 = NAND(g5314, g1514)
--	g2330 = NAND(I6134, I6135)
--	g6559 = NAND(g5814, g6109)
--	g3012 = NAND(I6758, I6759)
--	g9202 = NAND(I15881, I15882)
--	g3706 = NAND(g1556, g2510)
--	I9182 = NAND(g4231, I9181)
--	I9382 = NAND(g4062, I9381)
--	I10060 = NAND(g4910, g2226)
--	I10197 = NAND(g4724, I10196)
--	I6500 = NAND(g1913, I6499)
--	I10855 = NAND(g5521, I10854)
--	I8151 = NAND(g3229, I8150)
--	I13378 = NAND(g1472, I13376)
--	I9947 = NAND(g2128, I9946)
--	I11096 = NAND(g2734, I11094)
--	I10867 = NAND(g5480, I10866)
--	I5505 = NAND(g1532, g1528)
--	I13802 = NAND(g1061, I13800)
--	I10315 = NAND(g1041, I10313)
--	g5305 = NAND(g5009, g4335, g4328)
--	I6523 = NAND(g1919, I6522)
--	I10819 = NAND(g5567, I10818)
--	I12016 = NAND(g5874, I12015)
--	I10818 = NAND(g5567, g2039)
--	g5748 = NAND(I10306, I10307)
--	I11549 = NAND(g5984, g1045)
--	g9179 = NAND(I15818, I15819)
--	I7085 = NAND(g1753, g1918)
--	I7485 = NAND(g2989, g1708)
--	I6104 = NAND(g921, I6102)
--	I6499 = NAND(g1913, g1537)
--	g4256 = NAND(g3233, g1444)
--	I8134 = NAND(g1646, I8132)
--	g7503 = NAND(I13686, I13687)
--	I10094 = NAND(g2177, I10092)
--	I6273 = NAND(g840, g906)
--	g2367 = NAND(I6202, I6203)
--	g4700 = NAND(g2460, g4271)
--	I13002 = NAND(g7010, g1053)
--	I9233 = NAND(g4310, g2180)
--	I10019 = NAND(g2174, I10017)
--	g4263 = NAND(g3260, g1435)
--	I10196 = NAND(g4724, g1958)
--	I10018 = NAND(g4700, I10017)
--	g6282 = NAND(I11150, I11151)
--	I10866 = NAND(g5480, g2605)
--	I7270 = NAND(g955, I7268)
--	I10001 = NAND(g1929, I9999)
--	I7610 = NAND(g2471, I7609)
--	I9171 = NAND(g4244, I9169)
--	I10923 = NAND(g5525, g2752)
--	I7069 = NAND(g1639, I7068)
--	I10300 = NAND(g2562, I10298)
--	g7244 = NAND(g7050, g3757, g3739)
--	I7540 = NAND(g1715, I7538)
--	g7140 = NAND(I13003, I13004)
--	g5689 = NAND(I10197, I10198)
--	I9745 = NAND(g4826, g1549)
--	I9963 = NAND(g1938, g4869)
--	g7082 = NAND(I12853, I12854)
--	I6135 = NAND(g916, I6133)
--	g3678 = NAND(I7173, I7174)
--	I15881 = NAND(g9190, I15880)
--	I11080 = NAND(g2511, I11078)
--	I10854 = NAND(g5521, g2584)
--	I6916 = NAND(g2360, g1732)
--	g5564 = NAND(I10018, I10019)
--	I8658 = NAND(g2471, g2724)
--	I5696 = NAND(g1513, I5695)
--	I7510 = NAND(g2992, g1711)
--	I12853 = NAND(g6701, I12852)
--	g4474 = NAND(I8503, I8504)
--	I10314 = NAND(g5484, I10313)
--	I6102 = NAND(g849, g921)
--	I11843 = NAND(g6158, I11841)
--	I10307 = NAND(g3019, I10305)
--	g5589 = NAND(I10061, I10062)
--	I8132 = NAND(g3232, g1646)
--	I8680 = NAND(g2706, I8678)
--	g3602 = NAND(I7069, I7070)
--	I6752 = NAND(g1494, I6750)
--	I6917 = NAND(g2360, I6916)
--	g1775 = NAND(I5620, I5621)
--	I7215 = NAND(g815, I7214)
--	g3767 = NAND(I7240, I7241)
--	I5697 = NAND(g1524, I5695)
--	I8558 = NAND(g2502, g2790)
--	I12053 = NAND(g5939, I12051)
--	I6233 = NAND(g834, I6232)
--	I10335 = NAND(g5462, I10334)
--	g9205 = NAND(I15898, I15899)
--	I8511 = NAND(g2517, I8510)
--	I10993 = NAND(g2389, I10991)
--	I14839 = NAND(g1073, I14837)
--	g5538 = NAND(g5132, g1266)
--	I15897 = NAND(g9202, g9203)
--	I14838 = NAND(g8660, I14837)
--	g7237 = NAND(g7050, g3739)
--	I9070 = NAND(g4400, I9069)
--	g6153 = NAND(I10819, I10820)
--	g6680 = NAND(g5403, g6252)
--	g8239 = NAND(g8073, g8092)
--	I11171 = NAND(g5477, I11170)
--	I6171 = NAND(g843, I6170)
--	I10039 = NAND(g4893, I10038)
--	I10306 = NAND(g5470, I10305)
--	I10038 = NAND(g4893, g2202)
--	g3028 = NAND(I6775, I6776)
--	I11079 = NAND(g5697, I11078)
--	I7891 = NAND(g2979, g1499)
--	I10143 = NAND(g4707, I10142)
--	I13599 = NAND(g2551, I13598)
--	I11078 = NAND(g5697, g2511)
--	I13598 = NAND(g2551, g7244)
--	g5562 = NAND(I10010, I10011)
--	I10791 = NAND(g2170, I10789)
--	I15850 = NAND(g9154, I15848)
--	I8339 = NAND(g2966, I8338)
--	g5257 = NAND(I9768, I9769)
--	I6759 = NAND(g1983, I6757)
--	g5605 = NAND(I10093, I10094)
--	g3883 = NAND(g2276, g3188)
--	I11158 = NAND(g3052, I11156)
--	I6201 = NAND(g831, g891)
--	I9169 = NAND(g1935, g4244)
--	g5751 = NAND(I10321, I10322)
--	I9059 = NAND(g1504, I9057)
--	g6476 = NAND(g5939, g5269)
--	I11144 = NAND(g3062, I11142)
--	I9767 = NAND(g4832, g1114)
--	g6722 = NAND(I12079, I12080)
--	I10223 = NAND(g2522, g4895)
--	g6285 = NAND(I11171, I11172)
--	I12577 = NAND(g1049, I12575)
--	I6539 = NAND(g2555, I6538)
--	I10321 = NAND(g5459, I10320)
--	I13017 = NAND(g6941, I13016)
--	g6424 = NAND(I11550, I11551)
--	I10953 = NAND(g5565, I10952)
--	I15857 = NAND(g9165, I15855)
--	g6477 = NAND(g5269, g5918)
--	g4820 = NAND(I9170, I9171)
--	I10334 = NAND(g5462, g2573)
--	I13687 = NAND(g7237, I13685)
--	I11752 = NAND(g1486, I11750)
--	I7068 = NAND(g1639, g1643)
--	I12852 = NAND(g6701, g6695)
--	I7468 = NAND(g1704, I7466)
--	g6273 = NAND(I11095, I11096)
--	I9826 = NAND(g4729, g1509)
--	I8660 = NAND(g2724, I8658)
--	I10000 = NAND(g4839, I9999)
--	I10908 = NAND(g2605, I10906)
--	I11842 = NAND(g2548, I11841)
--	I7576 = NAND(g1718, I7574)
--	I7149 = NAND(g799, I7148)
--	I12576 = NAND(g6574, I12575)
--	I13016 = NAND(g6941, g1142)
--	g4294 = NAND(I8244, I8245)
--	I8679 = NAND(g2467, I8678)
--	I7241 = NAND(g2134, I7239)
--	I12052 = NAND(g5956, I12051)
--	I15856 = NAND(g9168, I15855)
--	I15880 = NAND(g9190, g9179)
--	I10992 = NAND(g5632, I10991)
--	I9827 = NAND(g4729, I9826)
--	g7069 = NAND(g5435, g6680)
--	I11124 = NAND(g2712, I11122)
--	I8560 = NAND(g2790, I8558)
--	g4954 = NAND(g4319, g2460)
--	g4810 = NAND(I9152, I9153)
--	g7540 = NAND(I13801, I13802)
--	g4363 = NAND(I8339, I8340)
--	I13686 = NAND(g1977, I13685)
--	I9196 = NAND(g1652, I9194)
--	I10835 = NAND(g5514, I10834)
--	g6178 = NAND(g2205, g5568)
--	I7893 = NAND(g1499, I7891)
--	I7186 = NAND(g2353, g1834)
--	I11875 = NAND(g6187, I11873)
--	g4912 = NAND(I9277, I9278)
--	g3890 = NAND(I7444, I7445)
--	I9994 = NAND(g4871, I9992)
--	g3011 = NAND(I6751, I6752)
--	I7939 = NAND(g1138, I7937)
--	I6203 = NAND(g891, I6201)
--	I9181 = NAND(g4231, g2007)
--	g5753 = NAND(I10335, I10336)
--	I8164 = NAND(g1943, g3231)
--	I9381 = NAND(g4062, g1908)
--	I15887 = NAND(g9192, g9191)
--	g7144 = NAND(I13017, I13018)
--	I10142 = NAND(g4707, g1916)
--	I6940 = NAND(g2161, I6939)
--	I7187 = NAND(g2353, I7186)
--	I7461 = NAND(g3815, I7459)
--	g5565 = NAND(g2044, g4933)
--	g5681 = NAND(g5132, g2043)
--	g6265 = NAND(I11079, I11080)
--	g5697 = NAND(g2044, g5005)
--	I11170 = NAND(g5477, g3038)
--	g6164 = NAND(I10848, I10849)
--	I8956 = NAND(g4246, I8955)
--	I6741 = NAND(g1970, I6739)
--	g6770 = NAND(I12180, I12181)
--	I13589 = NAND(g7234, I13587)
--	I13588 = NAND(g2556, I13587)
--	I8338 = NAND(g2966, g1698)
--	g3924 = NAND(I7568, I7569)
--	I10952 = NAND(g5565, g2340)
--	I6758 = NAND(g186, I6757)
--	I6066 = NAND(g883, I6064)
--	g7065 = NAND(I12833, I12834)
--	I11616 = NAND(g1519, I11614)
--	I10790 = NAND(g5512, I10789)
--	I9058 = NAND(g4059, I9057)
--	I10873 = NAND(g5516, g2595)
--	I8957 = NAND(g1110, I8955)
--	g3665 = NAND(I7157, I7158)
--	I6133 = NAND(g846, g916)
--	g6281 = NAND(I11143, I11144)
--	I6774 = NAND(g2386, g1134)
--	I11101 = NAND(g5491, g2712)
--	I11177 = NAND(g5466, g3019)
--	I10834 = NAND(g5514, g2584)
--	I6538 = NAND(g2555, g2557)
--	I9992 = NAND(g2145, g4871)
--	I11874 = NAND(g2543, I11873)
--	I15817 = NAND(g9151, g9148)
--	I12833 = NAND(g6722, I12832)
--	I10320 = NAND(g5459, g2573)
--	I10073 = NAND(g2253, I10071)
--	g8231 = NAND(I14473, I14474)
--	g5363 = NAND(I9827, I9828)
--	g3681 = NAND(g866, g2368)
--	I8504 = NAND(g2038, I8502)
--	g3914 = NAND(I7532, I7533)
--	I12951 = NAND(g7003, g1467)
--	g5568 = NAND(g2044, g4902, g4320)
--	I12033 = NAND(g5897, I12031)
--	I8470 = NAND(g2525, g2821)
--	I7512 = NAND(g1711, I7510)
--	g9203 = NAND(I15888, I15889)
--	I11185 = NAND(g5474, I11184)
--	g4244 = NAND(g3549, g3533)
--	I6257 = NAND(g837, g901)
--	I7148 = NAND(g799, g1974)
--	I9183 = NAND(g2007, I9181)
--	I9383 = NAND(g1908, I9381)
--	I14474 = NAND(g1069, I14472)
--	I8678 = NAND(g2467, g2706)
--	I10327 = NAND(g5467, g2562)
--	g7828 = NAND(I14245, I14246)
--	I8635 = NAND(g2481, g2743)
--	I6751 = NAND(g1733, I6750)
--	g6504 = NAND(g5269, g5874)
--	I13215 = NAND(g7082, I13213)
--	g2378 = NAND(I6233, I6234)
--	I10982 = NAND(g2210, I10980)
--	I7279 = NAND(g1898, I7277)
--	I9999 = NAND(g4839, g1929)
--	g4110 = NAND(I7938, I7939)
--	g4310 = NAND(g3666, g2460)
--	g4824 = NAND(I9182, I9183)
--	g5661 = NAND(I10143, I10144)
--	I8582 = NAND(g2498, I8581)
--	I7938 = NAND(g3614, I7937)
--	I5620 = NAND(g1092, I5619)
--	I10040 = NAND(g2202, I10038)
--	g8798 = NAND(g6984, g8644)
--	g4563 = NAND(I8659, I8660)
--	g6169 = NAND(I10867, I10868)
--	g6283 = NAND(I11157, I11158)
--	g4237 = NAND(I8151, I8152)
--	I11576 = NAND(g1122, I11574)
--	I8502 = NAND(g2986, g2038)
--	I10847 = NAND(g5490, g2595)
--	I8940 = NAND(g1545, I8938)
--	I10062 = NAND(g2226, I10060)
--	I11115 = NAND(g5481, g3062)
--	g5546 = NAND(I9964, I9965)
--	g7325 = NAND(I13396, I13397)
--	I5520 = NAND(g1087, I5519)
--	g6203 = NAND(I10953, I10954)
--	I11184 = NAND(g5474, g3029)
--	I7158 = NAND(g929, I7156)
--	I6924 = NAND(g1728, I6923)
--	I12832 = NAND(g6722, g6709)
--	I10072 = NAND(g4954, I10071)
--	g4836 = NAND(g4288, g1879)
--	g3894 = NAND(I7460, I7461)
--	g6188 = NAND(I10924, I10925)
--	I7174 = NAND(g2006, I7172)
--	I13214 = NAND(g7065, I13213)
--	I10820 = NAND(g2039, I10818)
--	I7239 = NAND(g1658, g2134)
--	I8165 = NAND(g1943, I8164)
--	I7180 = NAND(g2351, I7179)
--	I6103 = NAND(g849, I6102)
--	I8133 = NAND(g3232, I8132)
--	g1819 = NAND(I5696, I5697)
--	I12032 = NAND(g5918, I12031)
--	g5035 = NAND(I9382, I9383)
--	I9954 = NAND(g2131, I9953)
--	I8538 = NAND(g2798, I8536)
--	I15864 = NAND(g9171, I15862)
--	I12871 = NAND(g6618, I12869)
--	g6466 = NAND(I11615, I11616)
--	g7447 = NAND(I13599, I13600)
--	g6165 = NAND(I10855, I10856)
--	g6571 = NAND(I11758, I11759)
--	g5310 = NAND(g5009, g4335, g4963)
--	g4298 = NAND(I8254, I8255)
--	I10743 = NAND(g5550, g2100)
--	g5762 = NAND(I10360, I10361)
--	g3925 = NAND(I7575, I7576)
--	g5590 = NAND(g2044, g4906)
--	I11759 = NAND(g6118, I11757)
--	g5657 = NAND(g5021, g4381)
--	I11758 = NAND(g1758, I11757)
--	g6467 = NAND(g5956, g5269)
--	g5556 = NAND(I9986, I9987)
--	g4219 = NAND(I8120, I8121)
--	g2385 = NAND(I6258, I6259)
--	g7234 = NAND(g3757, g3739, g7050, g3770)
--	g4252 = NAND(g2276, g3313)
--	g3906 = NAND(I7504, I7505)
--	I6775 = NAND(g2386, I6774)
--	I7010 = NAND(g2295, I7009)
--	I10890 = NAND(g2259, I10888)
--	I8605 = NAND(g2487, g2764)
--	g6181 = NAND(I10907, I10908)
--	g4911 = NAND(g4320, g2044)
--	I9475 = NAND(g4038, g1942)
--	I6739 = NAND(g195, g1970)
--	I7172 = NAND(g1739, g2006)
--	I7278 = NAND(g2497, I7277)
--	I11135 = NAND(g5476, g3052)
--	I7618 = NAND(g1721, I7616)
--	g2801 = NAND(I6539, I6540)
--	g5557 = NAND(I9993, I9994)
--	g3907 = NAND(I7511, I7512)
--	I6501 = NAND(g1537, I6499)
--	I13004 = NAND(g1053, I13002)
--	I9276 = NAND(g2533, g4313)
--	g3656 = NAND(I7139, I7140)
--	g3915 = NAND(I7539, I7540)
--	g4399 = NAND(I8393, I8394)
--	I9986 = NAND(g4836, I9985)
--	I7567 = NAND(g2481, g3780)
--	I9277 = NAND(g2533, I9276)
--	I11163 = NAND(g5469, g3029)
--	I12551 = NAND(g6689, I12550)
--	g7121 = NAND(I12952, I12953)
--	I9987 = NAND(g2096, I9985)
--	g3899 = NAND(I7479, I7480)
--	I9547 = NAND(g1952, g4307)
--	I7179 = NAND(g2351, g795)
--	I8326 = NAND(g2011, g2721)
--	I12181 = NAND(g6163, I12179)
--	I10011 = NAND(g4821, I10009)
--	I7611 = NAND(g3771, I7609)
--	I10627 = NAND(g1514, I10625)
--	g4887 = NAND(I9234, I9235)
--	g4228 = NAND(g1408, g2665)
--	I10925 = NAND(g2752, I10923)
--	I6998 = NAND(g2242, I6996)
--	I8327 = NAND(g2011, I8326)
--	g6023 = NAND(I10626, I10627)
--	I7511 = NAND(g2992, I7510)
--	g2333 = NAND(g985, g990)
--	I8472 = NAND(g2821, I8470)
--	I7574 = NAND(g2999, g1718)
--	g9190 = NAND(I15849, I15850)
--	I12870 = NAND(g2536, I12869)
--	I6925 = NAND(g33, I6923)
--	I13395 = NAND(g7212, g1057)
--	g5540 = NAND(I9954, I9955)
--	I10626 = NAND(g5314, I10625)
--	I14245 = NAND(g7683, I14244)
--	I10299 = NAND(g5461, I10298)
--	g3895 = NAND(I7467, I7468)
--	I10298 = NAND(g5461, g2562)
--	g6472 = NAND(g5971, g5269)
--	I6906 = NAND(g1838, I6904)
--	I5599 = NAND(g1481, I5598)
--	I9194 = NAND(g4252, g1652)
--	I10856 = NAND(g2584, I10854)
--	I15882 = NAND(g9179, I15880)
--	I7139 = NAND(g2404, I7138)
--	I9071 = NAND(g1149, I9069)
--	I9242 = NAND(g2540, I9241)
--	g5291 = NAND(g4344, g5002, g4963)
--	I9948 = NAND(g4905, I9946)
--	I8581 = NAND(g2498, g2777)
--	I9955 = NAND(g4831, I9953)
--	g2751 = NAND(I6500, I6501)
--	I6876 = NAND(g1967, g1910)
--	I9769 = NAND(g1114, I9767)
--	I10080 = NAND(g2256, I10078)
--	I10924 = NAND(g5525, I10923)
--	I15849 = NAND(g9162, I15848)
--	g3286 = NAND(I6905, I6906)
--	I15848 = NAND(g9162, g9154)
--	I9993 = NAND(g2145, I9992)
--	I12597 = NAND(g6582, I12596)
--	I5695 = NAND(g1513, g1524)
--	I7444 = NAND(g2973, I7443)
--	I7269 = NAND(g2486, I7268)
--	I10198 = NAND(g1958, I10196)
--	g5594 = NAND(I10072, I10073)
--	I13785 = NAND(g7427, g1477)
--	I6877 = NAND(g1967, I6876)
--	I10868 = NAND(g2605, I10866)
--	g2474 = NAND(g1405, g1412)
--	I12854 = NAND(g6695, I12852)
--	I10225 = NAND(g4895, I10223)
--	I11151 = NAND(g3038, I11149)
--	I11172 = NAND(g3038, I11170)
--	I6064 = NAND(g852, g883)
--	g4893 = NAND(g2460, g4312)
--	g5550 = NAND(g1879, g4830)
--	I14244 = NAND(g7683, g1065)
--	g3900 = NAND(I7486, I7487)
--	g6163 = NAND(g5633, g3716)
--	I7436 = NAND(g2517, g3822)
--	I12550 = NAND(g6689, g1462)
--	g4821 = NAND(g4220, g3605)
--	I6844 = NAND(g2016, I6842)
--	I12596 = NAND(g6582, g1126)
--	I7422 = NAND(g2525, I7421)
--	I13377 = NAND(g7199, I13376)
--	I12180 = NAND(g1961, I12179)
--	I10010 = NAND(g1949, I10009)
--	g3886 = NAND(I7422, I7423)
--	I6814 = NAND(g210, I6813)
--	I10079 = NAND(g4911, I10078)
--	I7437 = NAND(g2517, I7436)
--	g3314 = NAND(I6917, I6918)
--	I10078 = NAND(g4911, g2256)
--	g5312 = NAND(g5009, g5002, g4963)
--	I10322 = NAND(g2573, I10320)
--	g2051 = NAND(g1444, g1450)
--	I10901 = NAND(g2752, I10899)
--	I6918 = NAND(g1732, I6916)
--	I9980 = NAND(g2092, I9978)
--	I9069 = NAND(g4400, g1149)
--	I8583 = NAND(g2777, I8581)
--	g4359 = NAND(I8327, I8328)
--	I10144 = NAND(g1916, I10142)
--	I11551 = NAND(g1045, I11549)
--	g3887 = NAND(I7429, I7430)
--	I7454 = NAND(g1106, I7452)
--	I10336 = NAND(g2573, I10334)
--	g6627 = NAND(I11874, I11875)
--	I7532 = NAND(g2487, I7531)
--	I10017 = NAND(g4700, g2174)
--	I5619 = NAND(g1092, g1130)
--	I13376 = NAND(g7199, g1472)
--	I11103 = NAND(g2712, I11101)
--	I11095 = NAND(g5515, I11094)
--	g8633 = NAND(g8176, g6232)
--	I8503 = NAND(g2986, I8502)
--	g4880 = NAND(g4287, g1879)
--	g5576 = NAND(g4894, g4888, g4884)
--	I10224 = NAND(g2522, I10223)
--	I7429 = NAND(g3222, I7428)
--	I8120 = NAND(g1904, I8119)
--	I12015 = NAND(g5874, g5847)
--	I5598 = NAND(g1481, g1489)
--	g6276 = NAND(I11116, I11117)
--	g4243 = NAND(I8165, I8166)
--	g5747 = NAND(I10299, I10300)
--	I6842 = NAND(g205, g2016)
--	I7138 = NAND(g2404, g2397)
--	I10954 = NAND(g2340, I10952)
--	I6941 = NAND(g2051, I6939)
--	g6503 = NAND(g5269, g5897)
--	I5519 = NAND(g1087, g1098)
--	I12179 = NAND(g1961, g6163)
--	g8681 = NAND(I14838, I14839)
--	I15899 = NAND(g9203, I15897)
--	I15898 = NAND(g9202, I15897)
--	I12953 = NAND(g1467, I12951)
--	I8244 = NAND(g2011, I8243)
--	g6277 = NAND(I11123, I11124)
--	I7575 = NAND(g2999, I7574)
--	I8340 = NAND(g1698, I8338)
--	g4090 = NAND(I7892, I7893)
--	I9768 = NAND(g4832, I9767)
--	g6516 = NAND(g5897, g5278)
--	g3129 = NAND(I6843, I6844)
--	g4456 = NAND(I8471, I8472)
--	I7539 = NAND(g2996, I7538)
--	g2995 = NAND(I6740, I6741)
--	g2294 = NAND(I6065, I6066)
--	g3221 = NAND(I6877, I6878)
--	I7268 = NAND(g2486, g955)
--	I5506 = NAND(g1532, I5505)
--	I7452 = NAND(g3226, g1106)
--	g6709 = NAND(I12052, I12053)
--	I6540 = NAND(g2557, I6538)
--	I10093 = NAND(g4881, I10092)
--	I9195 = NAND(g4252, I9194)
--	I7086 = NAND(g1753, I7085)
--	I7486 = NAND(g2989, I7485)
--	g6435 = NAND(I11575, I11576)
--	g6482 = NAND(g5269, g5847)
--	I7504 = NAND(g2498, I7503)
--	I10875 = NAND(g2595, I10873)
--	I7070 = NAND(g1643, I7068)
--	I14837 = NAND(g8660, g1073)
--	g4686 = NAND(I8956, I8957)
--	I11094 = NAND(g5515, g2734)
--	I5507 = NAND(g1528, I5505)
--	I11150 = NAND(g5473, I11149)
--	I13801 = NAND(g7429, I13800)
--	I9692 = NAND(g5096, I9691)
--	g7444 = NAND(I13588, I13589)
--	I13018 = NAND(g1142, I13016)
--	I6259 = NAND(g901, I6257)
--	I7087 = NAND(g1918, I7085)
--	I7487 = NAND(g1708, I7485)
--	I6923 = NAND(g1728, g33)
--	g3818 = NAND(I7278, I7279)
--	I8394 = NAND(g1925, I8392)
--	I9979 = NAND(g4880, I9978)
--	g3893 = NAND(I7453, I7454)
--	I7445 = NAND(g1701, I7443)
--	I7173 = NAND(g1739, I7172)
--	I8471 = NAND(g2525, I8470)
--	I9828 = NAND(g1509, I9826)
--	g5595 = NAND(I10079, I10080)
--	I8955 = NAND(g4246, g1110)
--	g9192 = NAND(I15863, I15864)
--	I8254 = NAND(g2454, I8253)
--	I10836 = NAND(g2584, I10834)
--	I9746 = NAND(g4826, I9745)
--	I7459 = NAND(g2506, g3815)
--	I11102 = NAND(g5491, I11101)
--	I11157 = NAND(g5482, I11156)
--	g3939 = NAND(I7617, I7618)
--	I8150 = NAND(g3229, g38)
--	g3083 = NAND(I6814, I6815)
--	I9953 = NAND(g2131, g4831)
--	g4879 = NAND(g2595, g2584, g4270, g4281)
--	I10313 = NAND(g5484, g1041)
--	I6065 = NAND(g852, I6064)
--	I10305 = NAND(g5470, g3019)
--	I10900 = NAND(g5520, I10899)
--	I9747 = NAND(g1549, I9745)
--	g8627 = NAND(g6232, g8091)
--	I11550 = NAND(g5984, I11549)
--	I9241 = NAND(g2540, g4305)
--	g5512 = NAND(g1879, g4877)
--	I7188 = NAND(g1834, I7186)
--	I10874 = NAND(g5516, I10873)
--	I7216 = NAND(g2091, I7214)
--	I12952 = NAND(g7003, I12951)
--	I7428 = NAND(g3222, g1541)
--	I10009 = NAND(g1949, g4821)
--	I7430 = NAND(g1541, I7428)
--	I11156 = NAND(g5482, g3052)
--	I9152 = NAND(g3883, I9151)
--	I5621 = NAND(g1130, I5619)
--	I6815 = NAND(g2052, I6813)
--	g4905 = NAND(g4282, g3533)
--	g3811 = NAND(I7269, I7270)
--	g3315 = NAND(I6924, I6925)
--	I10907 = NAND(g5492, I10906)
--	I7609 = NAND(g2471, g3771)
--	I12834 = NAND(g6709, I12832)
--	I8392 = NAND(g2949, g1925)
--	I9170 = NAND(g1935, I9169)
--	I15889 = NAND(g9191, I15887)
--	
--	g4884 = NOR(g4492, g4476, g4456, g4294)
--	g8656 = NOR(g8199, I14758, I14759)
--	g3260 = NOR(g1728, g2490)
--	g5615 = NOR(g4714, g3002)
--	g8236 = NOR(g8199, I14495, I14496)
--	g4160 = NOR(g1231, g2834)
--	g7406 = NOR(g7191, g1600)
--	g6259 = NOR(g3002, g5312)
--	g6465 = NOR(g5403, g5802, g5769, g5790)
--	g3515 = NOR(g1388, g2262, g2230, g2214)
--	g8812 = NOR(g8443, g8421, I15086)
--	g3528 = NOR(g2343, g1391)
--	g8073 = NOR(g7658, g7654)
--	g3555 = NOR(g2359, g1398)
--	g8819 = NOR(g8443, g8421, I15113)
--	g8694 = NOR(g7658, g8613, g7634)
--	g8806 = NOR(g8443, g8421, I15044)
--	g8230 = NOR(g8199, I14467, I14468)
--	g8807 = NOR(g8443, g8421, I15055)
--	g4888 = NOR(g4548, g4528, g4513, g4502)
--	g8859 = NOR(g8493, g8239, I15165)
--	g7326 = NOR(g7194, g6999)
--	g8699 = NOR(g7658, g8613, g7634)
--	g8855 = NOR(g7658, g8613, g7634)
--	g8644 = NOR(g4146, g8128)
--	g6193 = NOR(g1926, g5310)
--	g8818 = NOR(g8443, g8421, I15102)
--	g3885 = NOR(g3310, g3466)
--	g6174 = NOR(g1855, g5305)
--	g3233 = NOR(g1714, g1459)
--	g8811 = NOR(g8443, g8421, I15075)
--	g8629 = NOR(g6270, g8009)
--	g8279 = NOR(g7658, g7616, g8082, g7634)
--	g3504 = NOR(g1375, g2229, g2213, g2206)
--	g8625 = NOR(g1000, g6573, g1860, g8009)
--	g8232 = NOR(g8199, I14479, I14480)
--	g8659 = NOR(g8199, I14771, I14772)
--	g6209 = NOR(g2332, g5305)
--	g8630 = NOR(g6110, g7784, g3591, g1864)
--	g6184 = NOR(g875, g5291)
--	g8655 = NOR(g8199, I14753, I14754)
--	g5772 = NOR(g5428, g1888)
--	g2521 = NOR(g65, g62)
--	g7324 = NOR(g7189, g6994)
--	g5023 = NOR(g3894, g3889, g3886, g4359)
--	g8360 = NOR(g7658, g7616, g8082, g7634)
--	g8641 = NOR(g6559, g162, g7784, g3591)
--	g3505 = NOR(g2263, g1395)
--	g8658 = NOR(g8199, I14766, I14767)
--	g8680 = NOR(g8493, g8239, I14834)
--	g4894 = NOR(g4298, g4575, g4563)
--	g7314 = NOR(g7180, g6972)
--	g8092 = NOR(g7634, g7628, g7616, g7611)
--	g7322 = NOR(g7188, g6991)
--	g8523 = NOR(g7658, g7616, g8082, g7634)
--	g7312 = NOR(g7178, g6970)
--	g6452 = NOR(g6270, g2245)
--	g2014 = NOR(g1421, g1416)
--	g8862 = NOR(g8493, g8239, I15172)
--	g6185 = NOR(g5305, g1590)
--	g8679 = NOR(g8493, g8239, I14831)
--	g5039 = NOR(g3924, g3914, g3906, g3899)
--	g8805 = NOR(g8443, g8421, I15033)
--	g7152 = NOR(g6253, g7083, g5418)
--	g6664 = NOR(g5836, g1901, g1788)
--	g1980 = NOR(g1430, g1431)
--	g8233 = NOR(g8199, I14484, I14485)
--	g8706 = NOR(g7658, g8613, g7634)
--	g6910 = NOR(g1011, g1837, g6559, g1008)
--	g8707 = NOR(g7658, g8613, g7634)
--	g7328 = NOR(g7196, g7001)
--	g3516 = NOR(g2282, g1401)
--	g6197 = NOR(g875, g866, g1590, g5291)
--	g8635 = NOR(g1034, g8128)
--	g8801 = NOR(g8635, g3790)
--	g3310 = NOR(g936, g2557)
--	g7318 = NOR(g7185, g6979)
--	g7321 = NOR(g7187, g6990)
--	g3237 = NOR(g1444, g1838, g1454)
--	g8861 = NOR(g8493, g8239, I15169)
--	g4354 = NOR(g1424, g3541)
--	g8803 = NOR(g8443, g8421, I15021)
--	g4676 = NOR(g3885, g3094)
--	g8847 = NOR(g8493, g8239, I15147)
--	g4349 = NOR(g2496, g3310)
--	g3225 = NOR(g1021, g1025, g1889)
--	g7566 = NOR(g7421, g1597)
--	g8863 = NOR(g8493, g8239, I15175)
--	g1964 = NOR(g1428, g1429)
--	g7209 = NOR(g1789, g146, g6984)
--	g5614 = NOR(g3002, g1590, g4714)
--	g4318 = NOR(g3681, g1590)
--	g6214 = NOR(g878, g5284)
--	g4232 = NOR(g1934, g3591)
--	g6489 = NOR(g5802, g5769, g5790)
--	g3790 = NOR(g985, g990, g2295)
--	g5056 = NOR(g3556, g2872, g3938)
--	g8850 = NOR(g8493, g8239, I15152)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s13207 is
	port (
		CLK: in std_logic;
		G1: in std_logic;
		G9: in std_logic;
		G10: in std_logic;
		G11: in std_logic;
		G21: in std_logic;
		G22: in std_logic;
		G23: in std_logic;
		G24: in std_logic;
		G25: in std_logic;
		G26: in std_logic;
		G27: in std_logic;
		G28: in std_logic;
		G29: in std_logic;
		G30: in std_logic;
		G31: in std_logic;
		G32: in std_logic;
		G37: in std_logic;
		G41: in std_logic;
		G42: in std_logic;
		G43: in std_logic;
		G44: in std_logic;
		G45: in std_logic;
		G49: in std_logic;
		G633: in std_logic;
		G634: in std_logic;
		G635: in std_logic;
		G645: in std_logic;
		G647: in std_logic;
		G648: in std_logic;
		G690: in std_logic;
		G694: in std_logic;
		G698: in std_logic;
		G702: in std_logic;
		G722: in std_logic;
		G723: in std_logic;
		G751: in std_logic;
		G752: in std_logic;
		G753: in std_logic;
		G754: in std_logic;
		G755: in std_logic;
		G756: in std_logic;
		G757: in std_logic;
		G781: in std_logic;
		G786: in std_logic;
		G795: in std_logic;
		G929: in std_logic;
		G941: in std_logic;
		G955: in std_logic;
		G962: in std_logic;
		G1000: in std_logic;
		G1008: in std_logic;
		G1016: in std_logic;
		G1080: in std_logic;
		G1194: in std_logic;
		G1196: in std_logic;
		G1198: in std_logic;
		G1202: in std_logic;
		G1203: in std_logic;
		G1206: in std_logic;
		G1234: in std_logic;
		G1553: in std_logic;
		G1554: in std_logic;
		G206: out std_logic;
		G291: out std_logic;
		G372: out std_logic;
		G453: out std_logic;
		G534: out std_logic;
		G594: out std_logic;
		G785: out std_logic;
		G1006: out std_logic;
		G1015: out std_logic;
		G1017: out std_logic;
		G1193: out std_logic;
		G1195: out std_logic;
		G1197: out std_logic;
		G1201: out std_logic;
		G1205: out std_logic;
		G1246: out std_logic;
		G1724: out std_logic;
		G1783: out std_logic;
		G1798: out std_logic;
		G1804: out std_logic;
		G1810: out std_logic;
		G1817: out std_logic;
		G1824: out std_logic;
		G1829: out std_logic;
		G1870: out std_logic;
		G1871: out std_logic;
		G1894: out std_logic;
		G1911: out std_logic;
		G1944: out std_logic;
		G2662: out std_logic;
		G2844: out std_logic;
		G2888: out std_logic;
		G3077: out std_logic;
		G3096: out std_logic;
		G3130: out std_logic;
		G3159: out std_logic;
		G3191: out std_logic;
		G3829: out std_logic;
		G3854: out std_logic;
		G3856: out std_logic;
		G3857: out std_logic;
		G3859: out std_logic;
		G3860: out std_logic;
		G4267: out std_logic;
		G4316: out std_logic;
		G4370: out std_logic;
		G4371: out std_logic;
		G4372: out std_logic;
		G4373: out std_logic;
		G4655: out std_logic;
		G4657: out std_logic;
		G4660: out std_logic;
		G4661: out std_logic;
		G4663: out std_logic;
		G4664: out std_logic;
		G5143: out std_logic;
		G5164: out std_logic;
		G5571: out std_logic;
		G5669: out std_logic;
		G5678: out std_logic;
		G5682: out std_logic;
		G5684: out std_logic;
		G5687: out std_logic;
		G5729: out std_logic;
		G6207: out std_logic;
		G6212: out std_logic;
		G6223: out std_logic;
		G6236: out std_logic;
		G6269: out std_logic;
		G6288: out std_logic;
		G6289: out std_logic;
		G6290: out std_logic;
		G6291: out std_logic;
		G6292: out std_logic;
		G6293: out std_logic;
		G6294: out std_logic;
		G6295: out std_logic;
		G6296: out std_logic;
		G6297: out std_logic;
		G6298: out std_logic;
		G6299: out std_logic;
		G6300: out std_logic;
		G6301: out std_logic;
		G6302: out std_logic;
		G6303: out std_logic;
		G6304: out std_logic;
		G6305: out std_logic;
		G6306: out std_logic;
		G6307: out std_logic;
		G6308: out std_logic;
		G6376: out std_logic;
		G6425: out std_logic;
		G6648: out std_logic;
		G6653: out std_logic;
		G6675: out std_logic;
		G6849: out std_logic;
		G6850: out std_logic;
		G6895: out std_logic;
		G6909: out std_logic;
		G7048: out std_logic;
		G7063: out std_logic;
		G7103: out std_logic;
		G7283: out std_logic;
		G7284: out std_logic;
		G7285: out std_logic;
		G7286: out std_logic;
		G7287: out std_logic;
		G7288: out std_logic;
		G7289: out std_logic;
		G7290: out std_logic;
		G7291: out std_logic;
		G7292: out std_logic;
		G7293: out std_logic;
		G7294: out std_logic;
		G7295: out std_logic;
		G7298: out std_logic;
		G7423: out std_logic;
		G7424: out std_logic;
		G7425: out std_logic;
		G7474: out std_logic;
		G7504: out std_logic;
		G7505: out std_logic;
		G7506: out std_logic;
		G7507: out std_logic;
		G7508: out std_logic;
		G7514: out std_logic;
		G7729: out std_logic;
		G7730: out std_logic;
		G7731: out std_logic;
		G7732: out std_logic;
		G7763: out std_logic;
		G8216: out std_logic;
		G8217: out std_logic;
		G8218: out std_logic;
		G8219: out std_logic;
		G8234: out std_logic;
		G8661: out std_logic;
		G8663: out std_logic;
		G8872: out std_logic;
		G8958: out std_logic;
		G9128: out std_logic;
		G9132: out std_logic;
		G9204: out std_logic;
		G9280: out std_logic;
		G9297: out std_logic;
		G9299: out std_logic;
		G9305: out std_logic;
		G9308: out std_logic;
		G9310: out std_logic;
		G9312: out std_logic;
		G9314: out std_logic;
		G9378: out std_logic
	);
end entity;

architecture RTL of s13207 is
	attribute dont_touch: boolean;

	signal G2: std_logic; attribute dont_touch of G2: signal is true;
	signal G3: std_logic; attribute dont_touch of G3: signal is true;
	signal G4: std_logic; attribute dont_touch of G4: signal is true;
	signal G5: std_logic; attribute dont_touch of G5: signal is true;
	signal G6: std_logic; attribute dont_touch of G6: signal is true;
	signal G7: std_logic; attribute dont_touch of G7: signal is true;
	signal G8: std_logic; attribute dont_touch of G8: signal is true;
	signal G12: std_logic; attribute dont_touch of G12: signal is true;
	signal G13: std_logic; attribute dont_touch of G13: signal is true;
	signal G16: std_logic; attribute dont_touch of G16: signal is true;
	signal G20: std_logic; attribute dont_touch of G20: signal is true;
	signal G33: std_logic; attribute dont_touch of G33: signal is true;
	signal G38: std_logic; attribute dont_touch of G38: signal is true;
	signal G46: std_logic; attribute dont_touch of G46: signal is true;
	signal G47: std_logic; attribute dont_touch of G47: signal is true;
	signal G48: std_logic; attribute dont_touch of G48: signal is true;
	signal G52: std_logic; attribute dont_touch of G52: signal is true;
	signal G55: std_logic; attribute dont_touch of G55: signal is true;
	signal G58: std_logic; attribute dont_touch of G58: signal is true;
	signal G62: std_logic; attribute dont_touch of G62: signal is true;
	signal G65: std_logic; attribute dont_touch of G65: signal is true;
	signal G68: std_logic; attribute dont_touch of G68: signal is true;
	signal G71: std_logic; attribute dont_touch of G71: signal is true;
	signal G74: std_logic; attribute dont_touch of G74: signal is true;
	signal G77: std_logic; attribute dont_touch of G77: signal is true;
	signal G80: std_logic; attribute dont_touch of G80: signal is true;
	signal G83: std_logic; attribute dont_touch of G83: signal is true;
	signal G86: std_logic; attribute dont_touch of G86: signal is true;
	signal G89: std_logic; attribute dont_touch of G89: signal is true;
	signal G92: std_logic; attribute dont_touch of G92: signal is true;
	signal G93: std_logic; attribute dont_touch of G93: signal is true;
	signal G94: std_logic; attribute dont_touch of G94: signal is true;
	signal G95: std_logic; attribute dont_touch of G95: signal is true;
	signal G98: std_logic; attribute dont_touch of G98: signal is true;
	signal G99: std_logic; attribute dont_touch of G99: signal is true;
	signal G100: std_logic; attribute dont_touch of G100: signal is true;
	signal G103: std_logic; attribute dont_touch of G103: signal is true;
	signal G104: std_logic; attribute dont_touch of G104: signal is true;
	signal G105: std_logic; attribute dont_touch of G105: signal is true;
	signal G108: std_logic; attribute dont_touch of G108: signal is true;
	signal G109: std_logic; attribute dont_touch of G109: signal is true;
	signal G110: std_logic; attribute dont_touch of G110: signal is true;
	signal G113: std_logic; attribute dont_touch of G113: signal is true;
	signal G114: std_logic; attribute dont_touch of G114: signal is true;
	signal G117: std_logic; attribute dont_touch of G117: signal is true;
	signal G118: std_logic; attribute dont_touch of G118: signal is true;
	signal G121: std_logic; attribute dont_touch of G121: signal is true;
	signal G122: std_logic; attribute dont_touch of G122: signal is true;
	signal G125: std_logic; attribute dont_touch of G125: signal is true;
	signal G126: std_logic; attribute dont_touch of G126: signal is true;
	signal G129: std_logic; attribute dont_touch of G129: signal is true;
	signal G130: std_logic; attribute dont_touch of G130: signal is true;
	signal G133: std_logic; attribute dont_touch of G133: signal is true;
	signal G134: std_logic; attribute dont_touch of G134: signal is true;
	signal G137: std_logic; attribute dont_touch of G137: signal is true;
	signal G138: std_logic; attribute dont_touch of G138: signal is true;
	signal G141: std_logic; attribute dont_touch of G141: signal is true;
	signal G142: std_logic; attribute dont_touch of G142: signal is true;
	signal G145: std_logic; attribute dont_touch of G145: signal is true;
	signal G146: std_logic; attribute dont_touch of G146: signal is true;
	signal G150: std_logic; attribute dont_touch of G150: signal is true;
	signal G154: std_logic; attribute dont_touch of G154: signal is true;
	signal G158: std_logic; attribute dont_touch of G158: signal is true;
	signal G162: std_logic; attribute dont_touch of G162: signal is true;
	signal G168: std_logic; attribute dont_touch of G168: signal is true;
	signal G172: std_logic; attribute dont_touch of G172: signal is true;
	signal G173: std_logic; attribute dont_touch of G173: signal is true;
	signal G174: std_logic; attribute dont_touch of G174: signal is true;
	signal G179: std_logic; attribute dont_touch of G179: signal is true;
	signal G180: std_logic; attribute dont_touch of G180: signal is true;
	signal G181: std_logic; attribute dont_touch of G181: signal is true;
	signal G182: std_logic; attribute dont_touch of G182: signal is true;
	signal G183: std_logic; attribute dont_touch of G183: signal is true;
	signal G184: std_logic; attribute dont_touch of G184: signal is true;
	signal G185: std_logic; attribute dont_touch of G185: signal is true;
	signal G186: std_logic; attribute dont_touch of G186: signal is true;
	signal G187: std_logic; attribute dont_touch of G187: signal is true;
	signal G190: std_logic; attribute dont_touch of G190: signal is true;
	signal G195: std_logic; attribute dont_touch of G195: signal is true;
	signal G196: std_logic; attribute dont_touch of G196: signal is true;
	signal G199: std_logic; attribute dont_touch of G199: signal is true;
	signal G200: std_logic; attribute dont_touch of G200: signal is true;
	signal G201: std_logic; attribute dont_touch of G201: signal is true;
	signal G202: std_logic; attribute dont_touch of G202: signal is true;
	signal G205: std_logic; attribute dont_touch of G205: signal is true;
	signal G207: std_logic; attribute dont_touch of G207: signal is true;
	signal G210: std_logic; attribute dont_touch of G210: signal is true;
	signal G211: std_logic; attribute dont_touch of G211: signal is true;
	signal G212: std_logic; attribute dont_touch of G212: signal is true;
	signal G213: std_logic; attribute dont_touch of G213: signal is true;
	signal G214: std_logic; attribute dont_touch of G214: signal is true;
	signal G215: std_logic; attribute dont_touch of G215: signal is true;
	signal G216: std_logic; attribute dont_touch of G216: signal is true;
	signal G219: std_logic; attribute dont_touch of G219: signal is true;
	signal G222: std_logic; attribute dont_touch of G222: signal is true;
	signal G225: std_logic; attribute dont_touch of G225: signal is true;
	signal G228: std_logic; attribute dont_touch of G228: signal is true;
	signal G231: std_logic; attribute dont_touch of G231: signal is true;
	signal G232: std_logic; attribute dont_touch of G232: signal is true;
	signal G233: std_logic; attribute dont_touch of G233: signal is true;
	signal G234: std_logic; attribute dont_touch of G234: signal is true;
	signal G235: std_logic; attribute dont_touch of G235: signal is true;
	signal G236: std_logic; attribute dont_touch of G236: signal is true;
	signal G237: std_logic; attribute dont_touch of G237: signal is true;
	signal G240: std_logic; attribute dont_touch of G240: signal is true;
	signal G243: std_logic; attribute dont_touch of G243: signal is true;
	signal G246: std_logic; attribute dont_touch of G246: signal is true;
	signal G249: std_logic; attribute dont_touch of G249: signal is true;
	signal G252: std_logic; attribute dont_touch of G252: signal is true;
	signal G255: std_logic; attribute dont_touch of G255: signal is true;
	signal G258: std_logic; attribute dont_touch of G258: signal is true;
	signal G261: std_logic; attribute dont_touch of G261: signal is true;
	signal G264: std_logic; attribute dont_touch of G264: signal is true;
	signal G267: std_logic; attribute dont_touch of G267: signal is true;
	signal G270: std_logic; attribute dont_touch of G270: signal is true;
	signal G273: std_logic; attribute dont_touch of G273: signal is true;
	signal G274: std_logic; attribute dont_touch of G274: signal is true;
	signal G275: std_logic; attribute dont_touch of G275: signal is true;
	signal G278: std_logic; attribute dont_touch of G278: signal is true;
	signal G281: std_logic; attribute dont_touch of G281: signal is true;
	signal G284: std_logic; attribute dont_touch of G284: signal is true;
	signal G287: std_logic; attribute dont_touch of G287: signal is true;
	signal G290: std_logic; attribute dont_touch of G290: signal is true;
	signal G292: std_logic; attribute dont_touch of G292: signal is true;
	signal G293: std_logic; attribute dont_touch of G293: signal is true;
	signal G294: std_logic; attribute dont_touch of G294: signal is true;
	signal G295: std_logic; attribute dont_touch of G295: signal is true;
	signal G296: std_logic; attribute dont_touch of G296: signal is true;
	signal G297: std_logic; attribute dont_touch of G297: signal is true;
	signal G300: std_logic; attribute dont_touch of G300: signal is true;
	signal G303: std_logic; attribute dont_touch of G303: signal is true;
	signal G306: std_logic; attribute dont_touch of G306: signal is true;
	signal G309: std_logic; attribute dont_touch of G309: signal is true;
	signal G312: std_logic; attribute dont_touch of G312: signal is true;
	signal G313: std_logic; attribute dont_touch of G313: signal is true;
	signal G314: std_logic; attribute dont_touch of G314: signal is true;
	signal G315: std_logic; attribute dont_touch of G315: signal is true;
	signal G316: std_logic; attribute dont_touch of G316: signal is true;
	signal G317: std_logic; attribute dont_touch of G317: signal is true;
	signal G318: std_logic; attribute dont_touch of G318: signal is true;
	signal G321: std_logic; attribute dont_touch of G321: signal is true;
	signal G324: std_logic; attribute dont_touch of G324: signal is true;
	signal G327: std_logic; attribute dont_touch of G327: signal is true;
	signal G330: std_logic; attribute dont_touch of G330: signal is true;
	signal G333: std_logic; attribute dont_touch of G333: signal is true;
	signal G336: std_logic; attribute dont_touch of G336: signal is true;
	signal G339: std_logic; attribute dont_touch of G339: signal is true;
	signal G342: std_logic; attribute dont_touch of G342: signal is true;
	signal G345: std_logic; attribute dont_touch of G345: signal is true;
	signal G348: std_logic; attribute dont_touch of G348: signal is true;
	signal G351: std_logic; attribute dont_touch of G351: signal is true;
	signal G354: std_logic; attribute dont_touch of G354: signal is true;
	signal G355: std_logic; attribute dont_touch of G355: signal is true;
	signal G356: std_logic; attribute dont_touch of G356: signal is true;
	signal G359: std_logic; attribute dont_touch of G359: signal is true;
	signal G362: std_logic; attribute dont_touch of G362: signal is true;
	signal G365: std_logic; attribute dont_touch of G365: signal is true;
	signal G368: std_logic; attribute dont_touch of G368: signal is true;
	signal G371: std_logic; attribute dont_touch of G371: signal is true;
	signal G373: std_logic; attribute dont_touch of G373: signal is true;
	signal G374: std_logic; attribute dont_touch of G374: signal is true;
	signal G375: std_logic; attribute dont_touch of G375: signal is true;
	signal G376: std_logic; attribute dont_touch of G376: signal is true;
	signal G377: std_logic; attribute dont_touch of G377: signal is true;
	signal G378: std_logic; attribute dont_touch of G378: signal is true;
	signal G381: std_logic; attribute dont_touch of G381: signal is true;
	signal G384: std_logic; attribute dont_touch of G384: signal is true;
	signal G387: std_logic; attribute dont_touch of G387: signal is true;
	signal G390: std_logic; attribute dont_touch of G390: signal is true;
	signal G393: std_logic; attribute dont_touch of G393: signal is true;
	signal G394: std_logic; attribute dont_touch of G394: signal is true;
	signal G395: std_logic; attribute dont_touch of G395: signal is true;
	signal G396: std_logic; attribute dont_touch of G396: signal is true;
	signal G397: std_logic; attribute dont_touch of G397: signal is true;
	signal G398: std_logic; attribute dont_touch of G398: signal is true;
	signal G399: std_logic; attribute dont_touch of G399: signal is true;
	signal G402: std_logic; attribute dont_touch of G402: signal is true;
	signal G405: std_logic; attribute dont_touch of G405: signal is true;
	signal G408: std_logic; attribute dont_touch of G408: signal is true;
	signal G411: std_logic; attribute dont_touch of G411: signal is true;
	signal G414: std_logic; attribute dont_touch of G414: signal is true;
	signal G417: std_logic; attribute dont_touch of G417: signal is true;
	signal G420: std_logic; attribute dont_touch of G420: signal is true;
	signal G423: std_logic; attribute dont_touch of G423: signal is true;
	signal G426: std_logic; attribute dont_touch of G426: signal is true;
	signal G429: std_logic; attribute dont_touch of G429: signal is true;
	signal G432: std_logic; attribute dont_touch of G432: signal is true;
	signal G435: std_logic; attribute dont_touch of G435: signal is true;
	signal G436: std_logic; attribute dont_touch of G436: signal is true;
	signal G437: std_logic; attribute dont_touch of G437: signal is true;
	signal G440: std_logic; attribute dont_touch of G440: signal is true;
	signal G443: std_logic; attribute dont_touch of G443: signal is true;
	signal G446: std_logic; attribute dont_touch of G446: signal is true;
	signal G449: std_logic; attribute dont_touch of G449: signal is true;
	signal G452: std_logic; attribute dont_touch of G452: signal is true;
	signal G454: std_logic; attribute dont_touch of G454: signal is true;
	signal G455: std_logic; attribute dont_touch of G455: signal is true;
	signal G456: std_logic; attribute dont_touch of G456: signal is true;
	signal G457: std_logic; attribute dont_touch of G457: signal is true;
	signal G458: std_logic; attribute dont_touch of G458: signal is true;
	signal G459: std_logic; attribute dont_touch of G459: signal is true;
	signal G462: std_logic; attribute dont_touch of G462: signal is true;
	signal G465: std_logic; attribute dont_touch of G465: signal is true;
	signal G468: std_logic; attribute dont_touch of G468: signal is true;
	signal G471: std_logic; attribute dont_touch of G471: signal is true;
	signal G474: std_logic; attribute dont_touch of G474: signal is true;
	signal G475: std_logic; attribute dont_touch of G475: signal is true;
	signal G476: std_logic; attribute dont_touch of G476: signal is true;
	signal G477: std_logic; attribute dont_touch of G477: signal is true;
	signal G478: std_logic; attribute dont_touch of G478: signal is true;
	signal G479: std_logic; attribute dont_touch of G479: signal is true;
	signal G480: std_logic; attribute dont_touch of G480: signal is true;
	signal G483: std_logic; attribute dont_touch of G483: signal is true;
	signal G486: std_logic; attribute dont_touch of G486: signal is true;
	signal G489: std_logic; attribute dont_touch of G489: signal is true;
	signal G492: std_logic; attribute dont_touch of G492: signal is true;
	signal G495: std_logic; attribute dont_touch of G495: signal is true;
	signal G498: std_logic; attribute dont_touch of G498: signal is true;
	signal G501: std_logic; attribute dont_touch of G501: signal is true;
	signal G504: std_logic; attribute dont_touch of G504: signal is true;
	signal G507: std_logic; attribute dont_touch of G507: signal is true;
	signal G510: std_logic; attribute dont_touch of G510: signal is true;
	signal G513: std_logic; attribute dont_touch of G513: signal is true;
	signal G516: std_logic; attribute dont_touch of G516: signal is true;
	signal G517: std_logic; attribute dont_touch of G517: signal is true;
	signal G518: std_logic; attribute dont_touch of G518: signal is true;
	signal G521: std_logic; attribute dont_touch of G521: signal is true;
	signal G524: std_logic; attribute dont_touch of G524: signal is true;
	signal G527: std_logic; attribute dont_touch of G527: signal is true;
	signal G530: std_logic; attribute dont_touch of G530: signal is true;
	signal G533: std_logic; attribute dont_touch of G533: signal is true;
	signal G535: std_logic; attribute dont_touch of G535: signal is true;
	signal G536: std_logic; attribute dont_touch of G536: signal is true;
	signal G539: std_logic; attribute dont_touch of G539: signal is true;
	signal G540: std_logic; attribute dont_touch of G540: signal is true;
	signal G543: std_logic; attribute dont_touch of G543: signal is true;
	signal G544: std_logic; attribute dont_touch of G544: signal is true;
	signal G547: std_logic; attribute dont_touch of G547: signal is true;
	signal G550: std_logic; attribute dont_touch of G550: signal is true;
	signal G553: std_logic; attribute dont_touch of G553: signal is true;
	signal G556: std_logic; attribute dont_touch of G556: signal is true;
	signal G557: std_logic; attribute dont_touch of G557: signal is true;
	signal G560: std_logic; attribute dont_touch of G560: signal is true;
	signal G563: std_logic; attribute dont_touch of G563: signal is true;
	signal G566: std_logic; attribute dont_touch of G566: signal is true;
	signal G567: std_logic; attribute dont_touch of G567: signal is true;
	signal G570: std_logic; attribute dont_touch of G570: signal is true;
	signal G573: std_logic; attribute dont_touch of G573: signal is true;
	signal G576: std_logic; attribute dont_touch of G576: signal is true;
	signal G579: std_logic; attribute dont_touch of G579: signal is true;
	signal G580: std_logic; attribute dont_touch of G580: signal is true;
	signal G583: std_logic; attribute dont_touch of G583: signal is true;
	signal G584: std_logic; attribute dont_touch of G584: signal is true;
	signal G587: std_logic; attribute dont_touch of G587: signal is true;
	signal G588: std_logic; attribute dont_touch of G588: signal is true;
	signal G591: std_logic; attribute dont_touch of G591: signal is true;
	signal G595: std_logic; attribute dont_touch of G595: signal is true;
	signal G596: std_logic; attribute dont_touch of G596: signal is true;
	signal G597: std_logic; attribute dont_touch of G597: signal is true;
	signal G598: std_logic; attribute dont_touch of G598: signal is true;
	signal G599: std_logic; attribute dont_touch of G599: signal is true;
	signal G600: std_logic; attribute dont_touch of G600: signal is true;
	signal G601: std_logic; attribute dont_touch of G601: signal is true;
	signal G602: std_logic; attribute dont_touch of G602: signal is true;
	signal G603: std_logic; attribute dont_touch of G603: signal is true;
	signal G604: std_logic; attribute dont_touch of G604: signal is true;
	signal G605: std_logic; attribute dont_touch of G605: signal is true;
	signal G606: std_logic; attribute dont_touch of G606: signal is true;
	signal G607: std_logic; attribute dont_touch of G607: signal is true;
	signal G608: std_logic; attribute dont_touch of G608: signal is true;
	signal G609: std_logic; attribute dont_touch of G609: signal is true;
	signal G610: std_logic; attribute dont_touch of G610: signal is true;
	signal G611: std_logic; attribute dont_touch of G611: signal is true;
	signal G612: std_logic; attribute dont_touch of G612: signal is true;
	signal G613: std_logic; attribute dont_touch of G613: signal is true;
	signal G614: std_logic; attribute dont_touch of G614: signal is true;
	signal G615: std_logic; attribute dont_touch of G615: signal is true;
	signal G616: std_logic; attribute dont_touch of G616: signal is true;
	signal G617: std_logic; attribute dont_touch of G617: signal is true;
	signal G618: std_logic; attribute dont_touch of G618: signal is true;
	signal G619: std_logic; attribute dont_touch of G619: signal is true;
	signal G620: std_logic; attribute dont_touch of G620: signal is true;
	signal G621: std_logic; attribute dont_touch of G621: signal is true;
	signal G622: std_logic; attribute dont_touch of G622: signal is true;
	signal G623: std_logic; attribute dont_touch of G623: signal is true;
	signal G624: std_logic; attribute dont_touch of G624: signal is true;
	signal G625: std_logic; attribute dont_touch of G625: signal is true;
	signal G626: std_logic; attribute dont_touch of G626: signal is true;
	signal G627: std_logic; attribute dont_touch of G627: signal is true;
	signal G628: std_logic; attribute dont_touch of G628: signal is true;
	signal G629: std_logic; attribute dont_touch of G629: signal is true;
	signal G630: std_logic; attribute dont_touch of G630: signal is true;
	signal G631: std_logic; attribute dont_touch of G631: signal is true;
	signal G632: std_logic; attribute dont_touch of G632: signal is true;
	signal G636: std_logic; attribute dont_touch of G636: signal is true;
	signal G639: std_logic; attribute dont_touch of G639: signal is true;
	signal G642: std_logic; attribute dont_touch of G642: signal is true;
	signal G646: std_logic; attribute dont_touch of G646: signal is true;
	signal G649: std_logic; attribute dont_touch of G649: signal is true;
	signal G652: std_logic; attribute dont_touch of G652: signal is true;
	signal G655: std_logic; attribute dont_touch of G655: signal is true;
	signal G658: std_logic; attribute dont_touch of G658: signal is true;
	signal G661: std_logic; attribute dont_touch of G661: signal is true;
	signal G665: std_logic; attribute dont_touch of G665: signal is true;
	signal G669: std_logic; attribute dont_touch of G669: signal is true;
	signal G673: std_logic; attribute dont_touch of G673: signal is true;
	signal G677: std_logic; attribute dont_touch of G677: signal is true;
	signal G681: std_logic; attribute dont_touch of G681: signal is true;
	signal G685: std_logic; attribute dont_touch of G685: signal is true;
	signal G689: std_logic; attribute dont_touch of G689: signal is true;
	signal G691: std_logic; attribute dont_touch of G691: signal is true;
	signal G695: std_logic; attribute dont_touch of G695: signal is true;
	signal G699: std_logic; attribute dont_touch of G699: signal is true;
	signal G703: std_logic; attribute dont_touch of G703: signal is true;
	signal G706: std_logic; attribute dont_touch of G706: signal is true;
	signal G710: std_logic; attribute dont_touch of G710: signal is true;
	signal G714: std_logic; attribute dont_touch of G714: signal is true;
	signal G718: std_logic; attribute dont_touch of G718: signal is true;
	signal G724: std_logic; attribute dont_touch of G724: signal is true;
	signal G727: std_logic; attribute dont_touch of G727: signal is true;
	signal G730: std_logic; attribute dont_touch of G730: signal is true;
	signal G734: std_logic; attribute dont_touch of G734: signal is true;
	signal G738: std_logic; attribute dont_touch of G738: signal is true;
	signal G741: std_logic; attribute dont_touch of G741: signal is true;
	signal G746: std_logic; attribute dont_touch of G746: signal is true;
	signal G758: std_logic; attribute dont_touch of G758: signal is true;
	signal G759: std_logic; attribute dont_touch of G759: signal is true;
	signal G760: std_logic; attribute dont_touch of G760: signal is true;
	signal G761: std_logic; attribute dont_touch of G761: signal is true;
	signal G762: std_logic; attribute dont_touch of G762: signal is true;
	signal G763: std_logic; attribute dont_touch of G763: signal is true;
	signal G764: std_logic; attribute dont_touch of G764: signal is true;
	signal G765: std_logic; attribute dont_touch of G765: signal is true;
	signal G766: std_logic; attribute dont_touch of G766: signal is true;
	signal G767: std_logic; attribute dont_touch of G767: signal is true;
	signal G768: std_logic; attribute dont_touch of G768: signal is true;
	signal G769: std_logic; attribute dont_touch of G769: signal is true;
	signal G770: std_logic; attribute dont_touch of G770: signal is true;
	signal G771: std_logic; attribute dont_touch of G771: signal is true;
	signal G772: std_logic; attribute dont_touch of G772: signal is true;
	signal G773: std_logic; attribute dont_touch of G773: signal is true;
	signal G774: std_logic; attribute dont_touch of G774: signal is true;
	signal G775: std_logic; attribute dont_touch of G775: signal is true;
	signal G778: std_logic; attribute dont_touch of G778: signal is true;
	signal G782: std_logic; attribute dont_touch of G782: signal is true;
	signal G789: std_logic; attribute dont_touch of G789: signal is true;
	signal G792: std_logic; attribute dont_touch of G792: signal is true;
	signal G799: std_logic; attribute dont_touch of G799: signal is true;
	signal G803: std_logic; attribute dont_touch of G803: signal is true;
	signal G806: std_logic; attribute dont_touch of G806: signal is true;
	signal G809: std_logic; attribute dont_touch of G809: signal is true;
	signal G812: std_logic; attribute dont_touch of G812: signal is true;
	signal G815: std_logic; attribute dont_touch of G815: signal is true;
	signal G819: std_logic; attribute dont_touch of G819: signal is true;
	signal G822: std_logic; attribute dont_touch of G822: signal is true;
	signal G825: std_logic; attribute dont_touch of G825: signal is true;
	signal G828: std_logic; attribute dont_touch of G828: signal is true;
	signal G831: std_logic; attribute dont_touch of G831: signal is true;
	signal G834: std_logic; attribute dont_touch of G834: signal is true;
	signal G837: std_logic; attribute dont_touch of G837: signal is true;
	signal G840: std_logic; attribute dont_touch of G840: signal is true;
	signal G843: std_logic; attribute dont_touch of G843: signal is true;
	signal G846: std_logic; attribute dont_touch of G846: signal is true;
	signal G849: std_logic; attribute dont_touch of G849: signal is true;
	signal G852: std_logic; attribute dont_touch of G852: signal is true;
	signal G855: std_logic; attribute dont_touch of G855: signal is true;
	signal G859: std_logic; attribute dont_touch of G859: signal is true;
	signal G863: std_logic; attribute dont_touch of G863: signal is true;
	signal G866: std_logic; attribute dont_touch of G866: signal is true;
	signal G871: std_logic; attribute dont_touch of G871: signal is true;
	signal G874: std_logic; attribute dont_touch of G874: signal is true;
	signal G875: std_logic; attribute dont_touch of G875: signal is true;
	signal G878: std_logic; attribute dont_touch of G878: signal is true;
	signal G883: std_logic; attribute dont_touch of G883: signal is true;
	signal G887: std_logic; attribute dont_touch of G887: signal is true;
	signal G888: std_logic; attribute dont_touch of G888: signal is true;
	signal G889: std_logic; attribute dont_touch of G889: signal is true;
	signal G890: std_logic; attribute dont_touch of G890: signal is true;
	signal G891: std_logic; attribute dont_touch of G891: signal is true;
	signal G896: std_logic; attribute dont_touch of G896: signal is true;
	signal G901: std_logic; attribute dont_touch of G901: signal is true;
	signal G906: std_logic; attribute dont_touch of G906: signal is true;
	signal G911: std_logic; attribute dont_touch of G911: signal is true;
	signal G916: std_logic; attribute dont_touch of G916: signal is true;
	signal G921: std_logic; attribute dont_touch of G921: signal is true;
	signal G926: std_logic; attribute dont_touch of G926: signal is true;
	signal G933: std_logic; attribute dont_touch of G933: signal is true;
	signal G936: std_logic; attribute dont_touch of G936: signal is true;
	signal G940: std_logic; attribute dont_touch of G940: signal is true;
	signal G942: std_logic; attribute dont_touch of G942: signal is true;
	signal G943: std_logic; attribute dont_touch of G943: signal is true;
	signal G944: std_logic; attribute dont_touch of G944: signal is true;
	signal G945: std_logic; attribute dont_touch of G945: signal is true;
	signal G948: std_logic; attribute dont_touch of G948: signal is true;
	signal G949: std_logic; attribute dont_touch of G949: signal is true;
	signal G950: std_logic; attribute dont_touch of G950: signal is true;
	signal G951: std_logic; attribute dont_touch of G951: signal is true;
	signal G952: std_logic; attribute dont_touch of G952: signal is true;
	signal G953: std_logic; attribute dont_touch of G953: signal is true;
	signal G954: std_logic; attribute dont_touch of G954: signal is true;
	signal G959: std_logic; attribute dont_touch of G959: signal is true;
	signal G963: std_logic; attribute dont_touch of G963: signal is true;
	signal G966: std_logic; attribute dont_touch of G966: signal is true;
	signal G969: std_logic; attribute dont_touch of G969: signal is true;
	signal G970: std_logic; attribute dont_touch of G970: signal is true;
	signal G971: std_logic; attribute dont_touch of G971: signal is true;
	signal G972: std_logic; attribute dont_touch of G972: signal is true;
	signal G973: std_logic; attribute dont_touch of G973: signal is true;
	signal G976: std_logic; attribute dont_touch of G976: signal is true;
	signal G979: std_logic; attribute dont_touch of G979: signal is true;
	signal G984: std_logic; attribute dont_touch of G984: signal is true;
	signal G985: std_logic; attribute dont_touch of G985: signal is true;
	signal G990: std_logic; attribute dont_touch of G990: signal is true;
	signal G995: std_logic; attribute dont_touch of G995: signal is true;
	signal G998: std_logic; attribute dont_touch of G998: signal is true;
	signal G999: std_logic; attribute dont_touch of G999: signal is true;
	signal G1004: std_logic; attribute dont_touch of G1004: signal is true;
	signal G1005: std_logic; attribute dont_touch of G1005: signal is true;
	signal G1007: std_logic; attribute dont_touch of G1007: signal is true;
	signal G1011: std_logic; attribute dont_touch of G1011: signal is true;
	signal G1012: std_logic; attribute dont_touch of G1012: signal is true;
	signal G1013: std_logic; attribute dont_touch of G1013: signal is true;
	signal G1014: std_logic; attribute dont_touch of G1014: signal is true;
	signal G1018: std_logic; attribute dont_touch of G1018: signal is true;
	signal G1021: std_logic; attribute dont_touch of G1021: signal is true;
	signal G1025: std_logic; attribute dont_touch of G1025: signal is true;
	signal G1029: std_logic; attribute dont_touch of G1029: signal is true;
	signal G1030: std_logic; attribute dont_touch of G1030: signal is true;
	signal G1033: std_logic; attribute dont_touch of G1033: signal is true;
	signal G1034: std_logic; attribute dont_touch of G1034: signal is true;
	signal G1037: std_logic; attribute dont_touch of G1037: signal is true;
	signal G1041: std_logic; attribute dont_touch of G1041: signal is true;
	signal G1045: std_logic; attribute dont_touch of G1045: signal is true;
	signal G1049: std_logic; attribute dont_touch of G1049: signal is true;
	signal G1053: std_logic; attribute dont_touch of G1053: signal is true;
	signal G1057: std_logic; attribute dont_touch of G1057: signal is true;
	signal G1061: std_logic; attribute dont_touch of G1061: signal is true;
	signal G1065: std_logic; attribute dont_touch of G1065: signal is true;
	signal G1069: std_logic; attribute dont_touch of G1069: signal is true;
	signal G1073: std_logic; attribute dont_touch of G1073: signal is true;
	signal G1077: std_logic; attribute dont_touch of G1077: signal is true;
	signal G1081: std_logic; attribute dont_touch of G1081: signal is true;
	signal G1084: std_logic; attribute dont_touch of G1084: signal is true;
	signal G1087: std_logic; attribute dont_touch of G1087: signal is true;
	signal G1092: std_logic; attribute dont_touch of G1092: signal is true;
	signal G1097: std_logic; attribute dont_touch of G1097: signal is true;
	signal G1098: std_logic; attribute dont_touch of G1098: signal is true;
	signal G1102: std_logic; attribute dont_touch of G1102: signal is true;
	signal G1106: std_logic; attribute dont_touch of G1106: signal is true;
	signal G1110: std_logic; attribute dont_touch of G1110: signal is true;
	signal G1114: std_logic; attribute dont_touch of G1114: signal is true;
	signal G1118: std_logic; attribute dont_touch of G1118: signal is true;
	signal G1122: std_logic; attribute dont_touch of G1122: signal is true;
	signal G1126: std_logic; attribute dont_touch of G1126: signal is true;
	signal G1130: std_logic; attribute dont_touch of G1130: signal is true;
	signal G1134: std_logic; attribute dont_touch of G1134: signal is true;
	signal G1138: std_logic; attribute dont_touch of G1138: signal is true;
	signal G1142: std_logic; attribute dont_touch of G1142: signal is true;
	signal G1146: std_logic; attribute dont_touch of G1146: signal is true;
	signal G1147: std_logic; attribute dont_touch of G1147: signal is true;
	signal G1148: std_logic; attribute dont_touch of G1148: signal is true;
	signal G1149: std_logic; attribute dont_touch of G1149: signal is true;
	signal G1153: std_logic; attribute dont_touch of G1153: signal is true;
	signal G1154: std_logic; attribute dont_touch of G1154: signal is true;
	signal G1155: std_logic; attribute dont_touch of G1155: signal is true;
	signal G1156: std_logic; attribute dont_touch of G1156: signal is true;
	signal G1157: std_logic; attribute dont_touch of G1157: signal is true;
	signal G1158: std_logic; attribute dont_touch of G1158: signal is true;
	signal G1159: std_logic; attribute dont_touch of G1159: signal is true;
	signal G1160: std_logic; attribute dont_touch of G1160: signal is true;
	signal G1163: std_logic; attribute dont_touch of G1163: signal is true;
	signal G1166: std_logic; attribute dont_touch of G1166: signal is true;
	signal G1167: std_logic; attribute dont_touch of G1167: signal is true;
	signal G1170: std_logic; attribute dont_touch of G1170: signal is true;
	signal G1173: std_logic; attribute dont_touch of G1173: signal is true;
	signal G1176: std_logic; attribute dont_touch of G1176: signal is true;
	signal G1179: std_logic; attribute dont_touch of G1179: signal is true;
	signal G1182: std_logic; attribute dont_touch of G1182: signal is true;
	signal G1185: std_logic; attribute dont_touch of G1185: signal is true;
	signal G1186: std_logic; attribute dont_touch of G1186: signal is true;
	signal G1189: std_logic; attribute dont_touch of G1189: signal is true;
	signal G1190: std_logic; attribute dont_touch of G1190: signal is true;
	signal G1191: std_logic; attribute dont_touch of G1191: signal is true;
	signal G1192: std_logic; attribute dont_touch of G1192: signal is true;
	signal G1199: std_logic; attribute dont_touch of G1199: signal is true;
	signal G1200: std_logic; attribute dont_touch of G1200: signal is true;
	signal G1204: std_logic; attribute dont_touch of G1204: signal is true;
	signal G1207: std_logic; attribute dont_touch of G1207: signal is true;
	signal G1211: std_logic; attribute dont_touch of G1211: signal is true;
	signal G1214: std_logic; attribute dont_touch of G1214: signal is true;
	signal G1217: std_logic; attribute dont_touch of G1217: signal is true;
	signal G1220: std_logic; attribute dont_touch of G1220: signal is true;
	signal G1223: std_logic; attribute dont_touch of G1223: signal is true;
	signal G1224: std_logic; attribute dont_touch of G1224: signal is true;
	signal G1225: std_logic; attribute dont_touch of G1225: signal is true;
	signal G1226: std_logic; attribute dont_touch of G1226: signal is true;
	signal G1227: std_logic; attribute dont_touch of G1227: signal is true;
	signal G1228: std_logic; attribute dont_touch of G1228: signal is true;
	signal G1229: std_logic; attribute dont_touch of G1229: signal is true;
	signal G1230: std_logic; attribute dont_touch of G1230: signal is true;
	signal G1231: std_logic; attribute dont_touch of G1231: signal is true;
	signal G1235: std_logic; attribute dont_touch of G1235: signal is true;
	signal G1236: std_logic; attribute dont_touch of G1236: signal is true;
	signal G1240: std_logic; attribute dont_touch of G1240: signal is true;
	signal G1243: std_logic; attribute dont_touch of G1243: signal is true;
	signal G1244: std_logic; attribute dont_touch of G1244: signal is true;
	signal G1245: std_logic; attribute dont_touch of G1245: signal is true;
	signal G1247: std_logic; attribute dont_touch of G1247: signal is true;
	signal G1250: std_logic; attribute dont_touch of G1250: signal is true;
	signal G1251: std_logic; attribute dont_touch of G1251: signal is true;
	signal G1252: std_logic; attribute dont_touch of G1252: signal is true;
	signal G1253: std_logic; attribute dont_touch of G1253: signal is true;
	signal G1254: std_logic; attribute dont_touch of G1254: signal is true;
	signal G1257: std_logic; attribute dont_touch of G1257: signal is true;
	signal G1260: std_logic; attribute dont_touch of G1260: signal is true;
	signal G1263: std_logic; attribute dont_touch of G1263: signal is true;
	signal G1266: std_logic; attribute dont_touch of G1266: signal is true;
	signal G1267: std_logic; attribute dont_touch of G1267: signal is true;
	signal G1268: std_logic; attribute dont_touch of G1268: signal is true;
	signal G1269: std_logic; attribute dont_touch of G1269: signal is true;
	signal G1270: std_logic; attribute dont_touch of G1270: signal is true;
	signal G1271: std_logic; attribute dont_touch of G1271: signal is true;
	signal G1272: std_logic; attribute dont_touch of G1272: signal is true;
	signal G1276: std_logic; attribute dont_touch of G1276: signal is true;
	signal G1280: std_logic; attribute dont_touch of G1280: signal is true;
	signal G1284: std_logic; attribute dont_touch of G1284: signal is true;
	signal G1288: std_logic; attribute dont_touch of G1288: signal is true;
	signal G1292: std_logic; attribute dont_touch of G1292: signal is true;
	signal G1296: std_logic; attribute dont_touch of G1296: signal is true;
	signal G1300: std_logic; attribute dont_touch of G1300: signal is true;
	signal G1304: std_logic; attribute dont_touch of G1304: signal is true;
	signal G1307: std_logic; attribute dont_touch of G1307: signal is true;
	signal G1308: std_logic; attribute dont_touch of G1308: signal is true;
	signal G1309: std_logic; attribute dont_touch of G1309: signal is true;
	signal G1310: std_logic; attribute dont_touch of G1310: signal is true;
	signal G1311: std_logic; attribute dont_touch of G1311: signal is true;
	signal G1312: std_logic; attribute dont_touch of G1312: signal is true;
	signal G1313: std_logic; attribute dont_touch of G1313: signal is true;
	signal G1317: std_logic; attribute dont_touch of G1317: signal is true;
	signal G1318: std_logic; attribute dont_touch of G1318: signal is true;
	signal G1319: std_logic; attribute dont_touch of G1319: signal is true;
	signal G1320: std_logic; attribute dont_touch of G1320: signal is true;
	signal G1321: std_logic; attribute dont_touch of G1321: signal is true;
	signal G1322: std_logic; attribute dont_touch of G1322: signal is true;
	signal G1323: std_logic; attribute dont_touch of G1323: signal is true;
	signal G1324: std_logic; attribute dont_touch of G1324: signal is true;
	signal G1325: std_logic; attribute dont_touch of G1325: signal is true;
	signal G1326: std_logic; attribute dont_touch of G1326: signal is true;
	signal G1327: std_logic; attribute dont_touch of G1327: signal is true;
	signal G1328: std_logic; attribute dont_touch of G1328: signal is true;
	signal G1329: std_logic; attribute dont_touch of G1329: signal is true;
	signal G1330: std_logic; attribute dont_touch of G1330: signal is true;
	signal G1333: std_logic; attribute dont_touch of G1333: signal is true;
	signal G1336: std_logic; attribute dont_touch of G1336: signal is true;
	signal G1339: std_logic; attribute dont_touch of G1339: signal is true;
	signal G1342: std_logic; attribute dont_touch of G1342: signal is true;
	signal G1345: std_logic; attribute dont_touch of G1345: signal is true;
	signal G1348: std_logic; attribute dont_touch of G1348: signal is true;
	signal G1351: std_logic; attribute dont_touch of G1351: signal is true;
	signal G1354: std_logic; attribute dont_touch of G1354: signal is true;
	signal G1357: std_logic; attribute dont_touch of G1357: signal is true;
	signal G1360: std_logic; attribute dont_touch of G1360: signal is true;
	signal G1363: std_logic; attribute dont_touch of G1363: signal is true;
	signal G1364: std_logic; attribute dont_touch of G1364: signal is true;
	signal G1365: std_logic; attribute dont_touch of G1365: signal is true;
	signal G1366: std_logic; attribute dont_touch of G1366: signal is true;
	signal G1367: std_logic; attribute dont_touch of G1367: signal is true;
	signal G1368: std_logic; attribute dont_touch of G1368: signal is true;
	signal G1369: std_logic; attribute dont_touch of G1369: signal is true;
	signal G1370: std_logic; attribute dont_touch of G1370: signal is true;
	signal G1371: std_logic; attribute dont_touch of G1371: signal is true;
	signal G1372: std_logic; attribute dont_touch of G1372: signal is true;
	signal G1373: std_logic; attribute dont_touch of G1373: signal is true;
	signal G1374: std_logic; attribute dont_touch of G1374: signal is true;
	signal G1375: std_logic; attribute dont_touch of G1375: signal is true;
	signal G1376: std_logic; attribute dont_touch of G1376: signal is true;
	signal G1377: std_logic; attribute dont_touch of G1377: signal is true;
	signal G1378: std_logic; attribute dont_touch of G1378: signal is true;
	signal G1379: std_logic; attribute dont_touch of G1379: signal is true;
	signal G1380: std_logic; attribute dont_touch of G1380: signal is true;
	signal G1381: std_logic; attribute dont_touch of G1381: signal is true;
	signal G1382: std_logic; attribute dont_touch of G1382: signal is true;
	signal G1383: std_logic; attribute dont_touch of G1383: signal is true;
	signal G1384: std_logic; attribute dont_touch of G1384: signal is true;
	signal G1385: std_logic; attribute dont_touch of G1385: signal is true;
	signal G1386: std_logic; attribute dont_touch of G1386: signal is true;
	signal G1387: std_logic; attribute dont_touch of G1387: signal is true;
	signal G1388: std_logic; attribute dont_touch of G1388: signal is true;
	signal G1389: std_logic; attribute dont_touch of G1389: signal is true;
	signal G1390: std_logic; attribute dont_touch of G1390: signal is true;
	signal G1391: std_logic; attribute dont_touch of G1391: signal is true;
	signal G1392: std_logic; attribute dont_touch of G1392: signal is true;
	signal G1393: std_logic; attribute dont_touch of G1393: signal is true;
	signal G1394: std_logic; attribute dont_touch of G1394: signal is true;
	signal G1395: std_logic; attribute dont_touch of G1395: signal is true;
	signal G1396: std_logic; attribute dont_touch of G1396: signal is true;
	signal G1397: std_logic; attribute dont_touch of G1397: signal is true;
	signal G1398: std_logic; attribute dont_touch of G1398: signal is true;
	signal G1399: std_logic; attribute dont_touch of G1399: signal is true;
	signal G1400: std_logic; attribute dont_touch of G1400: signal is true;
	signal G1401: std_logic; attribute dont_touch of G1401: signal is true;
	signal G1402: std_logic; attribute dont_touch of G1402: signal is true;
	signal G1403: std_logic; attribute dont_touch of G1403: signal is true;
	signal G1404: std_logic; attribute dont_touch of G1404: signal is true;
	signal G1405: std_logic; attribute dont_touch of G1405: signal is true;
	signal G1408: std_logic; attribute dont_touch of G1408: signal is true;
	signal G1409: std_logic; attribute dont_touch of G1409: signal is true;
	signal G1412: std_logic; attribute dont_touch of G1412: signal is true;
	signal G1415: std_logic; attribute dont_touch of G1415: signal is true;
	signal G1416: std_logic; attribute dont_touch of G1416: signal is true;
	signal G1421: std_logic; attribute dont_touch of G1421: signal is true;
	signal G1424: std_logic; attribute dont_touch of G1424: signal is true;
	signal G1428: std_logic; attribute dont_touch of G1428: signal is true;
	signal G1429: std_logic; attribute dont_touch of G1429: signal is true;
	signal G1430: std_logic; attribute dont_touch of G1430: signal is true;
	signal G1431: std_logic; attribute dont_touch of G1431: signal is true;
	signal G1432: std_logic; attribute dont_touch of G1432: signal is true;
	signal G1435: std_logic; attribute dont_touch of G1435: signal is true;
	signal G1439: std_logic; attribute dont_touch of G1439: signal is true;
	signal G1443: std_logic; attribute dont_touch of G1443: signal is true;
	signal G1444: std_logic; attribute dont_touch of G1444: signal is true;
	signal G1450: std_logic; attribute dont_touch of G1450: signal is true;
	signal G1454: std_logic; attribute dont_touch of G1454: signal is true;
	signal G1459: std_logic; attribute dont_touch of G1459: signal is true;
	signal G1460: std_logic; attribute dont_touch of G1460: signal is true;
	signal G1461: std_logic; attribute dont_touch of G1461: signal is true;
	signal G1462: std_logic; attribute dont_touch of G1462: signal is true;
	signal G1467: std_logic; attribute dont_touch of G1467: signal is true;
	signal G1472: std_logic; attribute dont_touch of G1472: signal is true;
	signal G1477: std_logic; attribute dont_touch of G1477: signal is true;
	signal G1481: std_logic; attribute dont_touch of G1481: signal is true;
	signal G1486: std_logic; attribute dont_touch of G1486: signal is true;
	signal G1489: std_logic; attribute dont_touch of G1489: signal is true;
	signal G1494: std_logic; attribute dont_touch of G1494: signal is true;
	signal G1499: std_logic; attribute dont_touch of G1499: signal is true;
	signal G1504: std_logic; attribute dont_touch of G1504: signal is true;
	signal G1509: std_logic; attribute dont_touch of G1509: signal is true;
	signal G1513: std_logic; attribute dont_touch of G1513: signal is true;
	signal G1514: std_logic; attribute dont_touch of G1514: signal is true;
	signal G1519: std_logic; attribute dont_touch of G1519: signal is true;
	signal G1524: std_logic; attribute dont_touch of G1524: signal is true;
	signal G1528: std_logic; attribute dont_touch of G1528: signal is true;
	signal G1532: std_logic; attribute dont_touch of G1532: signal is true;
	signal G1537: std_logic; attribute dont_touch of G1537: signal is true;
	signal G1541: std_logic; attribute dont_touch of G1541: signal is true;
	signal G1545: std_logic; attribute dont_touch of G1545: signal is true;
	signal G1549: std_logic; attribute dont_touch of G1549: signal is true;
	signal G1555: std_logic; attribute dont_touch of G1555: signal is true;
	signal G1556: std_logic; attribute dont_touch of G1556: signal is true;
	signal G1557: std_logic; attribute dont_touch of G1557: signal is true;
	signal G1558: std_logic; attribute dont_touch of G1558: signal is true;
	signal G1562: std_logic; attribute dont_touch of G1562: signal is true;
	signal G1563: std_logic; attribute dont_touch of G1563: signal is true;
	signal G1564: std_logic; attribute dont_touch of G1564: signal is true;
	signal G1565: std_logic; attribute dont_touch of G1565: signal is true;
	signal G1566: std_logic; attribute dont_touch of G1566: signal is true;
	signal G1567: std_logic; attribute dont_touch of G1567: signal is true;
	signal G1568: std_logic; attribute dont_touch of G1568: signal is true;
	signal G1569: std_logic; attribute dont_touch of G1569: signal is true;
	signal G1570: std_logic; attribute dont_touch of G1570: signal is true;
	signal G1571: std_logic; attribute dont_touch of G1571: signal is true;
	signal G1572: std_logic; attribute dont_touch of G1572: signal is true;
	signal G1573: std_logic; attribute dont_touch of G1573: signal is true;
	signal G1574: std_logic; attribute dont_touch of G1574: signal is true;
	signal G1575: std_logic; attribute dont_touch of G1575: signal is true;
	signal G1576: std_logic; attribute dont_touch of G1576: signal is true;
	signal G1577: std_logic; attribute dont_touch of G1577: signal is true;
	signal G1578: std_logic; attribute dont_touch of G1578: signal is true;
	signal G1579: std_logic; attribute dont_touch of G1579: signal is true;
	signal G1580: std_logic; attribute dont_touch of G1580: signal is true;
	signal G1581: std_logic; attribute dont_touch of G1581: signal is true;
	signal G1582: std_logic; attribute dont_touch of G1582: signal is true;
	signal G1583: std_logic; attribute dont_touch of G1583: signal is true;
	signal G1584: std_logic; attribute dont_touch of G1584: signal is true;
	signal G1585: std_logic; attribute dont_touch of G1585: signal is true;
	signal G1586: std_logic; attribute dont_touch of G1586: signal is true;
	signal G1587: std_logic; attribute dont_touch of G1587: signal is true;
	signal G1588: std_logic; attribute dont_touch of G1588: signal is true;
	signal G1589: std_logic; attribute dont_touch of G1589: signal is true;
	signal G1590: std_logic; attribute dont_touch of G1590: signal is true;
	signal G1597: std_logic; attribute dont_touch of G1597: signal is true;
	signal G1600: std_logic; attribute dont_touch of G1600: signal is true;
	signal G1603: std_logic; attribute dont_touch of G1603: signal is true;
	signal G1611: std_logic; attribute dont_touch of G1611: signal is true;
	signal G1612: std_logic; attribute dont_touch of G1612: signal is true;
	signal G1616: std_logic; attribute dont_touch of G1616: signal is true;
	signal G1637: std_logic; attribute dont_touch of G1637: signal is true;
	signal G1638: std_logic; attribute dont_touch of G1638: signal is true;
	signal G1639: std_logic; attribute dont_touch of G1639: signal is true;
	signal G1643: std_logic; attribute dont_touch of G1643: signal is true;
	signal G1646: std_logic; attribute dont_touch of G1646: signal is true;
	signal G1649: std_logic; attribute dont_touch of G1649: signal is true;
	signal G1652: std_logic; attribute dont_touch of G1652: signal is true;
	signal G1655: std_logic; attribute dont_touch of G1655: signal is true;
	signal G1658: std_logic; attribute dont_touch of G1658: signal is true;
	signal G1661: std_logic; attribute dont_touch of G1661: signal is true;
	signal G1662: std_logic; attribute dont_touch of G1662: signal is true;
	signal G1663: std_logic; attribute dont_touch of G1663: signal is true;
	signal G1664: std_logic; attribute dont_touch of G1664: signal is true;
	signal G1665: std_logic; attribute dont_touch of G1665: signal is true;
	signal G1666: std_logic; attribute dont_touch of G1666: signal is true;
	signal G1667: std_logic; attribute dont_touch of G1667: signal is true;
	signal G1670: std_logic; attribute dont_touch of G1670: signal is true;
	signal G1671: std_logic; attribute dont_touch of G1671: signal is true;
	signal G1672: std_logic; attribute dont_touch of G1672: signal is true;
	signal G1673: std_logic; attribute dont_touch of G1673: signal is true;
	signal G1674: std_logic; attribute dont_touch of G1674: signal is true;
	signal G1675: std_logic; attribute dont_touch of G1675: signal is true;
	signal G1676: std_logic; attribute dont_touch of G1676: signal is true;
	signal G1677: std_logic; attribute dont_touch of G1677: signal is true;
	signal G1678: std_logic; attribute dont_touch of G1678: signal is true;
	signal G1679: std_logic; attribute dont_touch of G1679: signal is true;
	signal G1680: std_logic; attribute dont_touch of G1680: signal is true;
	signal G1681: std_logic; attribute dont_touch of G1681: signal is true;
	signal G1682: std_logic; attribute dont_touch of G1682: signal is true;
	signal G1683: std_logic; attribute dont_touch of G1683: signal is true;
	signal G1684: std_logic; attribute dont_touch of G1684: signal is true;
	signal G1685: std_logic; attribute dont_touch of G1685: signal is true;
	signal G1686: std_logic; attribute dont_touch of G1686: signal is true;
	signal G1687: std_logic; attribute dont_touch of G1687: signal is true;
	signal G1688: std_logic; attribute dont_touch of G1688: signal is true;
	signal G1689: std_logic; attribute dont_touch of G1689: signal is true;
	signal G1690: std_logic; attribute dont_touch of G1690: signal is true;
	signal G1694: std_logic; attribute dont_touch of G1694: signal is true;
	signal G1695: std_logic; attribute dont_touch of G1695: signal is true;
	signal G1698: std_logic; attribute dont_touch of G1698: signal is true;
	signal G1701: std_logic; attribute dont_touch of G1701: signal is true;
	signal G1704: std_logic; attribute dont_touch of G1704: signal is true;
	signal G1707: std_logic; attribute dont_touch of G1707: signal is true;
	signal G1708: std_logic; attribute dont_touch of G1708: signal is true;
	signal G1711: std_logic; attribute dont_touch of G1711: signal is true;
	signal G1714: std_logic; attribute dont_touch of G1714: signal is true;
	signal G1715: std_logic; attribute dont_touch of G1715: signal is true;
	signal G1718: std_logic; attribute dont_touch of G1718: signal is true;
	signal G1721: std_logic; attribute dont_touch of G1721: signal is true;
	signal G1725: std_logic; attribute dont_touch of G1725: signal is true;
	signal G1726: std_logic; attribute dont_touch of G1726: signal is true;
	signal G1727: std_logic; attribute dont_touch of G1727: signal is true;
	signal G1728: std_logic; attribute dont_touch of G1728: signal is true;
	signal G1732: std_logic; attribute dont_touch of G1732: signal is true;
	signal G1733: std_logic; attribute dont_touch of G1733: signal is true;
	signal G1736: std_logic; attribute dont_touch of G1736: signal is true;
	signal G1737: std_logic; attribute dont_touch of G1737: signal is true;
	signal G1738: std_logic; attribute dont_touch of G1738: signal is true;
	signal G1739: std_logic; attribute dont_touch of G1739: signal is true;
	signal G1742: std_logic; attribute dont_touch of G1742: signal is true;
	signal G1743: std_logic; attribute dont_touch of G1743: signal is true;
	signal G1744: std_logic; attribute dont_touch of G1744: signal is true;
	signal G1745: std_logic; attribute dont_touch of G1745: signal is true;
	signal G1746: std_logic; attribute dont_touch of G1746: signal is true;
	signal G1747: std_logic; attribute dont_touch of G1747: signal is true;
	signal G1748: std_logic; attribute dont_touch of G1748: signal is true;
	signal G1749: std_logic; attribute dont_touch of G1749: signal is true;
	signal G1750: std_logic; attribute dont_touch of G1750: signal is true;
	signal G1751: std_logic; attribute dont_touch of G1751: signal is true;
	signal G1752: std_logic; attribute dont_touch of G1752: signal is true;
	signal G1753: std_logic; attribute dont_touch of G1753: signal is true;
	signal G1756: std_logic; attribute dont_touch of G1756: signal is true;
	signal G1757: std_logic; attribute dont_touch of G1757: signal is true;
	signal G1758: std_logic; attribute dont_touch of G1758: signal is true;
	signal G1759: std_logic; attribute dont_touch of G1759: signal is true;
	signal G1760: std_logic; attribute dont_touch of G1760: signal is true;
	signal G1768: std_logic; attribute dont_touch of G1768: signal is true;
	signal G1769: std_logic; attribute dont_touch of G1769: signal is true;
	signal G1770: std_logic; attribute dont_touch of G1770: signal is true;
	signal G1771: std_logic; attribute dont_touch of G1771: signal is true;
	signal G1772: std_logic; attribute dont_touch of G1772: signal is true;
	signal G1773: std_logic; attribute dont_touch of G1773: signal is true;
	signal G1774: std_logic; attribute dont_touch of G1774: signal is true;
	signal G1775: std_logic; attribute dont_touch of G1775: signal is true;
	signal G1776: std_logic; attribute dont_touch of G1776: signal is true;
	signal G1777: std_logic; attribute dont_touch of G1777: signal is true;
	signal G1778: std_logic; attribute dont_touch of G1778: signal is true;
	signal G1779: std_logic; attribute dont_touch of G1779: signal is true;
	signal G1780: std_logic; attribute dont_touch of G1780: signal is true;
	signal G1781: std_logic; attribute dont_touch of G1781: signal is true;
	signal G1782: std_logic; attribute dont_touch of G1782: signal is true;
	signal G1784: std_logic; attribute dont_touch of G1784: signal is true;
	signal G1785: std_logic; attribute dont_touch of G1785: signal is true;
	signal G1786: std_logic; attribute dont_touch of G1786: signal is true;
	signal G1787: std_logic; attribute dont_touch of G1787: signal is true;
	signal G1788: std_logic; attribute dont_touch of G1788: signal is true;
	signal G1789: std_logic; attribute dont_touch of G1789: signal is true;
	signal G1792: std_logic; attribute dont_touch of G1792: signal is true;
	signal G1793: std_logic; attribute dont_touch of G1793: signal is true;
	signal G1794: std_logic; attribute dont_touch of G1794: signal is true;
	signal G1795: std_logic; attribute dont_touch of G1795: signal is true;
	signal G1796: std_logic; attribute dont_touch of G1796: signal is true;
	signal G1797: std_logic; attribute dont_touch of G1797: signal is true;
	signal G1799: std_logic; attribute dont_touch of G1799: signal is true;
	signal G1800: std_logic; attribute dont_touch of G1800: signal is true;
	signal G1801: std_logic; attribute dont_touch of G1801: signal is true;
	signal G1802: std_logic; attribute dont_touch of G1802: signal is true;
	signal G1803: std_logic; attribute dont_touch of G1803: signal is true;
	signal G1805: std_logic; attribute dont_touch of G1805: signal is true;
	signal G1806: std_logic; attribute dont_touch of G1806: signal is true;
	signal G1807: std_logic; attribute dont_touch of G1807: signal is true;
	signal G1808: std_logic; attribute dont_touch of G1808: signal is true;
	signal G1809: std_logic; attribute dont_touch of G1809: signal is true;
	signal G1811: std_logic; attribute dont_touch of G1811: signal is true;
	signal G1812: std_logic; attribute dont_touch of G1812: signal is true;
	signal G1813: std_logic; attribute dont_touch of G1813: signal is true;
	signal G1814: std_logic; attribute dont_touch of G1814: signal is true;
	signal G1815: std_logic; attribute dont_touch of G1815: signal is true;
	signal G1816: std_logic; attribute dont_touch of G1816: signal is true;
	signal G1818: std_logic; attribute dont_touch of G1818: signal is true;
	signal G1819: std_logic; attribute dont_touch of G1819: signal is true;
	signal G1820: std_logic; attribute dont_touch of G1820: signal is true;
	signal G1821: std_logic; attribute dont_touch of G1821: signal is true;
	signal G1822: std_logic; attribute dont_touch of G1822: signal is true;
	signal G1823: std_logic; attribute dont_touch of G1823: signal is true;
	signal G1825: std_logic; attribute dont_touch of G1825: signal is true;
	signal G1826: std_logic; attribute dont_touch of G1826: signal is true;
	signal G1827: std_logic; attribute dont_touch of G1827: signal is true;
	signal G1828: std_logic; attribute dont_touch of G1828: signal is true;
	signal G1830: std_logic; attribute dont_touch of G1830: signal is true;
	signal G1831: std_logic; attribute dont_touch of G1831: signal is true;
	signal G1832: std_logic; attribute dont_touch of G1832: signal is true;
	signal G1833: std_logic; attribute dont_touch of G1833: signal is true;
	signal G1834: std_logic; attribute dont_touch of G1834: signal is true;
	signal G1837: std_logic; attribute dont_touch of G1837: signal is true;
	signal G1838: std_logic; attribute dont_touch of G1838: signal is true;
	signal G1842: std_logic; attribute dont_touch of G1842: signal is true;
	signal G1843: std_logic; attribute dont_touch of G1843: signal is true;
	signal G1844: std_logic; attribute dont_touch of G1844: signal is true;
	signal G1847: std_logic; attribute dont_touch of G1847: signal is true;
	signal G1848: std_logic; attribute dont_touch of G1848: signal is true;
	signal G1849: std_logic; attribute dont_touch of G1849: signal is true;
	signal G1852: std_logic; attribute dont_touch of G1852: signal is true;
	signal G1853: std_logic; attribute dont_touch of G1853: signal is true;
	signal G1854: std_logic; attribute dont_touch of G1854: signal is true;
	signal G1855: std_logic; attribute dont_touch of G1855: signal is true;
	signal G1856: std_logic; attribute dont_touch of G1856: signal is true;
	signal G1857: std_logic; attribute dont_touch of G1857: signal is true;
	signal G1860: std_logic; attribute dont_touch of G1860: signal is true;
	signal G1863: std_logic; attribute dont_touch of G1863: signal is true;
	signal G1864: std_logic; attribute dont_touch of G1864: signal is true;
	signal G1865: std_logic; attribute dont_touch of G1865: signal is true;
	signal G1866: std_logic; attribute dont_touch of G1866: signal is true;
	signal G1867: std_logic; attribute dont_touch of G1867: signal is true;
	signal G1868: std_logic; attribute dont_touch of G1868: signal is true;
	signal G1869: std_logic; attribute dont_touch of G1869: signal is true;
	signal G1872: std_logic; attribute dont_touch of G1872: signal is true;
	signal G1876: std_logic; attribute dont_touch of G1876: signal is true;
	signal G1877: std_logic; attribute dont_touch of G1877: signal is true;
	signal G1878: std_logic; attribute dont_touch of G1878: signal is true;
	signal G1879: std_logic; attribute dont_touch of G1879: signal is true;
	signal G1886: std_logic; attribute dont_touch of G1886: signal is true;
	signal G1887: std_logic; attribute dont_touch of G1887: signal is true;
	signal G1888: std_logic; attribute dont_touch of G1888: signal is true;
	signal G1889: std_logic; attribute dont_touch of G1889: signal is true;
	signal G1895: std_logic; attribute dont_touch of G1895: signal is true;
	signal G1896: std_logic; attribute dont_touch of G1896: signal is true;
	signal G1897: std_logic; attribute dont_touch of G1897: signal is true;
	signal G1898: std_logic; attribute dont_touch of G1898: signal is true;
	signal G1901: std_logic; attribute dont_touch of G1901: signal is true;
	signal G1904: std_logic; attribute dont_touch of G1904: signal is true;
	signal G1907: std_logic; attribute dont_touch of G1907: signal is true;
	signal G1908: std_logic; attribute dont_touch of G1908: signal is true;
	signal G1909: std_logic; attribute dont_touch of G1909: signal is true;
	signal G1910: std_logic; attribute dont_touch of G1910: signal is true;
	signal G1912: std_logic; attribute dont_touch of G1912: signal is true;
	signal G1913: std_logic; attribute dont_touch of G1913: signal is true;
	signal G1916: std_logic; attribute dont_touch of G1916: signal is true;
	signal G1917: std_logic; attribute dont_touch of G1917: signal is true;
	signal G1918: std_logic; attribute dont_touch of G1918: signal is true;
	signal G1919: std_logic; attribute dont_touch of G1919: signal is true;
	signal G1922: std_logic; attribute dont_touch of G1922: signal is true;
	signal G1923: std_logic; attribute dont_touch of G1923: signal is true;
	signal G1924: std_logic; attribute dont_touch of G1924: signal is true;
	signal G1925: std_logic; attribute dont_touch of G1925: signal is true;
	signal G1926: std_logic; attribute dont_touch of G1926: signal is true;
	signal G1929: std_logic; attribute dont_touch of G1929: signal is true;
	signal G1933: std_logic; attribute dont_touch of G1933: signal is true;
	signal G1934: std_logic; attribute dont_touch of G1934: signal is true;
	signal G1935: std_logic; attribute dont_touch of G1935: signal is true;
	signal G1938: std_logic; attribute dont_touch of G1938: signal is true;
	signal G1941: std_logic; attribute dont_touch of G1941: signal is true;
	signal G1942: std_logic; attribute dont_touch of G1942: signal is true;
	signal G1943: std_logic; attribute dont_touch of G1943: signal is true;
	signal G1945: std_logic; attribute dont_touch of G1945: signal is true;
	signal G1948: std_logic; attribute dont_touch of G1948: signal is true;
	signal G1949: std_logic; attribute dont_touch of G1949: signal is true;
	signal G1952: std_logic; attribute dont_touch of G1952: signal is true;
	signal G1955: std_logic; attribute dont_touch of G1955: signal is true;
	signal G1958: std_logic; attribute dont_touch of G1958: signal is true;
	signal G1959: std_logic; attribute dont_touch of G1959: signal is true;
	signal G1960: std_logic; attribute dont_touch of G1960: signal is true;
	signal G1961: std_logic; attribute dont_touch of G1961: signal is true;
	signal G1964: std_logic; attribute dont_touch of G1964: signal is true;
	signal G1967: std_logic; attribute dont_touch of G1967: signal is true;
	signal G1970: std_logic; attribute dont_touch of G1970: signal is true;
	signal G1974: std_logic; attribute dont_touch of G1974: signal is true;
	signal G1975: std_logic; attribute dont_touch of G1975: signal is true;
	signal G1976: std_logic; attribute dont_touch of G1976: signal is true;
	signal G1977: std_logic; attribute dont_touch of G1977: signal is true;
	signal G1980: std_logic; attribute dont_touch of G1980: signal is true;
	signal G1983: std_logic; attribute dont_touch of G1983: signal is true;
	signal G1987: std_logic; attribute dont_touch of G1987: signal is true;
	signal G2006: std_logic; attribute dont_touch of G2006: signal is true;
	signal G2007: std_logic; attribute dont_touch of G2007: signal is true;
	signal G2011: std_logic; attribute dont_touch of G2011: signal is true;
	signal G2014: std_logic; attribute dont_touch of G2014: signal is true;
	signal G2015: std_logic; attribute dont_touch of G2015: signal is true;
	signal G2016: std_logic; attribute dont_touch of G2016: signal is true;
	signal G2020: std_logic; attribute dont_touch of G2020: signal is true;
	signal G2038: std_logic; attribute dont_touch of G2038: signal is true;
	signal G2039: std_logic; attribute dont_touch of G2039: signal is true;
	signal G2043: std_logic; attribute dont_touch of G2043: signal is true;
	signal G2044: std_logic; attribute dont_touch of G2044: signal is true;
	signal G2051: std_logic; attribute dont_touch of G2051: signal is true;
	signal G2052: std_logic; attribute dont_touch of G2052: signal is true;
	signal G2057: std_logic; attribute dont_touch of G2057: signal is true;
	signal G2073: std_logic; attribute dont_touch of G2073: signal is true;
	signal G2074: std_logic; attribute dont_touch of G2074: signal is true;
	signal G2091: std_logic; attribute dont_touch of G2091: signal is true;
	signal G2092: std_logic; attribute dont_touch of G2092: signal is true;
	signal G2096: std_logic; attribute dont_touch of G2096: signal is true;
	signal G2100: std_logic; attribute dont_touch of G2100: signal is true;
	signal G2104: std_logic; attribute dont_touch of G2104: signal is true;
	signal G2105: std_logic; attribute dont_touch of G2105: signal is true;
	signal G2106: std_logic; attribute dont_touch of G2106: signal is true;
	signal G2128: std_logic; attribute dont_touch of G2128: signal is true;
	signal G2131: std_logic; attribute dont_touch of G2131: signal is true;
	signal G2134: std_logic; attribute dont_touch of G2134: signal is true;
	signal G2137: std_logic; attribute dont_touch of G2137: signal is true;
	signal G2145: std_logic; attribute dont_touch of G2145: signal is true;
	signal G2148: std_logic; attribute dont_touch of G2148: signal is true;
	signal G2149: std_logic; attribute dont_touch of G2149: signal is true;
	signal G2157: std_logic; attribute dont_touch of G2157: signal is true;
	signal G2161: std_logic; attribute dont_touch of G2161: signal is true;
	signal G2162: std_logic; attribute dont_touch of G2162: signal is true;
	signal G2170: std_logic; attribute dont_touch of G2170: signal is true;
	signal G2174: std_logic; attribute dont_touch of G2174: signal is true;
	signal G2177: std_logic; attribute dont_touch of G2177: signal is true;
	signal G2180: std_logic; attribute dont_touch of G2180: signal is true;
	signal G2183: std_logic; attribute dont_touch of G2183: signal is true;
	signal G2184: std_logic; attribute dont_touch of G2184: signal is true;
	signal G2185: std_logic; attribute dont_touch of G2185: signal is true;
	signal G2202: std_logic; attribute dont_touch of G2202: signal is true;
	signal G2205: std_logic; attribute dont_touch of G2205: signal is true;
	signal G2206: std_logic; attribute dont_touch of G2206: signal is true;
	signal G2207: std_logic; attribute dont_touch of G2207: signal is true;
	signal G2208: std_logic; attribute dont_touch of G2208: signal is true;
	signal G2209: std_logic; attribute dont_touch of G2209: signal is true;
	signal G2210: std_logic; attribute dont_touch of G2210: signal is true;
	signal G2213: std_logic; attribute dont_touch of G2213: signal is true;
	signal G2214: std_logic; attribute dont_touch of G2214: signal is true;
	signal G2215: std_logic; attribute dont_touch of G2215: signal is true;
	signal G2216: std_logic; attribute dont_touch of G2216: signal is true;
	signal G2221: std_logic; attribute dont_touch of G2221: signal is true;
	signal G2222: std_logic; attribute dont_touch of G2222: signal is true;
	signal G2223: std_logic; attribute dont_touch of G2223: signal is true;
	signal G2224: std_logic; attribute dont_touch of G2224: signal is true;
	signal G2225: std_logic; attribute dont_touch of G2225: signal is true;
	signal G2226: std_logic; attribute dont_touch of G2226: signal is true;
	signal G2229: std_logic; attribute dont_touch of G2229: signal is true;
	signal G2230: std_logic; attribute dont_touch of G2230: signal is true;
	signal G2231: std_logic; attribute dont_touch of G2231: signal is true;
	signal G2232: std_logic; attribute dont_touch of G2232: signal is true;
	signal G2233: std_logic; attribute dont_touch of G2233: signal is true;
	signal G2234: std_logic; attribute dont_touch of G2234: signal is true;
	signal G2235: std_logic; attribute dont_touch of G2235: signal is true;
	signal G2236: std_logic; attribute dont_touch of G2236: signal is true;
	signal G2237: std_logic; attribute dont_touch of G2237: signal is true;
	signal G2238: std_logic; attribute dont_touch of G2238: signal is true;
	signal G2239: std_logic; attribute dont_touch of G2239: signal is true;
	signal G2240: std_logic; attribute dont_touch of G2240: signal is true;
	signal G2241: std_logic; attribute dont_touch of G2241: signal is true;
	signal G2242: std_logic; attribute dont_touch of G2242: signal is true;
	signal G2245: std_logic; attribute dont_touch of G2245: signal is true;
	signal G2246: std_logic; attribute dont_touch of G2246: signal is true;
	signal G2253: std_logic; attribute dont_touch of G2253: signal is true;
	signal G2256: std_logic; attribute dont_touch of G2256: signal is true;
	signal G2259: std_logic; attribute dont_touch of G2259: signal is true;
	signal G2262: std_logic; attribute dont_touch of G2262: signal is true;
	signal G2263: std_logic; attribute dont_touch of G2263: signal is true;
	signal G2264: std_logic; attribute dont_touch of G2264: signal is true;
	signal G2265: std_logic; attribute dont_touch of G2265: signal is true;
	signal G2266: std_logic; attribute dont_touch of G2266: signal is true;
	signal G2267: std_logic; attribute dont_touch of G2267: signal is true;
	signal G2268: std_logic; attribute dont_touch of G2268: signal is true;
	signal G2269: std_logic; attribute dont_touch of G2269: signal is true;
	signal G2270: std_logic; attribute dont_touch of G2270: signal is true;
	signal G2271: std_logic; attribute dont_touch of G2271: signal is true;
	signal G2272: std_logic; attribute dont_touch of G2272: signal is true;
	signal G2273: std_logic; attribute dont_touch of G2273: signal is true;
	signal G2274: std_logic; attribute dont_touch of G2274: signal is true;
	signal G2275: std_logic; attribute dont_touch of G2275: signal is true;
	signal G2276: std_logic; attribute dont_touch of G2276: signal is true;
	signal G2282: std_logic; attribute dont_touch of G2282: signal is true;
	signal G2283: std_logic; attribute dont_touch of G2283: signal is true;
	signal G2284: std_logic; attribute dont_touch of G2284: signal is true;
	signal G2285: std_logic; attribute dont_touch of G2285: signal is true;
	signal G2286: std_logic; attribute dont_touch of G2286: signal is true;
	signal G2287: std_logic; attribute dont_touch of G2287: signal is true;
	signal G2288: std_logic; attribute dont_touch of G2288: signal is true;
	signal G2289: std_logic; attribute dont_touch of G2289: signal is true;
	signal G2290: std_logic; attribute dont_touch of G2290: signal is true;
	signal G2291: std_logic; attribute dont_touch of G2291: signal is true;
	signal G2292: std_logic; attribute dont_touch of G2292: signal is true;
	signal G2293: std_logic; attribute dont_touch of G2293: signal is true;
	signal G2294: std_logic; attribute dont_touch of G2294: signal is true;
	signal G2295: std_logic; attribute dont_touch of G2295: signal is true;
	signal G2298: std_logic; attribute dont_touch of G2298: signal is true;
	signal G2306: std_logic; attribute dont_touch of G2306: signal is true;
	signal G2307: std_logic; attribute dont_touch of G2307: signal is true;
	signal G2308: std_logic; attribute dont_touch of G2308: signal is true;
	signal G2309: std_logic; attribute dont_touch of G2309: signal is true;
	signal G2310: std_logic; attribute dont_touch of G2310: signal is true;
	signal G2311: std_logic; attribute dont_touch of G2311: signal is true;
	signal G2312: std_logic; attribute dont_touch of G2312: signal is true;
	signal G2313: std_logic; attribute dont_touch of G2313: signal is true;
	signal G2314: std_logic; attribute dont_touch of G2314: signal is true;
	signal G2315: std_logic; attribute dont_touch of G2315: signal is true;
	signal G2316: std_logic; attribute dont_touch of G2316: signal is true;
	signal G2323: std_logic; attribute dont_touch of G2323: signal is true;
	signal G2324: std_logic; attribute dont_touch of G2324: signal is true;
	signal G2325: std_logic; attribute dont_touch of G2325: signal is true;
	signal G2326: std_logic; attribute dont_touch of G2326: signal is true;
	signal G2327: std_logic; attribute dont_touch of G2327: signal is true;
	signal G2328: std_logic; attribute dont_touch of G2328: signal is true;
	signal G2329: std_logic; attribute dont_touch of G2329: signal is true;
	signal G2330: std_logic; attribute dont_touch of G2330: signal is true;
	signal G2331: std_logic; attribute dont_touch of G2331: signal is true;
	signal G2332: std_logic; attribute dont_touch of G2332: signal is true;
	signal G2333: std_logic; attribute dont_touch of G2333: signal is true;
	signal G2334: std_logic; attribute dont_touch of G2334: signal is true;
	signal G2340: std_logic; attribute dont_touch of G2340: signal is true;
	signal G2343: std_logic; attribute dont_touch of G2343: signal is true;
	signal G2344: std_logic; attribute dont_touch of G2344: signal is true;
	signal G2345: std_logic; attribute dont_touch of G2345: signal is true;
	signal G2346: std_logic; attribute dont_touch of G2346: signal is true;
	signal G2347: std_logic; attribute dont_touch of G2347: signal is true;
	signal G2348: std_logic; attribute dont_touch of G2348: signal is true;
	signal G2349: std_logic; attribute dont_touch of G2349: signal is true;
	signal G2350: std_logic; attribute dont_touch of G2350: signal is true;
	signal G2351: std_logic; attribute dont_touch of G2351: signal is true;
	signal G2352: std_logic; attribute dont_touch of G2352: signal is true;
	signal G2353: std_logic; attribute dont_touch of G2353: signal is true;
	signal G2354: std_logic; attribute dont_touch of G2354: signal is true;
	signal G2359: std_logic; attribute dont_touch of G2359: signal is true;
	signal G2360: std_logic; attribute dont_touch of G2360: signal is true;
	signal G2361: std_logic; attribute dont_touch of G2361: signal is true;
	signal G2362: std_logic; attribute dont_touch of G2362: signal is true;
	signal G2363: std_logic; attribute dont_touch of G2363: signal is true;
	signal G2364: std_logic; attribute dont_touch of G2364: signal is true;
	signal G2365: std_logic; attribute dont_touch of G2365: signal is true;
	signal G2366: std_logic; attribute dont_touch of G2366: signal is true;
	signal G2367: std_logic; attribute dont_touch of G2367: signal is true;
	signal G2368: std_logic; attribute dont_touch of G2368: signal is true;
	signal G2371: std_logic; attribute dont_touch of G2371: signal is true;
	signal G2372: std_logic; attribute dont_touch of G2372: signal is true;
	signal G2373: std_logic; attribute dont_touch of G2373: signal is true;
	signal G2374: std_logic; attribute dont_touch of G2374: signal is true;
	signal G2375: std_logic; attribute dont_touch of G2375: signal is true;
	signal G2376: std_logic; attribute dont_touch of G2376: signal is true;
	signal G2377: std_logic; attribute dont_touch of G2377: signal is true;
	signal G2378: std_logic; attribute dont_touch of G2378: signal is true;
	signal G2379: std_logic; attribute dont_touch of G2379: signal is true;
	signal G2380: std_logic; attribute dont_touch of G2380: signal is true;
	signal G2381: std_logic; attribute dont_touch of G2381: signal is true;
	signal G2382: std_logic; attribute dont_touch of G2382: signal is true;
	signal G2383: std_logic; attribute dont_touch of G2383: signal is true;
	signal G2384: std_logic; attribute dont_touch of G2384: signal is true;
	signal G2385: std_logic; attribute dont_touch of G2385: signal is true;
	signal G2386: std_logic; attribute dont_touch of G2386: signal is true;
	signal G2389: std_logic; attribute dont_touch of G2389: signal is true;
	signal G2392: std_logic; attribute dont_touch of G2392: signal is true;
	signal G2393: std_logic; attribute dont_touch of G2393: signal is true;
	signal G2394: std_logic; attribute dont_touch of G2394: signal is true;
	signal G2395: std_logic; attribute dont_touch of G2395: signal is true;
	signal G2396: std_logic; attribute dont_touch of G2396: signal is true;
	signal G2397: std_logic; attribute dont_touch of G2397: signal is true;
	signal G2401: std_logic; attribute dont_touch of G2401: signal is true;
	signal G2402: std_logic; attribute dont_touch of G2402: signal is true;
	signal G2403: std_logic; attribute dont_touch of G2403: signal is true;
	signal G2404: std_logic; attribute dont_touch of G2404: signal is true;
	signal G2407: std_logic; attribute dont_touch of G2407: signal is true;
	signal G2424: std_logic; attribute dont_touch of G2424: signal is true;
	signal G2452: std_logic; attribute dont_touch of G2452: signal is true;
	signal G2453: std_logic; attribute dont_touch of G2453: signal is true;
	signal G2454: std_logic; attribute dont_touch of G2454: signal is true;
	signal G2457: std_logic; attribute dont_touch of G2457: signal is true;
	signal G2458: std_logic; attribute dont_touch of G2458: signal is true;
	signal G2459: std_logic; attribute dont_touch of G2459: signal is true;
	signal G2460: std_logic; attribute dont_touch of G2460: signal is true;
	signal G2467: std_logic; attribute dont_touch of G2467: signal is true;
	signal G2470: std_logic; attribute dont_touch of G2470: signal is true;
	signal G2471: std_logic; attribute dont_touch of G2471: signal is true;
	signal G2474: std_logic; attribute dont_touch of G2474: signal is true;
	signal G2477: std_logic; attribute dont_touch of G2477: signal is true;
	signal G2478: std_logic; attribute dont_touch of G2478: signal is true;
	signal G2479: std_logic; attribute dont_touch of G2479: signal is true;
	signal G2480: std_logic; attribute dont_touch of G2480: signal is true;
	signal G2481: std_logic; attribute dont_touch of G2481: signal is true;
	signal G2484: std_logic; attribute dont_touch of G2484: signal is true;
	signal G2485: std_logic; attribute dont_touch of G2485: signal is true;
	signal G2486: std_logic; attribute dont_touch of G2486: signal is true;
	signal G2487: std_logic; attribute dont_touch of G2487: signal is true;
	signal G2490: std_logic; attribute dont_touch of G2490: signal is true;
	signal G2494: std_logic; attribute dont_touch of G2494: signal is true;
	signal G2495: std_logic; attribute dont_touch of G2495: signal is true;
	signal G2496: std_logic; attribute dont_touch of G2496: signal is true;
	signal G2497: std_logic; attribute dont_touch of G2497: signal is true;
	signal G2498: std_logic; attribute dont_touch of G2498: signal is true;
	signal G2501: std_logic; attribute dont_touch of G2501: signal is true;
	signal G2502: std_logic; attribute dont_touch of G2502: signal is true;
	signal G2505: std_logic; attribute dont_touch of G2505: signal is true;
	signal G2506: std_logic; attribute dont_touch of G2506: signal is true;
	signal G2509: std_logic; attribute dont_touch of G2509: signal is true;
	signal G2510: std_logic; attribute dont_touch of G2510: signal is true;
	signal G2511: std_logic; attribute dont_touch of G2511: signal is true;
	signal G2514: std_logic; attribute dont_touch of G2514: signal is true;
	signal G2517: std_logic; attribute dont_touch of G2517: signal is true;
	signal G2520: std_logic; attribute dont_touch of G2520: signal is true;
	signal G2521: std_logic; attribute dont_touch of G2521: signal is true;
	signal G2522: std_logic; attribute dont_touch of G2522: signal is true;
	signal G2525: std_logic; attribute dont_touch of G2525: signal is true;
	signal G2528: std_logic; attribute dont_touch of G2528: signal is true;
	signal G2532: std_logic; attribute dont_touch of G2532: signal is true;
	signal G2533: std_logic; attribute dont_touch of G2533: signal is true;
	signal G2536: std_logic; attribute dont_touch of G2536: signal is true;
	signal G2539: std_logic; attribute dont_touch of G2539: signal is true;
	signal G2540: std_logic; attribute dont_touch of G2540: signal is true;
	signal G2543: std_logic; attribute dont_touch of G2543: signal is true;
	signal G2546: std_logic; attribute dont_touch of G2546: signal is true;
	signal G2547: std_logic; attribute dont_touch of G2547: signal is true;
	signal G2548: std_logic; attribute dont_touch of G2548: signal is true;
	signal G2551: std_logic; attribute dont_touch of G2551: signal is true;
	signal G2554: std_logic; attribute dont_touch of G2554: signal is true;
	signal G2555: std_logic; attribute dont_touch of G2555: signal is true;
	signal G2556: std_logic; attribute dont_touch of G2556: signal is true;
	signal G2557: std_logic; attribute dont_touch of G2557: signal is true;
	signal G2561: std_logic; attribute dont_touch of G2561: signal is true;
	signal G2562: std_logic; attribute dont_touch of G2562: signal is true;
	signal G2573: std_logic; attribute dont_touch of G2573: signal is true;
	signal G2584: std_logic; attribute dont_touch of G2584: signal is true;
	signal G2595: std_logic; attribute dont_touch of G2595: signal is true;
	signal G2605: std_logic; attribute dont_touch of G2605: signal is true;
	signal G2614: std_logic; attribute dont_touch of G2614: signal is true;
	signal G2615: std_logic; attribute dont_touch of G2615: signal is true;
	signal G2616: std_logic; attribute dont_touch of G2616: signal is true;
	signal G2617: std_logic; attribute dont_touch of G2617: signal is true;
	signal G2618: std_logic; attribute dont_touch of G2618: signal is true;
	signal G2621: std_logic; attribute dont_touch of G2621: signal is true;
	signal G2622: std_logic; attribute dont_touch of G2622: signal is true;
	signal G2623: std_logic; attribute dont_touch of G2623: signal is true;
	signal G2624: std_logic; attribute dont_touch of G2624: signal is true;
	signal G2625: std_logic; attribute dont_touch of G2625: signal is true;
	signal G2626: std_logic; attribute dont_touch of G2626: signal is true;
	signal G2627: std_logic; attribute dont_touch of G2627: signal is true;
	signal G2628: std_logic; attribute dont_touch of G2628: signal is true;
	signal G2629: std_logic; attribute dont_touch of G2629: signal is true;
	signal G2630: std_logic; attribute dont_touch of G2630: signal is true;
	signal G2631: std_logic; attribute dont_touch of G2631: signal is true;
	signal G2632: std_logic; attribute dont_touch of G2632: signal is true;
	signal G2633: std_logic; attribute dont_touch of G2633: signal is true;
	signal G2634: std_logic; attribute dont_touch of G2634: signal is true;
	signal G2635: std_logic; attribute dont_touch of G2635: signal is true;
	signal G2636: std_logic; attribute dont_touch of G2636: signal is true;
	signal G2637: std_logic; attribute dont_touch of G2637: signal is true;
	signal G2638: std_logic; attribute dont_touch of G2638: signal is true;
	signal G2639: std_logic; attribute dont_touch of G2639: signal is true;
	signal G2640: std_logic; attribute dont_touch of G2640: signal is true;
	signal G2641: std_logic; attribute dont_touch of G2641: signal is true;
	signal G2642: std_logic; attribute dont_touch of G2642: signal is true;
	signal G2643: std_logic; attribute dont_touch of G2643: signal is true;
	signal G2644: std_logic; attribute dont_touch of G2644: signal is true;
	signal G2645: std_logic; attribute dont_touch of G2645: signal is true;
	signal G2646: std_logic; attribute dont_touch of G2646: signal is true;
	signal G2647: std_logic; attribute dont_touch of G2647: signal is true;
	signal G2648: std_logic; attribute dont_touch of G2648: signal is true;
	signal G2649: std_logic; attribute dont_touch of G2649: signal is true;
	signal G2650: std_logic; attribute dont_touch of G2650: signal is true;
	signal G2651: std_logic; attribute dont_touch of G2651: signal is true;
	signal G2652: std_logic; attribute dont_touch of G2652: signal is true;
	signal G2653: std_logic; attribute dont_touch of G2653: signal is true;
	signal G2654: std_logic; attribute dont_touch of G2654: signal is true;
	signal G2655: std_logic; attribute dont_touch of G2655: signal is true;
	signal G2659: std_logic; attribute dont_touch of G2659: signal is true;
	signal G2660: std_logic; attribute dont_touch of G2660: signal is true;
	signal G2661: std_logic; attribute dont_touch of G2661: signal is true;
	signal G2663: std_logic; attribute dont_touch of G2663: signal is true;
	signal G2664: std_logic; attribute dont_touch of G2664: signal is true;
	signal G2665: std_logic; attribute dont_touch of G2665: signal is true;
	signal G2668: std_logic; attribute dont_touch of G2668: signal is true;
	signal G2671: std_logic; attribute dont_touch of G2671: signal is true;
	signal G2672: std_logic; attribute dont_touch of G2672: signal is true;
	signal G2673: std_logic; attribute dont_touch of G2673: signal is true;
	signal G2674: std_logic; attribute dont_touch of G2674: signal is true;
	signal G2677: std_logic; attribute dont_touch of G2677: signal is true;
	signal G2680: std_logic; attribute dont_touch of G2680: signal is true;
	signal G2683: std_logic; attribute dont_touch of G2683: signal is true;
	signal G2686: std_logic; attribute dont_touch of G2686: signal is true;
	signal G2689: std_logic; attribute dont_touch of G2689: signal is true;
	signal G2692: std_logic; attribute dont_touch of G2692: signal is true;
	signal G2695: std_logic; attribute dont_touch of G2695: signal is true;
	signal G2698: std_logic; attribute dont_touch of G2698: signal is true;
	signal G2699: std_logic; attribute dont_touch of G2699: signal is true;
	signal G2700: std_logic; attribute dont_touch of G2700: signal is true;
	signal G2703: std_logic; attribute dont_touch of G2703: signal is true;
	signal G2706: std_logic; attribute dont_touch of G2706: signal is true;
	signal G2709: std_logic; attribute dont_touch of G2709: signal is true;
	signal G2712: std_logic; attribute dont_touch of G2712: signal is true;
	signal G2721: std_logic; attribute dont_touch of G2721: signal is true;
	signal G2724: std_logic; attribute dont_touch of G2724: signal is true;
	signal G2727: std_logic; attribute dont_touch of G2727: signal is true;
	signal G2728: std_logic; attribute dont_touch of G2728: signal is true;
	signal G2734: std_logic; attribute dont_touch of G2734: signal is true;
	signal G2743: std_logic; attribute dont_touch of G2743: signal is true;
	signal G2746: std_logic; attribute dont_touch of G2746: signal is true;
	signal G2751: std_logic; attribute dont_touch of G2751: signal is true;
	signal G2752: std_logic; attribute dont_touch of G2752: signal is true;
	signal G2761: std_logic; attribute dont_touch of G2761: signal is true;
	signal G2764: std_logic; attribute dont_touch of G2764: signal is true;
	signal G2767: std_logic; attribute dont_touch of G2767: signal is true;
	signal G2768: std_logic; attribute dont_touch of G2768: signal is true;
	signal G2769: std_logic; attribute dont_touch of G2769: signal is true;
	signal G2770: std_logic; attribute dont_touch of G2770: signal is true;
	signal G2774: std_logic; attribute dont_touch of G2774: signal is true;
	signal G2777: std_logic; attribute dont_touch of G2777: signal is true;
	signal G2780: std_logic; attribute dont_touch of G2780: signal is true;
	signal G2781: std_logic; attribute dont_touch of G2781: signal is true;
	signal G2782: std_logic; attribute dont_touch of G2782: signal is true;
	signal G2783: std_logic; attribute dont_touch of G2783: signal is true;
	signal G2784: std_logic; attribute dont_touch of G2784: signal is true;
	signal G2787: std_logic; attribute dont_touch of G2787: signal is true;
	signal G2790: std_logic; attribute dont_touch of G2790: signal is true;
	signal G2793: std_logic; attribute dont_touch of G2793: signal is true;
	signal G2794: std_logic; attribute dont_touch of G2794: signal is true;
	signal G2795: std_logic; attribute dont_touch of G2795: signal is true;
	signal G2798: std_logic; attribute dont_touch of G2798: signal is true;
	signal G2801: std_logic; attribute dont_touch of G2801: signal is true;
	signal G2804: std_logic; attribute dont_touch of G2804: signal is true;
	signal G2807: std_logic; attribute dont_touch of G2807: signal is true;
	signal G2810: std_logic; attribute dont_touch of G2810: signal is true;
	signal G2816: std_logic; attribute dont_touch of G2816: signal is true;
	signal G2817: std_logic; attribute dont_touch of G2817: signal is true;
	signal G2818: std_logic; attribute dont_touch of G2818: signal is true;
	signal G2821: std_logic; attribute dont_touch of G2821: signal is true;
	signal G2824: std_logic; attribute dont_touch of G2824: signal is true;
	signal G2825: std_logic; attribute dont_touch of G2825: signal is true;
	signal G2826: std_logic; attribute dont_touch of G2826: signal is true;
	signal G2827: std_logic; attribute dont_touch of G2827: signal is true;
	signal G2828: std_logic; attribute dont_touch of G2828: signal is true;
	signal G2829: std_logic; attribute dont_touch of G2829: signal is true;
	signal G2832: std_logic; attribute dont_touch of G2832: signal is true;
	signal G2833: std_logic; attribute dont_touch of G2833: signal is true;
	signal G2834: std_logic; attribute dont_touch of G2834: signal is true;
	signal G2837: std_logic; attribute dont_touch of G2837: signal is true;
	signal G2840: std_logic; attribute dont_touch of G2840: signal is true;
	signal G2841: std_logic; attribute dont_touch of G2841: signal is true;
	signal G2842: std_logic; attribute dont_touch of G2842: signal is true;
	signal G2843: std_logic; attribute dont_touch of G2843: signal is true;
	signal G2845: std_logic; attribute dont_touch of G2845: signal is true;
	signal G2862: std_logic; attribute dont_touch of G2862: signal is true;
	signal G2863: std_logic; attribute dont_touch of G2863: signal is true;
	signal G2866: std_logic; attribute dont_touch of G2866: signal is true;
	signal G2867: std_logic; attribute dont_touch of G2867: signal is true;
	signal G2868: std_logic; attribute dont_touch of G2868: signal is true;
	signal G2869: std_logic; attribute dont_touch of G2869: signal is true;
	signal G2870: std_logic; attribute dont_touch of G2870: signal is true;
	signal G2871: std_logic; attribute dont_touch of G2871: signal is true;
	signal G2872: std_logic; attribute dont_touch of G2872: signal is true;
	signal G2873: std_logic; attribute dont_touch of G2873: signal is true;
	signal G2876: std_logic; attribute dont_touch of G2876: signal is true;
	signal G2877: std_logic; attribute dont_touch of G2877: signal is true;
	signal G2878: std_logic; attribute dont_touch of G2878: signal is true;
	signal G2879: std_logic; attribute dont_touch of G2879: signal is true;
	signal G2880: std_logic; attribute dont_touch of G2880: signal is true;
	signal G2881: std_logic; attribute dont_touch of G2881: signal is true;
	signal G2882: std_logic; attribute dont_touch of G2882: signal is true;
	signal G2883: std_logic; attribute dont_touch of G2883: signal is true;
	signal G2884: std_logic; attribute dont_touch of G2884: signal is true;
	signal G2885: std_logic; attribute dont_touch of G2885: signal is true;
	signal G2886: std_logic; attribute dont_touch of G2886: signal is true;
	signal G2887: std_logic; attribute dont_touch of G2887: signal is true;
	signal G2889: std_logic; attribute dont_touch of G2889: signal is true;
	signal G2890: std_logic; attribute dont_touch of G2890: signal is true;
	signal G2891: std_logic; attribute dont_touch of G2891: signal is true;
	signal G2892: std_logic; attribute dont_touch of G2892: signal is true;
	signal G2893: std_logic; attribute dont_touch of G2893: signal is true;
	signal G2894: std_logic; attribute dont_touch of G2894: signal is true;
	signal G2895: std_logic; attribute dont_touch of G2895: signal is true;
	signal G2896: std_logic; attribute dont_touch of G2896: signal is true;
	signal G2897: std_logic; attribute dont_touch of G2897: signal is true;
	signal G2898: std_logic; attribute dont_touch of G2898: signal is true;
	signal G2899: std_logic; attribute dont_touch of G2899: signal is true;
	signal G2900: std_logic; attribute dont_touch of G2900: signal is true;
	signal G2901: std_logic; attribute dont_touch of G2901: signal is true;
	signal G2902: std_logic; attribute dont_touch of G2902: signal is true;
	signal G2903: std_logic; attribute dont_touch of G2903: signal is true;
	signal G2904: std_logic; attribute dont_touch of G2904: signal is true;
	signal G2905: std_logic; attribute dont_touch of G2905: signal is true;
	signal G2906: std_logic; attribute dont_touch of G2906: signal is true;
	signal G2907: std_logic; attribute dont_touch of G2907: signal is true;
	signal G2908: std_logic; attribute dont_touch of G2908: signal is true;
	signal G2909: std_logic; attribute dont_touch of G2909: signal is true;
	signal G2910: std_logic; attribute dont_touch of G2910: signal is true;
	signal G2911: std_logic; attribute dont_touch of G2911: signal is true;
	signal G2912: std_logic; attribute dont_touch of G2912: signal is true;
	signal G2913: std_logic; attribute dont_touch of G2913: signal is true;
	signal G2914: std_logic; attribute dont_touch of G2914: signal is true;
	signal G2915: std_logic; attribute dont_touch of G2915: signal is true;
	signal G2916: std_logic; attribute dont_touch of G2916: signal is true;
	signal G2917: std_logic; attribute dont_touch of G2917: signal is true;
	signal G2918: std_logic; attribute dont_touch of G2918: signal is true;
	signal G2919: std_logic; attribute dont_touch of G2919: signal is true;
	signal G2920: std_logic; attribute dont_touch of G2920: signal is true;
	signal G2921: std_logic; attribute dont_touch of G2921: signal is true;
	signal G2922: std_logic; attribute dont_touch of G2922: signal is true;
	signal G2923: std_logic; attribute dont_touch of G2923: signal is true;
	signal G2924: std_logic; attribute dont_touch of G2924: signal is true;
	signal G2925: std_logic; attribute dont_touch of G2925: signal is true;
	signal G2926: std_logic; attribute dont_touch of G2926: signal is true;
	signal G2927: std_logic; attribute dont_touch of G2927: signal is true;
	signal G2928: std_logic; attribute dont_touch of G2928: signal is true;
	signal G2929: std_logic; attribute dont_touch of G2929: signal is true;
	signal G2930: std_logic; attribute dont_touch of G2930: signal is true;
	signal G2931: std_logic; attribute dont_touch of G2931: signal is true;
	signal G2932: std_logic; attribute dont_touch of G2932: signal is true;
	signal G2933: std_logic; attribute dont_touch of G2933: signal is true;
	signal G2934: std_logic; attribute dont_touch of G2934: signal is true;
	signal G2935: std_logic; attribute dont_touch of G2935: signal is true;
	signal G2936: std_logic; attribute dont_touch of G2936: signal is true;
	signal G2937: std_logic; attribute dont_touch of G2937: signal is true;
	signal G2938: std_logic; attribute dont_touch of G2938: signal is true;
	signal G2939: std_logic; attribute dont_touch of G2939: signal is true;
	signal G2940: std_logic; attribute dont_touch of G2940: signal is true;
	signal G2941: std_logic; attribute dont_touch of G2941: signal is true;
	signal G2942: std_logic; attribute dont_touch of G2942: signal is true;
	signal G2943: std_logic; attribute dont_touch of G2943: signal is true;
	signal G2944: std_logic; attribute dont_touch of G2944: signal is true;
	signal G2945: std_logic; attribute dont_touch of G2945: signal is true;
	signal G2946: std_logic; attribute dont_touch of G2946: signal is true;
	signal G2947: std_logic; attribute dont_touch of G2947: signal is true;
	signal G2948: std_logic; attribute dont_touch of G2948: signal is true;
	signal G2949: std_logic; attribute dont_touch of G2949: signal is true;
	signal G2952: std_logic; attribute dont_touch of G2952: signal is true;
	signal G2953: std_logic; attribute dont_touch of G2953: signal is true;
	signal G2954: std_logic; attribute dont_touch of G2954: signal is true;
	signal G2955: std_logic; attribute dont_touch of G2955: signal is true;
	signal G2956: std_logic; attribute dont_touch of G2956: signal is true;
	signal G2957: std_logic; attribute dont_touch of G2957: signal is true;
	signal G2958: std_logic; attribute dont_touch of G2958: signal is true;
	signal G2959: std_logic; attribute dont_touch of G2959: signal is true;
	signal G2960: std_logic; attribute dont_touch of G2960: signal is true;
	signal G2961: std_logic; attribute dont_touch of G2961: signal is true;
	signal G2962: std_logic; attribute dont_touch of G2962: signal is true;
	signal G2963: std_logic; attribute dont_touch of G2963: signal is true;
	signal G2964: std_logic; attribute dont_touch of G2964: signal is true;
	signal G2965: std_logic; attribute dont_touch of G2965: signal is true;
	signal G2966: std_logic; attribute dont_touch of G2966: signal is true;
	signal G2969: std_logic; attribute dont_touch of G2969: signal is true;
	signal G2970: std_logic; attribute dont_touch of G2970: signal is true;
	signal G2971: std_logic; attribute dont_touch of G2971: signal is true;
	signal G2972: std_logic; attribute dont_touch of G2972: signal is true;
	signal G2973: std_logic; attribute dont_touch of G2973: signal is true;
	signal G2976: std_logic; attribute dont_touch of G2976: signal is true;
	signal G2979: std_logic; attribute dont_touch of G2979: signal is true;
	signal G2982: std_logic; attribute dont_touch of G2982: signal is true;
	signal G2985: std_logic; attribute dont_touch of G2985: signal is true;
	signal G2986: std_logic; attribute dont_touch of G2986: signal is true;
	signal G2989: std_logic; attribute dont_touch of G2989: signal is true;
	signal G2992: std_logic; attribute dont_touch of G2992: signal is true;
	signal G2995: std_logic; attribute dont_touch of G2995: signal is true;
	signal G2996: std_logic; attribute dont_touch of G2996: signal is true;
	signal G2999: std_logic; attribute dont_touch of G2999: signal is true;
	signal G3002: std_logic; attribute dont_touch of G3002: signal is true;
	signal G3008: std_logic; attribute dont_touch of G3008: signal is true;
	signal G3011: std_logic; attribute dont_touch of G3011: signal is true;
	signal G3012: std_logic; attribute dont_touch of G3012: signal is true;
	signal G3013: std_logic; attribute dont_touch of G3013: signal is true;
	signal G3014: std_logic; attribute dont_touch of G3014: signal is true;
	signal G3018: std_logic; attribute dont_touch of G3018: signal is true;
	signal G3019: std_logic; attribute dont_touch of G3019: signal is true;
	signal G3028: std_logic; attribute dont_touch of G3028: signal is true;
	signal G3029: std_logic; attribute dont_touch of G3029: signal is true;
	signal G3038: std_logic; attribute dont_touch of G3038: signal is true;
	signal G3047: std_logic; attribute dont_touch of G3047: signal is true;
	signal G3048: std_logic; attribute dont_touch of G3048: signal is true;
	signal G3049: std_logic; attribute dont_touch of G3049: signal is true;
	signal G3050: std_logic; attribute dont_touch of G3050: signal is true;
	signal G3051: std_logic; attribute dont_touch of G3051: signal is true;
	signal G3052: std_logic; attribute dont_touch of G3052: signal is true;
	signal G3061: std_logic; attribute dont_touch of G3061: signal is true;
	signal G3062: std_logic; attribute dont_touch of G3062: signal is true;
	signal G3071: std_logic; attribute dont_touch of G3071: signal is true;
	signal G3074: std_logic; attribute dont_touch of G3074: signal is true;
	signal G3075: std_logic; attribute dont_touch of G3075: signal is true;
	signal G3076: std_logic; attribute dont_touch of G3076: signal is true;
	signal G3078: std_logic; attribute dont_touch of G3078: signal is true;
	signal G3079: std_logic; attribute dont_touch of G3079: signal is true;
	signal G3080: std_logic; attribute dont_touch of G3080: signal is true;
	signal G3081: std_logic; attribute dont_touch of G3081: signal is true;
	signal G3082: std_logic; attribute dont_touch of G3082: signal is true;
	signal G3083: std_logic; attribute dont_touch of G3083: signal is true;
	signal G3084: std_logic; attribute dont_touch of G3084: signal is true;
	signal G3085: std_logic; attribute dont_touch of G3085: signal is true;
	signal G3086: std_logic; attribute dont_touch of G3086: signal is true;
	signal G3091: std_logic; attribute dont_touch of G3091: signal is true;
	signal G3092: std_logic; attribute dont_touch of G3092: signal is true;
	signal G3093: std_logic; attribute dont_touch of G3093: signal is true;
	signal G3094: std_logic; attribute dont_touch of G3094: signal is true;
	signal G3095: std_logic; attribute dont_touch of G3095: signal is true;
	signal G3097: std_logic; attribute dont_touch of G3097: signal is true;
	signal G3124: std_logic; attribute dont_touch of G3124: signal is true;
	signal G3128: std_logic; attribute dont_touch of G3128: signal is true;
	signal G3129: std_logic; attribute dont_touch of G3129: signal is true;
	signal G3131: std_logic; attribute dont_touch of G3131: signal is true;
	signal G3158: std_logic; attribute dont_touch of G3158: signal is true;
	signal G3160: std_logic; attribute dont_touch of G3160: signal is true;
	signal G3187: std_logic; attribute dont_touch of G3187: signal is true;
	signal G3188: std_logic; attribute dont_touch of G3188: signal is true;
	signal G3189: std_logic; attribute dont_touch of G3189: signal is true;
	signal G3190: std_logic; attribute dont_touch of G3190: signal is true;
	signal G3192: std_logic; attribute dont_touch of G3192: signal is true;
	signal G3219: std_logic; attribute dont_touch of G3219: signal is true;
	signal G3220: std_logic; attribute dont_touch of G3220: signal is true;
	signal G3221: std_logic; attribute dont_touch of G3221: signal is true;
	signal G3222: std_logic; attribute dont_touch of G3222: signal is true;
	signal G3225: std_logic; attribute dont_touch of G3225: signal is true;
	signal G3226: std_logic; attribute dont_touch of G3226: signal is true;
	signal G3229: std_logic; attribute dont_touch of G3229: signal is true;
	signal G3230: std_logic; attribute dont_touch of G3230: signal is true;
	signal G3231: std_logic; attribute dont_touch of G3231: signal is true;
	signal G3232: std_logic; attribute dont_touch of G3232: signal is true;
	signal G3233: std_logic; attribute dont_touch of G3233: signal is true;
	signal G3237: std_logic; attribute dont_touch of G3237: signal is true;
	signal G3238: std_logic; attribute dont_touch of G3238: signal is true;
	signal G3258: std_logic; attribute dont_touch of G3258: signal is true;
	signal G3259: std_logic; attribute dont_touch of G3259: signal is true;
	signal G3260: std_logic; attribute dont_touch of G3260: signal is true;
	signal G3264: std_logic; attribute dont_touch of G3264: signal is true;
	signal G3285: std_logic; attribute dont_touch of G3285: signal is true;
	signal G3286: std_logic; attribute dont_touch of G3286: signal is true;
	signal G3287: std_logic; attribute dont_touch of G3287: signal is true;
	signal G3310: std_logic; attribute dont_touch of G3310: signal is true;
	signal G3313: std_logic; attribute dont_touch of G3313: signal is true;
	signal G3314: std_logic; attribute dont_touch of G3314: signal is true;
	signal G3315: std_logic; attribute dont_touch of G3315: signal is true;
	signal G3316: std_logic; attribute dont_touch of G3316: signal is true;
	signal G3338: std_logic; attribute dont_touch of G3338: signal is true;
	signal G3339: std_logic; attribute dont_touch of G3339: signal is true;
	signal G3340: std_logic; attribute dont_touch of G3340: signal is true;
	signal G3341: std_logic; attribute dont_touch of G3341: signal is true;
	signal G3358: std_logic; attribute dont_touch of G3358: signal is true;
	signal G3359: std_logic; attribute dont_touch of G3359: signal is true;
	signal G3390: std_logic; attribute dont_touch of G3390: signal is true;
	signal G3398: std_logic; attribute dont_touch of G3398: signal is true;
	signal G3429: std_logic; attribute dont_touch of G3429: signal is true;
	signal G3430: std_logic; attribute dont_touch of G3430: signal is true;
	signal G3461: std_logic; attribute dont_touch of G3461: signal is true;
	signal G3462: std_logic; attribute dont_touch of G3462: signal is true;
	signal G3465: std_logic; attribute dont_touch of G3465: signal is true;
	signal G3466: std_logic; attribute dont_touch of G3466: signal is true;
	signal G3485: std_logic; attribute dont_touch of G3485: signal is true;
	signal G3488: std_logic; attribute dont_touch of G3488: signal is true;
	signal G3491: std_logic; attribute dont_touch of G3491: signal is true;
	signal G3492: std_logic; attribute dont_touch of G3492: signal is true;
	signal G3495: std_logic; attribute dont_touch of G3495: signal is true;
	signal G3496: std_logic; attribute dont_touch of G3496: signal is true;
	signal G3497: std_logic; attribute dont_touch of G3497: signal is true;
	signal G3498: std_logic; attribute dont_touch of G3498: signal is true;
	signal G3499: std_logic; attribute dont_touch of G3499: signal is true;
	signal G3500: std_logic; attribute dont_touch of G3500: signal is true;
	signal G3501: std_logic; attribute dont_touch of G3501: signal is true;
	signal G3502: std_logic; attribute dont_touch of G3502: signal is true;
	signal G3503: std_logic; attribute dont_touch of G3503: signal is true;
	signal G3504: std_logic; attribute dont_touch of G3504: signal is true;
	signal G3505: std_logic; attribute dont_touch of G3505: signal is true;
	signal G3506: std_logic; attribute dont_touch of G3506: signal is true;
	signal G3509: std_logic; attribute dont_touch of G3509: signal is true;
	signal G3510: std_logic; attribute dont_touch of G3510: signal is true;
	signal G3511: std_logic; attribute dont_touch of G3511: signal is true;
	signal G3512: std_logic; attribute dont_touch of G3512: signal is true;
	signal G3513: std_logic; attribute dont_touch of G3513: signal is true;
	signal G3514: std_logic; attribute dont_touch of G3514: signal is true;
	signal G3515: std_logic; attribute dont_touch of G3515: signal is true;
	signal G3516: std_logic; attribute dont_touch of G3516: signal is true;
	signal G3517: std_logic; attribute dont_touch of G3517: signal is true;
	signal G3518: std_logic; attribute dont_touch of G3518: signal is true;
	signal G3519: std_logic; attribute dont_touch of G3519: signal is true;
	signal G3520: std_logic; attribute dont_touch of G3520: signal is true;
	signal G3521: std_logic; attribute dont_touch of G3521: signal is true;
	signal G3522: std_logic; attribute dont_touch of G3522: signal is true;
	signal G3523: std_logic; attribute dont_touch of G3523: signal is true;
	signal G3524: std_logic; attribute dont_touch of G3524: signal is true;
	signal G3525: std_logic; attribute dont_touch of G3525: signal is true;
	signal G3526: std_logic; attribute dont_touch of G3526: signal is true;
	signal G3527: std_logic; attribute dont_touch of G3527: signal is true;
	signal G3528: std_logic; attribute dont_touch of G3528: signal is true;
	signal G3529: std_logic; attribute dont_touch of G3529: signal is true;
	signal G3530: std_logic; attribute dont_touch of G3530: signal is true;
	signal G3531: std_logic; attribute dont_touch of G3531: signal is true;
	signal G3532: std_logic; attribute dont_touch of G3532: signal is true;
	signal G3533: std_logic; attribute dont_touch of G3533: signal is true;
	signal G3539: std_logic; attribute dont_touch of G3539: signal is true;
	signal G3540: std_logic; attribute dont_touch of G3540: signal is true;
	signal G3541: std_logic; attribute dont_touch of G3541: signal is true;
	signal G3542: std_logic; attribute dont_touch of G3542: signal is true;
	signal G3545: std_logic; attribute dont_touch of G3545: signal is true;
	signal G3546: std_logic; attribute dont_touch of G3546: signal is true;
	signal G3547: std_logic; attribute dont_touch of G3547: signal is true;
	signal G3548: std_logic; attribute dont_touch of G3548: signal is true;
	signal G3549: std_logic; attribute dont_touch of G3549: signal is true;
	signal G3555: std_logic; attribute dont_touch of G3555: signal is true;
	signal G3556: std_logic; attribute dont_touch of G3556: signal is true;
	signal G3557: std_logic; attribute dont_touch of G3557: signal is true;
	signal G3560: std_logic; attribute dont_touch of G3560: signal is true;
	signal G3561: std_logic; attribute dont_touch of G3561: signal is true;
	signal G3562: std_logic; attribute dont_touch of G3562: signal is true;
	signal G3563: std_logic; attribute dont_touch of G3563: signal is true;
	signal G3567: std_logic; attribute dont_touch of G3567: signal is true;
	signal G3568: std_logic; attribute dont_touch of G3568: signal is true;
	signal G3573: std_logic; attribute dont_touch of G3573: signal is true;
	signal G3574: std_logic; attribute dont_touch of G3574: signal is true;
	signal G3577: std_logic; attribute dont_touch of G3577: signal is true;
	signal G3578: std_logic; attribute dont_touch of G3578: signal is true;
	signal G3579: std_logic; attribute dont_touch of G3579: signal is true;
	signal G3582: std_logic; attribute dont_touch of G3582: signal is true;
	signal G3583: std_logic; attribute dont_touch of G3583: signal is true;
	signal G3587: std_logic; attribute dont_touch of G3587: signal is true;
	signal G3588: std_logic; attribute dont_touch of G3588: signal is true;
	signal G3589: std_logic; attribute dont_touch of G3589: signal is true;
	signal G3590: std_logic; attribute dont_touch of G3590: signal is true;
	signal G3591: std_logic; attribute dont_touch of G3591: signal is true;
	signal G3602: std_logic; attribute dont_touch of G3602: signal is true;
	signal G3603: std_logic; attribute dont_touch of G3603: signal is true;
	signal G3604: std_logic; attribute dont_touch of G3604: signal is true;
	signal G3605: std_logic; attribute dont_touch of G3605: signal is true;
	signal G3610: std_logic; attribute dont_touch of G3610: signal is true;
	signal G3611: std_logic; attribute dont_touch of G3611: signal is true;
	signal G3612: std_logic; attribute dont_touch of G3612: signal is true;
	signal G3613: std_logic; attribute dont_touch of G3613: signal is true;
	signal G3614: std_logic; attribute dont_touch of G3614: signal is true;
	signal G3617: std_logic; attribute dont_touch of G3617: signal is true;
	signal G3629: std_logic; attribute dont_touch of G3629: signal is true;
	signal G3630: std_logic; attribute dont_touch of G3630: signal is true;
	signal G3631: std_logic; attribute dont_touch of G3631: signal is true;
	signal G3632: std_logic; attribute dont_touch of G3632: signal is true;
	signal G3633: std_logic; attribute dont_touch of G3633: signal is true;
	signal G3634: std_logic; attribute dont_touch of G3634: signal is true;
	signal G3635: std_logic; attribute dont_touch of G3635: signal is true;
	signal G3639: std_logic; attribute dont_touch of G3639: signal is true;
	signal G3640: std_logic; attribute dont_touch of G3640: signal is true;
	signal G3641: std_logic; attribute dont_touch of G3641: signal is true;
	signal G3642: std_logic; attribute dont_touch of G3642: signal is true;
	signal G3643: std_logic; attribute dont_touch of G3643: signal is true;
	signal G3644: std_logic; attribute dont_touch of G3644: signal is true;
	signal G3647: std_logic; attribute dont_touch of G3647: signal is true;
	signal G3648: std_logic; attribute dont_touch of G3648: signal is true;
	signal G3649: std_logic; attribute dont_touch of G3649: signal is true;
	signal G3650: std_logic; attribute dont_touch of G3650: signal is true;
	signal G3651: std_logic; attribute dont_touch of G3651: signal is true;
	signal G3652: std_logic; attribute dont_touch of G3652: signal is true;
	signal G3653: std_logic; attribute dont_touch of G3653: signal is true;
	signal G3654: std_logic; attribute dont_touch of G3654: signal is true;
	signal G3655: std_logic; attribute dont_touch of G3655: signal is true;
	signal G3656: std_logic; attribute dont_touch of G3656: signal is true;
	signal G3657: std_logic; attribute dont_touch of G3657: signal is true;
	signal G3658: std_logic; attribute dont_touch of G3658: signal is true;
	signal G3659: std_logic; attribute dont_touch of G3659: signal is true;
	signal G3665: std_logic; attribute dont_touch of G3665: signal is true;
	signal G3666: std_logic; attribute dont_touch of G3666: signal is true;
	signal G3674: std_logic; attribute dont_touch of G3674: signal is true;
	signal G3675: std_logic; attribute dont_touch of G3675: signal is true;
	signal G3676: std_logic; attribute dont_touch of G3676: signal is true;
	signal G3677: std_logic; attribute dont_touch of G3677: signal is true;
	signal G3678: std_logic; attribute dont_touch of G3678: signal is true;
	signal G3679: std_logic; attribute dont_touch of G3679: signal is true;
	signal G3680: std_logic; attribute dont_touch of G3680: signal is true;
	signal G3681: std_logic; attribute dont_touch of G3681: signal is true;
	signal G3684: std_logic; attribute dont_touch of G3684: signal is true;
	signal G3691: std_logic; attribute dont_touch of G3691: signal is true;
	signal G3692: std_logic; attribute dont_touch of G3692: signal is true;
	signal G3693: std_logic; attribute dont_touch of G3693: signal is true;
	signal G3694: std_logic; attribute dont_touch of G3694: signal is true;
	signal G3700: std_logic; attribute dont_touch of G3700: signal is true;
	signal G3705: std_logic; attribute dont_touch of G3705: signal is true;
	signal G3706: std_logic; attribute dont_touch of G3706: signal is true;
	signal G3707: std_logic; attribute dont_touch of G3707: signal is true;
	signal G3712: std_logic; attribute dont_touch of G3712: signal is true;
	signal G3716: std_logic; attribute dont_touch of G3716: signal is true;
	signal G3721: std_logic; attribute dont_touch of G3721: signal is true;
	signal G3722: std_logic; attribute dont_touch of G3722: signal is true;
	signal G3723: std_logic; attribute dont_touch of G3723: signal is true;
	signal G3728: std_logic; attribute dont_touch of G3728: signal is true;
	signal G3732: std_logic; attribute dont_touch of G3732: signal is true;
	signal G3735: std_logic; attribute dont_touch of G3735: signal is true;
	signal G3739: std_logic; attribute dont_touch of G3739: signal is true;
	signal G3743: std_logic; attribute dont_touch of G3743: signal is true;
	signal G3746: std_logic; attribute dont_touch of G3746: signal is true;
	signal G3750: std_logic; attribute dont_touch of G3750: signal is true;
	signal G3753: std_logic; attribute dont_touch of G3753: signal is true;
	signal G3754: std_logic; attribute dont_touch of G3754: signal is true;
	signal G3757: std_logic; attribute dont_touch of G3757: signal is true;
	signal G3760: std_logic; attribute dont_touch of G3760: signal is true;
	signal G3761: std_logic; attribute dont_touch of G3761: signal is true;
	signal G3764: std_logic; attribute dont_touch of G3764: signal is true;
	signal G3767: std_logic; attribute dont_touch of G3767: signal is true;
	signal G3768: std_logic; attribute dont_touch of G3768: signal is true;
	signal G3769: std_logic; attribute dont_touch of G3769: signal is true;
	signal G3770: std_logic; attribute dont_touch of G3770: signal is true;
	signal G3771: std_logic; attribute dont_touch of G3771: signal is true;
	signal G3774: std_logic; attribute dont_touch of G3774: signal is true;
	signal G3777: std_logic; attribute dont_touch of G3777: signal is true;
	signal G3778: std_logic; attribute dont_touch of G3778: signal is true;
	signal G3779: std_logic; attribute dont_touch of G3779: signal is true;
	signal G3780: std_logic; attribute dont_touch of G3780: signal is true;
	signal G3783: std_logic; attribute dont_touch of G3783: signal is true;
	signal G3784: std_logic; attribute dont_touch of G3784: signal is true;
	signal G3787: std_logic; attribute dont_touch of G3787: signal is true;
	signal G3790: std_logic; attribute dont_touch of G3790: signal is true;
	signal G3798: std_logic; attribute dont_touch of G3798: signal is true;
	signal G3801: std_logic; attribute dont_touch of G3801: signal is true;
	signal G3802: std_logic; attribute dont_touch of G3802: signal is true;
	signal G3805: std_logic; attribute dont_touch of G3805: signal is true;
	signal G3808: std_logic; attribute dont_touch of G3808: signal is true;
	signal G3811: std_logic; attribute dont_touch of G3811: signal is true;
	signal G3812: std_logic; attribute dont_touch of G3812: signal is true;
	signal G3815: std_logic; attribute dont_touch of G3815: signal is true;
	signal G3818: std_logic; attribute dont_touch of G3818: signal is true;
	signal G3819: std_logic; attribute dont_touch of G3819: signal is true;
	signal G3822: std_logic; attribute dont_touch of G3822: signal is true;
	signal G3825: std_logic; attribute dont_touch of G3825: signal is true;
	signal G3828: std_logic; attribute dont_touch of G3828: signal is true;
	signal G3830: std_logic; attribute dont_touch of G3830: signal is true;
	signal G3831: std_logic; attribute dont_touch of G3831: signal is true;
	signal G3832: std_logic; attribute dont_touch of G3832: signal is true;
	signal G3833: std_logic; attribute dont_touch of G3833: signal is true;
	signal G3834: std_logic; attribute dont_touch of G3834: signal is true;
	signal G3835: std_logic; attribute dont_touch of G3835: signal is true;
	signal G3836: std_logic; attribute dont_touch of G3836: signal is true;
	signal G3837: std_logic; attribute dont_touch of G3837: signal is true;
	signal G3838: std_logic; attribute dont_touch of G3838: signal is true;
	signal G3839: std_logic; attribute dont_touch of G3839: signal is true;
	signal G3840: std_logic; attribute dont_touch of G3840: signal is true;
	signal G3841: std_logic; attribute dont_touch of G3841: signal is true;
	signal G3842: std_logic; attribute dont_touch of G3842: signal is true;
	signal G3843: std_logic; attribute dont_touch of G3843: signal is true;
	signal G3844: std_logic; attribute dont_touch of G3844: signal is true;
	signal G3845: std_logic; attribute dont_touch of G3845: signal is true;
	signal G3846: std_logic; attribute dont_touch of G3846: signal is true;
	signal G3847: std_logic; attribute dont_touch of G3847: signal is true;
	signal G3848: std_logic; attribute dont_touch of G3848: signal is true;
	signal G3849: std_logic; attribute dont_touch of G3849: signal is true;
	signal G3850: std_logic; attribute dont_touch of G3850: signal is true;
	signal G3851: std_logic; attribute dont_touch of G3851: signal is true;
	signal G3852: std_logic; attribute dont_touch of G3852: signal is true;
	signal G3853: std_logic; attribute dont_touch of G3853: signal is true;
	signal G3855: std_logic; attribute dont_touch of G3855: signal is true;
	signal G3858: std_logic; attribute dont_touch of G3858: signal is true;
	signal G3861: std_logic; attribute dont_touch of G3861: signal is true;
	signal G3862: std_logic; attribute dont_touch of G3862: signal is true;
	signal G3863: std_logic; attribute dont_touch of G3863: signal is true;
	signal G3864: std_logic; attribute dont_touch of G3864: signal is true;
	signal G3865: std_logic; attribute dont_touch of G3865: signal is true;
	signal G3866: std_logic; attribute dont_touch of G3866: signal is true;
	signal G3867: std_logic; attribute dont_touch of G3867: signal is true;
	signal G3868: std_logic; attribute dont_touch of G3868: signal is true;
	signal G3869: std_logic; attribute dont_touch of G3869: signal is true;
	signal G3870: std_logic; attribute dont_touch of G3870: signal is true;
	signal G3871: std_logic; attribute dont_touch of G3871: signal is true;
	signal G3872: std_logic; attribute dont_touch of G3872: signal is true;
	signal G3873: std_logic; attribute dont_touch of G3873: signal is true;
	signal G3874: std_logic; attribute dont_touch of G3874: signal is true;
	signal G3875: std_logic; attribute dont_touch of G3875: signal is true;
	signal G3876: std_logic; attribute dont_touch of G3876: signal is true;
	signal G3877: std_logic; attribute dont_touch of G3877: signal is true;
	signal G3878: std_logic; attribute dont_touch of G3878: signal is true;
	signal G3879: std_logic; attribute dont_touch of G3879: signal is true;
	signal G3880: std_logic; attribute dont_touch of G3880: signal is true;
	signal G3881: std_logic; attribute dont_touch of G3881: signal is true;
	signal G3882: std_logic; attribute dont_touch of G3882: signal is true;
	signal G3883: std_logic; attribute dont_touch of G3883: signal is true;
	signal G3884: std_logic; attribute dont_touch of G3884: signal is true;
	signal G3885: std_logic; attribute dont_touch of G3885: signal is true;
	signal G3886: std_logic; attribute dont_touch of G3886: signal is true;
	signal G3887: std_logic; attribute dont_touch of G3887: signal is true;
	signal G3888: std_logic; attribute dont_touch of G3888: signal is true;
	signal G3889: std_logic; attribute dont_touch of G3889: signal is true;
	signal G3890: std_logic; attribute dont_touch of G3890: signal is true;
	signal G3891: std_logic; attribute dont_touch of G3891: signal is true;
	signal G3892: std_logic; attribute dont_touch of G3892: signal is true;
	signal G3893: std_logic; attribute dont_touch of G3893: signal is true;
	signal G3894: std_logic; attribute dont_touch of G3894: signal is true;
	signal G3895: std_logic; attribute dont_touch of G3895: signal is true;
	signal G3896: std_logic; attribute dont_touch of G3896: signal is true;
	signal G3897: std_logic; attribute dont_touch of G3897: signal is true;
	signal G3898: std_logic; attribute dont_touch of G3898: signal is true;
	signal G3899: std_logic; attribute dont_touch of G3899: signal is true;
	signal G3900: std_logic; attribute dont_touch of G3900: signal is true;
	signal G3901: std_logic; attribute dont_touch of G3901: signal is true;
	signal G3902: std_logic; attribute dont_touch of G3902: signal is true;
	signal G3903: std_logic; attribute dont_touch of G3903: signal is true;
	signal G3904: std_logic; attribute dont_touch of G3904: signal is true;
	signal G3905: std_logic; attribute dont_touch of G3905: signal is true;
	signal G3906: std_logic; attribute dont_touch of G3906: signal is true;
	signal G3907: std_logic; attribute dont_touch of G3907: signal is true;
	signal G3908: std_logic; attribute dont_touch of G3908: signal is true;
	signal G3909: std_logic; attribute dont_touch of G3909: signal is true;
	signal G3910: std_logic; attribute dont_touch of G3910: signal is true;
	signal G3911: std_logic; attribute dont_touch of G3911: signal is true;
	signal G3912: std_logic; attribute dont_touch of G3912: signal is true;
	signal G3913: std_logic; attribute dont_touch of G3913: signal is true;
	signal G3914: std_logic; attribute dont_touch of G3914: signal is true;
	signal G3915: std_logic; attribute dont_touch of G3915: signal is true;
	signal G3916: std_logic; attribute dont_touch of G3916: signal is true;
	signal G3917: std_logic; attribute dont_touch of G3917: signal is true;
	signal G3918: std_logic; attribute dont_touch of G3918: signal is true;
	signal G3919: std_logic; attribute dont_touch of G3919: signal is true;
	signal G3920: std_logic; attribute dont_touch of G3920: signal is true;
	signal G3921: std_logic; attribute dont_touch of G3921: signal is true;
	signal G3922: std_logic; attribute dont_touch of G3922: signal is true;
	signal G3923: std_logic; attribute dont_touch of G3923: signal is true;
	signal G3924: std_logic; attribute dont_touch of G3924: signal is true;
	signal G3925: std_logic; attribute dont_touch of G3925: signal is true;
	signal G3926: std_logic; attribute dont_touch of G3926: signal is true;
	signal G3927: std_logic; attribute dont_touch of G3927: signal is true;
	signal G3928: std_logic; attribute dont_touch of G3928: signal is true;
	signal G3929: std_logic; attribute dont_touch of G3929: signal is true;
	signal G3930: std_logic; attribute dont_touch of G3930: signal is true;
	signal G3931: std_logic; attribute dont_touch of G3931: signal is true;
	signal G3932: std_logic; attribute dont_touch of G3932: signal is true;
	signal G3933: std_logic; attribute dont_touch of G3933: signal is true;
	signal G3934: std_logic; attribute dont_touch of G3934: signal is true;
	signal G3935: std_logic; attribute dont_touch of G3935: signal is true;
	signal G3936: std_logic; attribute dont_touch of G3936: signal is true;
	signal G3937: std_logic; attribute dont_touch of G3937: signal is true;
	signal G3938: std_logic; attribute dont_touch of G3938: signal is true;
	signal G3939: std_logic; attribute dont_touch of G3939: signal is true;
	signal G3940: std_logic; attribute dont_touch of G3940: signal is true;
	signal G3941: std_logic; attribute dont_touch of G3941: signal is true;
	signal G3942: std_logic; attribute dont_touch of G3942: signal is true;
	signal G3943: std_logic; attribute dont_touch of G3943: signal is true;
	signal G3944: std_logic; attribute dont_touch of G3944: signal is true;
	signal G3945: std_logic; attribute dont_touch of G3945: signal is true;
	signal G3946: std_logic; attribute dont_touch of G3946: signal is true;
	signal G3947: std_logic; attribute dont_touch of G3947: signal is true;
	signal G3948: std_logic; attribute dont_touch of G3948: signal is true;
	signal G3949: std_logic; attribute dont_touch of G3949: signal is true;
	signal G3950: std_logic; attribute dont_touch of G3950: signal is true;
	signal G3951: std_logic; attribute dont_touch of G3951: signal is true;
	signal G3952: std_logic; attribute dont_touch of G3952: signal is true;
	signal G3953: std_logic; attribute dont_touch of G3953: signal is true;
	signal G3954: std_logic; attribute dont_touch of G3954: signal is true;
	signal G3955: std_logic; attribute dont_touch of G3955: signal is true;
	signal G3956: std_logic; attribute dont_touch of G3956: signal is true;
	signal G3957: std_logic; attribute dont_touch of G3957: signal is true;
	signal G3958: std_logic; attribute dont_touch of G3958: signal is true;
	signal G3959: std_logic; attribute dont_touch of G3959: signal is true;
	signal G3960: std_logic; attribute dont_touch of G3960: signal is true;
	signal G3961: std_logic; attribute dont_touch of G3961: signal is true;
	signal G3962: std_logic; attribute dont_touch of G3962: signal is true;
	signal G3963: std_logic; attribute dont_touch of G3963: signal is true;
	signal G3964: std_logic; attribute dont_touch of G3964: signal is true;
	signal G3965: std_logic; attribute dont_touch of G3965: signal is true;
	signal G3966: std_logic; attribute dont_touch of G3966: signal is true;
	signal G3967: std_logic; attribute dont_touch of G3967: signal is true;
	signal G3968: std_logic; attribute dont_touch of G3968: signal is true;
	signal G3969: std_logic; attribute dont_touch of G3969: signal is true;
	signal G3970: std_logic; attribute dont_touch of G3970: signal is true;
	signal G3971: std_logic; attribute dont_touch of G3971: signal is true;
	signal G3972: std_logic; attribute dont_touch of G3972: signal is true;
	signal G3973: std_logic; attribute dont_touch of G3973: signal is true;
	signal G3974: std_logic; attribute dont_touch of G3974: signal is true;
	signal G3975: std_logic; attribute dont_touch of G3975: signal is true;
	signal G3976: std_logic; attribute dont_touch of G3976: signal is true;
	signal G3977: std_logic; attribute dont_touch of G3977: signal is true;
	signal G3978: std_logic; attribute dont_touch of G3978: signal is true;
	signal G3979: std_logic; attribute dont_touch of G3979: signal is true;
	signal G3980: std_logic; attribute dont_touch of G3980: signal is true;
	signal G3981: std_logic; attribute dont_touch of G3981: signal is true;
	signal G3982: std_logic; attribute dont_touch of G3982: signal is true;
	signal G3983: std_logic; attribute dont_touch of G3983: signal is true;
	signal G3984: std_logic; attribute dont_touch of G3984: signal is true;
	signal G3985: std_logic; attribute dont_touch of G3985: signal is true;
	signal G3986: std_logic; attribute dont_touch of G3986: signal is true;
	signal G3987: std_logic; attribute dont_touch of G3987: signal is true;
	signal G3988: std_logic; attribute dont_touch of G3988: signal is true;
	signal G3989: std_logic; attribute dont_touch of G3989: signal is true;
	signal G3990: std_logic; attribute dont_touch of G3990: signal is true;
	signal G3991: std_logic; attribute dont_touch of G3991: signal is true;
	signal G3992: std_logic; attribute dont_touch of G3992: signal is true;
	signal G3993: std_logic; attribute dont_touch of G3993: signal is true;
	signal G3994: std_logic; attribute dont_touch of G3994: signal is true;
	signal G3995: std_logic; attribute dont_touch of G3995: signal is true;
	signal G3996: std_logic; attribute dont_touch of G3996: signal is true;
	signal G3997: std_logic; attribute dont_touch of G3997: signal is true;
	signal G3998: std_logic; attribute dont_touch of G3998: signal is true;
	signal G3999: std_logic; attribute dont_touch of G3999: signal is true;
	signal G4000: std_logic; attribute dont_touch of G4000: signal is true;
	signal G4001: std_logic; attribute dont_touch of G4001: signal is true;
	signal G4002: std_logic; attribute dont_touch of G4002: signal is true;
	signal G4003: std_logic; attribute dont_touch of G4003: signal is true;
	signal G4004: std_logic; attribute dont_touch of G4004: signal is true;
	signal G4005: std_logic; attribute dont_touch of G4005: signal is true;
	signal G4006: std_logic; attribute dont_touch of G4006: signal is true;
	signal G4007: std_logic; attribute dont_touch of G4007: signal is true;
	signal G4008: std_logic; attribute dont_touch of G4008: signal is true;
	signal G4009: std_logic; attribute dont_touch of G4009: signal is true;
	signal G4010: std_logic; attribute dont_touch of G4010: signal is true;
	signal G4011: std_logic; attribute dont_touch of G4011: signal is true;
	signal G4012: std_logic; attribute dont_touch of G4012: signal is true;
	signal G4013: std_logic; attribute dont_touch of G4013: signal is true;
	signal G4014: std_logic; attribute dont_touch of G4014: signal is true;
	signal G4015: std_logic; attribute dont_touch of G4015: signal is true;
	signal G4016: std_logic; attribute dont_touch of G4016: signal is true;
	signal G4017: std_logic; attribute dont_touch of G4017: signal is true;
	signal G4018: std_logic; attribute dont_touch of G4018: signal is true;
	signal G4019: std_logic; attribute dont_touch of G4019: signal is true;
	signal G4020: std_logic; attribute dont_touch of G4020: signal is true;
	signal G4021: std_logic; attribute dont_touch of G4021: signal is true;
	signal G4022: std_logic; attribute dont_touch of G4022: signal is true;
	signal G4023: std_logic; attribute dont_touch of G4023: signal is true;
	signal G4024: std_logic; attribute dont_touch of G4024: signal is true;
	signal G4025: std_logic; attribute dont_touch of G4025: signal is true;
	signal G4026: std_logic; attribute dont_touch of G4026: signal is true;
	signal G4027: std_logic; attribute dont_touch of G4027: signal is true;
	signal G4028: std_logic; attribute dont_touch of G4028: signal is true;
	signal G4029: std_logic; attribute dont_touch of G4029: signal is true;
	signal G4030: std_logic; attribute dont_touch of G4030: signal is true;
	signal G4031: std_logic; attribute dont_touch of G4031: signal is true;
	signal G4032: std_logic; attribute dont_touch of G4032: signal is true;
	signal G4033: std_logic; attribute dont_touch of G4033: signal is true;
	signal G4034: std_logic; attribute dont_touch of G4034: signal is true;
	signal G4035: std_logic; attribute dont_touch of G4035: signal is true;
	signal G4036: std_logic; attribute dont_touch of G4036: signal is true;
	signal G4037: std_logic; attribute dont_touch of G4037: signal is true;
	signal G4038: std_logic; attribute dont_touch of G4038: signal is true;
	signal G4041: std_logic; attribute dont_touch of G4041: signal is true;
	signal G4044: std_logic; attribute dont_touch of G4044: signal is true;
	signal G4047: std_logic; attribute dont_touch of G4047: signal is true;
	signal G4048: std_logic; attribute dont_touch of G4048: signal is true;
	signal G4049: std_logic; attribute dont_touch of G4049: signal is true;
	signal G4050: std_logic; attribute dont_touch of G4050: signal is true;
	signal G4051: std_logic; attribute dont_touch of G4051: signal is true;
	signal G4052: std_logic; attribute dont_touch of G4052: signal is true;
	signal G4053: std_logic; attribute dont_touch of G4053: signal is true;
	signal G4054: std_logic; attribute dont_touch of G4054: signal is true;
	signal G4055: std_logic; attribute dont_touch of G4055: signal is true;
	signal G4056: std_logic; attribute dont_touch of G4056: signal is true;
	signal G4057: std_logic; attribute dont_touch of G4057: signal is true;
	signal G4058: std_logic; attribute dont_touch of G4058: signal is true;
	signal G4059: std_logic; attribute dont_touch of G4059: signal is true;
	signal G4062: std_logic; attribute dont_touch of G4062: signal is true;
	signal G4065: std_logic; attribute dont_touch of G4065: signal is true;
	signal G4066: std_logic; attribute dont_touch of G4066: signal is true;
	signal G4067: std_logic; attribute dont_touch of G4067: signal is true;
	signal G4068: std_logic; attribute dont_touch of G4068: signal is true;
	signal G4069: std_logic; attribute dont_touch of G4069: signal is true;
	signal G4070: std_logic; attribute dont_touch of G4070: signal is true;
	signal G4071: std_logic; attribute dont_touch of G4071: signal is true;
	signal G4072: std_logic; attribute dont_touch of G4072: signal is true;
	signal G4073: std_logic; attribute dont_touch of G4073: signal is true;
	signal G4074: std_logic; attribute dont_touch of G4074: signal is true;
	signal G4075: std_logic; attribute dont_touch of G4075: signal is true;
	signal G4076: std_logic; attribute dont_touch of G4076: signal is true;
	signal G4077: std_logic; attribute dont_touch of G4077: signal is true;
	signal G4078: std_logic; attribute dont_touch of G4078: signal is true;
	signal G4079: std_logic; attribute dont_touch of G4079: signal is true;
	signal G4080: std_logic; attribute dont_touch of G4080: signal is true;
	signal G4081: std_logic; attribute dont_touch of G4081: signal is true;
	signal G4082: std_logic; attribute dont_touch of G4082: signal is true;
	signal G4083: std_logic; attribute dont_touch of G4083: signal is true;
	signal G4084: std_logic; attribute dont_touch of G4084: signal is true;
	signal G4085: std_logic; attribute dont_touch of G4085: signal is true;
	signal G4086: std_logic; attribute dont_touch of G4086: signal is true;
	signal G4087: std_logic; attribute dont_touch of G4087: signal is true;
	signal G4088: std_logic; attribute dont_touch of G4088: signal is true;
	signal G4089: std_logic; attribute dont_touch of G4089: signal is true;
	signal G4090: std_logic; attribute dont_touch of G4090: signal is true;
	signal G4091: std_logic; attribute dont_touch of G4091: signal is true;
	signal G4092: std_logic; attribute dont_touch of G4092: signal is true;
	signal G4093: std_logic; attribute dont_touch of G4093: signal is true;
	signal G4094: std_logic; attribute dont_touch of G4094: signal is true;
	signal G4095: std_logic; attribute dont_touch of G4095: signal is true;
	signal G4096: std_logic; attribute dont_touch of G4096: signal is true;
	signal G4097: std_logic; attribute dont_touch of G4097: signal is true;
	signal G4098: std_logic; attribute dont_touch of G4098: signal is true;
	signal G4099: std_logic; attribute dont_touch of G4099: signal is true;
	signal G4100: std_logic; attribute dont_touch of G4100: signal is true;
	signal G4101: std_logic; attribute dont_touch of G4101: signal is true;
	signal G4102: std_logic; attribute dont_touch of G4102: signal is true;
	signal G4103: std_logic; attribute dont_touch of G4103: signal is true;
	signal G4104: std_logic; attribute dont_touch of G4104: signal is true;
	signal G4105: std_logic; attribute dont_touch of G4105: signal is true;
	signal G4106: std_logic; attribute dont_touch of G4106: signal is true;
	signal G4107: std_logic; attribute dont_touch of G4107: signal is true;
	signal G4108: std_logic; attribute dont_touch of G4108: signal is true;
	signal G4109: std_logic; attribute dont_touch of G4109: signal is true;
	signal G4110: std_logic; attribute dont_touch of G4110: signal is true;
	signal G4111: std_logic; attribute dont_touch of G4111: signal is true;
	signal G4112: std_logic; attribute dont_touch of G4112: signal is true;
	signal G4113: std_logic; attribute dont_touch of G4113: signal is true;
	signal G4114: std_logic; attribute dont_touch of G4114: signal is true;
	signal G4115: std_logic; attribute dont_touch of G4115: signal is true;
	signal G4116: std_logic; attribute dont_touch of G4116: signal is true;
	signal G4117: std_logic; attribute dont_touch of G4117: signal is true;
	signal G4118: std_logic; attribute dont_touch of G4118: signal is true;
	signal G4119: std_logic; attribute dont_touch of G4119: signal is true;
	signal G4120: std_logic; attribute dont_touch of G4120: signal is true;
	signal G4121: std_logic; attribute dont_touch of G4121: signal is true;
	signal G4122: std_logic; attribute dont_touch of G4122: signal is true;
	signal G4123: std_logic; attribute dont_touch of G4123: signal is true;
	signal G4124: std_logic; attribute dont_touch of G4124: signal is true;
	signal G4125: std_logic; attribute dont_touch of G4125: signal is true;
	signal G4126: std_logic; attribute dont_touch of G4126: signal is true;
	signal G4127: std_logic; attribute dont_touch of G4127: signal is true;
	signal G4128: std_logic; attribute dont_touch of G4128: signal is true;
	signal G4129: std_logic; attribute dont_touch of G4129: signal is true;
	signal G4130: std_logic; attribute dont_touch of G4130: signal is true;
	signal G4131: std_logic; attribute dont_touch of G4131: signal is true;
	signal G4132: std_logic; attribute dont_touch of G4132: signal is true;
	signal G4133: std_logic; attribute dont_touch of G4133: signal is true;
	signal G4134: std_logic; attribute dont_touch of G4134: signal is true;
	signal G4135: std_logic; attribute dont_touch of G4135: signal is true;
	signal G4138: std_logic; attribute dont_touch of G4138: signal is true;
	signal G4139: std_logic; attribute dont_touch of G4139: signal is true;
	signal G4142: std_logic; attribute dont_touch of G4142: signal is true;
	signal G4145: std_logic; attribute dont_touch of G4145: signal is true;
	signal G4146: std_logic; attribute dont_touch of G4146: signal is true;
	signal G4147: std_logic; attribute dont_touch of G4147: signal is true;
	signal G4150: std_logic; attribute dont_touch of G4150: signal is true;
	signal G4153: std_logic; attribute dont_touch of G4153: signal is true;
	signal G4154: std_logic; attribute dont_touch of G4154: signal is true;
	signal G4155: std_logic; attribute dont_touch of G4155: signal is true;
	signal G4158: std_logic; attribute dont_touch of G4158: signal is true;
	signal G4159: std_logic; attribute dont_touch of G4159: signal is true;
	signal G4160: std_logic; attribute dont_touch of G4160: signal is true;
	signal G4163: std_logic; attribute dont_touch of G4163: signal is true;
	signal G4166: std_logic; attribute dont_touch of G4166: signal is true;
	signal G4167: std_logic; attribute dont_touch of G4167: signal is true;
	signal G4168: std_logic; attribute dont_touch of G4168: signal is true;
	signal G4169: std_logic; attribute dont_touch of G4169: signal is true;
	signal G4172: std_logic; attribute dont_touch of G4172: signal is true;
	signal G4175: std_logic; attribute dont_touch of G4175: signal is true;
	signal G4176: std_logic; attribute dont_touch of G4176: signal is true;
	signal G4179: std_logic; attribute dont_touch of G4179: signal is true;
	signal G4180: std_logic; attribute dont_touch of G4180: signal is true;
	signal G4181: std_logic; attribute dont_touch of G4181: signal is true;
	signal G4182: std_logic; attribute dont_touch of G4182: signal is true;
	signal G4185: std_logic; attribute dont_touch of G4185: signal is true;
	signal G4186: std_logic; attribute dont_touch of G4186: signal is true;
	signal G4187: std_logic; attribute dont_touch of G4187: signal is true;
	signal G4190: std_logic; attribute dont_touch of G4190: signal is true;
	signal G4191: std_logic; attribute dont_touch of G4191: signal is true;
	signal G4192: std_logic; attribute dont_touch of G4192: signal is true;
	signal G4193: std_logic; attribute dont_touch of G4193: signal is true;
	signal G4194: std_logic; attribute dont_touch of G4194: signal is true;
	signal G4195: std_logic; attribute dont_touch of G4195: signal is true;
	signal G4196: std_logic; attribute dont_touch of G4196: signal is true;
	signal G4197: std_logic; attribute dont_touch of G4197: signal is true;
	signal G4198: std_logic; attribute dont_touch of G4198: signal is true;
	signal G4199: std_logic; attribute dont_touch of G4199: signal is true;
	signal G4200: std_logic; attribute dont_touch of G4200: signal is true;
	signal G4201: std_logic; attribute dont_touch of G4201: signal is true;
	signal G4202: std_logic; attribute dont_touch of G4202: signal is true;
	signal G4216: std_logic; attribute dont_touch of G4216: signal is true;
	signal G4219: std_logic; attribute dont_touch of G4219: signal is true;
	signal G4220: std_logic; attribute dont_touch of G4220: signal is true;
	signal G4224: std_logic; attribute dont_touch of G4224: signal is true;
	signal G4225: std_logic; attribute dont_touch of G4225: signal is true;
	signal G4226: std_logic; attribute dont_touch of G4226: signal is true;
	signal G4227: std_logic; attribute dont_touch of G4227: signal is true;
	signal G4228: std_logic; attribute dont_touch of G4228: signal is true;
	signal G4229: std_logic; attribute dont_touch of G4229: signal is true;
	signal G4230: std_logic; attribute dont_touch of G4230: signal is true;
	signal G4231: std_logic; attribute dont_touch of G4231: signal is true;
	signal G4232: std_logic; attribute dont_touch of G4232: signal is true;
	signal G4235: std_logic; attribute dont_touch of G4235: signal is true;
	signal G4236: std_logic; attribute dont_touch of G4236: signal is true;
	signal G4237: std_logic; attribute dont_touch of G4237: signal is true;
	signal G4238: std_logic; attribute dont_touch of G4238: signal is true;
	signal G4239: std_logic; attribute dont_touch of G4239: signal is true;
	signal G4242: std_logic; attribute dont_touch of G4242: signal is true;
	signal G4243: std_logic; attribute dont_touch of G4243: signal is true;
	signal G4244: std_logic; attribute dont_touch of G4244: signal is true;
	signal G4245: std_logic; attribute dont_touch of G4245: signal is true;
	signal G4246: std_logic; attribute dont_touch of G4246: signal is true;
	signal G4249: std_logic; attribute dont_touch of G4249: signal is true;
	signal G4250: std_logic; attribute dont_touch of G4250: signal is true;
	signal G4251: std_logic; attribute dont_touch of G4251: signal is true;
	signal G4252: std_logic; attribute dont_touch of G4252: signal is true;
	signal G4253: std_logic; attribute dont_touch of G4253: signal is true;
	signal G4254: std_logic; attribute dont_touch of G4254: signal is true;
	signal G4255: std_logic; attribute dont_touch of G4255: signal is true;
	signal G4256: std_logic; attribute dont_touch of G4256: signal is true;
	signal G4257: std_logic; attribute dont_touch of G4257: signal is true;
	signal G4258: std_logic; attribute dont_touch of G4258: signal is true;
	signal G4259: std_logic; attribute dont_touch of G4259: signal is true;
	signal G4263: std_logic; attribute dont_touch of G4263: signal is true;
	signal G4264: std_logic; attribute dont_touch of G4264: signal is true;
	signal G4265: std_logic; attribute dont_touch of G4265: signal is true;
	signal G4266: std_logic; attribute dont_touch of G4266: signal is true;
	signal G4268: std_logic; attribute dont_touch of G4268: signal is true;
	signal G4269: std_logic; attribute dont_touch of G4269: signal is true;
	signal G4270: std_logic; attribute dont_touch of G4270: signal is true;
	signal G4271: std_logic; attribute dont_touch of G4271: signal is true;
	signal G4272: std_logic; attribute dont_touch of G4272: signal is true;
	signal G4273: std_logic; attribute dont_touch of G4273: signal is true;
	signal G4274: std_logic; attribute dont_touch of G4274: signal is true;
	signal G4275: std_logic; attribute dont_touch of G4275: signal is true;
	signal G4276: std_logic; attribute dont_touch of G4276: signal is true;
	signal G4279: std_logic; attribute dont_touch of G4279: signal is true;
	signal G4280: std_logic; attribute dont_touch of G4280: signal is true;
	signal G4281: std_logic; attribute dont_touch of G4281: signal is true;
	signal G4282: std_logic; attribute dont_touch of G4282: signal is true;
	signal G4283: std_logic; attribute dont_touch of G4283: signal is true;
	signal G4284: std_logic; attribute dont_touch of G4284: signal is true;
	signal G4285: std_logic; attribute dont_touch of G4285: signal is true;
	signal G4286: std_logic; attribute dont_touch of G4286: signal is true;
	signal G4287: std_logic; attribute dont_touch of G4287: signal is true;
	signal G4288: std_logic; attribute dont_touch of G4288: signal is true;
	signal G4294: std_logic; attribute dont_touch of G4294: signal is true;
	signal G4295: std_logic; attribute dont_touch of G4295: signal is true;
	signal G4296: std_logic; attribute dont_touch of G4296: signal is true;
	signal G4297: std_logic; attribute dont_touch of G4297: signal is true;
	signal G4298: std_logic; attribute dont_touch of G4298: signal is true;
	signal G4299: std_logic; attribute dont_touch of G4299: signal is true;
	signal G4300: std_logic; attribute dont_touch of G4300: signal is true;
	signal G4301: std_logic; attribute dont_touch of G4301: signal is true;
	signal G4302: std_logic; attribute dont_touch of G4302: signal is true;
	signal G4303: std_logic; attribute dont_touch of G4303: signal is true;
	signal G4304: std_logic; attribute dont_touch of G4304: signal is true;
	signal G4305: std_logic; attribute dont_touch of G4305: signal is true;
	signal G4306: std_logic; attribute dont_touch of G4306: signal is true;
	signal G4307: std_logic; attribute dont_touch of G4307: signal is true;
	signal G4308: std_logic; attribute dont_touch of G4308: signal is true;
	signal G4309: std_logic; attribute dont_touch of G4309: signal is true;
	signal G4310: std_logic; attribute dont_touch of G4310: signal is true;
	signal G4311: std_logic; attribute dont_touch of G4311: signal is true;
	signal G4312: std_logic; attribute dont_touch of G4312: signal is true;
	signal G4313: std_logic; attribute dont_touch of G4313: signal is true;
	signal G4314: std_logic; attribute dont_touch of G4314: signal is true;
	signal G4315: std_logic; attribute dont_touch of G4315: signal is true;
	signal G4317: std_logic; attribute dont_touch of G4317: signal is true;
	signal G4318: std_logic; attribute dont_touch of G4318: signal is true;
	signal G4319: std_logic; attribute dont_touch of G4319: signal is true;
	signal G4320: std_logic; attribute dont_touch of G4320: signal is true;
	signal G4327: std_logic; attribute dont_touch of G4327: signal is true;
	signal G4328: std_logic; attribute dont_touch of G4328: signal is true;
	signal G4332: std_logic; attribute dont_touch of G4332: signal is true;
	signal G4333: std_logic; attribute dont_touch of G4333: signal is true;
	signal G4334: std_logic; attribute dont_touch of G4334: signal is true;
	signal G4335: std_logic; attribute dont_touch of G4335: signal is true;
	signal G4341: std_logic; attribute dont_touch of G4341: signal is true;
	signal G4342: std_logic; attribute dont_touch of G4342: signal is true;
	signal G4343: std_logic; attribute dont_touch of G4343: signal is true;
	signal G4344: std_logic; attribute dont_touch of G4344: signal is true;
	signal G4349: std_logic; attribute dont_touch of G4349: signal is true;
	signal G4350: std_logic; attribute dont_touch of G4350: signal is true;
	signal G4351: std_logic; attribute dont_touch of G4351: signal is true;
	signal G4352: std_logic; attribute dont_touch of G4352: signal is true;
	signal G4353: std_logic; attribute dont_touch of G4353: signal is true;
	signal G4354: std_logic; attribute dont_touch of G4354: signal is true;
	signal G4355: std_logic; attribute dont_touch of G4355: signal is true;
	signal G4356: std_logic; attribute dont_touch of G4356: signal is true;
	signal G4357: std_logic; attribute dont_touch of G4357: signal is true;
	signal G4358: std_logic; attribute dont_touch of G4358: signal is true;
	signal G4359: std_logic; attribute dont_touch of G4359: signal is true;
	signal G4360: std_logic; attribute dont_touch of G4360: signal is true;
	signal G4361: std_logic; attribute dont_touch of G4361: signal is true;
	signal G4362: std_logic; attribute dont_touch of G4362: signal is true;
	signal G4363: std_logic; attribute dont_touch of G4363: signal is true;
	signal G4364: std_logic; attribute dont_touch of G4364: signal is true;
	signal G4365: std_logic; attribute dont_touch of G4365: signal is true;
	signal G4366: std_logic; attribute dont_touch of G4366: signal is true;
	signal G4367: std_logic; attribute dont_touch of G4367: signal is true;
	signal G4368: std_logic; attribute dont_touch of G4368: signal is true;
	signal G4369: std_logic; attribute dont_touch of G4369: signal is true;
	signal G4374: std_logic; attribute dont_touch of G4374: signal is true;
	signal G4375: std_logic; attribute dont_touch of G4375: signal is true;
	signal G4376: std_logic; attribute dont_touch of G4376: signal is true;
	signal G4377: std_logic; attribute dont_touch of G4377: signal is true;
	signal G4378: std_logic; attribute dont_touch of G4378: signal is true;
	signal G4379: std_logic; attribute dont_touch of G4379: signal is true;
	signal G4380: std_logic; attribute dont_touch of G4380: signal is true;
	signal G4381: std_logic; attribute dont_touch of G4381: signal is true;
	signal G4382: std_logic; attribute dont_touch of G4382: signal is true;
	signal G4383: std_logic; attribute dont_touch of G4383: signal is true;
	signal G4384: std_logic; attribute dont_touch of G4384: signal is true;
	signal G4385: std_logic; attribute dont_touch of G4385: signal is true;
	signal G4386: std_logic; attribute dont_touch of G4386: signal is true;
	signal G4387: std_logic; attribute dont_touch of G4387: signal is true;
	signal G4388: std_logic; attribute dont_touch of G4388: signal is true;
	signal G4389: std_logic; attribute dont_touch of G4389: signal is true;
	signal G4390: std_logic; attribute dont_touch of G4390: signal is true;
	signal G4391: std_logic; attribute dont_touch of G4391: signal is true;
	signal G4392: std_logic; attribute dont_touch of G4392: signal is true;
	signal G4393: std_logic; attribute dont_touch of G4393: signal is true;
	signal G4394: std_logic; attribute dont_touch of G4394: signal is true;
	signal G4395: std_logic; attribute dont_touch of G4395: signal is true;
	signal G4396: std_logic; attribute dont_touch of G4396: signal is true;
	signal G4397: std_logic; attribute dont_touch of G4397: signal is true;
	signal G4398: std_logic; attribute dont_touch of G4398: signal is true;
	signal G4399: std_logic; attribute dont_touch of G4399: signal is true;
	signal G4400: std_logic; attribute dont_touch of G4400: signal is true;
	signal G4403: std_logic; attribute dont_touch of G4403: signal is true;
	signal G4407: std_logic; attribute dont_touch of G4407: signal is true;
	signal G4408: std_logic; attribute dont_touch of G4408: signal is true;
	signal G4409: std_logic; attribute dont_touch of G4409: signal is true;
	signal G4410: std_logic; attribute dont_touch of G4410: signal is true;
	signal G4411: std_logic; attribute dont_touch of G4411: signal is true;
	signal G4412: std_logic; attribute dont_touch of G4412: signal is true;
	signal G4413: std_logic; attribute dont_touch of G4413: signal is true;
	signal G4414: std_logic; attribute dont_touch of G4414: signal is true;
	signal G4417: std_logic; attribute dont_touch of G4417: signal is true;
	signal G4420: std_logic; attribute dont_touch of G4420: signal is true;
	signal G4421: std_logic; attribute dont_touch of G4421: signal is true;
	signal G4422: std_logic; attribute dont_touch of G4422: signal is true;
	signal G4423: std_logic; attribute dont_touch of G4423: signal is true;
	signal G4424: std_logic; attribute dont_touch of G4424: signal is true;
	signal G4425: std_logic; attribute dont_touch of G4425: signal is true;
	signal G4426: std_logic; attribute dont_touch of G4426: signal is true;
	signal G4427: std_logic; attribute dont_touch of G4427: signal is true;
	signal G4430: std_logic; attribute dont_touch of G4430: signal is true;
	signal G4433: std_logic; attribute dont_touch of G4433: signal is true;
	signal G4434: std_logic; attribute dont_touch of G4434: signal is true;
	signal G4435: std_logic; attribute dont_touch of G4435: signal is true;
	signal G4436: std_logic; attribute dont_touch of G4436: signal is true;
	signal G4437: std_logic; attribute dont_touch of G4437: signal is true;
	signal G4438: std_logic; attribute dont_touch of G4438: signal is true;
	signal G4443: std_logic; attribute dont_touch of G4443: signal is true;
	signal G4444: std_logic; attribute dont_touch of G4444: signal is true;
	signal G4445: std_logic; attribute dont_touch of G4445: signal is true;
	signal G4448: std_logic; attribute dont_touch of G4448: signal is true;
	signal G4451: std_logic; attribute dont_touch of G4451: signal is true;
	signal G4452: std_logic; attribute dont_touch of G4452: signal is true;
	signal G4453: std_logic; attribute dont_touch of G4453: signal is true;
	signal G4454: std_logic; attribute dont_touch of G4454: signal is true;
	signal G4455: std_logic; attribute dont_touch of G4455: signal is true;
	signal G4456: std_logic; attribute dont_touch of G4456: signal is true;
	signal G4457: std_logic; attribute dont_touch of G4457: signal is true;
	signal G4462: std_logic; attribute dont_touch of G4462: signal is true;
	signal G4463: std_logic; attribute dont_touch of G4463: signal is true;
	signal G4464: std_logic; attribute dont_touch of G4464: signal is true;
	signal G4465: std_logic; attribute dont_touch of G4465: signal is true;
	signal G4466: std_logic; attribute dont_touch of G4466: signal is true;
	signal G4469: std_logic; attribute dont_touch of G4469: signal is true;
	signal G4472: std_logic; attribute dont_touch of G4472: signal is true;
	signal G4473: std_logic; attribute dont_touch of G4473: signal is true;
	signal G4474: std_logic; attribute dont_touch of G4474: signal is true;
	signal G4475: std_logic; attribute dont_touch of G4475: signal is true;
	signal G4476: std_logic; attribute dont_touch of G4476: signal is true;
	signal G4477: std_logic; attribute dont_touch of G4477: signal is true;
	signal G4482: std_logic; attribute dont_touch of G4482: signal is true;
	signal G4483: std_logic; attribute dont_touch of G4483: signal is true;
	signal G4486: std_logic; attribute dont_touch of G4486: signal is true;
	signal G4489: std_logic; attribute dont_touch of G4489: signal is true;
	signal G4490: std_logic; attribute dont_touch of G4490: signal is true;
	signal G4491: std_logic; attribute dont_touch of G4491: signal is true;
	signal G4492: std_logic; attribute dont_touch of G4492: signal is true;
	signal G4493: std_logic; attribute dont_touch of G4493: signal is true;
	signal G4494: std_logic; attribute dont_touch of G4494: signal is true;
	signal G4497: std_logic; attribute dont_touch of G4497: signal is true;
	signal G4500: std_logic; attribute dont_touch of G4500: signal is true;
	signal G4501: std_logic; attribute dont_touch of G4501: signal is true;
	signal G4502: std_logic; attribute dont_touch of G4502: signal is true;
	signal G4503: std_logic; attribute dont_touch of G4503: signal is true;
	signal G4504: std_logic; attribute dont_touch of G4504: signal is true;
	signal G4507: std_logic; attribute dont_touch of G4507: signal is true;
	signal G4510: std_logic; attribute dont_touch of G4510: signal is true;
	signal G4511: std_logic; attribute dont_touch of G4511: signal is true;
	signal G4512: std_logic; attribute dont_touch of G4512: signal is true;
	signal G4513: std_logic; attribute dont_touch of G4513: signal is true;
	signal G4514: std_logic; attribute dont_touch of G4514: signal is true;
	signal G4517: std_logic; attribute dont_touch of G4517: signal is true;
	signal G4521: std_logic; attribute dont_touch of G4521: signal is true;
	signal G4522: std_logic; attribute dont_touch of G4522: signal is true;
	signal G4523: std_logic; attribute dont_touch of G4523: signal is true;
	signal G4524: std_logic; attribute dont_touch of G4524: signal is true;
	signal G4525: std_logic; attribute dont_touch of G4525: signal is true;
	signal G4526: std_logic; attribute dont_touch of G4526: signal is true;
	signal G4527: std_logic; attribute dont_touch of G4527: signal is true;
	signal G4528: std_logic; attribute dont_touch of G4528: signal is true;
	signal G4529: std_logic; attribute dont_touch of G4529: signal is true;
	signal G4532: std_logic; attribute dont_touch of G4532: signal is true;
	signal G4535: std_logic; attribute dont_touch of G4535: signal is true;
	signal G4536: std_logic; attribute dont_touch of G4536: signal is true;
	signal G4537: std_logic; attribute dont_touch of G4537: signal is true;
	signal G4538: std_logic; attribute dont_touch of G4538: signal is true;
	signal G4539: std_logic; attribute dont_touch of G4539: signal is true;
	signal G4540: std_logic; attribute dont_touch of G4540: signal is true;
	signal G4541: std_logic; attribute dont_touch of G4541: signal is true;
	signal G4542: std_logic; attribute dont_touch of G4542: signal is true;
	signal G4543: std_logic; attribute dont_touch of G4543: signal is true;
	signal G4544: std_logic; attribute dont_touch of G4544: signal is true;
	signal G4545: std_logic; attribute dont_touch of G4545: signal is true;
	signal G4546: std_logic; attribute dont_touch of G4546: signal is true;
	signal G4547: std_logic; attribute dont_touch of G4547: signal is true;
	signal G4548: std_logic; attribute dont_touch of G4548: signal is true;
	signal G4549: std_logic; attribute dont_touch of G4549: signal is true;
	signal G4552: std_logic; attribute dont_touch of G4552: signal is true;
	signal G4553: std_logic; attribute dont_touch of G4553: signal is true;
	signal G4554: std_logic; attribute dont_touch of G4554: signal is true;
	signal G4555: std_logic; attribute dont_touch of G4555: signal is true;
	signal G4556: std_logic; attribute dont_touch of G4556: signal is true;
	signal G4557: std_logic; attribute dont_touch of G4557: signal is true;
	signal G4558: std_logic; attribute dont_touch of G4558: signal is true;
	signal G4559: std_logic; attribute dont_touch of G4559: signal is true;
	signal G4560: std_logic; attribute dont_touch of G4560: signal is true;
	signal G4561: std_logic; attribute dont_touch of G4561: signal is true;
	signal G4562: std_logic; attribute dont_touch of G4562: signal is true;
	signal G4563: std_logic; attribute dont_touch of G4563: signal is true;
	signal G4564: std_logic; attribute dont_touch of G4564: signal is true;
	signal G4565: std_logic; attribute dont_touch of G4565: signal is true;
	signal G4566: std_logic; attribute dont_touch of G4566: signal is true;
	signal G4567: std_logic; attribute dont_touch of G4567: signal is true;
	signal G4568: std_logic; attribute dont_touch of G4568: signal is true;
	signal G4569: std_logic; attribute dont_touch of G4569: signal is true;
	signal G4570: std_logic; attribute dont_touch of G4570: signal is true;
	signal G4571: std_logic; attribute dont_touch of G4571: signal is true;
	signal G4572: std_logic; attribute dont_touch of G4572: signal is true;
	signal G4573: std_logic; attribute dont_touch of G4573: signal is true;
	signal G4574: std_logic; attribute dont_touch of G4574: signal is true;
	signal G4575: std_logic; attribute dont_touch of G4575: signal is true;
	signal G4576: std_logic; attribute dont_touch of G4576: signal is true;
	signal G4577: std_logic; attribute dont_touch of G4577: signal is true;
	signal G4578: std_logic; attribute dont_touch of G4578: signal is true;
	signal G4579: std_logic; attribute dont_touch of G4579: signal is true;
	signal G4580: std_logic; attribute dont_touch of G4580: signal is true;
	signal G4581: std_logic; attribute dont_touch of G4581: signal is true;
	signal G4582: std_logic; attribute dont_touch of G4582: signal is true;
	signal G4583: std_logic; attribute dont_touch of G4583: signal is true;
	signal G4584: std_logic; attribute dont_touch of G4584: signal is true;
	signal G4585: std_logic; attribute dont_touch of G4585: signal is true;
	signal G4586: std_logic; attribute dont_touch of G4586: signal is true;
	signal G4587: std_logic; attribute dont_touch of G4587: signal is true;
	signal G4588: std_logic; attribute dont_touch of G4588: signal is true;
	signal G4589: std_logic; attribute dont_touch of G4589: signal is true;
	signal G4590: std_logic; attribute dont_touch of G4590: signal is true;
	signal G4591: std_logic; attribute dont_touch of G4591: signal is true;
	signal G4592: std_logic; attribute dont_touch of G4592: signal is true;
	signal G4593: std_logic; attribute dont_touch of G4593: signal is true;
	signal G4594: std_logic; attribute dont_touch of G4594: signal is true;
	signal G4595: std_logic; attribute dont_touch of G4595: signal is true;
	signal G4596: std_logic; attribute dont_touch of G4596: signal is true;
	signal G4597: std_logic; attribute dont_touch of G4597: signal is true;
	signal G4598: std_logic; attribute dont_touch of G4598: signal is true;
	signal G4599: std_logic; attribute dont_touch of G4599: signal is true;
	signal G4600: std_logic; attribute dont_touch of G4600: signal is true;
	signal G4601: std_logic; attribute dont_touch of G4601: signal is true;
	signal G4602: std_logic; attribute dont_touch of G4602: signal is true;
	signal G4603: std_logic; attribute dont_touch of G4603: signal is true;
	signal G4604: std_logic; attribute dont_touch of G4604: signal is true;
	signal G4605: std_logic; attribute dont_touch of G4605: signal is true;
	signal G4606: std_logic; attribute dont_touch of G4606: signal is true;
	signal G4607: std_logic; attribute dont_touch of G4607: signal is true;
	signal G4608: std_logic; attribute dont_touch of G4608: signal is true;
	signal G4609: std_logic; attribute dont_touch of G4609: signal is true;
	signal G4610: std_logic; attribute dont_touch of G4610: signal is true;
	signal G4611: std_logic; attribute dont_touch of G4611: signal is true;
	signal G4612: std_logic; attribute dont_touch of G4612: signal is true;
	signal G4613: std_logic; attribute dont_touch of G4613: signal is true;
	signal G4614: std_logic; attribute dont_touch of G4614: signal is true;
	signal G4615: std_logic; attribute dont_touch of G4615: signal is true;
	signal G4616: std_logic; attribute dont_touch of G4616: signal is true;
	signal G4617: std_logic; attribute dont_touch of G4617: signal is true;
	signal G4618: std_logic; attribute dont_touch of G4618: signal is true;
	signal G4619: std_logic; attribute dont_touch of G4619: signal is true;
	signal G4620: std_logic; attribute dont_touch of G4620: signal is true;
	signal G4621: std_logic; attribute dont_touch of G4621: signal is true;
	signal G4622: std_logic; attribute dont_touch of G4622: signal is true;
	signal G4623: std_logic; attribute dont_touch of G4623: signal is true;
	signal G4624: std_logic; attribute dont_touch of G4624: signal is true;
	signal G4625: std_logic; attribute dont_touch of G4625: signal is true;
	signal G4626: std_logic; attribute dont_touch of G4626: signal is true;
	signal G4627: std_logic; attribute dont_touch of G4627: signal is true;
	signal G4628: std_logic; attribute dont_touch of G4628: signal is true;
	signal G4629: std_logic; attribute dont_touch of G4629: signal is true;
	signal G4630: std_logic; attribute dont_touch of G4630: signal is true;
	signal G4631: std_logic; attribute dont_touch of G4631: signal is true;
	signal G4632: std_logic; attribute dont_touch of G4632: signal is true;
	signal G4633: std_logic; attribute dont_touch of G4633: signal is true;
	signal G4634: std_logic; attribute dont_touch of G4634: signal is true;
	signal G4635: std_logic; attribute dont_touch of G4635: signal is true;
	signal G4636: std_logic; attribute dont_touch of G4636: signal is true;
	signal G4637: std_logic; attribute dont_touch of G4637: signal is true;
	signal G4638: std_logic; attribute dont_touch of G4638: signal is true;
	signal G4639: std_logic; attribute dont_touch of G4639: signal is true;
	signal G4640: std_logic; attribute dont_touch of G4640: signal is true;
	signal G4641: std_logic; attribute dont_touch of G4641: signal is true;
	signal G4642: std_logic; attribute dont_touch of G4642: signal is true;
	signal G4643: std_logic; attribute dont_touch of G4643: signal is true;
	signal G4644: std_logic; attribute dont_touch of G4644: signal is true;
	signal G4645: std_logic; attribute dont_touch of G4645: signal is true;
	signal G4646: std_logic; attribute dont_touch of G4646: signal is true;
	signal G4647: std_logic; attribute dont_touch of G4647: signal is true;
	signal G4648: std_logic; attribute dont_touch of G4648: signal is true;
	signal G4649: std_logic; attribute dont_touch of G4649: signal is true;
	signal G4650: std_logic; attribute dont_touch of G4650: signal is true;
	signal G4651: std_logic; attribute dont_touch of G4651: signal is true;
	signal G4652: std_logic; attribute dont_touch of G4652: signal is true;
	signal G4653: std_logic; attribute dont_touch of G4653: signal is true;
	signal G4654: std_logic; attribute dont_touch of G4654: signal is true;
	signal G4656: std_logic; attribute dont_touch of G4656: signal is true;
	signal G4658: std_logic; attribute dont_touch of G4658: signal is true;
	signal G4659: std_logic; attribute dont_touch of G4659: signal is true;
	signal G4662: std_logic; attribute dont_touch of G4662: signal is true;
	signal G4665: std_logic; attribute dont_touch of G4665: signal is true;
	signal G4666: std_logic; attribute dont_touch of G4666: signal is true;
	signal G4667: std_logic; attribute dont_touch of G4667: signal is true;
	signal G4668: std_logic; attribute dont_touch of G4668: signal is true;
	signal G4669: std_logic; attribute dont_touch of G4669: signal is true;
	signal G4670: std_logic; attribute dont_touch of G4670: signal is true;
	signal G4673: std_logic; attribute dont_touch of G4673: signal is true;
	signal G4676: std_logic; attribute dont_touch of G4676: signal is true;
	signal G4677: std_logic; attribute dont_touch of G4677: signal is true;
	signal G4678: std_logic; attribute dont_touch of G4678: signal is true;
	signal G4679: std_logic; attribute dont_touch of G4679: signal is true;
	signal G4680: std_logic; attribute dont_touch of G4680: signal is true;
	signal G4681: std_logic; attribute dont_touch of G4681: signal is true;
	signal G4684: std_logic; attribute dont_touch of G4684: signal is true;
	signal G4685: std_logic; attribute dont_touch of G4685: signal is true;
	signal G4686: std_logic; attribute dont_touch of G4686: signal is true;
	signal G4687: std_logic; attribute dont_touch of G4687: signal is true;
	signal G4688: std_logic; attribute dont_touch of G4688: signal is true;
	signal G4689: std_logic; attribute dont_touch of G4689: signal is true;
	signal G4690: std_logic; attribute dont_touch of G4690: signal is true;
	signal G4691: std_logic; attribute dont_touch of G4691: signal is true;
	signal G4692: std_logic; attribute dont_touch of G4692: signal is true;
	signal G4693: std_logic; attribute dont_touch of G4693: signal is true;
	signal G4694: std_logic; attribute dont_touch of G4694: signal is true;
	signal G4695: std_logic; attribute dont_touch of G4695: signal is true;
	signal G4696: std_logic; attribute dont_touch of G4696: signal is true;
	signal G4697: std_logic; attribute dont_touch of G4697: signal is true;
	signal G4698: std_logic; attribute dont_touch of G4698: signal is true;
	signal G4699: std_logic; attribute dont_touch of G4699: signal is true;
	signal G4700: std_logic; attribute dont_touch of G4700: signal is true;
	signal G4701: std_logic; attribute dont_touch of G4701: signal is true;
	signal G4702: std_logic; attribute dont_touch of G4702: signal is true;
	signal G4703: std_logic; attribute dont_touch of G4703: signal is true;
	signal G4704: std_logic; attribute dont_touch of G4704: signal is true;
	signal G4705: std_logic; attribute dont_touch of G4705: signal is true;
	signal G4706: std_logic; attribute dont_touch of G4706: signal is true;
	signal G4707: std_logic; attribute dont_touch of G4707: signal is true;
	signal G4710: std_logic; attribute dont_touch of G4710: signal is true;
	signal G4711: std_logic; attribute dont_touch of G4711: signal is true;
	signal G4712: std_logic; attribute dont_touch of G4712: signal is true;
	signal G4713: std_logic; attribute dont_touch of G4713: signal is true;
	signal G4714: std_logic; attribute dont_touch of G4714: signal is true;
	signal G4718: std_logic; attribute dont_touch of G4718: signal is true;
	signal G4719: std_logic; attribute dont_touch of G4719: signal is true;
	signal G4720: std_logic; attribute dont_touch of G4720: signal is true;
	signal G4721: std_logic; attribute dont_touch of G4721: signal is true;
	signal G4724: std_logic; attribute dont_touch of G4724: signal is true;
	signal G4727: std_logic; attribute dont_touch of G4727: signal is true;
	signal G4728: std_logic; attribute dont_touch of G4728: signal is true;
	signal G4729: std_logic; attribute dont_touch of G4729: signal is true;
	signal G4732: std_logic; attribute dont_touch of G4732: signal is true;
	signal G4733: std_logic; attribute dont_touch of G4733: signal is true;
	signal G4734: std_logic; attribute dont_touch of G4734: signal is true;
	signal G4735: std_logic; attribute dont_touch of G4735: signal is true;
	signal G4736: std_logic; attribute dont_touch of G4736: signal is true;
	signal G4737: std_logic; attribute dont_touch of G4737: signal is true;
	signal G4738: std_logic; attribute dont_touch of G4738: signal is true;
	signal G4739: std_logic; attribute dont_touch of G4739: signal is true;
	signal G4740: std_logic; attribute dont_touch of G4740: signal is true;
	signal G4741: std_logic; attribute dont_touch of G4741: signal is true;
	signal G4742: std_logic; attribute dont_touch of G4742: signal is true;
	signal G4743: std_logic; attribute dont_touch of G4743: signal is true;
	signal G4744: std_logic; attribute dont_touch of G4744: signal is true;
	signal G4745: std_logic; attribute dont_touch of G4745: signal is true;
	signal G4746: std_logic; attribute dont_touch of G4746: signal is true;
	signal G4747: std_logic; attribute dont_touch of G4747: signal is true;
	signal G4748: std_logic; attribute dont_touch of G4748: signal is true;
	signal G4776: std_logic; attribute dont_touch of G4776: signal is true;
	signal G4777: std_logic; attribute dont_touch of G4777: signal is true;
	signal G4778: std_logic; attribute dont_touch of G4778: signal is true;
	signal G4779: std_logic; attribute dont_touch of G4779: signal is true;
	signal G4780: std_logic; attribute dont_touch of G4780: signal is true;
	signal G4781: std_logic; attribute dont_touch of G4781: signal is true;
	signal G4782: std_logic; attribute dont_touch of G4782: signal is true;
	signal G4783: std_logic; attribute dont_touch of G4783: signal is true;
	signal G4784: std_logic; attribute dont_touch of G4784: signal is true;
	signal G4785: std_logic; attribute dont_touch of G4785: signal is true;
	signal G4786: std_logic; attribute dont_touch of G4786: signal is true;
	signal G4787: std_logic; attribute dont_touch of G4787: signal is true;
	signal G4788: std_logic; attribute dont_touch of G4788: signal is true;
	signal G4789: std_logic; attribute dont_touch of G4789: signal is true;
	signal G4790: std_logic; attribute dont_touch of G4790: signal is true;
	signal G4791: std_logic; attribute dont_touch of G4791: signal is true;
	signal G4792: std_logic; attribute dont_touch of G4792: signal is true;
	signal G4793: std_logic; attribute dont_touch of G4793: signal is true;
	signal G4794: std_logic; attribute dont_touch of G4794: signal is true;
	signal G4795: std_logic; attribute dont_touch of G4795: signal is true;
	signal G4796: std_logic; attribute dont_touch of G4796: signal is true;
	signal G4797: std_logic; attribute dont_touch of G4797: signal is true;
	signal G4798: std_logic; attribute dont_touch of G4798: signal is true;
	signal G4799: std_logic; attribute dont_touch of G4799: signal is true;
	signal G4800: std_logic; attribute dont_touch of G4800: signal is true;
	signal G4801: std_logic; attribute dont_touch of G4801: signal is true;
	signal G4802: std_logic; attribute dont_touch of G4802: signal is true;
	signal G4803: std_logic; attribute dont_touch of G4803: signal is true;
	signal G4804: std_logic; attribute dont_touch of G4804: signal is true;
	signal G4805: std_logic; attribute dont_touch of G4805: signal is true;
	signal G4806: std_logic; attribute dont_touch of G4806: signal is true;
	signal G4807: std_logic; attribute dont_touch of G4807: signal is true;
	signal G4808: std_logic; attribute dont_touch of G4808: signal is true;
	signal G4809: std_logic; attribute dont_touch of G4809: signal is true;
	signal G4810: std_logic; attribute dont_touch of G4810: signal is true;
	signal G4811: std_logic; attribute dont_touch of G4811: signal is true;
	signal G4812: std_logic; attribute dont_touch of G4812: signal is true;
	signal G4813: std_logic; attribute dont_touch of G4813: signal is true;
	signal G4814: std_logic; attribute dont_touch of G4814: signal is true;
	signal G4819: std_logic; attribute dont_touch of G4819: signal is true;
	signal G4820: std_logic; attribute dont_touch of G4820: signal is true;
	signal G4821: std_logic; attribute dont_touch of G4821: signal is true;
	signal G4822: std_logic; attribute dont_touch of G4822: signal is true;
	signal G4823: std_logic; attribute dont_touch of G4823: signal is true;
	signal G4824: std_logic; attribute dont_touch of G4824: signal is true;
	signal G4825: std_logic; attribute dont_touch of G4825: signal is true;
	signal G4826: std_logic; attribute dont_touch of G4826: signal is true;
	signal G4829: std_logic; attribute dont_touch of G4829: signal is true;
	signal G4830: std_logic; attribute dont_touch of G4830: signal is true;
	signal G4831: std_logic; attribute dont_touch of G4831: signal is true;
	signal G4832: std_logic; attribute dont_touch of G4832: signal is true;
	signal G4835: std_logic; attribute dont_touch of G4835: signal is true;
	signal G4836: std_logic; attribute dont_touch of G4836: signal is true;
	signal G4837: std_logic; attribute dont_touch of G4837: signal is true;
	signal G4838: std_logic; attribute dont_touch of G4838: signal is true;
	signal G4839: std_logic; attribute dont_touch of G4839: signal is true;
	signal G4840: std_logic; attribute dont_touch of G4840: signal is true;
	signal G4841: std_logic; attribute dont_touch of G4841: signal is true;
	signal G4867: std_logic; attribute dont_touch of G4867: signal is true;
	signal G4868: std_logic; attribute dont_touch of G4868: signal is true;
	signal G4869: std_logic; attribute dont_touch of G4869: signal is true;
	signal G4870: std_logic; attribute dont_touch of G4870: signal is true;
	signal G4871: std_logic; attribute dont_touch of G4871: signal is true;
	signal G4872: std_logic; attribute dont_touch of G4872: signal is true;
	signal G4873: std_logic; attribute dont_touch of G4873: signal is true;
	signal G4876: std_logic; attribute dont_touch of G4876: signal is true;
	signal G4877: std_logic; attribute dont_touch of G4877: signal is true;
	signal G4878: std_logic; attribute dont_touch of G4878: signal is true;
	signal G4879: std_logic; attribute dont_touch of G4879: signal is true;
	signal G4880: std_logic; attribute dont_touch of G4880: signal is true;
	signal G4881: std_logic; attribute dont_touch of G4881: signal is true;
	signal G4882: std_logic; attribute dont_touch of G4882: signal is true;
	signal G4883: std_logic; attribute dont_touch of G4883: signal is true;
	signal G4884: std_logic; attribute dont_touch of G4884: signal is true;
	signal G4885: std_logic; attribute dont_touch of G4885: signal is true;
	signal G4886: std_logic; attribute dont_touch of G4886: signal is true;
	signal G4887: std_logic; attribute dont_touch of G4887: signal is true;
	signal G4888: std_logic; attribute dont_touch of G4888: signal is true;
	signal G4889: std_logic; attribute dont_touch of G4889: signal is true;
	signal G4890: std_logic; attribute dont_touch of G4890: signal is true;
	signal G4891: std_logic; attribute dont_touch of G4891: signal is true;
	signal G4892: std_logic; attribute dont_touch of G4892: signal is true;
	signal G4893: std_logic; attribute dont_touch of G4893: signal is true;
	signal G4894: std_logic; attribute dont_touch of G4894: signal is true;
	signal G4895: std_logic; attribute dont_touch of G4895: signal is true;
	signal G4898: std_logic; attribute dont_touch of G4898: signal is true;
	signal G4899: std_logic; attribute dont_touch of G4899: signal is true;
	signal G4900: std_logic; attribute dont_touch of G4900: signal is true;
	signal G4901: std_logic; attribute dont_touch of G4901: signal is true;
	signal G4902: std_logic; attribute dont_touch of G4902: signal is true;
	signal G4903: std_logic; attribute dont_touch of G4903: signal is true;
	signal G4904: std_logic; attribute dont_touch of G4904: signal is true;
	signal G4905: std_logic; attribute dont_touch of G4905: signal is true;
	signal G4906: std_logic; attribute dont_touch of G4906: signal is true;
	signal G4907: std_logic; attribute dont_touch of G4907: signal is true;
	signal G4908: std_logic; attribute dont_touch of G4908: signal is true;
	signal G4909: std_logic; attribute dont_touch of G4909: signal is true;
	signal G4910: std_logic; attribute dont_touch of G4910: signal is true;
	signal G4911: std_logic; attribute dont_touch of G4911: signal is true;
	signal G4912: std_logic; attribute dont_touch of G4912: signal is true;
	signal G4913: std_logic; attribute dont_touch of G4913: signal is true;
	signal G4914: std_logic; attribute dont_touch of G4914: signal is true;
	signal G4915: std_logic; attribute dont_touch of G4915: signal is true;
	signal G4916: std_logic; attribute dont_touch of G4916: signal is true;
	signal G4917: std_logic; attribute dont_touch of G4917: signal is true;
	signal G4918: std_logic; attribute dont_touch of G4918: signal is true;
	signal G4919: std_logic; attribute dont_touch of G4919: signal is true;
	signal G4920: std_logic; attribute dont_touch of G4920: signal is true;
	signal G4921: std_logic; attribute dont_touch of G4921: signal is true;
	signal G4922: std_logic; attribute dont_touch of G4922: signal is true;
	signal G4923: std_logic; attribute dont_touch of G4923: signal is true;
	signal G4924: std_logic; attribute dont_touch of G4924: signal is true;
	signal G4925: std_logic; attribute dont_touch of G4925: signal is true;
	signal G4926: std_logic; attribute dont_touch of G4926: signal is true;
	signal G4927: std_logic; attribute dont_touch of G4927: signal is true;
	signal G4928: std_logic; attribute dont_touch of G4928: signal is true;
	signal G4929: std_logic; attribute dont_touch of G4929: signal is true;
	signal G4930: std_logic; attribute dont_touch of G4930: signal is true;
	signal G4931: std_logic; attribute dont_touch of G4931: signal is true;
	signal G4932: std_logic; attribute dont_touch of G4932: signal is true;
	signal G4933: std_logic; attribute dont_touch of G4933: signal is true;
	signal G4934: std_logic; attribute dont_touch of G4934: signal is true;
	signal G4935: std_logic; attribute dont_touch of G4935: signal is true;
	signal G4936: std_logic; attribute dont_touch of G4936: signal is true;
	signal G4937: std_logic; attribute dont_touch of G4937: signal is true;
	signal G4938: std_logic; attribute dont_touch of G4938: signal is true;
	signal G4954: std_logic; attribute dont_touch of G4954: signal is true;
	signal G4955: std_logic; attribute dont_touch of G4955: signal is true;
	signal G4956: std_logic; attribute dont_touch of G4956: signal is true;
	signal G4957: std_logic; attribute dont_touch of G4957: signal is true;
	signal G4958: std_logic; attribute dont_touch of G4958: signal is true;
	signal G4959: std_logic; attribute dont_touch of G4959: signal is true;
	signal G4960: std_logic; attribute dont_touch of G4960: signal is true;
	signal G4961: std_logic; attribute dont_touch of G4961: signal is true;
	signal G4962: std_logic; attribute dont_touch of G4962: signal is true;
	signal G4963: std_logic; attribute dont_touch of G4963: signal is true;
	signal G4968: std_logic; attribute dont_touch of G4968: signal is true;
	signal G4969: std_logic; attribute dont_touch of G4969: signal is true;
	signal G5000: std_logic; attribute dont_touch of G5000: signal is true;
	signal G5001: std_logic; attribute dont_touch of G5001: signal is true;
	signal G5002: std_logic; attribute dont_touch of G5002: signal is true;
	signal G5005: std_logic; attribute dont_touch of G5005: signal is true;
	signal G5006: std_logic; attribute dont_touch of G5006: signal is true;
	signal G5007: std_logic; attribute dont_touch of G5007: signal is true;
	signal G5008: std_logic; attribute dont_touch of G5008: signal is true;
	signal G5009: std_logic; attribute dont_touch of G5009: signal is true;
	signal G5013: std_logic; attribute dont_touch of G5013: signal is true;
	signal G5014: std_logic; attribute dont_touch of G5014: signal is true;
	signal G5015: std_logic; attribute dont_touch of G5015: signal is true;
	signal G5016: std_logic; attribute dont_touch of G5016: signal is true;
	signal G5017: std_logic; attribute dont_touch of G5017: signal is true;
	signal G5018: std_logic; attribute dont_touch of G5018: signal is true;
	signal G5019: std_logic; attribute dont_touch of G5019: signal is true;
	signal G5020: std_logic; attribute dont_touch of G5020: signal is true;
	signal G5021: std_logic; attribute dont_touch of G5021: signal is true;
	signal G5022: std_logic; attribute dont_touch of G5022: signal is true;
	signal G5023: std_logic; attribute dont_touch of G5023: signal is true;
	signal G5024: std_logic; attribute dont_touch of G5024: signal is true;
	signal G5025: std_logic; attribute dont_touch of G5025: signal is true;
	signal G5026: std_logic; attribute dont_touch of G5026: signal is true;
	signal G5027: std_logic; attribute dont_touch of G5027: signal is true;
	signal G5028: std_logic; attribute dont_touch of G5028: signal is true;
	signal G5029: std_logic; attribute dont_touch of G5029: signal is true;
	signal G5030: std_logic; attribute dont_touch of G5030: signal is true;
	signal G5031: std_logic; attribute dont_touch of G5031: signal is true;
	signal G5032: std_logic; attribute dont_touch of G5032: signal is true;
	signal G5033: std_logic; attribute dont_touch of G5033: signal is true;
	signal G5034: std_logic; attribute dont_touch of G5034: signal is true;
	signal G5035: std_logic; attribute dont_touch of G5035: signal is true;
	signal G5036: std_logic; attribute dont_touch of G5036: signal is true;
	signal G5037: std_logic; attribute dont_touch of G5037: signal is true;
	signal G5038: std_logic; attribute dont_touch of G5038: signal is true;
	signal G5039: std_logic; attribute dont_touch of G5039: signal is true;
	signal G5040: std_logic; attribute dont_touch of G5040: signal is true;
	signal G5041: std_logic; attribute dont_touch of G5041: signal is true;
	signal G5042: std_logic; attribute dont_touch of G5042: signal is true;
	signal G5043: std_logic; attribute dont_touch of G5043: signal is true;
	signal G5044: std_logic; attribute dont_touch of G5044: signal is true;
	signal G5045: std_logic; attribute dont_touch of G5045: signal is true;
	signal G5046: std_logic; attribute dont_touch of G5046: signal is true;
	signal G5047: std_logic; attribute dont_touch of G5047: signal is true;
	signal G5048: std_logic; attribute dont_touch of G5048: signal is true;
	signal G5049: std_logic; attribute dont_touch of G5049: signal is true;
	signal G5050: std_logic; attribute dont_touch of G5050: signal is true;
	signal G5051: std_logic; attribute dont_touch of G5051: signal is true;
	signal G5052: std_logic; attribute dont_touch of G5052: signal is true;
	signal G5053: std_logic; attribute dont_touch of G5053: signal is true;
	signal G5054: std_logic; attribute dont_touch of G5054: signal is true;
	signal G5055: std_logic; attribute dont_touch of G5055: signal is true;
	signal G5056: std_logic; attribute dont_touch of G5056: signal is true;
	signal G5057: std_logic; attribute dont_touch of G5057: signal is true;
	signal G5058: std_logic; attribute dont_touch of G5058: signal is true;
	signal G5059: std_logic; attribute dont_touch of G5059: signal is true;
	signal G5060: std_logic; attribute dont_touch of G5060: signal is true;
	signal G5061: std_logic; attribute dont_touch of G5061: signal is true;
	signal G5062: std_logic; attribute dont_touch of G5062: signal is true;
	signal G5063: std_logic; attribute dont_touch of G5063: signal is true;
	signal G5064: std_logic; attribute dont_touch of G5064: signal is true;
	signal G5065: std_logic; attribute dont_touch of G5065: signal is true;
	signal G5066: std_logic; attribute dont_touch of G5066: signal is true;
	signal G5067: std_logic; attribute dont_touch of G5067: signal is true;
	signal G5068: std_logic; attribute dont_touch of G5068: signal is true;
	signal G5069: std_logic; attribute dont_touch of G5069: signal is true;
	signal G5070: std_logic; attribute dont_touch of G5070: signal is true;
	signal G5071: std_logic; attribute dont_touch of G5071: signal is true;
	signal G5072: std_logic; attribute dont_touch of G5072: signal is true;
	signal G5073: std_logic; attribute dont_touch of G5073: signal is true;
	signal G5074: std_logic; attribute dont_touch of G5074: signal is true;
	signal G5075: std_logic; attribute dont_touch of G5075: signal is true;
	signal G5076: std_logic; attribute dont_touch of G5076: signal is true;
	signal G5077: std_logic; attribute dont_touch of G5077: signal is true;
	signal G5078: std_logic; attribute dont_touch of G5078: signal is true;
	signal G5079: std_logic; attribute dont_touch of G5079: signal is true;
	signal G5080: std_logic; attribute dont_touch of G5080: signal is true;
	signal G5081: std_logic; attribute dont_touch of G5081: signal is true;
	signal G5082: std_logic; attribute dont_touch of G5082: signal is true;
	signal G5083: std_logic; attribute dont_touch of G5083: signal is true;
	signal G5084: std_logic; attribute dont_touch of G5084: signal is true;
	signal G5085: std_logic; attribute dont_touch of G5085: signal is true;
	signal G5086: std_logic; attribute dont_touch of G5086: signal is true;
	signal G5087: std_logic; attribute dont_touch of G5087: signal is true;
	signal G5088: std_logic; attribute dont_touch of G5088: signal is true;
	signal G5089: std_logic; attribute dont_touch of G5089: signal is true;
	signal G5090: std_logic; attribute dont_touch of G5090: signal is true;
	signal G5091: std_logic; attribute dont_touch of G5091: signal is true;
	signal G5092: std_logic; attribute dont_touch of G5092: signal is true;
	signal G5093: std_logic; attribute dont_touch of G5093: signal is true;
	signal G5094: std_logic; attribute dont_touch of G5094: signal is true;
	signal G5095: std_logic; attribute dont_touch of G5095: signal is true;
	signal G5096: std_logic; attribute dont_touch of G5096: signal is true;
	signal G5099: std_logic; attribute dont_touch of G5099: signal is true;
	signal G5100: std_logic; attribute dont_touch of G5100: signal is true;
	signal G5101: std_logic; attribute dont_touch of G5101: signal is true;
	signal G5104: std_logic; attribute dont_touch of G5104: signal is true;
	signal G5105: std_logic; attribute dont_touch of G5105: signal is true;
	signal G5106: std_logic; attribute dont_touch of G5106: signal is true;
	signal G5107: std_logic; attribute dont_touch of G5107: signal is true;
	signal G5108: std_logic; attribute dont_touch of G5108: signal is true;
	signal G5109: std_logic; attribute dont_touch of G5109: signal is true;
	signal G5112: std_logic; attribute dont_touch of G5112: signal is true;
	signal G5113: std_logic; attribute dont_touch of G5113: signal is true;
	signal G5114: std_logic; attribute dont_touch of G5114: signal is true;
	signal G5115: std_logic; attribute dont_touch of G5115: signal is true;
	signal G5116: std_logic; attribute dont_touch of G5116: signal is true;
	signal G5117: std_logic; attribute dont_touch of G5117: signal is true;
	signal G5118: std_logic; attribute dont_touch of G5118: signal is true;
	signal G5119: std_logic; attribute dont_touch of G5119: signal is true;
	signal G5120: std_logic; attribute dont_touch of G5120: signal is true;
	signal G5121: std_logic; attribute dont_touch of G5121: signal is true;
	signal G5122: std_logic; attribute dont_touch of G5122: signal is true;
	signal G5123: std_logic; attribute dont_touch of G5123: signal is true;
	signal G5124: std_logic; attribute dont_touch of G5124: signal is true;
	signal G5125: std_logic; attribute dont_touch of G5125: signal is true;
	signal G5126: std_logic; attribute dont_touch of G5126: signal is true;
	signal G5127: std_logic; attribute dont_touch of G5127: signal is true;
	signal G5128: std_logic; attribute dont_touch of G5128: signal is true;
	signal G5129: std_logic; attribute dont_touch of G5129: signal is true;
	signal G5132: std_logic; attribute dont_touch of G5132: signal is true;
	signal G5137: std_logic; attribute dont_touch of G5137: signal is true;
	signal G5138: std_logic; attribute dont_touch of G5138: signal is true;
	signal G5139: std_logic; attribute dont_touch of G5139: signal is true;
	signal G5140: std_logic; attribute dont_touch of G5140: signal is true;
	signal G5141: std_logic; attribute dont_touch of G5141: signal is true;
	signal G5142: std_logic; attribute dont_touch of G5142: signal is true;
	signal G5144: std_logic; attribute dont_touch of G5144: signal is true;
	signal G5145: std_logic; attribute dont_touch of G5145: signal is true;
	signal G5146: std_logic; attribute dont_touch of G5146: signal is true;
	signal G5147: std_logic; attribute dont_touch of G5147: signal is true;
	signal G5148: std_logic; attribute dont_touch of G5148: signal is true;
	signal G5149: std_logic; attribute dont_touch of G5149: signal is true;
	signal G5150: std_logic; attribute dont_touch of G5150: signal is true;
	signal G5151: std_logic; attribute dont_touch of G5151: signal is true;
	signal G5152: std_logic; attribute dont_touch of G5152: signal is true;
	signal G5153: std_logic; attribute dont_touch of G5153: signal is true;
	signal G5154: std_logic; attribute dont_touch of G5154: signal is true;
	signal G5155: std_logic; attribute dont_touch of G5155: signal is true;
	signal G5156: std_logic; attribute dont_touch of G5156: signal is true;
	signal G5157: std_logic; attribute dont_touch of G5157: signal is true;
	signal G5158: std_logic; attribute dont_touch of G5158: signal is true;
	signal G5159: std_logic; attribute dont_touch of G5159: signal is true;
	signal G5160: std_logic; attribute dont_touch of G5160: signal is true;
	signal G5161: std_logic; attribute dont_touch of G5161: signal is true;
	signal G5162: std_logic; attribute dont_touch of G5162: signal is true;
	signal G5163: std_logic; attribute dont_touch of G5163: signal is true;
	signal G5165: std_logic; attribute dont_touch of G5165: signal is true;
	signal G5166: std_logic; attribute dont_touch of G5166: signal is true;
	signal G5167: std_logic; attribute dont_touch of G5167: signal is true;
	signal G5168: std_logic; attribute dont_touch of G5168: signal is true;
	signal G5169: std_logic; attribute dont_touch of G5169: signal is true;
	signal G5170: std_logic; attribute dont_touch of G5170: signal is true;
	signal G5171: std_logic; attribute dont_touch of G5171: signal is true;
	signal G5172: std_logic; attribute dont_touch of G5172: signal is true;
	signal G5173: std_logic; attribute dont_touch of G5173: signal is true;
	signal G5174: std_logic; attribute dont_touch of G5174: signal is true;
	signal G5175: std_logic; attribute dont_touch of G5175: signal is true;
	signal G5176: std_logic; attribute dont_touch of G5176: signal is true;
	signal G5177: std_logic; attribute dont_touch of G5177: signal is true;
	signal G5178: std_logic; attribute dont_touch of G5178: signal is true;
	signal G5179: std_logic; attribute dont_touch of G5179: signal is true;
	signal G5180: std_logic; attribute dont_touch of G5180: signal is true;
	signal G5181: std_logic; attribute dont_touch of G5181: signal is true;
	signal G5182: std_logic; attribute dont_touch of G5182: signal is true;
	signal G5183: std_logic; attribute dont_touch of G5183: signal is true;
	signal G5184: std_logic; attribute dont_touch of G5184: signal is true;
	signal G5185: std_logic; attribute dont_touch of G5185: signal is true;
	signal G5186: std_logic; attribute dont_touch of G5186: signal is true;
	signal G5187: std_logic; attribute dont_touch of G5187: signal is true;
	signal G5188: std_logic; attribute dont_touch of G5188: signal is true;
	signal G5189: std_logic; attribute dont_touch of G5189: signal is true;
	signal G5190: std_logic; attribute dont_touch of G5190: signal is true;
	signal G5191: std_logic; attribute dont_touch of G5191: signal is true;
	signal G5192: std_logic; attribute dont_touch of G5192: signal is true;
	signal G5193: std_logic; attribute dont_touch of G5193: signal is true;
	signal G5194: std_logic; attribute dont_touch of G5194: signal is true;
	signal G5195: std_logic; attribute dont_touch of G5195: signal is true;
	signal G5196: std_logic; attribute dont_touch of G5196: signal is true;
	signal G5197: std_logic; attribute dont_touch of G5197: signal is true;
	signal G5198: std_logic; attribute dont_touch of G5198: signal is true;
	signal G5199: std_logic; attribute dont_touch of G5199: signal is true;
	signal G5200: std_logic; attribute dont_touch of G5200: signal is true;
	signal G5201: std_logic; attribute dont_touch of G5201: signal is true;
	signal G5202: std_logic; attribute dont_touch of G5202: signal is true;
	signal G5203: std_logic; attribute dont_touch of G5203: signal is true;
	signal G5204: std_logic; attribute dont_touch of G5204: signal is true;
	signal G5205: std_logic; attribute dont_touch of G5205: signal is true;
	signal G5206: std_logic; attribute dont_touch of G5206: signal is true;
	signal G5207: std_logic; attribute dont_touch of G5207: signal is true;
	signal G5208: std_logic; attribute dont_touch of G5208: signal is true;
	signal G5209: std_logic; attribute dont_touch of G5209: signal is true;
	signal G5210: std_logic; attribute dont_touch of G5210: signal is true;
	signal G5211: std_logic; attribute dont_touch of G5211: signal is true;
	signal G5212: std_logic; attribute dont_touch of G5212: signal is true;
	signal G5213: std_logic; attribute dont_touch of G5213: signal is true;
	signal G5214: std_logic; attribute dont_touch of G5214: signal is true;
	signal G5215: std_logic; attribute dont_touch of G5215: signal is true;
	signal G5216: std_logic; attribute dont_touch of G5216: signal is true;
	signal G5217: std_logic; attribute dont_touch of G5217: signal is true;
	signal G5218: std_logic; attribute dont_touch of G5218: signal is true;
	signal G5219: std_logic; attribute dont_touch of G5219: signal is true;
	signal G5220: std_logic; attribute dont_touch of G5220: signal is true;
	signal G5221: std_logic; attribute dont_touch of G5221: signal is true;
	signal G5222: std_logic; attribute dont_touch of G5222: signal is true;
	signal G5223: std_logic; attribute dont_touch of G5223: signal is true;
	signal G5224: std_logic; attribute dont_touch of G5224: signal is true;
	signal G5227: std_logic; attribute dont_touch of G5227: signal is true;
	signal G5228: std_logic; attribute dont_touch of G5228: signal is true;
	signal G5229: std_logic; attribute dont_touch of G5229: signal is true;
	signal G5230: std_logic; attribute dont_touch of G5230: signal is true;
	signal G5231: std_logic; attribute dont_touch of G5231: signal is true;
	signal G5232: std_logic; attribute dont_touch of G5232: signal is true;
	signal G5233: std_logic; attribute dont_touch of G5233: signal is true;
	signal G5234: std_logic; attribute dont_touch of G5234: signal is true;
	signal G5235: std_logic; attribute dont_touch of G5235: signal is true;
	signal G5236: std_logic; attribute dont_touch of G5236: signal is true;
	signal G5237: std_logic; attribute dont_touch of G5237: signal is true;
	signal G5238: std_logic; attribute dont_touch of G5238: signal is true;
	signal G5239: std_logic; attribute dont_touch of G5239: signal is true;
	signal G5240: std_logic; attribute dont_touch of G5240: signal is true;
	signal G5241: std_logic; attribute dont_touch of G5241: signal is true;
	signal G5242: std_logic; attribute dont_touch of G5242: signal is true;
	signal G5243: std_logic; attribute dont_touch of G5243: signal is true;
	signal G5244: std_logic; attribute dont_touch of G5244: signal is true;
	signal G5245: std_logic; attribute dont_touch of G5245: signal is true;
	signal G5246: std_logic; attribute dont_touch of G5246: signal is true;
	signal G5253: std_logic; attribute dont_touch of G5253: signal is true;
	signal G5254: std_logic; attribute dont_touch of G5254: signal is true;
	signal G5255: std_logic; attribute dont_touch of G5255: signal is true;
	signal G5256: std_logic; attribute dont_touch of G5256: signal is true;
	signal G5257: std_logic; attribute dont_touch of G5257: signal is true;
	signal G5258: std_logic; attribute dont_touch of G5258: signal is true;
	signal G5259: std_logic; attribute dont_touch of G5259: signal is true;
	signal G5260: std_logic; attribute dont_touch of G5260: signal is true;
	signal G5261: std_logic; attribute dont_touch of G5261: signal is true;
	signal G5264: std_logic; attribute dont_touch of G5264: signal is true;
	signal G5265: std_logic; attribute dont_touch of G5265: signal is true;
	signal G5266: std_logic; attribute dont_touch of G5266: signal is true;
	signal G5267: std_logic; attribute dont_touch of G5267: signal is true;
	signal G5268: std_logic; attribute dont_touch of G5268: signal is true;
	signal G5269: std_logic; attribute dont_touch of G5269: signal is true;
	signal G5278: std_logic; attribute dont_touch of G5278: signal is true;
	signal G5284: std_logic; attribute dont_touch of G5284: signal is true;
	signal G5285: std_logic; attribute dont_touch of G5285: signal is true;
	signal G5286: std_logic; attribute dont_touch of G5286: signal is true;
	signal G5287: std_logic; attribute dont_touch of G5287: signal is true;
	signal G5291: std_logic; attribute dont_touch of G5291: signal is true;
	signal G5294: std_logic; attribute dont_touch of G5294: signal is true;
	signal G5298: std_logic; attribute dont_touch of G5298: signal is true;
	signal G5299: std_logic; attribute dont_touch of G5299: signal is true;
	signal G5302: std_logic; attribute dont_touch of G5302: signal is true;
	signal G5305: std_logic; attribute dont_touch of G5305: signal is true;
	signal G5309: std_logic; attribute dont_touch of G5309: signal is true;
	signal G5310: std_logic; attribute dont_touch of G5310: signal is true;
	signal G5311: std_logic; attribute dont_touch of G5311: signal is true;
	signal G5312: std_logic; attribute dont_touch of G5312: signal is true;
	signal G5313: std_logic; attribute dont_touch of G5313: signal is true;
	signal G5314: std_logic; attribute dont_touch of G5314: signal is true;
	signal G5317: std_logic; attribute dont_touch of G5317: signal is true;
	signal G5334: std_logic; attribute dont_touch of G5334: signal is true;
	signal G5335: std_logic; attribute dont_touch of G5335: signal is true;
	signal G5343: std_logic; attribute dont_touch of G5343: signal is true;
	signal G5344: std_logic; attribute dont_touch of G5344: signal is true;
	signal G5345: std_logic; attribute dont_touch of G5345: signal is true;
	signal G5362: std_logic; attribute dont_touch of G5362: signal is true;
	signal G5363: std_logic; attribute dont_touch of G5363: signal is true;
	signal G5364: std_logic; attribute dont_touch of G5364: signal is true;
	signal G5367: std_logic; attribute dont_touch of G5367: signal is true;
	signal G5384: std_logic; attribute dont_touch of G5384: signal is true;
	signal G5395: std_logic; attribute dont_touch of G5395: signal is true;
	signal G5396: std_logic; attribute dont_touch of G5396: signal is true;
	signal G5397: std_logic; attribute dont_touch of G5397: signal is true;
	signal G5401: std_logic; attribute dont_touch of G5401: signal is true;
	signal G5402: std_logic; attribute dont_touch of G5402: signal is true;
	signal G5403: std_logic; attribute dont_touch of G5403: signal is true;
	signal G5412: std_logic; attribute dont_touch of G5412: signal is true;
	signal G5417: std_logic; attribute dont_touch of G5417: signal is true;
	signal G5418: std_logic; attribute dont_touch of G5418: signal is true;
	signal G5425: std_logic; attribute dont_touch of G5425: signal is true;
	signal G5426: std_logic; attribute dont_touch of G5426: signal is true;
	signal G5427: std_logic; attribute dont_touch of G5427: signal is true;
	signal G5428: std_logic; attribute dont_touch of G5428: signal is true;
	signal G5432: std_logic; attribute dont_touch of G5432: signal is true;
	signal G5433: std_logic; attribute dont_touch of G5433: signal is true;
	signal G5434: std_logic; attribute dont_touch of G5434: signal is true;
	signal G5435: std_logic; attribute dont_touch of G5435: signal is true;
	signal G5436: std_logic; attribute dont_touch of G5436: signal is true;
	signal G5437: std_logic; attribute dont_touch of G5437: signal is true;
	signal G5438: std_logic; attribute dont_touch of G5438: signal is true;
	signal G5439: std_logic; attribute dont_touch of G5439: signal is true;
	signal G5440: std_logic; attribute dont_touch of G5440: signal is true;
	signal G5441: std_logic; attribute dont_touch of G5441: signal is true;
	signal G5442: std_logic; attribute dont_touch of G5442: signal is true;
	signal G5443: std_logic; attribute dont_touch of G5443: signal is true;
	signal G5444: std_logic; attribute dont_touch of G5444: signal is true;
	signal G5445: std_logic; attribute dont_touch of G5445: signal is true;
	signal G5448: std_logic; attribute dont_touch of G5448: signal is true;
	signal G5452: std_logic; attribute dont_touch of G5452: signal is true;
	signal G5453: std_logic; attribute dont_touch of G5453: signal is true;
	signal G5458: std_logic; attribute dont_touch of G5458: signal is true;
	signal G5459: std_logic; attribute dont_touch of G5459: signal is true;
	signal G5460: std_logic; attribute dont_touch of G5460: signal is true;
	signal G5461: std_logic; attribute dont_touch of G5461: signal is true;
	signal G5462: std_logic; attribute dont_touch of G5462: signal is true;
	signal G5463: std_logic; attribute dont_touch of G5463: signal is true;
	signal G5466: std_logic; attribute dont_touch of G5466: signal is true;
	signal G5467: std_logic; attribute dont_touch of G5467: signal is true;
	signal G5468: std_logic; attribute dont_touch of G5468: signal is true;
	signal G5469: std_logic; attribute dont_touch of G5469: signal is true;
	signal G5470: std_logic; attribute dont_touch of G5470: signal is true;
	signal G5471: std_logic; attribute dont_touch of G5471: signal is true;
	signal G5472: std_logic; attribute dont_touch of G5472: signal is true;
	signal G5473: std_logic; attribute dont_touch of G5473: signal is true;
	signal G5474: std_logic; attribute dont_touch of G5474: signal is true;
	signal G5475: std_logic; attribute dont_touch of G5475: signal is true;
	signal G5476: std_logic; attribute dont_touch of G5476: signal is true;
	signal G5477: std_logic; attribute dont_touch of G5477: signal is true;
	signal G5478: std_logic; attribute dont_touch of G5478: signal is true;
	signal G5479: std_logic; attribute dont_touch of G5479: signal is true;
	signal G5480: std_logic; attribute dont_touch of G5480: signal is true;
	signal G5481: std_logic; attribute dont_touch of G5481: signal is true;
	signal G5482: std_logic; attribute dont_touch of G5482: signal is true;
	signal G5483: std_logic; attribute dont_touch of G5483: signal is true;
	signal G5484: std_logic; attribute dont_touch of G5484: signal is true;
	signal G5487: std_logic; attribute dont_touch of G5487: signal is true;
	signal G5488: std_logic; attribute dont_touch of G5488: signal is true;
	signal G5489: std_logic; attribute dont_touch of G5489: signal is true;
	signal G5490: std_logic; attribute dont_touch of G5490: signal is true;
	signal G5491: std_logic; attribute dont_touch of G5491: signal is true;
	signal G5492: std_logic; attribute dont_touch of G5492: signal is true;
	signal G5493: std_logic; attribute dont_touch of G5493: signal is true;
	signal G5494: std_logic; attribute dont_touch of G5494: signal is true;
	signal G5511: std_logic; attribute dont_touch of G5511: signal is true;
	signal G5512: std_logic; attribute dont_touch of G5512: signal is true;
	signal G5513: std_logic; attribute dont_touch of G5513: signal is true;
	signal G5514: std_logic; attribute dont_touch of G5514: signal is true;
	signal G5515: std_logic; attribute dont_touch of G5515: signal is true;
	signal G5516: std_logic; attribute dont_touch of G5516: signal is true;
	signal G5517: std_logic; attribute dont_touch of G5517: signal is true;
	signal G5518: std_logic; attribute dont_touch of G5518: signal is true;
	signal G5519: std_logic; attribute dont_touch of G5519: signal is true;
	signal G5520: std_logic; attribute dont_touch of G5520: signal is true;
	signal G5521: std_logic; attribute dont_touch of G5521: signal is true;
	signal G5522: std_logic; attribute dont_touch of G5522: signal is true;
	signal G5523: std_logic; attribute dont_touch of G5523: signal is true;
	signal G5524: std_logic; attribute dont_touch of G5524: signal is true;
	signal G5525: std_logic; attribute dont_touch of G5525: signal is true;
	signal G5526: std_logic; attribute dont_touch of G5526: signal is true;
	signal G5529: std_logic; attribute dont_touch of G5529: signal is true;
	signal G5537: std_logic; attribute dont_touch of G5537: signal is true;
	signal G5538: std_logic; attribute dont_touch of G5538: signal is true;
	signal G5539: std_logic; attribute dont_touch of G5539: signal is true;
	signal G5540: std_logic; attribute dont_touch of G5540: signal is true;
	signal G5541: std_logic; attribute dont_touch of G5541: signal is true;
	signal G5542: std_logic; attribute dont_touch of G5542: signal is true;
	signal G5545: std_logic; attribute dont_touch of G5545: signal is true;
	signal G5546: std_logic; attribute dont_touch of G5546: signal is true;
	signal G5547: std_logic; attribute dont_touch of G5547: signal is true;
	signal G5548: std_logic; attribute dont_touch of G5548: signal is true;
	signal G5549: std_logic; attribute dont_touch of G5549: signal is true;
	signal G5550: std_logic; attribute dont_touch of G5550: signal is true;
	signal G5551: std_logic; attribute dont_touch of G5551: signal is true;
	signal G5552: std_logic; attribute dont_touch of G5552: signal is true;
	signal G5555: std_logic; attribute dont_touch of G5555: signal is true;
	signal G5556: std_logic; attribute dont_touch of G5556: signal is true;
	signal G5557: std_logic; attribute dont_touch of G5557: signal is true;
	signal G5558: std_logic; attribute dont_touch of G5558: signal is true;
	signal G5559: std_logic; attribute dont_touch of G5559: signal is true;
	signal G5560: std_logic; attribute dont_touch of G5560: signal is true;
	signal G5561: std_logic; attribute dont_touch of G5561: signal is true;
	signal G5562: std_logic; attribute dont_touch of G5562: signal is true;
	signal G5563: std_logic; attribute dont_touch of G5563: signal is true;
	signal G5564: std_logic; attribute dont_touch of G5564: signal is true;
	signal G5565: std_logic; attribute dont_touch of G5565: signal is true;
	signal G5566: std_logic; attribute dont_touch of G5566: signal is true;
	signal G5567: std_logic; attribute dont_touch of G5567: signal is true;
	signal G5568: std_logic; attribute dont_touch of G5568: signal is true;
	signal G5569: std_logic; attribute dont_touch of G5569: signal is true;
	signal G5570: std_logic; attribute dont_touch of G5570: signal is true;
	signal G5572: std_logic; attribute dont_touch of G5572: signal is true;
	signal G5573: std_logic; attribute dont_touch of G5573: signal is true;
	signal G5574: std_logic; attribute dont_touch of G5574: signal is true;
	signal G5575: std_logic; attribute dont_touch of G5575: signal is true;
	signal G5576: std_logic; attribute dont_touch of G5576: signal is true;
	signal G5577: std_logic; attribute dont_touch of G5577: signal is true;
	signal G5578: std_logic; attribute dont_touch of G5578: signal is true;
	signal G5579: std_logic; attribute dont_touch of G5579: signal is true;
	signal G5580: std_logic; attribute dont_touch of G5580: signal is true;
	signal G5581: std_logic; attribute dont_touch of G5581: signal is true;
	signal G5582: std_logic; attribute dont_touch of G5582: signal is true;
	signal G5583: std_logic; attribute dont_touch of G5583: signal is true;
	signal G5584: std_logic; attribute dont_touch of G5584: signal is true;
	signal G5585: std_logic; attribute dont_touch of G5585: signal is true;
	signal G5586: std_logic; attribute dont_touch of G5586: signal is true;
	signal G5587: std_logic; attribute dont_touch of G5587: signal is true;
	signal G5588: std_logic; attribute dont_touch of G5588: signal is true;
	signal G5589: std_logic; attribute dont_touch of G5589: signal is true;
	signal G5590: std_logic; attribute dont_touch of G5590: signal is true;
	signal G5591: std_logic; attribute dont_touch of G5591: signal is true;
	signal G5592: std_logic; attribute dont_touch of G5592: signal is true;
	signal G5593: std_logic; attribute dont_touch of G5593: signal is true;
	signal G5594: std_logic; attribute dont_touch of G5594: signal is true;
	signal G5595: std_logic; attribute dont_touch of G5595: signal is true;
	signal G5596: std_logic; attribute dont_touch of G5596: signal is true;
	signal G5597: std_logic; attribute dont_touch of G5597: signal is true;
	signal G5598: std_logic; attribute dont_touch of G5598: signal is true;
	signal G5599: std_logic; attribute dont_touch of G5599: signal is true;
	signal G5600: std_logic; attribute dont_touch of G5600: signal is true;
	signal G5603: std_logic; attribute dont_touch of G5603: signal is true;
	signal G5604: std_logic; attribute dont_touch of G5604: signal is true;
	signal G5605: std_logic; attribute dont_touch of G5605: signal is true;
	signal G5606: std_logic; attribute dont_touch of G5606: signal is true;
	signal G5607: std_logic; attribute dont_touch of G5607: signal is true;
	signal G5608: std_logic; attribute dont_touch of G5608: signal is true;
	signal G5609: std_logic; attribute dont_touch of G5609: signal is true;
	signal G5610: std_logic; attribute dont_touch of G5610: signal is true;
	signal G5611: std_logic; attribute dont_touch of G5611: signal is true;
	signal G5612: std_logic; attribute dont_touch of G5612: signal is true;
	signal G5613: std_logic; attribute dont_touch of G5613: signal is true;
	signal G5614: std_logic; attribute dont_touch of G5614: signal is true;
	signal G5615: std_logic; attribute dont_touch of G5615: signal is true;
	signal G5616: std_logic; attribute dont_touch of G5616: signal is true;
	signal G5617: std_logic; attribute dont_touch of G5617: signal is true;
	signal G5618: std_logic; attribute dont_touch of G5618: signal is true;
	signal G5621: std_logic; attribute dont_touch of G5621: signal is true;
	signal G5622: std_logic; attribute dont_touch of G5622: signal is true;
	signal G5623: std_logic; attribute dont_touch of G5623: signal is true;
	signal G5624: std_logic; attribute dont_touch of G5624: signal is true;
	signal G5625: std_logic; attribute dont_touch of G5625: signal is true;
	signal G5626: std_logic; attribute dont_touch of G5626: signal is true;
	signal G5627: std_logic; attribute dont_touch of G5627: signal is true;
	signal G5628: std_logic; attribute dont_touch of G5628: signal is true;
	signal G5631: std_logic; attribute dont_touch of G5631: signal is true;
	signal G5632: std_logic; attribute dont_touch of G5632: signal is true;
	signal G5633: std_logic; attribute dont_touch of G5633: signal is true;
	signal G5638: std_logic; attribute dont_touch of G5638: signal is true;
	signal G5639: std_logic; attribute dont_touch of G5639: signal is true;
	signal G5642: std_logic; attribute dont_touch of G5642: signal is true;
	signal G5643: std_logic; attribute dont_touch of G5643: signal is true;
	signal G5644: std_logic; attribute dont_touch of G5644: signal is true;
	signal G5645: std_logic; attribute dont_touch of G5645: signal is true;
	signal G5648: std_logic; attribute dont_touch of G5648: signal is true;
	signal G5649: std_logic; attribute dont_touch of G5649: signal is true;
	signal G5652: std_logic; attribute dont_touch of G5652: signal is true;
	signal G5653: std_logic; attribute dont_touch of G5653: signal is true;
	signal G5654: std_logic; attribute dont_touch of G5654: signal is true;
	signal G5657: std_logic; attribute dont_touch of G5657: signal is true;
	signal G5658: std_logic; attribute dont_touch of G5658: signal is true;
	signal G5661: std_logic; attribute dont_touch of G5661: signal is true;
	signal G5662: std_logic; attribute dont_touch of G5662: signal is true;
	signal G5665: std_logic; attribute dont_touch of G5665: signal is true;
	signal G5668: std_logic; attribute dont_touch of G5668: signal is true;
	signal G5670: std_logic; attribute dont_touch of G5670: signal is true;
	signal G5671: std_logic; attribute dont_touch of G5671: signal is true;
	signal G5672: std_logic; attribute dont_touch of G5672: signal is true;
	signal G5673: std_logic; attribute dont_touch of G5673: signal is true;
	signal G5674: std_logic; attribute dont_touch of G5674: signal is true;
	signal G5677: std_logic; attribute dont_touch of G5677: signal is true;
	signal G5679: std_logic; attribute dont_touch of G5679: signal is true;
	signal G5680: std_logic; attribute dont_touch of G5680: signal is true;
	signal G5681: std_logic; attribute dont_touch of G5681: signal is true;
	signal G5683: std_logic; attribute dont_touch of G5683: signal is true;
	signal G5685: std_logic; attribute dont_touch of G5685: signal is true;
	signal G5686: std_logic; attribute dont_touch of G5686: signal is true;
	signal G5688: std_logic; attribute dont_touch of G5688: signal is true;
	signal G5689: std_logic; attribute dont_touch of G5689: signal is true;
	signal G5690: std_logic; attribute dont_touch of G5690: signal is true;
	signal G5693: std_logic; attribute dont_touch of G5693: signal is true;
	signal G5696: std_logic; attribute dont_touch of G5696: signal is true;
	signal G5697: std_logic; attribute dont_touch of G5697: signal is true;
	signal G5698: std_logic; attribute dont_touch of G5698: signal is true;
	signal G5699: std_logic; attribute dont_touch of G5699: signal is true;
	signal G5700: std_logic; attribute dont_touch of G5700: signal is true;
	signal G5701: std_logic; attribute dont_touch of G5701: signal is true;
	signal G5704: std_logic; attribute dont_touch of G5704: signal is true;
	signal G5705: std_logic; attribute dont_touch of G5705: signal is true;
	signal G5706: std_logic; attribute dont_touch of G5706: signal is true;
	signal G5707: std_logic; attribute dont_touch of G5707: signal is true;
	signal G5708: std_logic; attribute dont_touch of G5708: signal is true;
	signal G5709: std_logic; attribute dont_touch of G5709: signal is true;
	signal G5710: std_logic; attribute dont_touch of G5710: signal is true;
	signal G5711: std_logic; attribute dont_touch of G5711: signal is true;
	signal G5712: std_logic; attribute dont_touch of G5712: signal is true;
	signal G5713: std_logic; attribute dont_touch of G5713: signal is true;
	signal G5714: std_logic; attribute dont_touch of G5714: signal is true;
	signal G5715: std_logic; attribute dont_touch of G5715: signal is true;
	signal G5716: std_logic; attribute dont_touch of G5716: signal is true;
	signal G5717: std_logic; attribute dont_touch of G5717: signal is true;
	signal G5718: std_logic; attribute dont_touch of G5718: signal is true;
	signal G5719: std_logic; attribute dont_touch of G5719: signal is true;
	signal G5722: std_logic; attribute dont_touch of G5722: signal is true;
	signal G5723: std_logic; attribute dont_touch of G5723: signal is true;
	signal G5724: std_logic; attribute dont_touch of G5724: signal is true;
	signal G5725: std_logic; attribute dont_touch of G5725: signal is true;
	signal G5726: std_logic; attribute dont_touch of G5726: signal is true;
	signal G5730: std_logic; attribute dont_touch of G5730: signal is true;
	signal G5731: std_logic; attribute dont_touch of G5731: signal is true;
	signal G5732: std_logic; attribute dont_touch of G5732: signal is true;
	signal G5733: std_logic; attribute dont_touch of G5733: signal is true;
	signal G5734: std_logic; attribute dont_touch of G5734: signal is true;
	signal G5735: std_logic; attribute dont_touch of G5735: signal is true;
	signal G5736: std_logic; attribute dont_touch of G5736: signal is true;
	signal G5737: std_logic; attribute dont_touch of G5737: signal is true;
	signal G5738: std_logic; attribute dont_touch of G5738: signal is true;
	signal G5739: std_logic; attribute dont_touch of G5739: signal is true;
	signal G5740: std_logic; attribute dont_touch of G5740: signal is true;
	signal G5741: std_logic; attribute dont_touch of G5741: signal is true;
	signal G5742: std_logic; attribute dont_touch of G5742: signal is true;
	signal G5743: std_logic; attribute dont_touch of G5743: signal is true;
	signal G5744: std_logic; attribute dont_touch of G5744: signal is true;
	signal G5745: std_logic; attribute dont_touch of G5745: signal is true;
	signal G5746: std_logic; attribute dont_touch of G5746: signal is true;
	signal G5747: std_logic; attribute dont_touch of G5747: signal is true;
	signal G5748: std_logic; attribute dont_touch of G5748: signal is true;
	signal G5749: std_logic; attribute dont_touch of G5749: signal is true;
	signal G5750: std_logic; attribute dont_touch of G5750: signal is true;
	signal G5751: std_logic; attribute dont_touch of G5751: signal is true;
	signal G5752: std_logic; attribute dont_touch of G5752: signal is true;
	signal G5753: std_logic; attribute dont_touch of G5753: signal is true;
	signal G5754: std_logic; attribute dont_touch of G5754: signal is true;
	signal G5755: std_logic; attribute dont_touch of G5755: signal is true;
	signal G5756: std_logic; attribute dont_touch of G5756: signal is true;
	signal G5757: std_logic; attribute dont_touch of G5757: signal is true;
	signal G5758: std_logic; attribute dont_touch of G5758: signal is true;
	signal G5759: std_logic; attribute dont_touch of G5759: signal is true;
	signal G5760: std_logic; attribute dont_touch of G5760: signal is true;
	signal G5761: std_logic; attribute dont_touch of G5761: signal is true;
	signal G5762: std_logic; attribute dont_touch of G5762: signal is true;
	signal G5763: std_logic; attribute dont_touch of G5763: signal is true;
	signal G5764: std_logic; attribute dont_touch of G5764: signal is true;
	signal G5765: std_logic; attribute dont_touch of G5765: signal is true;
	signal G5766: std_logic; attribute dont_touch of G5766: signal is true;
	signal G5767: std_logic; attribute dont_touch of G5767: signal is true;
	signal G5768: std_logic; attribute dont_touch of G5768: signal is true;
	signal G5769: std_logic; attribute dont_touch of G5769: signal is true;
	signal G5772: std_logic; attribute dont_touch of G5772: signal is true;
	signal G5779: std_logic; attribute dont_touch of G5779: signal is true;
	signal G5780: std_logic; attribute dont_touch of G5780: signal is true;
	signal G5781: std_logic; attribute dont_touch of G5781: signal is true;
	signal G5782: std_logic; attribute dont_touch of G5782: signal is true;
	signal G5783: std_logic; attribute dont_touch of G5783: signal is true;
	signal G5784: std_logic; attribute dont_touch of G5784: signal is true;
	signal G5785: std_logic; attribute dont_touch of G5785: signal is true;
	signal G5786: std_logic; attribute dont_touch of G5786: signal is true;
	signal G5787: std_logic; attribute dont_touch of G5787: signal is true;
	signal G5788: std_logic; attribute dont_touch of G5788: signal is true;
	signal G5789: std_logic; attribute dont_touch of G5789: signal is true;
	signal G5790: std_logic; attribute dont_touch of G5790: signal is true;
	signal G5793: std_logic; attribute dont_touch of G5793: signal is true;
	signal G5794: std_logic; attribute dont_touch of G5794: signal is true;
	signal G5795: std_logic; attribute dont_touch of G5795: signal is true;
	signal G5796: std_logic; attribute dont_touch of G5796: signal is true;
	signal G5797: std_logic; attribute dont_touch of G5797: signal is true;
	signal G5798: std_logic; attribute dont_touch of G5798: signal is true;
	signal G5799: std_logic; attribute dont_touch of G5799: signal is true;
	signal G5800: std_logic; attribute dont_touch of G5800: signal is true;
	signal G5801: std_logic; attribute dont_touch of G5801: signal is true;
	signal G5802: std_logic; attribute dont_touch of G5802: signal is true;
	signal G5805: std_logic; attribute dont_touch of G5805: signal is true;
	signal G5806: std_logic; attribute dont_touch of G5806: signal is true;
	signal G5807: std_logic; attribute dont_touch of G5807: signal is true;
	signal G5808: std_logic; attribute dont_touch of G5808: signal is true;
	signal G5809: std_logic; attribute dont_touch of G5809: signal is true;
	signal G5810: std_logic; attribute dont_touch of G5810: signal is true;
	signal G5811: std_logic; attribute dont_touch of G5811: signal is true;
	signal G5812: std_logic; attribute dont_touch of G5812: signal is true;
	signal G5813: std_logic; attribute dont_touch of G5813: signal is true;
	signal G5814: std_logic; attribute dont_touch of G5814: signal is true;
	signal G5817: std_logic; attribute dont_touch of G5817: signal is true;
	signal G5818: std_logic; attribute dont_touch of G5818: signal is true;
	signal G5819: std_logic; attribute dont_touch of G5819: signal is true;
	signal G5820: std_logic; attribute dont_touch of G5820: signal is true;
	signal G5821: std_logic; attribute dont_touch of G5821: signal is true;
	signal G5822: std_logic; attribute dont_touch of G5822: signal is true;
	signal G5823: std_logic; attribute dont_touch of G5823: signal is true;
	signal G5824: std_logic; attribute dont_touch of G5824: signal is true;
	signal G5825: std_logic; attribute dont_touch of G5825: signal is true;
	signal G5826: std_logic; attribute dont_touch of G5826: signal is true;
	signal G5827: std_logic; attribute dont_touch of G5827: signal is true;
	signal G5828: std_logic; attribute dont_touch of G5828: signal is true;
	signal G5829: std_logic; attribute dont_touch of G5829: signal is true;
	signal G5830: std_logic; attribute dont_touch of G5830: signal is true;
	signal G5831: std_logic; attribute dont_touch of G5831: signal is true;
	signal G5832: std_logic; attribute dont_touch of G5832: signal is true;
	signal G5833: std_logic; attribute dont_touch of G5833: signal is true;
	signal G5834: std_logic; attribute dont_touch of G5834: signal is true;
	signal G5835: std_logic; attribute dont_touch of G5835: signal is true;
	signal G5836: std_logic; attribute dont_touch of G5836: signal is true;
	signal G5839: std_logic; attribute dont_touch of G5839: signal is true;
	signal G5840: std_logic; attribute dont_touch of G5840: signal is true;
	signal G5841: std_logic; attribute dont_touch of G5841: signal is true;
	signal G5842: std_logic; attribute dont_touch of G5842: signal is true;
	signal G5843: std_logic; attribute dont_touch of G5843: signal is true;
	signal G5844: std_logic; attribute dont_touch of G5844: signal is true;
	signal G5845: std_logic; attribute dont_touch of G5845: signal is true;
	signal G5846: std_logic; attribute dont_touch of G5846: signal is true;
	signal G5847: std_logic; attribute dont_touch of G5847: signal is true;
	signal G5868: std_logic; attribute dont_touch of G5868: signal is true;
	signal G5871: std_logic; attribute dont_touch of G5871: signal is true;
	signal G5872: std_logic; attribute dont_touch of G5872: signal is true;
	signal G5873: std_logic; attribute dont_touch of G5873: signal is true;
	signal G5874: std_logic; attribute dont_touch of G5874: signal is true;
	signal G5894: std_logic; attribute dont_touch of G5894: signal is true;
	signal G5897: std_logic; attribute dont_touch of G5897: signal is true;
	signal G5916: std_logic; attribute dont_touch of G5916: signal is true;
	signal G5917: std_logic; attribute dont_touch of G5917: signal is true;
	signal G5918: std_logic; attribute dont_touch of G5918: signal is true;
	signal G5937: std_logic; attribute dont_touch of G5937: signal is true;
	signal G5938: std_logic; attribute dont_touch of G5938: signal is true;
	signal G5939: std_logic; attribute dont_touch of G5939: signal is true;
	signal G5956: std_logic; attribute dont_touch of G5956: signal is true;
	signal G5969: std_logic; attribute dont_touch of G5969: signal is true;
	signal G5970: std_logic; attribute dont_touch of G5970: signal is true;
	signal G5971: std_logic; attribute dont_touch of G5971: signal is true;
	signal G5984: std_logic; attribute dont_touch of G5984: signal is true;
	signal G5987: std_logic; attribute dont_touch of G5987: signal is true;
	signal G5988: std_logic; attribute dont_touch of G5988: signal is true;
	signal G6001: std_logic; attribute dont_touch of G6001: signal is true;
	signal G6002: std_logic; attribute dont_touch of G6002: signal is true;
	signal G6003: std_logic; attribute dont_touch of G6003: signal is true;
	signal G6004: std_logic; attribute dont_touch of G6004: signal is true;
	signal G6005: std_logic; attribute dont_touch of G6005: signal is true;
	signal G6006: std_logic; attribute dont_touch of G6006: signal is true;
	signal G6007: std_logic; attribute dont_touch of G6007: signal is true;
	signal G6008: std_logic; attribute dont_touch of G6008: signal is true;
	signal G6009: std_logic; attribute dont_touch of G6009: signal is true;
	signal G6010: std_logic; attribute dont_touch of G6010: signal is true;
	signal G6011: std_logic; attribute dont_touch of G6011: signal is true;
	signal G6012: std_logic; attribute dont_touch of G6012: signal is true;
	signal G6013: std_logic; attribute dont_touch of G6013: signal is true;
	signal G6014: std_logic; attribute dont_touch of G6014: signal is true;
	signal G6015: std_logic; attribute dont_touch of G6015: signal is true;
	signal G6018: std_logic; attribute dont_touch of G6018: signal is true;
	signal G6019: std_logic; attribute dont_touch of G6019: signal is true;
	signal G6020: std_logic; attribute dont_touch of G6020: signal is true;
	signal G6021: std_logic; attribute dont_touch of G6021: signal is true;
	signal G6022: std_logic; attribute dont_touch of G6022: signal is true;
	signal G6023: std_logic; attribute dont_touch of G6023: signal is true;
	signal G6024: std_logic; attribute dont_touch of G6024: signal is true;
	signal G6025: std_logic; attribute dont_touch of G6025: signal is true;
	signal G6026: std_logic; attribute dont_touch of G6026: signal is true;
	signal G6027: std_logic; attribute dont_touch of G6027: signal is true;
	signal G6028: std_logic; attribute dont_touch of G6028: signal is true;
	signal G6032: std_logic; attribute dont_touch of G6032: signal is true;
	signal G6033: std_logic; attribute dont_touch of G6033: signal is true;
	signal G6034: std_logic; attribute dont_touch of G6034: signal is true;
	signal G6035: std_logic; attribute dont_touch of G6035: signal is true;
	signal G6036: std_logic; attribute dont_touch of G6036: signal is true;
	signal G6037: std_logic; attribute dont_touch of G6037: signal is true;
	signal G6038: std_logic; attribute dont_touch of G6038: signal is true;
	signal G6039: std_logic; attribute dont_touch of G6039: signal is true;
	signal G6040: std_logic; attribute dont_touch of G6040: signal is true;
	signal G6041: std_logic; attribute dont_touch of G6041: signal is true;
	signal G6042: std_logic; attribute dont_touch of G6042: signal is true;
	signal G6043: std_logic; attribute dont_touch of G6043: signal is true;
	signal G6044: std_logic; attribute dont_touch of G6044: signal is true;
	signal G6045: std_logic; attribute dont_touch of G6045: signal is true;
	signal G6046: std_logic; attribute dont_touch of G6046: signal is true;
	signal G6047: std_logic; attribute dont_touch of G6047: signal is true;
	signal G6048: std_logic; attribute dont_touch of G6048: signal is true;
	signal G6049: std_logic; attribute dont_touch of G6049: signal is true;
	signal G6050: std_logic; attribute dont_touch of G6050: signal is true;
	signal G6051: std_logic; attribute dont_touch of G6051: signal is true;
	signal G6052: std_logic; attribute dont_touch of G6052: signal is true;
	signal G6053: std_logic; attribute dont_touch of G6053: signal is true;
	signal G6054: std_logic; attribute dont_touch of G6054: signal is true;
	signal G6055: std_logic; attribute dont_touch of G6055: signal is true;
	signal G6056: std_logic; attribute dont_touch of G6056: signal is true;
	signal G6057: std_logic; attribute dont_touch of G6057: signal is true;
	signal G6058: std_logic; attribute dont_touch of G6058: signal is true;
	signal G6059: std_logic; attribute dont_touch of G6059: signal is true;
	signal G6060: std_logic; attribute dont_touch of G6060: signal is true;
	signal G6061: std_logic; attribute dont_touch of G6061: signal is true;
	signal G6062: std_logic; attribute dont_touch of G6062: signal is true;
	signal G6063: std_logic; attribute dont_touch of G6063: signal is true;
	signal G6064: std_logic; attribute dont_touch of G6064: signal is true;
	signal G6065: std_logic; attribute dont_touch of G6065: signal is true;
	signal G6068: std_logic; attribute dont_touch of G6068: signal is true;
	signal G6069: std_logic; attribute dont_touch of G6069: signal is true;
	signal G6070: std_logic; attribute dont_touch of G6070: signal is true;
	signal G6071: std_logic; attribute dont_touch of G6071: signal is true;
	signal G6072: std_logic; attribute dont_touch of G6072: signal is true;
	signal G6073: std_logic; attribute dont_touch of G6073: signal is true;
	signal G6074: std_logic; attribute dont_touch of G6074: signal is true;
	signal G6075: std_logic; attribute dont_touch of G6075: signal is true;
	signal G6076: std_logic; attribute dont_touch of G6076: signal is true;
	signal G6083: std_logic; attribute dont_touch of G6083: signal is true;
	signal G6087: std_logic; attribute dont_touch of G6087: signal is true;
	signal G6088: std_logic; attribute dont_touch of G6088: signal is true;
	signal G6089: std_logic; attribute dont_touch of G6089: signal is true;
	signal G6090: std_logic; attribute dont_touch of G6090: signal is true;
	signal G6091: std_logic; attribute dont_touch of G6091: signal is true;
	signal G6092: std_logic; attribute dont_touch of G6092: signal is true;
	signal G6093: std_logic; attribute dont_touch of G6093: signal is true;
	signal G6094: std_logic; attribute dont_touch of G6094: signal is true;
	signal G6095: std_logic; attribute dont_touch of G6095: signal is true;
	signal G6096: std_logic; attribute dont_touch of G6096: signal is true;
	signal G6097: std_logic; attribute dont_touch of G6097: signal is true;
	signal G6098: std_logic; attribute dont_touch of G6098: signal is true;
	signal G6101: std_logic; attribute dont_touch of G6101: signal is true;
	signal G6102: std_logic; attribute dont_touch of G6102: signal is true;
	signal G6103: std_logic; attribute dont_touch of G6103: signal is true;
	signal G6104: std_logic; attribute dont_touch of G6104: signal is true;
	signal G6105: std_logic; attribute dont_touch of G6105: signal is true;
	signal G6106: std_logic; attribute dont_touch of G6106: signal is true;
	signal G6107: std_logic; attribute dont_touch of G6107: signal is true;
	signal G6108: std_logic; attribute dont_touch of G6108: signal is true;
	signal G6109: std_logic; attribute dont_touch of G6109: signal is true;
	signal G6110: std_logic; attribute dont_touch of G6110: signal is true;
	signal G6111: std_logic; attribute dont_touch of G6111: signal is true;
	signal G6112: std_logic; attribute dont_touch of G6112: signal is true;
	signal G6115: std_logic; attribute dont_touch of G6115: signal is true;
	signal G6116: std_logic; attribute dont_touch of G6116: signal is true;
	signal G6117: std_logic; attribute dont_touch of G6117: signal is true;
	signal G6118: std_logic; attribute dont_touch of G6118: signal is true;
	signal G6119: std_logic; attribute dont_touch of G6119: signal is true;
	signal G6120: std_logic; attribute dont_touch of G6120: signal is true;
	signal G6121: std_logic; attribute dont_touch of G6121: signal is true;
	signal G6122: std_logic; attribute dont_touch of G6122: signal is true;
	signal G6123: std_logic; attribute dont_touch of G6123: signal is true;
	signal G6124: std_logic; attribute dont_touch of G6124: signal is true;
	signal G6125: std_logic; attribute dont_touch of G6125: signal is true;
	signal G6129: std_logic; attribute dont_touch of G6129: signal is true;
	signal G6130: std_logic; attribute dont_touch of G6130: signal is true;
	signal G6131: std_logic; attribute dont_touch of G6131: signal is true;
	signal G6132: std_logic; attribute dont_touch of G6132: signal is true;
	signal G6133: std_logic; attribute dont_touch of G6133: signal is true;
	signal G6134: std_logic; attribute dont_touch of G6134: signal is true;
	signal G6135: std_logic; attribute dont_touch of G6135: signal is true;
	signal G6136: std_logic; attribute dont_touch of G6136: signal is true;
	signal G6137: std_logic; attribute dont_touch of G6137: signal is true;
	signal G6138: std_logic; attribute dont_touch of G6138: signal is true;
	signal G6139: std_logic; attribute dont_touch of G6139: signal is true;
	signal G6140: std_logic; attribute dont_touch of G6140: signal is true;
	signal G6141: std_logic; attribute dont_touch of G6141: signal is true;
	signal G6142: std_logic; attribute dont_touch of G6142: signal is true;
	signal G6143: std_logic; attribute dont_touch of G6143: signal is true;
	signal G6144: std_logic; attribute dont_touch of G6144: signal is true;
	signal G6145: std_logic; attribute dont_touch of G6145: signal is true;
	signal G6146: std_logic; attribute dont_touch of G6146: signal is true;
	signal G6147: std_logic; attribute dont_touch of G6147: signal is true;
	signal G6148: std_logic; attribute dont_touch of G6148: signal is true;
	signal G6149: std_logic; attribute dont_touch of G6149: signal is true;
	signal G6150: std_logic; attribute dont_touch of G6150: signal is true;
	signal G6151: std_logic; attribute dont_touch of G6151: signal is true;
	signal G6152: std_logic; attribute dont_touch of G6152: signal is true;
	signal G6153: std_logic; attribute dont_touch of G6153: signal is true;
	signal G6154: std_logic; attribute dont_touch of G6154: signal is true;
	signal G6155: std_logic; attribute dont_touch of G6155: signal is true;
	signal G6156: std_logic; attribute dont_touch of G6156: signal is true;
	signal G6157: std_logic; attribute dont_touch of G6157: signal is true;
	signal G6158: std_logic; attribute dont_touch of G6158: signal is true;
	signal G6159: std_logic; attribute dont_touch of G6159: signal is true;
	signal G6160: std_logic; attribute dont_touch of G6160: signal is true;
	signal G6161: std_logic; attribute dont_touch of G6161: signal is true;
	signal G6162: std_logic; attribute dont_touch of G6162: signal is true;
	signal G6163: std_logic; attribute dont_touch of G6163: signal is true;
	signal G6164: std_logic; attribute dont_touch of G6164: signal is true;
	signal G6165: std_logic; attribute dont_touch of G6165: signal is true;
	signal G6166: std_logic; attribute dont_touch of G6166: signal is true;
	signal G6167: std_logic; attribute dont_touch of G6167: signal is true;
	signal G6168: std_logic; attribute dont_touch of G6168: signal is true;
	signal G6169: std_logic; attribute dont_touch of G6169: signal is true;
	signal G6170: std_logic; attribute dont_touch of G6170: signal is true;
	signal G6171: std_logic; attribute dont_touch of G6171: signal is true;
	signal G6172: std_logic; attribute dont_touch of G6172: signal is true;
	signal G6173: std_logic; attribute dont_touch of G6173: signal is true;
	signal G6174: std_logic; attribute dont_touch of G6174: signal is true;
	signal G6175: std_logic; attribute dont_touch of G6175: signal is true;
	signal G6176: std_logic; attribute dont_touch of G6176: signal is true;
	signal G6177: std_logic; attribute dont_touch of G6177: signal is true;
	signal G6178: std_logic; attribute dont_touch of G6178: signal is true;
	signal G6179: std_logic; attribute dont_touch of G6179: signal is true;
	signal G6180: std_logic; attribute dont_touch of G6180: signal is true;
	signal G6181: std_logic; attribute dont_touch of G6181: signal is true;
	signal G6182: std_logic; attribute dont_touch of G6182: signal is true;
	signal G6183: std_logic; attribute dont_touch of G6183: signal is true;
	signal G6184: std_logic; attribute dont_touch of G6184: signal is true;
	signal G6185: std_logic; attribute dont_touch of G6185: signal is true;
	signal G6186: std_logic; attribute dont_touch of G6186: signal is true;
	signal G6187: std_logic; attribute dont_touch of G6187: signal is true;
	signal G6188: std_logic; attribute dont_touch of G6188: signal is true;
	signal G6189: std_logic; attribute dont_touch of G6189: signal is true;
	signal G6190: std_logic; attribute dont_touch of G6190: signal is true;
	signal G6193: std_logic; attribute dont_touch of G6193: signal is true;
	signal G6194: std_logic; attribute dont_touch of G6194: signal is true;
	signal G6195: std_logic; attribute dont_touch of G6195: signal is true;
	signal G6196: std_logic; attribute dont_touch of G6196: signal is true;
	signal G6197: std_logic; attribute dont_touch of G6197: signal is true;
	signal G6198: std_logic; attribute dont_touch of G6198: signal is true;
	signal G6201: std_logic; attribute dont_touch of G6201: signal is true;
	signal G6202: std_logic; attribute dont_touch of G6202: signal is true;
	signal G6203: std_logic; attribute dont_touch of G6203: signal is true;
	signal G6204: std_logic; attribute dont_touch of G6204: signal is true;
	signal G6205: std_logic; attribute dont_touch of G6205: signal is true;
	signal G6206: std_logic; attribute dont_touch of G6206: signal is true;
	signal G6208: std_logic; attribute dont_touch of G6208: signal is true;
	signal G6209: std_logic; attribute dont_touch of G6209: signal is true;
	signal G6210: std_logic; attribute dont_touch of G6210: signal is true;
	signal G6211: std_logic; attribute dont_touch of G6211: signal is true;
	signal G6213: std_logic; attribute dont_touch of G6213: signal is true;
	signal G6214: std_logic; attribute dont_touch of G6214: signal is true;
	signal G6215: std_logic; attribute dont_touch of G6215: signal is true;
	signal G6216: std_logic; attribute dont_touch of G6216: signal is true;
	signal G6217: std_logic; attribute dont_touch of G6217: signal is true;
	signal G6218: std_logic; attribute dont_touch of G6218: signal is true;
	signal G6219: std_logic; attribute dont_touch of G6219: signal is true;
	signal G6220: std_logic; attribute dont_touch of G6220: signal is true;
	signal G6221: std_logic; attribute dont_touch of G6221: signal is true;
	signal G6222: std_logic; attribute dont_touch of G6222: signal is true;
	signal G6224: std_logic; attribute dont_touch of G6224: signal is true;
	signal G6225: std_logic; attribute dont_touch of G6225: signal is true;
	signal G6226: std_logic; attribute dont_touch of G6226: signal is true;
	signal G6227: std_logic; attribute dont_touch of G6227: signal is true;
	signal G6228: std_logic; attribute dont_touch of G6228: signal is true;
	signal G6229: std_logic; attribute dont_touch of G6229: signal is true;
	signal G6230: std_logic; attribute dont_touch of G6230: signal is true;
	signal G6231: std_logic; attribute dont_touch of G6231: signal is true;
	signal G6232: std_logic; attribute dont_touch of G6232: signal is true;
	signal G6235: std_logic; attribute dont_touch of G6235: signal is true;
	signal G6237: std_logic; attribute dont_touch of G6237: signal is true;
	signal G6238: std_logic; attribute dont_touch of G6238: signal is true;
	signal G6239: std_logic; attribute dont_touch of G6239: signal is true;
	signal G6242: std_logic; attribute dont_touch of G6242: signal is true;
	signal G6243: std_logic; attribute dont_touch of G6243: signal is true;
	signal G6244: std_logic; attribute dont_touch of G6244: signal is true;
	signal G6245: std_logic; attribute dont_touch of G6245: signal is true;
	signal G6246: std_logic; attribute dont_touch of G6246: signal is true;
	signal G6249: std_logic; attribute dont_touch of G6249: signal is true;
	signal G6250: std_logic; attribute dont_touch of G6250: signal is true;
	signal G6251: std_logic; attribute dont_touch of G6251: signal is true;
	signal G6252: std_logic; attribute dont_touch of G6252: signal is true;
	signal G6253: std_logic; attribute dont_touch of G6253: signal is true;
	signal G6254: std_logic; attribute dont_touch of G6254: signal is true;
	signal G6255: std_logic; attribute dont_touch of G6255: signal is true;
	signal G6256: std_logic; attribute dont_touch of G6256: signal is true;
	signal G6257: std_logic; attribute dont_touch of G6257: signal is true;
	signal G6258: std_logic; attribute dont_touch of G6258: signal is true;
	signal G6259: std_logic; attribute dont_touch of G6259: signal is true;
	signal G6262: std_logic; attribute dont_touch of G6262: signal is true;
	signal G6263: std_logic; attribute dont_touch of G6263: signal is true;
	signal G6264: std_logic; attribute dont_touch of G6264: signal is true;
	signal G6265: std_logic; attribute dont_touch of G6265: signal is true;
	signal G6266: std_logic; attribute dont_touch of G6266: signal is true;
	signal G6267: std_logic; attribute dont_touch of G6267: signal is true;
	signal G6268: std_logic; attribute dont_touch of G6268: signal is true;
	signal G6270: std_logic; attribute dont_touch of G6270: signal is true;
	signal G6273: std_logic; attribute dont_touch of G6273: signal is true;
	signal G6274: std_logic; attribute dont_touch of G6274: signal is true;
	signal G6275: std_logic; attribute dont_touch of G6275: signal is true;
	signal G6276: std_logic; attribute dont_touch of G6276: signal is true;
	signal G6277: std_logic; attribute dont_touch of G6277: signal is true;
	signal G6278: std_logic; attribute dont_touch of G6278: signal is true;
	signal G6279: std_logic; attribute dont_touch of G6279: signal is true;
	signal G6280: std_logic; attribute dont_touch of G6280: signal is true;
	signal G6281: std_logic; attribute dont_touch of G6281: signal is true;
	signal G6282: std_logic; attribute dont_touch of G6282: signal is true;
	signal G6283: std_logic; attribute dont_touch of G6283: signal is true;
	signal G6284: std_logic; attribute dont_touch of G6284: signal is true;
	signal G6285: std_logic; attribute dont_touch of G6285: signal is true;
	signal G6286: std_logic; attribute dont_touch of G6286: signal is true;
	signal G6287: std_logic; attribute dont_touch of G6287: signal is true;
	signal G6309: std_logic; attribute dont_touch of G6309: signal is true;
	signal G6310: std_logic; attribute dont_touch of G6310: signal is true;
	signal G6311: std_logic; attribute dont_touch of G6311: signal is true;
	signal G6312: std_logic; attribute dont_touch of G6312: signal is true;
	signal G6313: std_logic; attribute dont_touch of G6313: signal is true;
	signal G6314: std_logic; attribute dont_touch of G6314: signal is true;
	signal G6315: std_logic; attribute dont_touch of G6315: signal is true;
	signal G6316: std_logic; attribute dont_touch of G6316: signal is true;
	signal G6317: std_logic; attribute dont_touch of G6317: signal is true;
	signal G6318: std_logic; attribute dont_touch of G6318: signal is true;
	signal G6319: std_logic; attribute dont_touch of G6319: signal is true;
	signal G6320: std_logic; attribute dont_touch of G6320: signal is true;
	signal G6321: std_logic; attribute dont_touch of G6321: signal is true;
	signal G6322: std_logic; attribute dont_touch of G6322: signal is true;
	signal G6323: std_logic; attribute dont_touch of G6323: signal is true;
	signal G6324: std_logic; attribute dont_touch of G6324: signal is true;
	signal G6325: std_logic; attribute dont_touch of G6325: signal is true;
	signal G6326: std_logic; attribute dont_touch of G6326: signal is true;
	signal G6327: std_logic; attribute dont_touch of G6327: signal is true;
	signal G6328: std_logic; attribute dont_touch of G6328: signal is true;
	signal G6329: std_logic; attribute dont_touch of G6329: signal is true;
	signal G6330: std_logic; attribute dont_touch of G6330: signal is true;
	signal G6331: std_logic; attribute dont_touch of G6331: signal is true;
	signal G6332: std_logic; attribute dont_touch of G6332: signal is true;
	signal G6333: std_logic; attribute dont_touch of G6333: signal is true;
	signal G6334: std_logic; attribute dont_touch of G6334: signal is true;
	signal G6335: std_logic; attribute dont_touch of G6335: signal is true;
	signal G6336: std_logic; attribute dont_touch of G6336: signal is true;
	signal G6337: std_logic; attribute dont_touch of G6337: signal is true;
	signal G6338: std_logic; attribute dont_touch of G6338: signal is true;
	signal G6339: std_logic; attribute dont_touch of G6339: signal is true;
	signal G6340: std_logic; attribute dont_touch of G6340: signal is true;
	signal G6341: std_logic; attribute dont_touch of G6341: signal is true;
	signal G6342: std_logic; attribute dont_touch of G6342: signal is true;
	signal G6343: std_logic; attribute dont_touch of G6343: signal is true;
	signal G6344: std_logic; attribute dont_touch of G6344: signal is true;
	signal G6345: std_logic; attribute dont_touch of G6345: signal is true;
	signal G6346: std_logic; attribute dont_touch of G6346: signal is true;
	signal G6347: std_logic; attribute dont_touch of G6347: signal is true;
	signal G6348: std_logic; attribute dont_touch of G6348: signal is true;
	signal G6349: std_logic; attribute dont_touch of G6349: signal is true;
	signal G6350: std_logic; attribute dont_touch of G6350: signal is true;
	signal G6351: std_logic; attribute dont_touch of G6351: signal is true;
	signal G6352: std_logic; attribute dont_touch of G6352: signal is true;
	signal G6353: std_logic; attribute dont_touch of G6353: signal is true;
	signal G6354: std_logic; attribute dont_touch of G6354: signal is true;
	signal G6355: std_logic; attribute dont_touch of G6355: signal is true;
	signal G6356: std_logic; attribute dont_touch of G6356: signal is true;
	signal G6357: std_logic; attribute dont_touch of G6357: signal is true;
	signal G6358: std_logic; attribute dont_touch of G6358: signal is true;
	signal G6359: std_logic; attribute dont_touch of G6359: signal is true;
	signal G6360: std_logic; attribute dont_touch of G6360: signal is true;
	signal G6361: std_logic; attribute dont_touch of G6361: signal is true;
	signal G6362: std_logic; attribute dont_touch of G6362: signal is true;
	signal G6363: std_logic; attribute dont_touch of G6363: signal is true;
	signal G6364: std_logic; attribute dont_touch of G6364: signal is true;
	signal G6365: std_logic; attribute dont_touch of G6365: signal is true;
	signal G6366: std_logic; attribute dont_touch of G6366: signal is true;
	signal G6367: std_logic; attribute dont_touch of G6367: signal is true;
	signal G6368: std_logic; attribute dont_touch of G6368: signal is true;
	signal G6369: std_logic; attribute dont_touch of G6369: signal is true;
	signal G6370: std_logic; attribute dont_touch of G6370: signal is true;
	signal G6371: std_logic; attribute dont_touch of G6371: signal is true;
	signal G6372: std_logic; attribute dont_touch of G6372: signal is true;
	signal G6373: std_logic; attribute dont_touch of G6373: signal is true;
	signal G6374: std_logic; attribute dont_touch of G6374: signal is true;
	signal G6375: std_logic; attribute dont_touch of G6375: signal is true;
	signal G6377: std_logic; attribute dont_touch of G6377: signal is true;
	signal G6378: std_logic; attribute dont_touch of G6378: signal is true;
	signal G6379: std_logic; attribute dont_touch of G6379: signal is true;
	signal G6380: std_logic; attribute dont_touch of G6380: signal is true;
	signal G6381: std_logic; attribute dont_touch of G6381: signal is true;
	signal G6382: std_logic; attribute dont_touch of G6382: signal is true;
	signal G6383: std_logic; attribute dont_touch of G6383: signal is true;
	signal G6384: std_logic; attribute dont_touch of G6384: signal is true;
	signal G6385: std_logic; attribute dont_touch of G6385: signal is true;
	signal G6386: std_logic; attribute dont_touch of G6386: signal is true;
	signal G6387: std_logic; attribute dont_touch of G6387: signal is true;
	signal G6388: std_logic; attribute dont_touch of G6388: signal is true;
	signal G6389: std_logic; attribute dont_touch of G6389: signal is true;
	signal G6390: std_logic; attribute dont_touch of G6390: signal is true;
	signal G6391: std_logic; attribute dont_touch of G6391: signal is true;
	signal G6392: std_logic; attribute dont_touch of G6392: signal is true;
	signal G6393: std_logic; attribute dont_touch of G6393: signal is true;
	signal G6394: std_logic; attribute dont_touch of G6394: signal is true;
	signal G6395: std_logic; attribute dont_touch of G6395: signal is true;
	signal G6396: std_logic; attribute dont_touch of G6396: signal is true;
	signal G6397: std_logic; attribute dont_touch of G6397: signal is true;
	signal G6398: std_logic; attribute dont_touch of G6398: signal is true;
	signal G6399: std_logic; attribute dont_touch of G6399: signal is true;
	signal G6400: std_logic; attribute dont_touch of G6400: signal is true;
	signal G6401: std_logic; attribute dont_touch of G6401: signal is true;
	signal G6402: std_logic; attribute dont_touch of G6402: signal is true;
	signal G6403: std_logic; attribute dont_touch of G6403: signal is true;
	signal G6404: std_logic; attribute dont_touch of G6404: signal is true;
	signal G6405: std_logic; attribute dont_touch of G6405: signal is true;
	signal G6406: std_logic; attribute dont_touch of G6406: signal is true;
	signal G6407: std_logic; attribute dont_touch of G6407: signal is true;
	signal G6408: std_logic; attribute dont_touch of G6408: signal is true;
	signal G6409: std_logic; attribute dont_touch of G6409: signal is true;
	signal G6410: std_logic; attribute dont_touch of G6410: signal is true;
	signal G6411: std_logic; attribute dont_touch of G6411: signal is true;
	signal G6412: std_logic; attribute dont_touch of G6412: signal is true;
	signal G6413: std_logic; attribute dont_touch of G6413: signal is true;
	signal G6414: std_logic; attribute dont_touch of G6414: signal is true;
	signal G6415: std_logic; attribute dont_touch of G6415: signal is true;
	signal G6416: std_logic; attribute dont_touch of G6416: signal is true;
	signal G6417: std_logic; attribute dont_touch of G6417: signal is true;
	signal G6418: std_logic; attribute dont_touch of G6418: signal is true;
	signal G6419: std_logic; attribute dont_touch of G6419: signal is true;
	signal G6420: std_logic; attribute dont_touch of G6420: signal is true;
	signal G6421: std_logic; attribute dont_touch of G6421: signal is true;
	signal G6422: std_logic; attribute dont_touch of G6422: signal is true;
	signal G6423: std_logic; attribute dont_touch of G6423: signal is true;
	signal G6424: std_logic; attribute dont_touch of G6424: signal is true;
	signal G6426: std_logic; attribute dont_touch of G6426: signal is true;
	signal G6427: std_logic; attribute dont_touch of G6427: signal is true;
	signal G6428: std_logic; attribute dont_touch of G6428: signal is true;
	signal G6429: std_logic; attribute dont_touch of G6429: signal is true;
	signal G6430: std_logic; attribute dont_touch of G6430: signal is true;
	signal G6431: std_logic; attribute dont_touch of G6431: signal is true;
	signal G6432: std_logic; attribute dont_touch of G6432: signal is true;
	signal G6433: std_logic; attribute dont_touch of G6433: signal is true;
	signal G6434: std_logic; attribute dont_touch of G6434: signal is true;
	signal G6435: std_logic; attribute dont_touch of G6435: signal is true;
	signal G6436: std_logic; attribute dont_touch of G6436: signal is true;
	signal G6437: std_logic; attribute dont_touch of G6437: signal is true;
	signal G6438: std_logic; attribute dont_touch of G6438: signal is true;
	signal G6439: std_logic; attribute dont_touch of G6439: signal is true;
	signal G6440: std_logic; attribute dont_touch of G6440: signal is true;
	signal G6441: std_logic; attribute dont_touch of G6441: signal is true;
	signal G6444: std_logic; attribute dont_touch of G6444: signal is true;
	signal G6445: std_logic; attribute dont_touch of G6445: signal is true;
	signal G6446: std_logic; attribute dont_touch of G6446: signal is true;
	signal G6447: std_logic; attribute dont_touch of G6447: signal is true;
	signal G6448: std_logic; attribute dont_touch of G6448: signal is true;
	signal G6449: std_logic; attribute dont_touch of G6449: signal is true;
	signal G6452: std_logic; attribute dont_touch of G6452: signal is true;
	signal G6456: std_logic; attribute dont_touch of G6456: signal is true;
	signal G6457: std_logic; attribute dont_touch of G6457: signal is true;
	signal G6458: std_logic; attribute dont_touch of G6458: signal is true;
	signal G6459: std_logic; attribute dont_touch of G6459: signal is true;
	signal G6460: std_logic; attribute dont_touch of G6460: signal is true;
	signal G6461: std_logic; attribute dont_touch of G6461: signal is true;
	signal G6462: std_logic; attribute dont_touch of G6462: signal is true;
	signal G6463: std_logic; attribute dont_touch of G6463: signal is true;
	signal G6464: std_logic; attribute dont_touch of G6464: signal is true;
	signal G6465: std_logic; attribute dont_touch of G6465: signal is true;
	signal G6466: std_logic; attribute dont_touch of G6466: signal is true;
	signal G6467: std_logic; attribute dont_touch of G6467: signal is true;
	signal G6468: std_logic; attribute dont_touch of G6468: signal is true;
	signal G6469: std_logic; attribute dont_touch of G6469: signal is true;
	signal G6470: std_logic; attribute dont_touch of G6470: signal is true;
	signal G6471: std_logic; attribute dont_touch of G6471: signal is true;
	signal G6472: std_logic; attribute dont_touch of G6472: signal is true;
	signal G6473: std_logic; attribute dont_touch of G6473: signal is true;
	signal G6474: std_logic; attribute dont_touch of G6474: signal is true;
	signal G6475: std_logic; attribute dont_touch of G6475: signal is true;
	signal G6476: std_logic; attribute dont_touch of G6476: signal is true;
	signal G6477: std_logic; attribute dont_touch of G6477: signal is true;
	signal G6478: std_logic; attribute dont_touch of G6478: signal is true;
	signal G6481: std_logic; attribute dont_touch of G6481: signal is true;
	signal G6482: std_logic; attribute dont_touch of G6482: signal is true;
	signal G6483: std_logic; attribute dont_touch of G6483: signal is true;
	signal G6486: std_logic; attribute dont_touch of G6486: signal is true;
	signal G6487: std_logic; attribute dont_touch of G6487: signal is true;
	signal G6488: std_logic; attribute dont_touch of G6488: signal is true;
	signal G6489: std_logic; attribute dont_touch of G6489: signal is true;
	signal G6490: std_logic; attribute dont_touch of G6490: signal is true;
	signal G6493: std_logic; attribute dont_touch of G6493: signal is true;
	signal G6496: std_logic; attribute dont_touch of G6496: signal is true;
	signal G6497: std_logic; attribute dont_touch of G6497: signal is true;
	signal G6498: std_logic; attribute dont_touch of G6498: signal is true;
	signal G6501: std_logic; attribute dont_touch of G6501: signal is true;
	signal G6502: std_logic; attribute dont_touch of G6502: signal is true;
	signal G6503: std_logic; attribute dont_touch of G6503: signal is true;
	signal G6504: std_logic; attribute dont_touch of G6504: signal is true;
	signal G6505: std_logic; attribute dont_touch of G6505: signal is true;
	signal G6506: std_logic; attribute dont_touch of G6506: signal is true;
	signal G6507: std_logic; attribute dont_touch of G6507: signal is true;
	signal G6508: std_logic; attribute dont_touch of G6508: signal is true;
	signal G6509: std_logic; attribute dont_touch of G6509: signal is true;
	signal G6510: std_logic; attribute dont_touch of G6510: signal is true;
	signal G6511: std_logic; attribute dont_touch of G6511: signal is true;
	signal G6514: std_logic; attribute dont_touch of G6514: signal is true;
	signal G6515: std_logic; attribute dont_touch of G6515: signal is true;
	signal G6516: std_logic; attribute dont_touch of G6516: signal is true;
	signal G6517: std_logic; attribute dont_touch of G6517: signal is true;
	signal G6520: std_logic; attribute dont_touch of G6520: signal is true;
	signal G6523: std_logic; attribute dont_touch of G6523: signal is true;
	signal G6524: std_logic; attribute dont_touch of G6524: signal is true;
	signal G6525: std_logic; attribute dont_touch of G6525: signal is true;
	signal G6538: std_logic; attribute dont_touch of G6538: signal is true;
	signal G6541: std_logic; attribute dont_touch of G6541: signal is true;
	signal G6542: std_logic; attribute dont_touch of G6542: signal is true;
	signal G6543: std_logic; attribute dont_touch of G6543: signal is true;
	signal G6552: std_logic; attribute dont_touch of G6552: signal is true;
	signal G6553: std_logic; attribute dont_touch of G6553: signal is true;
	signal G6554: std_logic; attribute dont_touch of G6554: signal is true;
	signal G6555: std_logic; attribute dont_touch of G6555: signal is true;
	signal G6556: std_logic; attribute dont_touch of G6556: signal is true;
	signal G6559: std_logic; attribute dont_touch of G6559: signal is true;
	signal G6562: std_logic; attribute dont_touch of G6562: signal is true;
	signal G6565: std_logic; attribute dont_touch of G6565: signal is true;
	signal G6566: std_logic; attribute dont_touch of G6566: signal is true;
	signal G6567: std_logic; attribute dont_touch of G6567: signal is true;
	signal G6568: std_logic; attribute dont_touch of G6568: signal is true;
	signal G6569: std_logic; attribute dont_touch of G6569: signal is true;
	signal G6570: std_logic; attribute dont_touch of G6570: signal is true;
	signal G6571: std_logic; attribute dont_touch of G6571: signal is true;
	signal G6572: std_logic; attribute dont_touch of G6572: signal is true;
	signal G6573: std_logic; attribute dont_touch of G6573: signal is true;
	signal G6574: std_logic; attribute dont_touch of G6574: signal is true;
	signal G6577: std_logic; attribute dont_touch of G6577: signal is true;
	signal G6578: std_logic; attribute dont_touch of G6578: signal is true;
	signal G6579: std_logic; attribute dont_touch of G6579: signal is true;
	signal G6580: std_logic; attribute dont_touch of G6580: signal is true;
	signal G6581: std_logic; attribute dont_touch of G6581: signal is true;
	signal G6582: std_logic; attribute dont_touch of G6582: signal is true;
	signal G6585: std_logic; attribute dont_touch of G6585: signal is true;
	signal G6586: std_logic; attribute dont_touch of G6586: signal is true;
	signal G6587: std_logic; attribute dont_touch of G6587: signal is true;
	signal G6588: std_logic; attribute dont_touch of G6588: signal is true;
	signal G6589: std_logic; attribute dont_touch of G6589: signal is true;
	signal G6590: std_logic; attribute dont_touch of G6590: signal is true;
	signal G6591: std_logic; attribute dont_touch of G6591: signal is true;
	signal G6592: std_logic; attribute dont_touch of G6592: signal is true;
	signal G6593: std_logic; attribute dont_touch of G6593: signal is true;
	signal G6594: std_logic; attribute dont_touch of G6594: signal is true;
	signal G6595: std_logic; attribute dont_touch of G6595: signal is true;
	signal G6596: std_logic; attribute dont_touch of G6596: signal is true;
	signal G6597: std_logic; attribute dont_touch of G6597: signal is true;
	signal G6598: std_logic; attribute dont_touch of G6598: signal is true;
	signal G6599: std_logic; attribute dont_touch of G6599: signal is true;
	signal G6600: std_logic; attribute dont_touch of G6600: signal is true;
	signal G6601: std_logic; attribute dont_touch of G6601: signal is true;
	signal G6602: std_logic; attribute dont_touch of G6602: signal is true;
	signal G6603: std_logic; attribute dont_touch of G6603: signal is true;
	signal G6604: std_logic; attribute dont_touch of G6604: signal is true;
	signal G6605: std_logic; attribute dont_touch of G6605: signal is true;
	signal G6606: std_logic; attribute dont_touch of G6606: signal is true;
	signal G6607: std_logic; attribute dont_touch of G6607: signal is true;
	signal G6610: std_logic; attribute dont_touch of G6610: signal is true;
	signal G6611: std_logic; attribute dont_touch of G6611: signal is true;
	signal G6612: std_logic; attribute dont_touch of G6612: signal is true;
	signal G6613: std_logic; attribute dont_touch of G6613: signal is true;
	signal G6614: std_logic; attribute dont_touch of G6614: signal is true;
	signal G6615: std_logic; attribute dont_touch of G6615: signal is true;
	signal G6616: std_logic; attribute dont_touch of G6616: signal is true;
	signal G6617: std_logic; attribute dont_touch of G6617: signal is true;
	signal G6618: std_logic; attribute dont_touch of G6618: signal is true;
	signal G6621: std_logic; attribute dont_touch of G6621: signal is true;
	signal G6622: std_logic; attribute dont_touch of G6622: signal is true;
	signal G6623: std_logic; attribute dont_touch of G6623: signal is true;
	signal G6624: std_logic; attribute dont_touch of G6624: signal is true;
	signal G6625: std_logic; attribute dont_touch of G6625: signal is true;
	signal G6626: std_logic; attribute dont_touch of G6626: signal is true;
	signal G6627: std_logic; attribute dont_touch of G6627: signal is true;
	signal G6628: std_logic; attribute dont_touch of G6628: signal is true;
	signal G6629: std_logic; attribute dont_touch of G6629: signal is true;
	signal G6630: std_logic; attribute dont_touch of G6630: signal is true;
	signal G6631: std_logic; attribute dont_touch of G6631: signal is true;
	signal G6632: std_logic; attribute dont_touch of G6632: signal is true;
	signal G6633: std_logic; attribute dont_touch of G6633: signal is true;
	signal G6634: std_logic; attribute dont_touch of G6634: signal is true;
	signal G6635: std_logic; attribute dont_touch of G6635: signal is true;
	signal G6636: std_logic; attribute dont_touch of G6636: signal is true;
	signal G6637: std_logic; attribute dont_touch of G6637: signal is true;
	signal G6638: std_logic; attribute dont_touch of G6638: signal is true;
	signal G6639: std_logic; attribute dont_touch of G6639: signal is true;
	signal G6640: std_logic; attribute dont_touch of G6640: signal is true;
	signal G6641: std_logic; attribute dont_touch of G6641: signal is true;
	signal G6642: std_logic; attribute dont_touch of G6642: signal is true;
	signal G6643: std_logic; attribute dont_touch of G6643: signal is true;
	signal G6644: std_logic; attribute dont_touch of G6644: signal is true;
	signal G6645: std_logic; attribute dont_touch of G6645: signal is true;
	signal G6646: std_logic; attribute dont_touch of G6646: signal is true;
	signal G6647: std_logic; attribute dont_touch of G6647: signal is true;
	signal G6649: std_logic; attribute dont_touch of G6649: signal is true;
	signal G6650: std_logic; attribute dont_touch of G6650: signal is true;
	signal G6651: std_logic; attribute dont_touch of G6651: signal is true;
	signal G6652: std_logic; attribute dont_touch of G6652: signal is true;
	signal G6654: std_logic; attribute dont_touch of G6654: signal is true;
	signal G6655: std_logic; attribute dont_touch of G6655: signal is true;
	signal G6656: std_logic; attribute dont_touch of G6656: signal is true;
	signal G6657: std_logic; attribute dont_touch of G6657: signal is true;
	signal G6658: std_logic; attribute dont_touch of G6658: signal is true;
	signal G6659: std_logic; attribute dont_touch of G6659: signal is true;
	signal G6660: std_logic; attribute dont_touch of G6660: signal is true;
	signal G6661: std_logic; attribute dont_touch of G6661: signal is true;
	signal G6662: std_logic; attribute dont_touch of G6662: signal is true;
	signal G6663: std_logic; attribute dont_touch of G6663: signal is true;
	signal G6664: std_logic; attribute dont_touch of G6664: signal is true;
	signal G6671: std_logic; attribute dont_touch of G6671: signal is true;
	signal G6672: std_logic; attribute dont_touch of G6672: signal is true;
	signal G6673: std_logic; attribute dont_touch of G6673: signal is true;
	signal G6674: std_logic; attribute dont_touch of G6674: signal is true;
	signal G6676: std_logic; attribute dont_touch of G6676: signal is true;
	signal G6677: std_logic; attribute dont_touch of G6677: signal is true;
	signal G6680: std_logic; attribute dont_touch of G6680: signal is true;
	signal G6681: std_logic; attribute dont_touch of G6681: signal is true;
	signal G6682: std_logic; attribute dont_touch of G6682: signal is true;
	signal G6683: std_logic; attribute dont_touch of G6683: signal is true;
	signal G6684: std_logic; attribute dont_touch of G6684: signal is true;
	signal G6685: std_logic; attribute dont_touch of G6685: signal is true;
	signal G6686: std_logic; attribute dont_touch of G6686: signal is true;
	signal G6687: std_logic; attribute dont_touch of G6687: signal is true;
	signal G6688: std_logic; attribute dont_touch of G6688: signal is true;
	signal G6689: std_logic; attribute dont_touch of G6689: signal is true;
	signal G6692: std_logic; attribute dont_touch of G6692: signal is true;
	signal G6693: std_logic; attribute dont_touch of G6693: signal is true;
	signal G6694: std_logic; attribute dont_touch of G6694: signal is true;
	signal G6695: std_logic; attribute dont_touch of G6695: signal is true;
	signal G6696: std_logic; attribute dont_touch of G6696: signal is true;
	signal G6697: std_logic; attribute dont_touch of G6697: signal is true;
	signal G6698: std_logic; attribute dont_touch of G6698: signal is true;
	signal G6699: std_logic; attribute dont_touch of G6699: signal is true;
	signal G6700: std_logic; attribute dont_touch of G6700: signal is true;
	signal G6701: std_logic; attribute dont_touch of G6701: signal is true;
	signal G6702: std_logic; attribute dont_touch of G6702: signal is true;
	signal G6703: std_logic; attribute dont_touch of G6703: signal is true;
	signal G6704: std_logic; attribute dont_touch of G6704: signal is true;
	signal G6705: std_logic; attribute dont_touch of G6705: signal is true;
	signal G6706: std_logic; attribute dont_touch of G6706: signal is true;
	signal G6707: std_logic; attribute dont_touch of G6707: signal is true;
	signal G6708: std_logic; attribute dont_touch of G6708: signal is true;
	signal G6709: std_logic; attribute dont_touch of G6709: signal is true;
	signal G6710: std_logic; attribute dont_touch of G6710: signal is true;
	signal G6711: std_logic; attribute dont_touch of G6711: signal is true;
	signal G6712: std_logic; attribute dont_touch of G6712: signal is true;
	signal G6713: std_logic; attribute dont_touch of G6713: signal is true;
	signal G6714: std_logic; attribute dont_touch of G6714: signal is true;
	signal G6715: std_logic; attribute dont_touch of G6715: signal is true;
	signal G6716: std_logic; attribute dont_touch of G6716: signal is true;
	signal G6717: std_logic; attribute dont_touch of G6717: signal is true;
	signal G6718: std_logic; attribute dont_touch of G6718: signal is true;
	signal G6719: std_logic; attribute dont_touch of G6719: signal is true;
	signal G6720: std_logic; attribute dont_touch of G6720: signal is true;
	signal G6721: std_logic; attribute dont_touch of G6721: signal is true;
	signal G6722: std_logic; attribute dont_touch of G6722: signal is true;
	signal G6723: std_logic; attribute dont_touch of G6723: signal is true;
	signal G6724: std_logic; attribute dont_touch of G6724: signal is true;
	signal G6725: std_logic; attribute dont_touch of G6725: signal is true;
	signal G6726: std_logic; attribute dont_touch of G6726: signal is true;
	signal G6727: std_logic; attribute dont_touch of G6727: signal is true;
	signal G6728: std_logic; attribute dont_touch of G6728: signal is true;
	signal G6729: std_logic; attribute dont_touch of G6729: signal is true;
	signal G6730: std_logic; attribute dont_touch of G6730: signal is true;
	signal G6731: std_logic; attribute dont_touch of G6731: signal is true;
	signal G6732: std_logic; attribute dont_touch of G6732: signal is true;
	signal G6733: std_logic; attribute dont_touch of G6733: signal is true;
	signal G6734: std_logic; attribute dont_touch of G6734: signal is true;
	signal G6735: std_logic; attribute dont_touch of G6735: signal is true;
	signal G6736: std_logic; attribute dont_touch of G6736: signal is true;
	signal G6737: std_logic; attribute dont_touch of G6737: signal is true;
	signal G6738: std_logic; attribute dont_touch of G6738: signal is true;
	signal G6739: std_logic; attribute dont_touch of G6739: signal is true;
	signal G6740: std_logic; attribute dont_touch of G6740: signal is true;
	signal G6741: std_logic; attribute dont_touch of G6741: signal is true;
	signal G6742: std_logic; attribute dont_touch of G6742: signal is true;
	signal G6743: std_logic; attribute dont_touch of G6743: signal is true;
	signal G6744: std_logic; attribute dont_touch of G6744: signal is true;
	signal G6745: std_logic; attribute dont_touch of G6745: signal is true;
	signal G6751: std_logic; attribute dont_touch of G6751: signal is true;
	signal G6752: std_logic; attribute dont_touch of G6752: signal is true;
	signal G6753: std_logic; attribute dont_touch of G6753: signal is true;
	signal G6754: std_logic; attribute dont_touch of G6754: signal is true;
	signal G6755: std_logic; attribute dont_touch of G6755: signal is true;
	signal G6756: std_logic; attribute dont_touch of G6756: signal is true;
	signal G6757: std_logic; attribute dont_touch of G6757: signal is true;
	signal G6758: std_logic; attribute dont_touch of G6758: signal is true;
	signal G6759: std_logic; attribute dont_touch of G6759: signal is true;
	signal G6760: std_logic; attribute dont_touch of G6760: signal is true;
	signal G6761: std_logic; attribute dont_touch of G6761: signal is true;
	signal G6762: std_logic; attribute dont_touch of G6762: signal is true;
	signal G6763: std_logic; attribute dont_touch of G6763: signal is true;
	signal G6764: std_logic; attribute dont_touch of G6764: signal is true;
	signal G6765: std_logic; attribute dont_touch of G6765: signal is true;
	signal G6766: std_logic; attribute dont_touch of G6766: signal is true;
	signal G6767: std_logic; attribute dont_touch of G6767: signal is true;
	signal G6768: std_logic; attribute dont_touch of G6768: signal is true;
	signal G6769: std_logic; attribute dont_touch of G6769: signal is true;
	signal G6770: std_logic; attribute dont_touch of G6770: signal is true;
	signal G6771: std_logic; attribute dont_touch of G6771: signal is true;
	signal G6772: std_logic; attribute dont_touch of G6772: signal is true;
	signal G6773: std_logic; attribute dont_touch of G6773: signal is true;
	signal G6774: std_logic; attribute dont_touch of G6774: signal is true;
	signal G6775: std_logic; attribute dont_touch of G6775: signal is true;
	signal G6776: std_logic; attribute dont_touch of G6776: signal is true;
	signal G6777: std_logic; attribute dont_touch of G6777: signal is true;
	signal G6778: std_logic; attribute dont_touch of G6778: signal is true;
	signal G6779: std_logic; attribute dont_touch of G6779: signal is true;
	signal G6780: std_logic; attribute dont_touch of G6780: signal is true;
	signal G6781: std_logic; attribute dont_touch of G6781: signal is true;
	signal G6782: std_logic; attribute dont_touch of G6782: signal is true;
	signal G6783: std_logic; attribute dont_touch of G6783: signal is true;
	signal G6784: std_logic; attribute dont_touch of G6784: signal is true;
	signal G6785: std_logic; attribute dont_touch of G6785: signal is true;
	signal G6786: std_logic; attribute dont_touch of G6786: signal is true;
	signal G6787: std_logic; attribute dont_touch of G6787: signal is true;
	signal G6788: std_logic; attribute dont_touch of G6788: signal is true;
	signal G6789: std_logic; attribute dont_touch of G6789: signal is true;
	signal G6790: std_logic; attribute dont_touch of G6790: signal is true;
	signal G6791: std_logic; attribute dont_touch of G6791: signal is true;
	signal G6792: std_logic; attribute dont_touch of G6792: signal is true;
	signal G6793: std_logic; attribute dont_touch of G6793: signal is true;
	signal G6794: std_logic; attribute dont_touch of G6794: signal is true;
	signal G6795: std_logic; attribute dont_touch of G6795: signal is true;
	signal G6796: std_logic; attribute dont_touch of G6796: signal is true;
	signal G6797: std_logic; attribute dont_touch of G6797: signal is true;
	signal G6798: std_logic; attribute dont_touch of G6798: signal is true;
	signal G6799: std_logic; attribute dont_touch of G6799: signal is true;
	signal G6800: std_logic; attribute dont_touch of G6800: signal is true;
	signal G6801: std_logic; attribute dont_touch of G6801: signal is true;
	signal G6802: std_logic; attribute dont_touch of G6802: signal is true;
	signal G6803: std_logic; attribute dont_touch of G6803: signal is true;
	signal G6804: std_logic; attribute dont_touch of G6804: signal is true;
	signal G6805: std_logic; attribute dont_touch of G6805: signal is true;
	signal G6806: std_logic; attribute dont_touch of G6806: signal is true;
	signal G6807: std_logic; attribute dont_touch of G6807: signal is true;
	signal G6808: std_logic; attribute dont_touch of G6808: signal is true;
	signal G6809: std_logic; attribute dont_touch of G6809: signal is true;
	signal G6810: std_logic; attribute dont_touch of G6810: signal is true;
	signal G6811: std_logic; attribute dont_touch of G6811: signal is true;
	signal G6812: std_logic; attribute dont_touch of G6812: signal is true;
	signal G6813: std_logic; attribute dont_touch of G6813: signal is true;
	signal G6814: std_logic; attribute dont_touch of G6814: signal is true;
	signal G6815: std_logic; attribute dont_touch of G6815: signal is true;
	signal G6816: std_logic; attribute dont_touch of G6816: signal is true;
	signal G6817: std_logic; attribute dont_touch of G6817: signal is true;
	signal G6818: std_logic; attribute dont_touch of G6818: signal is true;
	signal G6819: std_logic; attribute dont_touch of G6819: signal is true;
	signal G6820: std_logic; attribute dont_touch of G6820: signal is true;
	signal G6821: std_logic; attribute dont_touch of G6821: signal is true;
	signal G6822: std_logic; attribute dont_touch of G6822: signal is true;
	signal G6823: std_logic; attribute dont_touch of G6823: signal is true;
	signal G6824: std_logic; attribute dont_touch of G6824: signal is true;
	signal G6825: std_logic; attribute dont_touch of G6825: signal is true;
	signal G6826: std_logic; attribute dont_touch of G6826: signal is true;
	signal G6827: std_logic; attribute dont_touch of G6827: signal is true;
	signal G6828: std_logic; attribute dont_touch of G6828: signal is true;
	signal G6829: std_logic; attribute dont_touch of G6829: signal is true;
	signal G6830: std_logic; attribute dont_touch of G6830: signal is true;
	signal G6831: std_logic; attribute dont_touch of G6831: signal is true;
	signal G6832: std_logic; attribute dont_touch of G6832: signal is true;
	signal G6833: std_logic; attribute dont_touch of G6833: signal is true;
	signal G6834: std_logic; attribute dont_touch of G6834: signal is true;
	signal G6835: std_logic; attribute dont_touch of G6835: signal is true;
	signal G6836: std_logic; attribute dont_touch of G6836: signal is true;
	signal G6837: std_logic; attribute dont_touch of G6837: signal is true;
	signal G6838: std_logic; attribute dont_touch of G6838: signal is true;
	signal G6839: std_logic; attribute dont_touch of G6839: signal is true;
	signal G6840: std_logic; attribute dont_touch of G6840: signal is true;
	signal G6841: std_logic; attribute dont_touch of G6841: signal is true;
	signal G6842: std_logic; attribute dont_touch of G6842: signal is true;
	signal G6843: std_logic; attribute dont_touch of G6843: signal is true;
	signal G6844: std_logic; attribute dont_touch of G6844: signal is true;
	signal G6845: std_logic; attribute dont_touch of G6845: signal is true;
	signal G6846: std_logic; attribute dont_touch of G6846: signal is true;
	signal G6847: std_logic; attribute dont_touch of G6847: signal is true;
	signal G6848: std_logic; attribute dont_touch of G6848: signal is true;
	signal G6851: std_logic; attribute dont_touch of G6851: signal is true;
	signal G6852: std_logic; attribute dont_touch of G6852: signal is true;
	signal G6853: std_logic; attribute dont_touch of G6853: signal is true;
	signal G6854: std_logic; attribute dont_touch of G6854: signal is true;
	signal G6855: std_logic; attribute dont_touch of G6855: signal is true;
	signal G6856: std_logic; attribute dont_touch of G6856: signal is true;
	signal G6857: std_logic; attribute dont_touch of G6857: signal is true;
	signal G6858: std_logic; attribute dont_touch of G6858: signal is true;
	signal G6859: std_logic; attribute dont_touch of G6859: signal is true;
	signal G6860: std_logic; attribute dont_touch of G6860: signal is true;
	signal G6861: std_logic; attribute dont_touch of G6861: signal is true;
	signal G6862: std_logic; attribute dont_touch of G6862: signal is true;
	signal G6863: std_logic; attribute dont_touch of G6863: signal is true;
	signal G6864: std_logic; attribute dont_touch of G6864: signal is true;
	signal G6865: std_logic; attribute dont_touch of G6865: signal is true;
	signal G6866: std_logic; attribute dont_touch of G6866: signal is true;
	signal G6867: std_logic; attribute dont_touch of G6867: signal is true;
	signal G6868: std_logic; attribute dont_touch of G6868: signal is true;
	signal G6869: std_logic; attribute dont_touch of G6869: signal is true;
	signal G6870: std_logic; attribute dont_touch of G6870: signal is true;
	signal G6871: std_logic; attribute dont_touch of G6871: signal is true;
	signal G6872: std_logic; attribute dont_touch of G6872: signal is true;
	signal G6873: std_logic; attribute dont_touch of G6873: signal is true;
	signal G6874: std_logic; attribute dont_touch of G6874: signal is true;
	signal G6875: std_logic; attribute dont_touch of G6875: signal is true;
	signal G6876: std_logic; attribute dont_touch of G6876: signal is true;
	signal G6877: std_logic; attribute dont_touch of G6877: signal is true;
	signal G6878: std_logic; attribute dont_touch of G6878: signal is true;
	signal G6879: std_logic; attribute dont_touch of G6879: signal is true;
	signal G6880: std_logic; attribute dont_touch of G6880: signal is true;
	signal G6881: std_logic; attribute dont_touch of G6881: signal is true;
	signal G6882: std_logic; attribute dont_touch of G6882: signal is true;
	signal G6883: std_logic; attribute dont_touch of G6883: signal is true;
	signal G6884: std_logic; attribute dont_touch of G6884: signal is true;
	signal G6885: std_logic; attribute dont_touch of G6885: signal is true;
	signal G6886: std_logic; attribute dont_touch of G6886: signal is true;
	signal G6887: std_logic; attribute dont_touch of G6887: signal is true;
	signal G6888: std_logic; attribute dont_touch of G6888: signal is true;
	signal G6889: std_logic; attribute dont_touch of G6889: signal is true;
	signal G6890: std_logic; attribute dont_touch of G6890: signal is true;
	signal G6891: std_logic; attribute dont_touch of G6891: signal is true;
	signal G6892: std_logic; attribute dont_touch of G6892: signal is true;
	signal G6893: std_logic; attribute dont_touch of G6893: signal is true;
	signal G6894: std_logic; attribute dont_touch of G6894: signal is true;
	signal G6896: std_logic; attribute dont_touch of G6896: signal is true;
	signal G6897: std_logic; attribute dont_touch of G6897: signal is true;
	signal G6898: std_logic; attribute dont_touch of G6898: signal is true;
	signal G6899: std_logic; attribute dont_touch of G6899: signal is true;
	signal G6900: std_logic; attribute dont_touch of G6900: signal is true;
	signal G6901: std_logic; attribute dont_touch of G6901: signal is true;
	signal G6902: std_logic; attribute dont_touch of G6902: signal is true;
	signal G6903: std_logic; attribute dont_touch of G6903: signal is true;
	signal G6904: std_logic; attribute dont_touch of G6904: signal is true;
	signal G6905: std_logic; attribute dont_touch of G6905: signal is true;
	signal G6906: std_logic; attribute dont_touch of G6906: signal is true;
	signal G6907: std_logic; attribute dont_touch of G6907: signal is true;
	signal G6908: std_logic; attribute dont_touch of G6908: signal is true;
	signal G6910: std_logic; attribute dont_touch of G6910: signal is true;
	signal G6911: std_logic; attribute dont_touch of G6911: signal is true;
	signal G6912: std_logic; attribute dont_touch of G6912: signal is true;
	signal G6913: std_logic; attribute dont_touch of G6913: signal is true;
	signal G6914: std_logic; attribute dont_touch of G6914: signal is true;
	signal G6915: std_logic; attribute dont_touch of G6915: signal is true;
	signal G6916: std_logic; attribute dont_touch of G6916: signal is true;
	signal G6917: std_logic; attribute dont_touch of G6917: signal is true;
	signal G6918: std_logic; attribute dont_touch of G6918: signal is true;
	signal G6919: std_logic; attribute dont_touch of G6919: signal is true;
	signal G6920: std_logic; attribute dont_touch of G6920: signal is true;
	signal G6921: std_logic; attribute dont_touch of G6921: signal is true;
	signal G6922: std_logic; attribute dont_touch of G6922: signal is true;
	signal G6923: std_logic; attribute dont_touch of G6923: signal is true;
	signal G6924: std_logic; attribute dont_touch of G6924: signal is true;
	signal G6925: std_logic; attribute dont_touch of G6925: signal is true;
	signal G6926: std_logic; attribute dont_touch of G6926: signal is true;
	signal G6927: std_logic; attribute dont_touch of G6927: signal is true;
	signal G6928: std_logic; attribute dont_touch of G6928: signal is true;
	signal G6929: std_logic; attribute dont_touch of G6929: signal is true;
	signal G6930: std_logic; attribute dont_touch of G6930: signal is true;
	signal G6931: std_logic; attribute dont_touch of G6931: signal is true;
	signal G6932: std_logic; attribute dont_touch of G6932: signal is true;
	signal G6933: std_logic; attribute dont_touch of G6933: signal is true;
	signal G6934: std_logic; attribute dont_touch of G6934: signal is true;
	signal G6935: std_logic; attribute dont_touch of G6935: signal is true;
	signal G6936: std_logic; attribute dont_touch of G6936: signal is true;
	signal G6937: std_logic; attribute dont_touch of G6937: signal is true;
	signal G6938: std_logic; attribute dont_touch of G6938: signal is true;
	signal G6939: std_logic; attribute dont_touch of G6939: signal is true;
	signal G6940: std_logic; attribute dont_touch of G6940: signal is true;
	signal G6941: std_logic; attribute dont_touch of G6941: signal is true;
	signal G6944: std_logic; attribute dont_touch of G6944: signal is true;
	signal G6945: std_logic; attribute dont_touch of G6945: signal is true;
	signal G6946: std_logic; attribute dont_touch of G6946: signal is true;
	signal G6947: std_logic; attribute dont_touch of G6947: signal is true;
	signal G6948: std_logic; attribute dont_touch of G6948: signal is true;
	signal G6949: std_logic; attribute dont_touch of G6949: signal is true;
	signal G6950: std_logic; attribute dont_touch of G6950: signal is true;
	signal G6951: std_logic; attribute dont_touch of G6951: signal is true;
	signal G6952: std_logic; attribute dont_touch of G6952: signal is true;
	signal G6953: std_logic; attribute dont_touch of G6953: signal is true;
	signal G6954: std_logic; attribute dont_touch of G6954: signal is true;
	signal G6955: std_logic; attribute dont_touch of G6955: signal is true;
	signal G6956: std_logic; attribute dont_touch of G6956: signal is true;
	signal G6957: std_logic; attribute dont_touch of G6957: signal is true;
	signal G6958: std_logic; attribute dont_touch of G6958: signal is true;
	signal G6959: std_logic; attribute dont_touch of G6959: signal is true;
	signal G6960: std_logic; attribute dont_touch of G6960: signal is true;
	signal G6961: std_logic; attribute dont_touch of G6961: signal is true;
	signal G6962: std_logic; attribute dont_touch of G6962: signal is true;
	signal G6963: std_logic; attribute dont_touch of G6963: signal is true;
	signal G6964: std_logic; attribute dont_touch of G6964: signal is true;
	signal G6965: std_logic; attribute dont_touch of G6965: signal is true;
	signal G6966: std_logic; attribute dont_touch of G6966: signal is true;
	signal G6967: std_logic; attribute dont_touch of G6967: signal is true;
	signal G6968: std_logic; attribute dont_touch of G6968: signal is true;
	signal G6969: std_logic; attribute dont_touch of G6969: signal is true;
	signal G6970: std_logic; attribute dont_touch of G6970: signal is true;
	signal G6971: std_logic; attribute dont_touch of G6971: signal is true;
	signal G6972: std_logic; attribute dont_touch of G6972: signal is true;
	signal G6973: std_logic; attribute dont_touch of G6973: signal is true;
	signal G6974: std_logic; attribute dont_touch of G6974: signal is true;
	signal G6975: std_logic; attribute dont_touch of G6975: signal is true;
	signal G6976: std_logic; attribute dont_touch of G6976: signal is true;
	signal G6977: std_logic; attribute dont_touch of G6977: signal is true;
	signal G6978: std_logic; attribute dont_touch of G6978: signal is true;
	signal G6979: std_logic; attribute dont_touch of G6979: signal is true;
	signal G6980: std_logic; attribute dont_touch of G6980: signal is true;
	signal G6983: std_logic; attribute dont_touch of G6983: signal is true;
	signal G6984: std_logic; attribute dont_touch of G6984: signal is true;
	signal G6990: std_logic; attribute dont_touch of G6990: signal is true;
	signal G6991: std_logic; attribute dont_touch of G6991: signal is true;
	signal G6992: std_logic; attribute dont_touch of G6992: signal is true;
	signal G6993: std_logic; attribute dont_touch of G6993: signal is true;
	signal G6994: std_logic; attribute dont_touch of G6994: signal is true;
	signal G6995: std_logic; attribute dont_touch of G6995: signal is true;
	signal G6996: std_logic; attribute dont_touch of G6996: signal is true;
	signal G6997: std_logic; attribute dont_touch of G6997: signal is true;
	signal G6998: std_logic; attribute dont_touch of G6998: signal is true;
	signal G6999: std_logic; attribute dont_touch of G6999: signal is true;
	signal G7000: std_logic; attribute dont_touch of G7000: signal is true;
	signal G7001: std_logic; attribute dont_touch of G7001: signal is true;
	signal G7002: std_logic; attribute dont_touch of G7002: signal is true;
	signal G7003: std_logic; attribute dont_touch of G7003: signal is true;
	signal G7006: std_logic; attribute dont_touch of G7006: signal is true;
	signal G7007: std_logic; attribute dont_touch of G7007: signal is true;
	signal G7008: std_logic; attribute dont_touch of G7008: signal is true;
	signal G7009: std_logic; attribute dont_touch of G7009: signal is true;
	signal G7010: std_logic; attribute dont_touch of G7010: signal is true;
	signal G7013: std_logic; attribute dont_touch of G7013: signal is true;
	signal G7014: std_logic; attribute dont_touch of G7014: signal is true;
	signal G7015: std_logic; attribute dont_touch of G7015: signal is true;
	signal G7016: std_logic; attribute dont_touch of G7016: signal is true;
	signal G7017: std_logic; attribute dont_touch of G7017: signal is true;
	signal G7018: std_logic; attribute dont_touch of G7018: signal is true;
	signal G7019: std_logic; attribute dont_touch of G7019: signal is true;
	signal G7020: std_logic; attribute dont_touch of G7020: signal is true;
	signal G7021: std_logic; attribute dont_touch of G7021: signal is true;
	signal G7022: std_logic; attribute dont_touch of G7022: signal is true;
	signal G7023: std_logic; attribute dont_touch of G7023: signal is true;
	signal G7024: std_logic; attribute dont_touch of G7024: signal is true;
	signal G7025: std_logic; attribute dont_touch of G7025: signal is true;
	signal G7026: std_logic; attribute dont_touch of G7026: signal is true;
	signal G7027: std_logic; attribute dont_touch of G7027: signal is true;
	signal G7028: std_logic; attribute dont_touch of G7028: signal is true;
	signal G7029: std_logic; attribute dont_touch of G7029: signal is true;
	signal G7030: std_logic; attribute dont_touch of G7030: signal is true;
	signal G7031: std_logic; attribute dont_touch of G7031: signal is true;
	signal G7032: std_logic; attribute dont_touch of G7032: signal is true;
	signal G7033: std_logic; attribute dont_touch of G7033: signal is true;
	signal G7034: std_logic; attribute dont_touch of G7034: signal is true;
	signal G7035: std_logic; attribute dont_touch of G7035: signal is true;
	signal G7036: std_logic; attribute dont_touch of G7036: signal is true;
	signal G7037: std_logic; attribute dont_touch of G7037: signal is true;
	signal G7038: std_logic; attribute dont_touch of G7038: signal is true;
	signal G7039: std_logic; attribute dont_touch of G7039: signal is true;
	signal G7040: std_logic; attribute dont_touch of G7040: signal is true;
	signal G7041: std_logic; attribute dont_touch of G7041: signal is true;
	signal G7042: std_logic; attribute dont_touch of G7042: signal is true;
	signal G7043: std_logic; attribute dont_touch of G7043: signal is true;
	signal G7044: std_logic; attribute dont_touch of G7044: signal is true;
	signal G7045: std_logic; attribute dont_touch of G7045: signal is true;
	signal G7046: std_logic; attribute dont_touch of G7046: signal is true;
	signal G7047: std_logic; attribute dont_touch of G7047: signal is true;
	signal G7049: std_logic; attribute dont_touch of G7049: signal is true;
	signal G7050: std_logic; attribute dont_touch of G7050: signal is true;
	signal G7054: std_logic; attribute dont_touch of G7054: signal is true;
	signal G7055: std_logic; attribute dont_touch of G7055: signal is true;
	signal G7056: std_logic; attribute dont_touch of G7056: signal is true;
	signal G7057: std_logic; attribute dont_touch of G7057: signal is true;
	signal G7058: std_logic; attribute dont_touch of G7058: signal is true;
	signal G7059: std_logic; attribute dont_touch of G7059: signal is true;
	signal G7060: std_logic; attribute dont_touch of G7060: signal is true;
	signal G7061: std_logic; attribute dont_touch of G7061: signal is true;
	signal G7062: std_logic; attribute dont_touch of G7062: signal is true;
	signal G7064: std_logic; attribute dont_touch of G7064: signal is true;
	signal G7065: std_logic; attribute dont_touch of G7065: signal is true;
	signal G7066: std_logic; attribute dont_touch of G7066: signal is true;
	signal G7067: std_logic; attribute dont_touch of G7067: signal is true;
	signal G7068: std_logic; attribute dont_touch of G7068: signal is true;
	signal G7069: std_logic; attribute dont_touch of G7069: signal is true;
	signal G7070: std_logic; attribute dont_touch of G7070: signal is true;
	signal G7071: std_logic; attribute dont_touch of G7071: signal is true;
	signal G7077: std_logic; attribute dont_touch of G7077: signal is true;
	signal G7078: std_logic; attribute dont_touch of G7078: signal is true;
	signal G7079: std_logic; attribute dont_touch of G7079: signal is true;
	signal G7080: std_logic; attribute dont_touch of G7080: signal is true;
	signal G7081: std_logic; attribute dont_touch of G7081: signal is true;
	signal G7082: std_logic; attribute dont_touch of G7082: signal is true;
	signal G7083: std_logic; attribute dont_touch of G7083: signal is true;
	signal G7086: std_logic; attribute dont_touch of G7086: signal is true;
	signal G7087: std_logic; attribute dont_touch of G7087: signal is true;
	signal G7088: std_logic; attribute dont_touch of G7088: signal is true;
	signal G7089: std_logic; attribute dont_touch of G7089: signal is true;
	signal G7090: std_logic; attribute dont_touch of G7090: signal is true;
	signal G7091: std_logic; attribute dont_touch of G7091: signal is true;
	signal G7092: std_logic; attribute dont_touch of G7092: signal is true;
	signal G7093: std_logic; attribute dont_touch of G7093: signal is true;
	signal G7094: std_logic; attribute dont_touch of G7094: signal is true;
	signal G7095: std_logic; attribute dont_touch of G7095: signal is true;
	signal G7096: std_logic; attribute dont_touch of G7096: signal is true;
	signal G7097: std_logic; attribute dont_touch of G7097: signal is true;
	signal G7098: std_logic; attribute dont_touch of G7098: signal is true;
	signal G7099: std_logic; attribute dont_touch of G7099: signal is true;
	signal G7100: std_logic; attribute dont_touch of G7100: signal is true;
	signal G7101: std_logic; attribute dont_touch of G7101: signal is true;
	signal G7102: std_logic; attribute dont_touch of G7102: signal is true;
	signal G7104: std_logic; attribute dont_touch of G7104: signal is true;
	signal G7105: std_logic; attribute dont_touch of G7105: signal is true;
	signal G7106: std_logic; attribute dont_touch of G7106: signal is true;
	signal G7107: std_logic; attribute dont_touch of G7107: signal is true;
	signal G7108: std_logic; attribute dont_touch of G7108: signal is true;
	signal G7109: std_logic; attribute dont_touch of G7109: signal is true;
	signal G7110: std_logic; attribute dont_touch of G7110: signal is true;
	signal G7111: std_logic; attribute dont_touch of G7111: signal is true;
	signal G7112: std_logic; attribute dont_touch of G7112: signal is true;
	signal G7113: std_logic; attribute dont_touch of G7113: signal is true;
	signal G7114: std_logic; attribute dont_touch of G7114: signal is true;
	signal G7115: std_logic; attribute dont_touch of G7115: signal is true;
	signal G7116: std_logic; attribute dont_touch of G7116: signal is true;
	signal G7117: std_logic; attribute dont_touch of G7117: signal is true;
	signal G7118: std_logic; attribute dont_touch of G7118: signal is true;
	signal G7119: std_logic; attribute dont_touch of G7119: signal is true;
	signal G7120: std_logic; attribute dont_touch of G7120: signal is true;
	signal G7121: std_logic; attribute dont_touch of G7121: signal is true;
	signal G7122: std_logic; attribute dont_touch of G7122: signal is true;
	signal G7123: std_logic; attribute dont_touch of G7123: signal is true;
	signal G7124: std_logic; attribute dont_touch of G7124: signal is true;
	signal G7125: std_logic; attribute dont_touch of G7125: signal is true;
	signal G7126: std_logic; attribute dont_touch of G7126: signal is true;
	signal G7127: std_logic; attribute dont_touch of G7127: signal is true;
	signal G7128: std_logic; attribute dont_touch of G7128: signal is true;
	signal G7129: std_logic; attribute dont_touch of G7129: signal is true;
	signal G7130: std_logic; attribute dont_touch of G7130: signal is true;
	signal G7131: std_logic; attribute dont_touch of G7131: signal is true;
	signal G7132: std_logic; attribute dont_touch of G7132: signal is true;
	signal G7133: std_logic; attribute dont_touch of G7133: signal is true;
	signal G7134: std_logic; attribute dont_touch of G7134: signal is true;
	signal G7135: std_logic; attribute dont_touch of G7135: signal is true;
	signal G7136: std_logic; attribute dont_touch of G7136: signal is true;
	signal G7137: std_logic; attribute dont_touch of G7137: signal is true;
	signal G7138: std_logic; attribute dont_touch of G7138: signal is true;
	signal G7139: std_logic; attribute dont_touch of G7139: signal is true;
	signal G7140: std_logic; attribute dont_touch of G7140: signal is true;
	signal G7141: std_logic; attribute dont_touch of G7141: signal is true;
	signal G7142: std_logic; attribute dont_touch of G7142: signal is true;
	signal G7143: std_logic; attribute dont_touch of G7143: signal is true;
	signal G7144: std_logic; attribute dont_touch of G7144: signal is true;
	signal G7145: std_logic; attribute dont_touch of G7145: signal is true;
	signal G7146: std_logic; attribute dont_touch of G7146: signal is true;
	signal G7147: std_logic; attribute dont_touch of G7147: signal is true;
	signal G7148: std_logic; attribute dont_touch of G7148: signal is true;
	signal G7149: std_logic; attribute dont_touch of G7149: signal is true;
	signal G7150: std_logic; attribute dont_touch of G7150: signal is true;
	signal G7151: std_logic; attribute dont_touch of G7151: signal is true;
	signal G7152: std_logic; attribute dont_touch of G7152: signal is true;
	signal G7155: std_logic; attribute dont_touch of G7155: signal is true;
	signal G7156: std_logic; attribute dont_touch of G7156: signal is true;
	signal G7157: std_logic; attribute dont_touch of G7157: signal is true;
	signal G7158: std_logic; attribute dont_touch of G7158: signal is true;
	signal G7159: std_logic; attribute dont_touch of G7159: signal is true;
	signal G7160: std_logic; attribute dont_touch of G7160: signal is true;
	signal G7161: std_logic; attribute dont_touch of G7161: signal is true;
	signal G7162: std_logic; attribute dont_touch of G7162: signal is true;
	signal G7163: std_logic; attribute dont_touch of G7163: signal is true;
	signal G7164: std_logic; attribute dont_touch of G7164: signal is true;
	signal G7165: std_logic; attribute dont_touch of G7165: signal is true;
	signal G7166: std_logic; attribute dont_touch of G7166: signal is true;
	signal G7167: std_logic; attribute dont_touch of G7167: signal is true;
	signal G7168: std_logic; attribute dont_touch of G7168: signal is true;
	signal G7169: std_logic; attribute dont_touch of G7169: signal is true;
	signal G7170: std_logic; attribute dont_touch of G7170: signal is true;
	signal G7171: std_logic; attribute dont_touch of G7171: signal is true;
	signal G7172: std_logic; attribute dont_touch of G7172: signal is true;
	signal G7173: std_logic; attribute dont_touch of G7173: signal is true;
	signal G7174: std_logic; attribute dont_touch of G7174: signal is true;
	signal G7175: std_logic; attribute dont_touch of G7175: signal is true;
	signal G7176: std_logic; attribute dont_touch of G7176: signal is true;
	signal G7177: std_logic; attribute dont_touch of G7177: signal is true;
	signal G7178: std_logic; attribute dont_touch of G7178: signal is true;
	signal G7179: std_logic; attribute dont_touch of G7179: signal is true;
	signal G7180: std_logic; attribute dont_touch of G7180: signal is true;
	signal G7181: std_logic; attribute dont_touch of G7181: signal is true;
	signal G7182: std_logic; attribute dont_touch of G7182: signal is true;
	signal G7183: std_logic; attribute dont_touch of G7183: signal is true;
	signal G7184: std_logic; attribute dont_touch of G7184: signal is true;
	signal G7185: std_logic; attribute dont_touch of G7185: signal is true;
	signal G7186: std_logic; attribute dont_touch of G7186: signal is true;
	signal G7187: std_logic; attribute dont_touch of G7187: signal is true;
	signal G7188: std_logic; attribute dont_touch of G7188: signal is true;
	signal G7189: std_logic; attribute dont_touch of G7189: signal is true;
	signal G7190: std_logic; attribute dont_touch of G7190: signal is true;
	signal G7191: std_logic; attribute dont_touch of G7191: signal is true;
	signal G7192: std_logic; attribute dont_touch of G7192: signal is true;
	signal G7193: std_logic; attribute dont_touch of G7193: signal is true;
	signal G7194: std_logic; attribute dont_touch of G7194: signal is true;
	signal G7195: std_logic; attribute dont_touch of G7195: signal is true;
	signal G7196: std_logic; attribute dont_touch of G7196: signal is true;
	signal G7197: std_logic; attribute dont_touch of G7197: signal is true;
	signal G7198: std_logic; attribute dont_touch of G7198: signal is true;
	signal G7199: std_logic; attribute dont_touch of G7199: signal is true;
	signal G7202: std_logic; attribute dont_touch of G7202: signal is true;
	signal G7205: std_logic; attribute dont_touch of G7205: signal is true;
	signal G7206: std_logic; attribute dont_touch of G7206: signal is true;
	signal G7207: std_logic; attribute dont_touch of G7207: signal is true;
	signal G7208: std_logic; attribute dont_touch of G7208: signal is true;
	signal G7209: std_logic; attribute dont_touch of G7209: signal is true;
	signal G7210: std_logic; attribute dont_touch of G7210: signal is true;
	signal G7211: std_logic; attribute dont_touch of G7211: signal is true;
	signal G7212: std_logic; attribute dont_touch of G7212: signal is true;
	signal G7215: std_logic; attribute dont_touch of G7215: signal is true;
	signal G7216: std_logic; attribute dont_touch of G7216: signal is true;
	signal G7217: std_logic; attribute dont_touch of G7217: signal is true;
	signal G7220: std_logic; attribute dont_touch of G7220: signal is true;
	signal G7221: std_logic; attribute dont_touch of G7221: signal is true;
	signal G7222: std_logic; attribute dont_touch of G7222: signal is true;
	signal G7223: std_logic; attribute dont_touch of G7223: signal is true;
	signal G7224: std_logic; attribute dont_touch of G7224: signal is true;
	signal G7225: std_logic; attribute dont_touch of G7225: signal is true;
	signal G7226: std_logic; attribute dont_touch of G7226: signal is true;
	signal G7227: std_logic; attribute dont_touch of G7227: signal is true;
	signal G7228: std_logic; attribute dont_touch of G7228: signal is true;
	signal G7229: std_logic; attribute dont_touch of G7229: signal is true;
	signal G7230: std_logic; attribute dont_touch of G7230: signal is true;
	signal G7231: std_logic; attribute dont_touch of G7231: signal is true;
	signal G7232: std_logic; attribute dont_touch of G7232: signal is true;
	signal G7233: std_logic; attribute dont_touch of G7233: signal is true;
	signal G7234: std_logic; attribute dont_touch of G7234: signal is true;
	signal G7235: std_logic; attribute dont_touch of G7235: signal is true;
	signal G7236: std_logic; attribute dont_touch of G7236: signal is true;
	signal G7237: std_logic; attribute dont_touch of G7237: signal is true;
	signal G7238: std_logic; attribute dont_touch of G7238: signal is true;
	signal G7239: std_logic; attribute dont_touch of G7239: signal is true;
	signal G7240: std_logic; attribute dont_touch of G7240: signal is true;
	signal G7241: std_logic; attribute dont_touch of G7241: signal is true;
	signal G7242: std_logic; attribute dont_touch of G7242: signal is true;
	signal G7243: std_logic; attribute dont_touch of G7243: signal is true;
	signal G7244: std_logic; attribute dont_touch of G7244: signal is true;
	signal G7245: std_logic; attribute dont_touch of G7245: signal is true;
	signal G7246: std_logic; attribute dont_touch of G7246: signal is true;
	signal G7247: std_logic; attribute dont_touch of G7247: signal is true;
	signal G7248: std_logic; attribute dont_touch of G7248: signal is true;
	signal G7251: std_logic; attribute dont_touch of G7251: signal is true;
	signal G7252: std_logic; attribute dont_touch of G7252: signal is true;
	signal G7253: std_logic; attribute dont_touch of G7253: signal is true;
	signal G7254: std_logic; attribute dont_touch of G7254: signal is true;
	signal G7255: std_logic; attribute dont_touch of G7255: signal is true;
	signal G7256: std_logic; attribute dont_touch of G7256: signal is true;
	signal G7257: std_logic; attribute dont_touch of G7257: signal is true;
	signal G7258: std_logic; attribute dont_touch of G7258: signal is true;
	signal G7259: std_logic; attribute dont_touch of G7259: signal is true;
	signal G7260: std_logic; attribute dont_touch of G7260: signal is true;
	signal G7261: std_logic; attribute dont_touch of G7261: signal is true;
	signal G7262: std_logic; attribute dont_touch of G7262: signal is true;
	signal G7263: std_logic; attribute dont_touch of G7263: signal is true;
	signal G7264: std_logic; attribute dont_touch of G7264: signal is true;
	signal G7265: std_logic; attribute dont_touch of G7265: signal is true;
	signal G7266: std_logic; attribute dont_touch of G7266: signal is true;
	signal G7267: std_logic; attribute dont_touch of G7267: signal is true;
	signal G7268: std_logic; attribute dont_touch of G7268: signal is true;
	signal G7269: std_logic; attribute dont_touch of G7269: signal is true;
	signal G7270: std_logic; attribute dont_touch of G7270: signal is true;
	signal G7271: std_logic; attribute dont_touch of G7271: signal is true;
	signal G7272: std_logic; attribute dont_touch of G7272: signal is true;
	signal G7273: std_logic; attribute dont_touch of G7273: signal is true;
	signal G7274: std_logic; attribute dont_touch of G7274: signal is true;
	signal G7275: std_logic; attribute dont_touch of G7275: signal is true;
	signal G7276: std_logic; attribute dont_touch of G7276: signal is true;
	signal G7277: std_logic; attribute dont_touch of G7277: signal is true;
	signal G7278: std_logic; attribute dont_touch of G7278: signal is true;
	signal G7279: std_logic; attribute dont_touch of G7279: signal is true;
	signal G7280: std_logic; attribute dont_touch of G7280: signal is true;
	signal G7281: std_logic; attribute dont_touch of G7281: signal is true;
	signal G7282: std_logic; attribute dont_touch of G7282: signal is true;
	signal G7296: std_logic; attribute dont_touch of G7296: signal is true;
	signal G7297: std_logic; attribute dont_touch of G7297: signal is true;
	signal G7299: std_logic; attribute dont_touch of G7299: signal is true;
	signal G7300: std_logic; attribute dont_touch of G7300: signal is true;
	signal G7301: std_logic; attribute dont_touch of G7301: signal is true;
	signal G7302: std_logic; attribute dont_touch of G7302: signal is true;
	signal G7303: std_logic; attribute dont_touch of G7303: signal is true;
	signal G7304: std_logic; attribute dont_touch of G7304: signal is true;
	signal G7305: std_logic; attribute dont_touch of G7305: signal is true;
	signal G7306: std_logic; attribute dont_touch of G7306: signal is true;
	signal G7307: std_logic; attribute dont_touch of G7307: signal is true;
	signal G7308: std_logic; attribute dont_touch of G7308: signal is true;
	signal G7309: std_logic; attribute dont_touch of G7309: signal is true;
	signal G7310: std_logic; attribute dont_touch of G7310: signal is true;
	signal G7311: std_logic; attribute dont_touch of G7311: signal is true;
	signal G7312: std_logic; attribute dont_touch of G7312: signal is true;
	signal G7313: std_logic; attribute dont_touch of G7313: signal is true;
	signal G7314: std_logic; attribute dont_touch of G7314: signal is true;
	signal G7315: std_logic; attribute dont_touch of G7315: signal is true;
	signal G7316: std_logic; attribute dont_touch of G7316: signal is true;
	signal G7317: std_logic; attribute dont_touch of G7317: signal is true;
	signal G7318: std_logic; attribute dont_touch of G7318: signal is true;
	signal G7319: std_logic; attribute dont_touch of G7319: signal is true;
	signal G7320: std_logic; attribute dont_touch of G7320: signal is true;
	signal G7321: std_logic; attribute dont_touch of G7321: signal is true;
	signal G7322: std_logic; attribute dont_touch of G7322: signal is true;
	signal G7323: std_logic; attribute dont_touch of G7323: signal is true;
	signal G7324: std_logic; attribute dont_touch of G7324: signal is true;
	signal G7325: std_logic; attribute dont_touch of G7325: signal is true;
	signal G7326: std_logic; attribute dont_touch of G7326: signal is true;
	signal G7327: std_logic; attribute dont_touch of G7327: signal is true;
	signal G7328: std_logic; attribute dont_touch of G7328: signal is true;
	signal G7329: std_logic; attribute dont_touch of G7329: signal is true;
	signal G7330: std_logic; attribute dont_touch of G7330: signal is true;
	signal G7331: std_logic; attribute dont_touch of G7331: signal is true;
	signal G7332: std_logic; attribute dont_touch of G7332: signal is true;
	signal G7333: std_logic; attribute dont_touch of G7333: signal is true;
	signal G7334: std_logic; attribute dont_touch of G7334: signal is true;
	signal G7335: std_logic; attribute dont_touch of G7335: signal is true;
	signal G7336: std_logic; attribute dont_touch of G7336: signal is true;
	signal G7337: std_logic; attribute dont_touch of G7337: signal is true;
	signal G7338: std_logic; attribute dont_touch of G7338: signal is true;
	signal G7339: std_logic; attribute dont_touch of G7339: signal is true;
	signal G7340: std_logic; attribute dont_touch of G7340: signal is true;
	signal G7341: std_logic; attribute dont_touch of G7341: signal is true;
	signal G7342: std_logic; attribute dont_touch of G7342: signal is true;
	signal G7343: std_logic; attribute dont_touch of G7343: signal is true;
	signal G7344: std_logic; attribute dont_touch of G7344: signal is true;
	signal G7345: std_logic; attribute dont_touch of G7345: signal is true;
	signal G7346: std_logic; attribute dont_touch of G7346: signal is true;
	signal G7347: std_logic; attribute dont_touch of G7347: signal is true;
	signal G7348: std_logic; attribute dont_touch of G7348: signal is true;
	signal G7349: std_logic; attribute dont_touch of G7349: signal is true;
	signal G7350: std_logic; attribute dont_touch of G7350: signal is true;
	signal G7351: std_logic; attribute dont_touch of G7351: signal is true;
	signal G7352: std_logic; attribute dont_touch of G7352: signal is true;
	signal G7353: std_logic; attribute dont_touch of G7353: signal is true;
	signal G7354: std_logic; attribute dont_touch of G7354: signal is true;
	signal G7355: std_logic; attribute dont_touch of G7355: signal is true;
	signal G7356: std_logic; attribute dont_touch of G7356: signal is true;
	signal G7357: std_logic; attribute dont_touch of G7357: signal is true;
	signal G7358: std_logic; attribute dont_touch of G7358: signal is true;
	signal G7359: std_logic; attribute dont_touch of G7359: signal is true;
	signal G7360: std_logic; attribute dont_touch of G7360: signal is true;
	signal G7361: std_logic; attribute dont_touch of G7361: signal is true;
	signal G7362: std_logic; attribute dont_touch of G7362: signal is true;
	signal G7363: std_logic; attribute dont_touch of G7363: signal is true;
	signal G7364: std_logic; attribute dont_touch of G7364: signal is true;
	signal G7365: std_logic; attribute dont_touch of G7365: signal is true;
	signal G7366: std_logic; attribute dont_touch of G7366: signal is true;
	signal G7367: std_logic; attribute dont_touch of G7367: signal is true;
	signal G7405: std_logic; attribute dont_touch of G7405: signal is true;
	signal G7406: std_logic; attribute dont_touch of G7406: signal is true;
	signal G7411: std_logic; attribute dont_touch of G7411: signal is true;
	signal G7412: std_logic; attribute dont_touch of G7412: signal is true;
	signal G7413: std_logic; attribute dont_touch of G7413: signal is true;
	signal G7414: std_logic; attribute dont_touch of G7414: signal is true;
	signal G7415: std_logic; attribute dont_touch of G7415: signal is true;
	signal G7416: std_logic; attribute dont_touch of G7416: signal is true;
	signal G7417: std_logic; attribute dont_touch of G7417: signal is true;
	signal G7418: std_logic; attribute dont_touch of G7418: signal is true;
	signal G7419: std_logic; attribute dont_touch of G7419: signal is true;
	signal G7420: std_logic; attribute dont_touch of G7420: signal is true;
	signal G7421: std_logic; attribute dont_touch of G7421: signal is true;
	signal G7422: std_logic; attribute dont_touch of G7422: signal is true;
	signal G7426: std_logic; attribute dont_touch of G7426: signal is true;
	signal G7427: std_logic; attribute dont_touch of G7427: signal is true;
	signal G7428: std_logic; attribute dont_touch of G7428: signal is true;
	signal G7429: std_logic; attribute dont_touch of G7429: signal is true;
	signal G7432: std_logic; attribute dont_touch of G7432: signal is true;
	signal G7433: std_logic; attribute dont_touch of G7433: signal is true;
	signal G7434: std_logic; attribute dont_touch of G7434: signal is true;
	signal G7435: std_logic; attribute dont_touch of G7435: signal is true;
	signal G7436: std_logic; attribute dont_touch of G7436: signal is true;
	signal G7437: std_logic; attribute dont_touch of G7437: signal is true;
	signal G7438: std_logic; attribute dont_touch of G7438: signal is true;
	signal G7439: std_logic; attribute dont_touch of G7439: signal is true;
	signal G7440: std_logic; attribute dont_touch of G7440: signal is true;
	signal G7441: std_logic; attribute dont_touch of G7441: signal is true;
	signal G7442: std_logic; attribute dont_touch of G7442: signal is true;
	signal G7443: std_logic; attribute dont_touch of G7443: signal is true;
	signal G7444: std_logic; attribute dont_touch of G7444: signal is true;
	signal G7445: std_logic; attribute dont_touch of G7445: signal is true;
	signal G7446: std_logic; attribute dont_touch of G7446: signal is true;
	signal G7447: std_logic; attribute dont_touch of G7447: signal is true;
	signal G7448: std_logic; attribute dont_touch of G7448: signal is true;
	signal G7449: std_logic; attribute dont_touch of G7449: signal is true;
	signal G7450: std_logic; attribute dont_touch of G7450: signal is true;
	signal G7454: std_logic; attribute dont_touch of G7454: signal is true;
	signal G7455: std_logic; attribute dont_touch of G7455: signal is true;
	signal G7456: std_logic; attribute dont_touch of G7456: signal is true;
	signal G7459: std_logic; attribute dont_touch of G7459: signal is true;
	signal G7460: std_logic; attribute dont_touch of G7460: signal is true;
	signal G7463: std_logic; attribute dont_touch of G7463: signal is true;
	signal G7466: std_logic; attribute dont_touch of G7466: signal is true;
	signal G7467: std_logic; attribute dont_touch of G7467: signal is true;
	signal G7470: std_logic; attribute dont_touch of G7470: signal is true;
	signal G7471: std_logic; attribute dont_touch of G7471: signal is true;
	signal G7475: std_logic; attribute dont_touch of G7475: signal is true;
	signal G7476: std_logic; attribute dont_touch of G7476: signal is true;
	signal G7479: std_logic; attribute dont_touch of G7479: signal is true;
	signal G7480: std_logic; attribute dont_touch of G7480: signal is true;
	signal G7483: std_logic; attribute dont_touch of G7483: signal is true;
	signal G7486: std_logic; attribute dont_touch of G7486: signal is true;
	signal G7487: std_logic; attribute dont_touch of G7487: signal is true;
	signal G7488: std_logic; attribute dont_touch of G7488: signal is true;
	signal G7491: std_logic; attribute dont_touch of G7491: signal is true;
	signal G7492: std_logic; attribute dont_touch of G7492: signal is true;
	signal G7493: std_logic; attribute dont_touch of G7493: signal is true;
	signal G7494: std_logic; attribute dont_touch of G7494: signal is true;
	signal G7495: std_logic; attribute dont_touch of G7495: signal is true;
	signal G7496: std_logic; attribute dont_touch of G7496: signal is true;
	signal G7497: std_logic; attribute dont_touch of G7497: signal is true;
	signal G7498: std_logic; attribute dont_touch of G7498: signal is true;
	signal G7499: std_logic; attribute dont_touch of G7499: signal is true;
	signal G7500: std_logic; attribute dont_touch of G7500: signal is true;
	signal G7501: std_logic; attribute dont_touch of G7501: signal is true;
	signal G7502: std_logic; attribute dont_touch of G7502: signal is true;
	signal G7503: std_logic; attribute dont_touch of G7503: signal is true;
	signal G7509: std_logic; attribute dont_touch of G7509: signal is true;
	signal G7510: std_logic; attribute dont_touch of G7510: signal is true;
	signal G7511: std_logic; attribute dont_touch of G7511: signal is true;
	signal G7512: std_logic; attribute dont_touch of G7512: signal is true;
	signal G7513: std_logic; attribute dont_touch of G7513: signal is true;
	signal G7515: std_logic; attribute dont_touch of G7515: signal is true;
	signal G7516: std_logic; attribute dont_touch of G7516: signal is true;
	signal G7517: std_logic; attribute dont_touch of G7517: signal is true;
	signal G7518: std_logic; attribute dont_touch of G7518: signal is true;
	signal G7519: std_logic; attribute dont_touch of G7519: signal is true;
	signal G7520: std_logic; attribute dont_touch of G7520: signal is true;
	signal G7521: std_logic; attribute dont_touch of G7521: signal is true;
	signal G7522: std_logic; attribute dont_touch of G7522: signal is true;
	signal G7523: std_logic; attribute dont_touch of G7523: signal is true;
	signal G7524: std_logic; attribute dont_touch of G7524: signal is true;
	signal G7525: std_logic; attribute dont_touch of G7525: signal is true;
	signal G7526: std_logic; attribute dont_touch of G7526: signal is true;
	signal G7527: std_logic; attribute dont_touch of G7527: signal is true;
	signal G7528: std_logic; attribute dont_touch of G7528: signal is true;
	signal G7529: std_logic; attribute dont_touch of G7529: signal is true;
	signal G7530: std_logic; attribute dont_touch of G7530: signal is true;
	signal G7531: std_logic; attribute dont_touch of G7531: signal is true;
	signal G7532: std_logic; attribute dont_touch of G7532: signal is true;
	signal G7533: std_logic; attribute dont_touch of G7533: signal is true;
	signal G7534: std_logic; attribute dont_touch of G7534: signal is true;
	signal G7535: std_logic; attribute dont_touch of G7535: signal is true;
	signal G7536: std_logic; attribute dont_touch of G7536: signal is true;
	signal G7537: std_logic; attribute dont_touch of G7537: signal is true;
	signal G7538: std_logic; attribute dont_touch of G7538: signal is true;
	signal G7539: std_logic; attribute dont_touch of G7539: signal is true;
	signal G7540: std_logic; attribute dont_touch of G7540: signal is true;
	signal G7541: std_logic; attribute dont_touch of G7541: signal is true;
	signal G7542: std_logic; attribute dont_touch of G7542: signal is true;
	signal G7543: std_logic; attribute dont_touch of G7543: signal is true;
	signal G7544: std_logic; attribute dont_touch of G7544: signal is true;
	signal G7545: std_logic; attribute dont_touch of G7545: signal is true;
	signal G7546: std_logic; attribute dont_touch of G7546: signal is true;
	signal G7547: std_logic; attribute dont_touch of G7547: signal is true;
	signal G7548: std_logic; attribute dont_touch of G7548: signal is true;
	signal G7549: std_logic; attribute dont_touch of G7549: signal is true;
	signal G7550: std_logic; attribute dont_touch of G7550: signal is true;
	signal G7551: std_logic; attribute dont_touch of G7551: signal is true;
	signal G7552: std_logic; attribute dont_touch of G7552: signal is true;
	signal G7553: std_logic; attribute dont_touch of G7553: signal is true;
	signal G7554: std_logic; attribute dont_touch of G7554: signal is true;
	signal G7555: std_logic; attribute dont_touch of G7555: signal is true;
	signal G7556: std_logic; attribute dont_touch of G7556: signal is true;
	signal G7557: std_logic; attribute dont_touch of G7557: signal is true;
	signal G7558: std_logic; attribute dont_touch of G7558: signal is true;
	signal G7559: std_logic; attribute dont_touch of G7559: signal is true;
	signal G7560: std_logic; attribute dont_touch of G7560: signal is true;
	signal G7561: std_logic; attribute dont_touch of G7561: signal is true;
	signal G7562: std_logic; attribute dont_touch of G7562: signal is true;
	signal G7563: std_logic; attribute dont_touch of G7563: signal is true;
	signal G7564: std_logic; attribute dont_touch of G7564: signal is true;
	signal G7565: std_logic; attribute dont_touch of G7565: signal is true;
	signal G7566: std_logic; attribute dont_touch of G7566: signal is true;
	signal G7574: std_logic; attribute dont_touch of G7574: signal is true;
	signal G7575: std_logic; attribute dont_touch of G7575: signal is true;
	signal G7576: std_logic; attribute dont_touch of G7576: signal is true;
	signal G7577: std_logic; attribute dont_touch of G7577: signal is true;
	signal G7578: std_logic; attribute dont_touch of G7578: signal is true;
	signal G7579: std_logic; attribute dont_touch of G7579: signal is true;
	signal G7580: std_logic; attribute dont_touch of G7580: signal is true;
	signal G7581: std_logic; attribute dont_touch of G7581: signal is true;
	signal G7582: std_logic; attribute dont_touch of G7582: signal is true;
	signal G7583: std_logic; attribute dont_touch of G7583: signal is true;
	signal G7584: std_logic; attribute dont_touch of G7584: signal is true;
	signal G7585: std_logic; attribute dont_touch of G7585: signal is true;
	signal G7586: std_logic; attribute dont_touch of G7586: signal is true;
	signal G7587: std_logic; attribute dont_touch of G7587: signal is true;
	signal G7588: std_logic; attribute dont_touch of G7588: signal is true;
	signal G7589: std_logic; attribute dont_touch of G7589: signal is true;
	signal G7590: std_logic; attribute dont_touch of G7590: signal is true;
	signal G7591: std_logic; attribute dont_touch of G7591: signal is true;
	signal G7592: std_logic; attribute dont_touch of G7592: signal is true;
	signal G7593: std_logic; attribute dont_touch of G7593: signal is true;
	signal G7594: std_logic; attribute dont_touch of G7594: signal is true;
	signal G7595: std_logic; attribute dont_touch of G7595: signal is true;
	signal G7596: std_logic; attribute dont_touch of G7596: signal is true;
	signal G7597: std_logic; attribute dont_touch of G7597: signal is true;
	signal G7598: std_logic; attribute dont_touch of G7598: signal is true;
	signal G7599: std_logic; attribute dont_touch of G7599: signal is true;
	signal G7600: std_logic; attribute dont_touch of G7600: signal is true;
	signal G7601: std_logic; attribute dont_touch of G7601: signal is true;
	signal G7602: std_logic; attribute dont_touch of G7602: signal is true;
	signal G7603: std_logic; attribute dont_touch of G7603: signal is true;
	signal G7604: std_logic; attribute dont_touch of G7604: signal is true;
	signal G7605: std_logic; attribute dont_touch of G7605: signal is true;
	signal G7606: std_logic; attribute dont_touch of G7606: signal is true;
	signal G7607: std_logic; attribute dont_touch of G7607: signal is true;
	signal G7608: std_logic; attribute dont_touch of G7608: signal is true;
	signal G7609: std_logic; attribute dont_touch of G7609: signal is true;
	signal G7610: std_logic; attribute dont_touch of G7610: signal is true;
	signal G7611: std_logic; attribute dont_touch of G7611: signal is true;
	signal G7614: std_logic; attribute dont_touch of G7614: signal is true;
	signal G7615: std_logic; attribute dont_touch of G7615: signal is true;
	signal G7616: std_logic; attribute dont_touch of G7616: signal is true;
	signal G7625: std_logic; attribute dont_touch of G7625: signal is true;
	signal G7626: std_logic; attribute dont_touch of G7626: signal is true;
	signal G7627: std_logic; attribute dont_touch of G7627: signal is true;
	signal G7628: std_logic; attribute dont_touch of G7628: signal is true;
	signal G7631: std_logic; attribute dont_touch of G7631: signal is true;
	signal G7632: std_logic; attribute dont_touch of G7632: signal is true;
	signal G7633: std_logic; attribute dont_touch of G7633: signal is true;
	signal G7634: std_logic; attribute dont_touch of G7634: signal is true;
	signal G7652: std_logic; attribute dont_touch of G7652: signal is true;
	signal G7653: std_logic; attribute dont_touch of G7653: signal is true;
	signal G7654: std_logic; attribute dont_touch of G7654: signal is true;
	signal G7657: std_logic; attribute dont_touch of G7657: signal is true;
	signal G7658: std_logic; attribute dont_touch of G7658: signal is true;
	signal G7676: std_logic; attribute dont_touch of G7676: signal is true;
	signal G7677: std_logic; attribute dont_touch of G7677: signal is true;
	signal G7678: std_logic; attribute dont_touch of G7678: signal is true;
	signal G7679: std_logic; attribute dont_touch of G7679: signal is true;
	signal G7680: std_logic; attribute dont_touch of G7680: signal is true;
	signal G7681: std_logic; attribute dont_touch of G7681: signal is true;
	signal G7682: std_logic; attribute dont_touch of G7682: signal is true;
	signal G7683: std_logic; attribute dont_touch of G7683: signal is true;
	signal G7686: std_logic; attribute dont_touch of G7686: signal is true;
	signal G7687: std_logic; attribute dont_touch of G7687: signal is true;
	signal G7688: std_logic; attribute dont_touch of G7688: signal is true;
	signal G7689: std_logic; attribute dont_touch of G7689: signal is true;
	signal G7690: std_logic; attribute dont_touch of G7690: signal is true;
	signal G7691: std_logic; attribute dont_touch of G7691: signal is true;
	signal G7692: std_logic; attribute dont_touch of G7692: signal is true;
	signal G7693: std_logic; attribute dont_touch of G7693: signal is true;
	signal G7694: std_logic; attribute dont_touch of G7694: signal is true;
	signal G7695: std_logic; attribute dont_touch of G7695: signal is true;
	signal G7696: std_logic; attribute dont_touch of G7696: signal is true;
	signal G7697: std_logic; attribute dont_touch of G7697: signal is true;
	signal G7698: std_logic; attribute dont_touch of G7698: signal is true;
	signal G7699: std_logic; attribute dont_touch of G7699: signal is true;
	signal G7700: std_logic; attribute dont_touch of G7700: signal is true;
	signal G7701: std_logic; attribute dont_touch of G7701: signal is true;
	signal G7702: std_logic; attribute dont_touch of G7702: signal is true;
	signal G7703: std_logic; attribute dont_touch of G7703: signal is true;
	signal G7704: std_logic; attribute dont_touch of G7704: signal is true;
	signal G7705: std_logic; attribute dont_touch of G7705: signal is true;
	signal G7708: std_logic; attribute dont_touch of G7708: signal is true;
	signal G7709: std_logic; attribute dont_touch of G7709: signal is true;
	signal G7710: std_logic; attribute dont_touch of G7710: signal is true;
	signal G7711: std_logic; attribute dont_touch of G7711: signal is true;
	signal G7712: std_logic; attribute dont_touch of G7712: signal is true;
	signal G7713: std_logic; attribute dont_touch of G7713: signal is true;
	signal G7714: std_logic; attribute dont_touch of G7714: signal is true;
	signal G7715: std_logic; attribute dont_touch of G7715: signal is true;
	signal G7716: std_logic; attribute dont_touch of G7716: signal is true;
	signal G7717: std_logic; attribute dont_touch of G7717: signal is true;
	signal G7718: std_logic; attribute dont_touch of G7718: signal is true;
	signal G7719: std_logic; attribute dont_touch of G7719: signal is true;
	signal G7720: std_logic; attribute dont_touch of G7720: signal is true;
	signal G7721: std_logic; attribute dont_touch of G7721: signal is true;
	signal G7722: std_logic; attribute dont_touch of G7722: signal is true;
	signal G7723: std_logic; attribute dont_touch of G7723: signal is true;
	signal G7724: std_logic; attribute dont_touch of G7724: signal is true;
	signal G7725: std_logic; attribute dont_touch of G7725: signal is true;
	signal G7726: std_logic; attribute dont_touch of G7726: signal is true;
	signal G7727: std_logic; attribute dont_touch of G7727: signal is true;
	signal G7728: std_logic; attribute dont_touch of G7728: signal is true;
	signal G7733: std_logic; attribute dont_touch of G7733: signal is true;
	signal G7734: std_logic; attribute dont_touch of G7734: signal is true;
	signal G7735: std_logic; attribute dont_touch of G7735: signal is true;
	signal G7736: std_logic; attribute dont_touch of G7736: signal is true;
	signal G7737: std_logic; attribute dont_touch of G7737: signal is true;
	signal G7738: std_logic; attribute dont_touch of G7738: signal is true;
	signal G7739: std_logic; attribute dont_touch of G7739: signal is true;
	signal G7740: std_logic; attribute dont_touch of G7740: signal is true;
	signal G7741: std_logic; attribute dont_touch of G7741: signal is true;
	signal G7742: std_logic; attribute dont_touch of G7742: signal is true;
	signal G7743: std_logic; attribute dont_touch of G7743: signal is true;
	signal G7744: std_logic; attribute dont_touch of G7744: signal is true;
	signal G7745: std_logic; attribute dont_touch of G7745: signal is true;
	signal G7746: std_logic; attribute dont_touch of G7746: signal is true;
	signal G7747: std_logic; attribute dont_touch of G7747: signal is true;
	signal G7748: std_logic; attribute dont_touch of G7748: signal is true;
	signal G7749: std_logic; attribute dont_touch of G7749: signal is true;
	signal G7750: std_logic; attribute dont_touch of G7750: signal is true;
	signal G7751: std_logic; attribute dont_touch of G7751: signal is true;
	signal G7752: std_logic; attribute dont_touch of G7752: signal is true;
	signal G7753: std_logic; attribute dont_touch of G7753: signal is true;
	signal G7754: std_logic; attribute dont_touch of G7754: signal is true;
	signal G7755: std_logic; attribute dont_touch of G7755: signal is true;
	signal G7756: std_logic; attribute dont_touch of G7756: signal is true;
	signal G7757: std_logic; attribute dont_touch of G7757: signal is true;
	signal G7758: std_logic; attribute dont_touch of G7758: signal is true;
	signal G7759: std_logic; attribute dont_touch of G7759: signal is true;
	signal G7760: std_logic; attribute dont_touch of G7760: signal is true;
	signal G7761: std_logic; attribute dont_touch of G7761: signal is true;
	signal G7762: std_logic; attribute dont_touch of G7762: signal is true;
	signal G7764: std_logic; attribute dont_touch of G7764: signal is true;
	signal G7765: std_logic; attribute dont_touch of G7765: signal is true;
	signal G7766: std_logic; attribute dont_touch of G7766: signal is true;
	signal G7767: std_logic; attribute dont_touch of G7767: signal is true;
	signal G7768: std_logic; attribute dont_touch of G7768: signal is true;
	signal G7769: std_logic; attribute dont_touch of G7769: signal is true;
	signal G7770: std_logic; attribute dont_touch of G7770: signal is true;
	signal G7771: std_logic; attribute dont_touch of G7771: signal is true;
	signal G7772: std_logic; attribute dont_touch of G7772: signal is true;
	signal G7773: std_logic; attribute dont_touch of G7773: signal is true;
	signal G7774: std_logic; attribute dont_touch of G7774: signal is true;
	signal G7775: std_logic; attribute dont_touch of G7775: signal is true;
	signal G7776: std_logic; attribute dont_touch of G7776: signal is true;
	signal G7777: std_logic; attribute dont_touch of G7777: signal is true;
	signal G7778: std_logic; attribute dont_touch of G7778: signal is true;
	signal G7779: std_logic; attribute dont_touch of G7779: signal is true;
	signal G7780: std_logic; attribute dont_touch of G7780: signal is true;
	signal G7781: std_logic; attribute dont_touch of G7781: signal is true;
	signal G7782: std_logic; attribute dont_touch of G7782: signal is true;
	signal G7783: std_logic; attribute dont_touch of G7783: signal is true;
	signal G7784: std_logic; attribute dont_touch of G7784: signal is true;
	signal G7787: std_logic; attribute dont_touch of G7787: signal is true;
	signal G7788: std_logic; attribute dont_touch of G7788: signal is true;
	signal G7789: std_logic; attribute dont_touch of G7789: signal is true;
	signal G7790: std_logic; attribute dont_touch of G7790: signal is true;
	signal G7791: std_logic; attribute dont_touch of G7791: signal is true;
	signal G7792: std_logic; attribute dont_touch of G7792: signal is true;
	signal G7793: std_logic; attribute dont_touch of G7793: signal is true;
	signal G7810: std_logic; attribute dont_touch of G7810: signal is true;
	signal G7811: std_logic; attribute dont_touch of G7811: signal is true;
	signal G7825: std_logic; attribute dont_touch of G7825: signal is true;
	signal G7826: std_logic; attribute dont_touch of G7826: signal is true;
	signal G7827: std_logic; attribute dont_touch of G7827: signal is true;
	signal G7828: std_logic; attribute dont_touch of G7828: signal is true;
	signal G7829: std_logic; attribute dont_touch of G7829: signal is true;
	signal G7832: std_logic; attribute dont_touch of G7832: signal is true;
	signal G7833: std_logic; attribute dont_touch of G7833: signal is true;
	signal G7834: std_logic; attribute dont_touch of G7834: signal is true;
	signal G7835: std_logic; attribute dont_touch of G7835: signal is true;
	signal G7836: std_logic; attribute dont_touch of G7836: signal is true;
	signal G7837: std_logic; attribute dont_touch of G7837: signal is true;
	signal G7838: std_logic; attribute dont_touch of G7838: signal is true;
	signal G7855: std_logic; attribute dont_touch of G7855: signal is true;
	signal G7870: std_logic; attribute dont_touch of G7870: signal is true;
	signal G7887: std_logic; attribute dont_touch of G7887: signal is true;
	signal G7904: std_logic; attribute dont_touch of G7904: signal is true;
	signal G7905: std_logic; attribute dont_touch of G7905: signal is true;
	signal G7920: std_logic; attribute dont_touch of G7920: signal is true;
	signal G7937: std_logic; attribute dont_touch of G7937: signal is true;
	signal G7951: std_logic; attribute dont_touch of G7951: signal is true;
	signal G7966: std_logic; attribute dont_touch of G7966: signal is true;
	signal G7983: std_logic; attribute dont_touch of G7983: signal is true;
	signal G7992: std_logic; attribute dont_touch of G7992: signal is true;
	signal G7993: std_logic; attribute dont_touch of G7993: signal is true;
	signal G8008: std_logic; attribute dont_touch of G8008: signal is true;
	signal G8009: std_logic; attribute dont_touch of G8009: signal is true;
	signal G8012: std_logic; attribute dont_touch of G8012: signal is true;
	signal G8013: std_logic; attribute dont_touch of G8013: signal is true;
	signal G8014: std_logic; attribute dont_touch of G8014: signal is true;
	signal G8015: std_logic; attribute dont_touch of G8015: signal is true;
	signal G8016: std_logic; attribute dont_touch of G8016: signal is true;
	signal G8017: std_logic; attribute dont_touch of G8017: signal is true;
	signal G8018: std_logic; attribute dont_touch of G8018: signal is true;
	signal G8029: std_logic; attribute dont_touch of G8029: signal is true;
	signal G8038: std_logic; attribute dont_touch of G8038: signal is true;
	signal G8039: std_logic; attribute dont_touch of G8039: signal is true;
	signal G8040: std_logic; attribute dont_touch of G8040: signal is true;
	signal G8041: std_logic; attribute dont_touch of G8041: signal is true;
	signal G8042: std_logic; attribute dont_touch of G8042: signal is true;
	signal G8059: std_logic; attribute dont_touch of G8059: signal is true;
	signal G8060: std_logic; attribute dont_touch of G8060: signal is true;
	signal G8061: std_logic; attribute dont_touch of G8061: signal is true;
	signal G8062: std_logic; attribute dont_touch of G8062: signal is true;
	signal G8063: std_logic; attribute dont_touch of G8063: signal is true;
	signal G8064: std_logic; attribute dont_touch of G8064: signal is true;
	signal G8065: std_logic; attribute dont_touch of G8065: signal is true;
	signal G8066: std_logic; attribute dont_touch of G8066: signal is true;
	signal G8067: std_logic; attribute dont_touch of G8067: signal is true;
	signal G8068: std_logic; attribute dont_touch of G8068: signal is true;
	signal G8069: std_logic; attribute dont_touch of G8069: signal is true;
	signal G8070: std_logic; attribute dont_touch of G8070: signal is true;
	signal G8071: std_logic; attribute dont_touch of G8071: signal is true;
	signal G8072: std_logic; attribute dont_touch of G8072: signal is true;
	signal G8073: std_logic; attribute dont_touch of G8073: signal is true;
	signal G8074: std_logic; attribute dont_touch of G8074: signal is true;
	signal G8075: std_logic; attribute dont_touch of G8075: signal is true;
	signal G8076: std_logic; attribute dont_touch of G8076: signal is true;
	signal G8077: std_logic; attribute dont_touch of G8077: signal is true;
	signal G8078: std_logic; attribute dont_touch of G8078: signal is true;
	signal G8079: std_logic; attribute dont_touch of G8079: signal is true;
	signal G8080: std_logic; attribute dont_touch of G8080: signal is true;
	signal G8081: std_logic; attribute dont_touch of G8081: signal is true;
	signal G8082: std_logic; attribute dont_touch of G8082: signal is true;
	signal G8087: std_logic; attribute dont_touch of G8087: signal is true;
	signal G8088: std_logic; attribute dont_touch of G8088: signal is true;
	signal G8089: std_logic; attribute dont_touch of G8089: signal is true;
	signal G8090: std_logic; attribute dont_touch of G8090: signal is true;
	signal G8091: std_logic; attribute dont_touch of G8091: signal is true;
	signal G8092: std_logic; attribute dont_touch of G8092: signal is true;
	signal G8093: std_logic; attribute dont_touch of G8093: signal is true;
	signal G8094: std_logic; attribute dont_touch of G8094: signal is true;
	signal G8111: std_logic; attribute dont_touch of G8111: signal is true;
	signal G8128: std_logic; attribute dont_touch of G8128: signal is true;
	signal G8131: std_logic; attribute dont_touch of G8131: signal is true;
	signal G8145: std_logic; attribute dont_touch of G8145: signal is true;
	signal G8146: std_logic; attribute dont_touch of G8146: signal is true;
	signal G8147: std_logic; attribute dont_touch of G8147: signal is true;
	signal G8150: std_logic; attribute dont_touch of G8150: signal is true;
	signal G8151: std_logic; attribute dont_touch of G8151: signal is true;
	signal G8152: std_logic; attribute dont_touch of G8152: signal is true;
	signal G8153: std_logic; attribute dont_touch of G8153: signal is true;
	signal G8154: std_logic; attribute dont_touch of G8154: signal is true;
	signal G8155: std_logic; attribute dont_touch of G8155: signal is true;
	signal G8156: std_logic; attribute dont_touch of G8156: signal is true;
	signal G8172: std_logic; attribute dont_touch of G8172: signal is true;
	signal G8173: std_logic; attribute dont_touch of G8173: signal is true;
	signal G8174: std_logic; attribute dont_touch of G8174: signal is true;
	signal G8175: std_logic; attribute dont_touch of G8175: signal is true;
	signal G8176: std_logic; attribute dont_touch of G8176: signal is true;
	signal G8177: std_logic; attribute dont_touch of G8177: signal is true;
	signal G8178: std_logic; attribute dont_touch of G8178: signal is true;
	signal G8179: std_logic; attribute dont_touch of G8179: signal is true;
	signal G8180: std_logic; attribute dont_touch of G8180: signal is true;
	signal G8181: std_logic; attribute dont_touch of G8181: signal is true;
	signal G8198: std_logic; attribute dont_touch of G8198: signal is true;
	signal G8199: std_logic; attribute dont_touch of G8199: signal is true;
	signal G8220: std_logic; attribute dont_touch of G8220: signal is true;
	signal G8221: std_logic; attribute dont_touch of G8221: signal is true;
	signal G8222: std_logic; attribute dont_touch of G8222: signal is true;
	signal G8223: std_logic; attribute dont_touch of G8223: signal is true;
	signal G8224: std_logic; attribute dont_touch of G8224: signal is true;
	signal G8225: std_logic; attribute dont_touch of G8225: signal is true;
	signal G8226: std_logic; attribute dont_touch of G8226: signal is true;
	signal G8227: std_logic; attribute dont_touch of G8227: signal is true;
	signal G8228: std_logic; attribute dont_touch of G8228: signal is true;
	signal G8229: std_logic; attribute dont_touch of G8229: signal is true;
	signal G8230: std_logic; attribute dont_touch of G8230: signal is true;
	signal G8231: std_logic; attribute dont_touch of G8231: signal is true;
	signal G8232: std_logic; attribute dont_touch of G8232: signal is true;
	signal G8233: std_logic; attribute dont_touch of G8233: signal is true;
	signal G8235: std_logic; attribute dont_touch of G8235: signal is true;
	signal G8236: std_logic; attribute dont_touch of G8236: signal is true;
	signal G8237: std_logic; attribute dont_touch of G8237: signal is true;
	signal G8238: std_logic; attribute dont_touch of G8238: signal is true;
	signal G8239: std_logic; attribute dont_touch of G8239: signal is true;
	signal G8256: std_logic; attribute dont_touch of G8256: signal is true;
	signal G8257: std_logic; attribute dont_touch of G8257: signal is true;
	signal G8258: std_logic; attribute dont_touch of G8258: signal is true;
	signal G8259: std_logic; attribute dont_touch of G8259: signal is true;
	signal G8260: std_logic; attribute dont_touch of G8260: signal is true;
	signal G8261: std_logic; attribute dont_touch of G8261: signal is true;
	signal G8262: std_logic; attribute dont_touch of G8262: signal is true;
	signal G8263: std_logic; attribute dont_touch of G8263: signal is true;
	signal G8264: std_logic; attribute dont_touch of G8264: signal is true;
	signal G8265: std_logic; attribute dont_touch of G8265: signal is true;
	signal G8266: std_logic; attribute dont_touch of G8266: signal is true;
	signal G8267: std_logic; attribute dont_touch of G8267: signal is true;
	signal G8268: std_logic; attribute dont_touch of G8268: signal is true;
	signal G8269: std_logic; attribute dont_touch of G8269: signal is true;
	signal G8270: std_logic; attribute dont_touch of G8270: signal is true;
	signal G8271: std_logic; attribute dont_touch of G8271: signal is true;
	signal G8272: std_logic; attribute dont_touch of G8272: signal is true;
	signal G8273: std_logic; attribute dont_touch of G8273: signal is true;
	signal G8274: std_logic; attribute dont_touch of G8274: signal is true;
	signal G8275: std_logic; attribute dont_touch of G8275: signal is true;
	signal G8276: std_logic; attribute dont_touch of G8276: signal is true;
	signal G8277: std_logic; attribute dont_touch of G8277: signal is true;
	signal G8278: std_logic; attribute dont_touch of G8278: signal is true;
	signal G8279: std_logic; attribute dont_touch of G8279: signal is true;
	signal G8280: std_logic; attribute dont_touch of G8280: signal is true;
	signal G8281: std_logic; attribute dont_touch of G8281: signal is true;
	signal G8282: std_logic; attribute dont_touch of G8282: signal is true;
	signal G8283: std_logic; attribute dont_touch of G8283: signal is true;
	signal G8284: std_logic; attribute dont_touch of G8284: signal is true;
	signal G8285: std_logic; attribute dont_touch of G8285: signal is true;
	signal G8286: std_logic; attribute dont_touch of G8286: signal is true;
	signal G8287: std_logic; attribute dont_touch of G8287: signal is true;
	signal G8288: std_logic; attribute dont_touch of G8288: signal is true;
	signal G8289: std_logic; attribute dont_touch of G8289: signal is true;
	signal G8290: std_logic; attribute dont_touch of G8290: signal is true;
	signal G8291: std_logic; attribute dont_touch of G8291: signal is true;
	signal G8292: std_logic; attribute dont_touch of G8292: signal is true;
	signal G8293: std_logic; attribute dont_touch of G8293: signal is true;
	signal G8294: std_logic; attribute dont_touch of G8294: signal is true;
	signal G8295: std_logic; attribute dont_touch of G8295: signal is true;
	signal G8296: std_logic; attribute dont_touch of G8296: signal is true;
	signal G8297: std_logic; attribute dont_touch of G8297: signal is true;
	signal G8298: std_logic; attribute dont_touch of G8298: signal is true;
	signal G8299: std_logic; attribute dont_touch of G8299: signal is true;
	signal G8300: std_logic; attribute dont_touch of G8300: signal is true;
	signal G8301: std_logic; attribute dont_touch of G8301: signal is true;
	signal G8302: std_logic; attribute dont_touch of G8302: signal is true;
	signal G8303: std_logic; attribute dont_touch of G8303: signal is true;
	signal G8304: std_logic; attribute dont_touch of G8304: signal is true;
	signal G8305: std_logic; attribute dont_touch of G8305: signal is true;
	signal G8306: std_logic; attribute dont_touch of G8306: signal is true;
	signal G8307: std_logic; attribute dont_touch of G8307: signal is true;
	signal G8308: std_logic; attribute dont_touch of G8308: signal is true;
	signal G8309: std_logic; attribute dont_touch of G8309: signal is true;
	signal G8310: std_logic; attribute dont_touch of G8310: signal is true;
	signal G8311: std_logic; attribute dont_touch of G8311: signal is true;
	signal G8312: std_logic; attribute dont_touch of G8312: signal is true;
	signal G8313: std_logic; attribute dont_touch of G8313: signal is true;
	signal G8314: std_logic; attribute dont_touch of G8314: signal is true;
	signal G8315: std_logic; attribute dont_touch of G8315: signal is true;
	signal G8316: std_logic; attribute dont_touch of G8316: signal is true;
	signal G8317: std_logic; attribute dont_touch of G8317: signal is true;
	signal G8318: std_logic; attribute dont_touch of G8318: signal is true;
	signal G8319: std_logic; attribute dont_touch of G8319: signal is true;
	signal G8320: std_logic; attribute dont_touch of G8320: signal is true;
	signal G8321: std_logic; attribute dont_touch of G8321: signal is true;
	signal G8322: std_logic; attribute dont_touch of G8322: signal is true;
	signal G8323: std_logic; attribute dont_touch of G8323: signal is true;
	signal G8324: std_logic; attribute dont_touch of G8324: signal is true;
	signal G8325: std_logic; attribute dont_touch of G8325: signal is true;
	signal G8326: std_logic; attribute dont_touch of G8326: signal is true;
	signal G8327: std_logic; attribute dont_touch of G8327: signal is true;
	signal G8328: std_logic; attribute dont_touch of G8328: signal is true;
	signal G8329: std_logic; attribute dont_touch of G8329: signal is true;
	signal G8330: std_logic; attribute dont_touch of G8330: signal is true;
	signal G8331: std_logic; attribute dont_touch of G8331: signal is true;
	signal G8332: std_logic; attribute dont_touch of G8332: signal is true;
	signal G8333: std_logic; attribute dont_touch of G8333: signal is true;
	signal G8334: std_logic; attribute dont_touch of G8334: signal is true;
	signal G8335: std_logic; attribute dont_touch of G8335: signal is true;
	signal G8336: std_logic; attribute dont_touch of G8336: signal is true;
	signal G8337: std_logic; attribute dont_touch of G8337: signal is true;
	signal G8338: std_logic; attribute dont_touch of G8338: signal is true;
	signal G8339: std_logic; attribute dont_touch of G8339: signal is true;
	signal G8340: std_logic; attribute dont_touch of G8340: signal is true;
	signal G8341: std_logic; attribute dont_touch of G8341: signal is true;
	signal G8342: std_logic; attribute dont_touch of G8342: signal is true;
	signal G8359: std_logic; attribute dont_touch of G8359: signal is true;
	signal G8360: std_logic; attribute dont_touch of G8360: signal is true;
	signal G8361: std_logic; attribute dont_touch of G8361: signal is true;
	signal G8362: std_logic; attribute dont_touch of G8362: signal is true;
	signal G8363: std_logic; attribute dont_touch of G8363: signal is true;
	signal G8377: std_logic; attribute dont_touch of G8377: signal is true;
	signal G8378: std_logic; attribute dont_touch of G8378: signal is true;
	signal G8379: std_logic; attribute dont_touch of G8379: signal is true;
	signal G8380: std_logic; attribute dont_touch of G8380: signal is true;
	signal G8381: std_logic; attribute dont_touch of G8381: signal is true;
	signal G8382: std_logic; attribute dont_touch of G8382: signal is true;
	signal G8383: std_logic; attribute dont_touch of G8383: signal is true;
	signal G8384: std_logic; attribute dont_touch of G8384: signal is true;
	signal G8385: std_logic; attribute dont_touch of G8385: signal is true;
	signal G8386: std_logic; attribute dont_touch of G8386: signal is true;
	signal G8403: std_logic; attribute dont_touch of G8403: signal is true;
	signal G8404: std_logic; attribute dont_touch of G8404: signal is true;
	signal G8405: std_logic; attribute dont_touch of G8405: signal is true;
	signal G8406: std_logic; attribute dont_touch of G8406: signal is true;
	signal G8407: std_logic; attribute dont_touch of G8407: signal is true;
	signal G8421: std_logic; attribute dont_touch of G8421: signal is true;
	signal G8438: std_logic; attribute dont_touch of G8438: signal is true;
	signal G8439: std_logic; attribute dont_touch of G8439: signal is true;
	signal G8440: std_logic; attribute dont_touch of G8440: signal is true;
	signal G8441: std_logic; attribute dont_touch of G8441: signal is true;
	signal G8442: std_logic; attribute dont_touch of G8442: signal is true;
	signal G8443: std_logic; attribute dont_touch of G8443: signal is true;
	signal G8455: std_logic; attribute dont_touch of G8455: signal is true;
	signal G8456: std_logic; attribute dont_touch of G8456: signal is true;
	signal G8457: std_logic; attribute dont_touch of G8457: signal is true;
	signal G8458: std_logic; attribute dont_touch of G8458: signal is true;
	signal G8459: std_logic; attribute dont_touch of G8459: signal is true;
	signal G8460: std_logic; attribute dont_touch of G8460: signal is true;
	signal G8461: std_logic; attribute dont_touch of G8461: signal is true;
	signal G8462: std_logic; attribute dont_touch of G8462: signal is true;
	signal G8463: std_logic; attribute dont_touch of G8463: signal is true;
	signal G8464: std_logic; attribute dont_touch of G8464: signal is true;
	signal G8481: std_logic; attribute dont_touch of G8481: signal is true;
	signal G8482: std_logic; attribute dont_touch of G8482: signal is true;
	signal G8483: std_logic; attribute dont_touch of G8483: signal is true;
	signal G8493: std_logic; attribute dont_touch of G8493: signal is true;
	signal G8510: std_logic; attribute dont_touch of G8510: signal is true;
	signal G8511: std_logic; attribute dont_touch of G8511: signal is true;
	signal G8512: std_logic; attribute dont_touch of G8512: signal is true;
	signal G8513: std_logic; attribute dont_touch of G8513: signal is true;
	signal G8514: std_logic; attribute dont_touch of G8514: signal is true;
	signal G8523: std_logic; attribute dont_touch of G8523: signal is true;
	signal G8524: std_logic; attribute dont_touch of G8524: signal is true;
	signal G8541: std_logic; attribute dont_touch of G8541: signal is true;
	signal G8542: std_logic; attribute dont_touch of G8542: signal is true;
	signal G8543: std_logic; attribute dont_touch of G8543: signal is true;
	signal G8544: std_logic; attribute dont_touch of G8544: signal is true;
	signal G8545: std_logic; attribute dont_touch of G8545: signal is true;
	signal G8562: std_logic; attribute dont_touch of G8562: signal is true;
	signal G8563: std_logic; attribute dont_touch of G8563: signal is true;
	signal G8564: std_logic; attribute dont_touch of G8564: signal is true;
	signal G8581: std_logic; attribute dont_touch of G8581: signal is true;
	signal G8582: std_logic; attribute dont_touch of G8582: signal is true;
	signal G8583: std_logic; attribute dont_touch of G8583: signal is true;
	signal G8584: std_logic; attribute dont_touch of G8584: signal is true;
	signal G8585: std_logic; attribute dont_touch of G8585: signal is true;
	signal G8602: std_logic; attribute dont_touch of G8602: signal is true;
	signal G8603: std_logic; attribute dont_touch of G8603: signal is true;
	signal G8604: std_logic; attribute dont_touch of G8604: signal is true;
	signal G8605: std_logic; attribute dont_touch of G8605: signal is true;
	signal G8606: std_logic; attribute dont_touch of G8606: signal is true;
	signal G8607: std_logic; attribute dont_touch of G8607: signal is true;
	signal G8608: std_logic; attribute dont_touch of G8608: signal is true;
	signal G8609: std_logic; attribute dont_touch of G8609: signal is true;
	signal G8610: std_logic; attribute dont_touch of G8610: signal is true;
	signal G8611: std_logic; attribute dont_touch of G8611: signal is true;
	signal G8612: std_logic; attribute dont_touch of G8612: signal is true;
	signal G8613: std_logic; attribute dont_touch of G8613: signal is true;
	signal G8619: std_logic; attribute dont_touch of G8619: signal is true;
	signal G8620: std_logic; attribute dont_touch of G8620: signal is true;
	signal G8621: std_logic; attribute dont_touch of G8621: signal is true;
	signal G8622: std_logic; attribute dont_touch of G8622: signal is true;
	signal G8623: std_logic; attribute dont_touch of G8623: signal is true;
	signal G8624: std_logic; attribute dont_touch of G8624: signal is true;
	signal G8625: std_logic; attribute dont_touch of G8625: signal is true;
	signal G8626: std_logic; attribute dont_touch of G8626: signal is true;
	signal G8627: std_logic; attribute dont_touch of G8627: signal is true;
	signal G8628: std_logic; attribute dont_touch of G8628: signal is true;
	signal G8629: std_logic; attribute dont_touch of G8629: signal is true;
	signal G8630: std_logic; attribute dont_touch of G8630: signal is true;
	signal G8631: std_logic; attribute dont_touch of G8631: signal is true;
	signal G8632: std_logic; attribute dont_touch of G8632: signal is true;
	signal G8633: std_logic; attribute dont_touch of G8633: signal is true;
	signal G8634: std_logic; attribute dont_touch of G8634: signal is true;
	signal G8635: std_logic; attribute dont_touch of G8635: signal is true;
	signal G8636: std_logic; attribute dont_touch of G8636: signal is true;
	signal G8637: std_logic; attribute dont_touch of G8637: signal is true;
	signal G8638: std_logic; attribute dont_touch of G8638: signal is true;
	signal G8639: std_logic; attribute dont_touch of G8639: signal is true;
	signal G8640: std_logic; attribute dont_touch of G8640: signal is true;
	signal G8641: std_logic; attribute dont_touch of G8641: signal is true;
	signal G8642: std_logic; attribute dont_touch of G8642: signal is true;
	signal G8643: std_logic; attribute dont_touch of G8643: signal is true;
	signal G8644: std_logic; attribute dont_touch of G8644: signal is true;
	signal G8645: std_logic; attribute dont_touch of G8645: signal is true;
	signal G8646: std_logic; attribute dont_touch of G8646: signal is true;
	signal G8647: std_logic; attribute dont_touch of G8647: signal is true;
	signal G8648: std_logic; attribute dont_touch of G8648: signal is true;
	signal G8649: std_logic; attribute dont_touch of G8649: signal is true;
	signal G8650: std_logic; attribute dont_touch of G8650: signal is true;
	signal G8651: std_logic; attribute dont_touch of G8651: signal is true;
	signal G8652: std_logic; attribute dont_touch of G8652: signal is true;
	signal G8653: std_logic; attribute dont_touch of G8653: signal is true;
	signal G8654: std_logic; attribute dont_touch of G8654: signal is true;
	signal G8655: std_logic; attribute dont_touch of G8655: signal is true;
	signal G8656: std_logic; attribute dont_touch of G8656: signal is true;
	signal G8657: std_logic; attribute dont_touch of G8657: signal is true;
	signal G8658: std_logic; attribute dont_touch of G8658: signal is true;
	signal G8659: std_logic; attribute dont_touch of G8659: signal is true;
	signal G8660: std_logic; attribute dont_touch of G8660: signal is true;
	signal G8662: std_logic; attribute dont_touch of G8662: signal is true;
	signal G8664: std_logic; attribute dont_touch of G8664: signal is true;
	signal G8665: std_logic; attribute dont_touch of G8665: signal is true;
	signal G8666: std_logic; attribute dont_touch of G8666: signal is true;
	signal G8667: std_logic; attribute dont_touch of G8667: signal is true;
	signal G8668: std_logic; attribute dont_touch of G8668: signal is true;
	signal G8669: std_logic; attribute dont_touch of G8669: signal is true;
	signal G8670: std_logic; attribute dont_touch of G8670: signal is true;
	signal G8671: std_logic; attribute dont_touch of G8671: signal is true;
	signal G8672: std_logic; attribute dont_touch of G8672: signal is true;
	signal G8673: std_logic; attribute dont_touch of G8673: signal is true;
	signal G8674: std_logic; attribute dont_touch of G8674: signal is true;
	signal G8675: std_logic; attribute dont_touch of G8675: signal is true;
	signal G8676: std_logic; attribute dont_touch of G8676: signal is true;
	signal G8677: std_logic; attribute dont_touch of G8677: signal is true;
	signal G8678: std_logic; attribute dont_touch of G8678: signal is true;
	signal G8679: std_logic; attribute dont_touch of G8679: signal is true;
	signal G8680: std_logic; attribute dont_touch of G8680: signal is true;
	signal G8681: std_logic; attribute dont_touch of G8681: signal is true;
	signal G8682: std_logic; attribute dont_touch of G8682: signal is true;
	signal G8683: std_logic; attribute dont_touch of G8683: signal is true;
	signal G8684: std_logic; attribute dont_touch of G8684: signal is true;
	signal G8685: std_logic; attribute dont_touch of G8685: signal is true;
	signal G8686: std_logic; attribute dont_touch of G8686: signal is true;
	signal G8687: std_logic; attribute dont_touch of G8687: signal is true;
	signal G8688: std_logic; attribute dont_touch of G8688: signal is true;
	signal G8689: std_logic; attribute dont_touch of G8689: signal is true;
	signal G8690: std_logic; attribute dont_touch of G8690: signal is true;
	signal G8691: std_logic; attribute dont_touch of G8691: signal is true;
	signal G8692: std_logic; attribute dont_touch of G8692: signal is true;
	signal G8693: std_logic; attribute dont_touch of G8693: signal is true;
	signal G8694: std_logic; attribute dont_touch of G8694: signal is true;
	signal G8695: std_logic; attribute dont_touch of G8695: signal is true;
	signal G8696: std_logic; attribute dont_touch of G8696: signal is true;
	signal G8697: std_logic; attribute dont_touch of G8697: signal is true;
	signal G8698: std_logic; attribute dont_touch of G8698: signal is true;
	signal G8699: std_logic; attribute dont_touch of G8699: signal is true;
	signal G8700: std_logic; attribute dont_touch of G8700: signal is true;
	signal G8701: std_logic; attribute dont_touch of G8701: signal is true;
	signal G8702: std_logic; attribute dont_touch of G8702: signal is true;
	signal G8703: std_logic; attribute dont_touch of G8703: signal is true;
	signal G8704: std_logic; attribute dont_touch of G8704: signal is true;
	signal G8705: std_logic; attribute dont_touch of G8705: signal is true;
	signal G8706: std_logic; attribute dont_touch of G8706: signal is true;
	signal G8707: std_logic; attribute dont_touch of G8707: signal is true;
	signal G8708: std_logic; attribute dont_touch of G8708: signal is true;
	signal G8709: std_logic; attribute dont_touch of G8709: signal is true;
	signal G8710: std_logic; attribute dont_touch of G8710: signal is true;
	signal G8711: std_logic; attribute dont_touch of G8711: signal is true;
	signal G8712: std_logic; attribute dont_touch of G8712: signal is true;
	signal G8713: std_logic; attribute dont_touch of G8713: signal is true;
	signal G8714: std_logic; attribute dont_touch of G8714: signal is true;
	signal G8715: std_logic; attribute dont_touch of G8715: signal is true;
	signal G8716: std_logic; attribute dont_touch of G8716: signal is true;
	signal G8717: std_logic; attribute dont_touch of G8717: signal is true;
	signal G8718: std_logic; attribute dont_touch of G8718: signal is true;
	signal G8719: std_logic; attribute dont_touch of G8719: signal is true;
	signal G8720: std_logic; attribute dont_touch of G8720: signal is true;
	signal G8721: std_logic; attribute dont_touch of G8721: signal is true;
	signal G8722: std_logic; attribute dont_touch of G8722: signal is true;
	signal G8723: std_logic; attribute dont_touch of G8723: signal is true;
	signal G8724: std_logic; attribute dont_touch of G8724: signal is true;
	signal G8725: std_logic; attribute dont_touch of G8725: signal is true;
	signal G8726: std_logic; attribute dont_touch of G8726: signal is true;
	signal G8727: std_logic; attribute dont_touch of G8727: signal is true;
	signal G8728: std_logic; attribute dont_touch of G8728: signal is true;
	signal G8729: std_logic; attribute dont_touch of G8729: signal is true;
	signal G8730: std_logic; attribute dont_touch of G8730: signal is true;
	signal G8731: std_logic; attribute dont_touch of G8731: signal is true;
	signal G8732: std_logic; attribute dont_touch of G8732: signal is true;
	signal G8733: std_logic; attribute dont_touch of G8733: signal is true;
	signal G8734: std_logic; attribute dont_touch of G8734: signal is true;
	signal G8735: std_logic; attribute dont_touch of G8735: signal is true;
	signal G8736: std_logic; attribute dont_touch of G8736: signal is true;
	signal G8737: std_logic; attribute dont_touch of G8737: signal is true;
	signal G8738: std_logic; attribute dont_touch of G8738: signal is true;
	signal G8739: std_logic; attribute dont_touch of G8739: signal is true;
	signal G8740: std_logic; attribute dont_touch of G8740: signal is true;
	signal G8741: std_logic; attribute dont_touch of G8741: signal is true;
	signal G8742: std_logic; attribute dont_touch of G8742: signal is true;
	signal G8743: std_logic; attribute dont_touch of G8743: signal is true;
	signal G8744: std_logic; attribute dont_touch of G8744: signal is true;
	signal G8745: std_logic; attribute dont_touch of G8745: signal is true;
	signal G8746: std_logic; attribute dont_touch of G8746: signal is true;
	signal G8747: std_logic; attribute dont_touch of G8747: signal is true;
	signal G8748: std_logic; attribute dont_touch of G8748: signal is true;
	signal G8749: std_logic; attribute dont_touch of G8749: signal is true;
	signal G8750: std_logic; attribute dont_touch of G8750: signal is true;
	signal G8751: std_logic; attribute dont_touch of G8751: signal is true;
	signal G8752: std_logic; attribute dont_touch of G8752: signal is true;
	signal G8753: std_logic; attribute dont_touch of G8753: signal is true;
	signal G8754: std_logic; attribute dont_touch of G8754: signal is true;
	signal G8755: std_logic; attribute dont_touch of G8755: signal is true;
	signal G8756: std_logic; attribute dont_touch of G8756: signal is true;
	signal G8757: std_logic; attribute dont_touch of G8757: signal is true;
	signal G8758: std_logic; attribute dont_touch of G8758: signal is true;
	signal G8759: std_logic; attribute dont_touch of G8759: signal is true;
	signal G8760: std_logic; attribute dont_touch of G8760: signal is true;
	signal G8761: std_logic; attribute dont_touch of G8761: signal is true;
	signal G8762: std_logic; attribute dont_touch of G8762: signal is true;
	signal G8763: std_logic; attribute dont_touch of G8763: signal is true;
	signal G8764: std_logic; attribute dont_touch of G8764: signal is true;
	signal G8765: std_logic; attribute dont_touch of G8765: signal is true;
	signal G8766: std_logic; attribute dont_touch of G8766: signal is true;
	signal G8767: std_logic; attribute dont_touch of G8767: signal is true;
	signal G8768: std_logic; attribute dont_touch of G8768: signal is true;
	signal G8769: std_logic; attribute dont_touch of G8769: signal is true;
	signal G8770: std_logic; attribute dont_touch of G8770: signal is true;
	signal G8771: std_logic; attribute dont_touch of G8771: signal is true;
	signal G8772: std_logic; attribute dont_touch of G8772: signal is true;
	signal G8773: std_logic; attribute dont_touch of G8773: signal is true;
	signal G8774: std_logic; attribute dont_touch of G8774: signal is true;
	signal G8775: std_logic; attribute dont_touch of G8775: signal is true;
	signal G8776: std_logic; attribute dont_touch of G8776: signal is true;
	signal G8777: std_logic; attribute dont_touch of G8777: signal is true;
	signal G8778: std_logic; attribute dont_touch of G8778: signal is true;
	signal G8779: std_logic; attribute dont_touch of G8779: signal is true;
	signal G8780: std_logic; attribute dont_touch of G8780: signal is true;
	signal G8781: std_logic; attribute dont_touch of G8781: signal is true;
	signal G8782: std_logic; attribute dont_touch of G8782: signal is true;
	signal G8783: std_logic; attribute dont_touch of G8783: signal is true;
	signal G8784: std_logic; attribute dont_touch of G8784: signal is true;
	signal G8785: std_logic; attribute dont_touch of G8785: signal is true;
	signal G8786: std_logic; attribute dont_touch of G8786: signal is true;
	signal G8787: std_logic; attribute dont_touch of G8787: signal is true;
	signal G8788: std_logic; attribute dont_touch of G8788: signal is true;
	signal G8789: std_logic; attribute dont_touch of G8789: signal is true;
	signal G8790: std_logic; attribute dont_touch of G8790: signal is true;
	signal G8791: std_logic; attribute dont_touch of G8791: signal is true;
	signal G8792: std_logic; attribute dont_touch of G8792: signal is true;
	signal G8793: std_logic; attribute dont_touch of G8793: signal is true;
	signal G8794: std_logic; attribute dont_touch of G8794: signal is true;
	signal G8795: std_logic; attribute dont_touch of G8795: signal is true;
	signal G8796: std_logic; attribute dont_touch of G8796: signal is true;
	signal G8797: std_logic; attribute dont_touch of G8797: signal is true;
	signal G8798: std_logic; attribute dont_touch of G8798: signal is true;
	signal G8799: std_logic; attribute dont_touch of G8799: signal is true;
	signal G8800: std_logic; attribute dont_touch of G8800: signal is true;
	signal G8801: std_logic; attribute dont_touch of G8801: signal is true;
	signal G8802: std_logic; attribute dont_touch of G8802: signal is true;
	signal G8803: std_logic; attribute dont_touch of G8803: signal is true;
	signal G8804: std_logic; attribute dont_touch of G8804: signal is true;
	signal G8805: std_logic; attribute dont_touch of G8805: signal is true;
	signal G8806: std_logic; attribute dont_touch of G8806: signal is true;
	signal G8807: std_logic; attribute dont_touch of G8807: signal is true;
	signal G8808: std_logic; attribute dont_touch of G8808: signal is true;
	signal G8809: std_logic; attribute dont_touch of G8809: signal is true;
	signal G8810: std_logic; attribute dont_touch of G8810: signal is true;
	signal G8811: std_logic; attribute dont_touch of G8811: signal is true;
	signal G8812: std_logic; attribute dont_touch of G8812: signal is true;
	signal G8813: std_logic; attribute dont_touch of G8813: signal is true;
	signal G8814: std_logic; attribute dont_touch of G8814: signal is true;
	signal G8815: std_logic; attribute dont_touch of G8815: signal is true;
	signal G8816: std_logic; attribute dont_touch of G8816: signal is true;
	signal G8817: std_logic; attribute dont_touch of G8817: signal is true;
	signal G8818: std_logic; attribute dont_touch of G8818: signal is true;
	signal G8819: std_logic; attribute dont_touch of G8819: signal is true;
	signal G8820: std_logic; attribute dont_touch of G8820: signal is true;
	signal G8821: std_logic; attribute dont_touch of G8821: signal is true;
	signal G8822: std_logic; attribute dont_touch of G8822: signal is true;
	signal G8823: std_logic; attribute dont_touch of G8823: signal is true;
	signal G8824: std_logic; attribute dont_touch of G8824: signal is true;
	signal G8825: std_logic; attribute dont_touch of G8825: signal is true;
	signal G8826: std_logic; attribute dont_touch of G8826: signal is true;
	signal G8827: std_logic; attribute dont_touch of G8827: signal is true;
	signal G8828: std_logic; attribute dont_touch of G8828: signal is true;
	signal G8829: std_logic; attribute dont_touch of G8829: signal is true;
	signal G8830: std_logic; attribute dont_touch of G8830: signal is true;
	signal G8831: std_logic; attribute dont_touch of G8831: signal is true;
	signal G8832: std_logic; attribute dont_touch of G8832: signal is true;
	signal G8833: std_logic; attribute dont_touch of G8833: signal is true;
	signal G8834: std_logic; attribute dont_touch of G8834: signal is true;
	signal G8835: std_logic; attribute dont_touch of G8835: signal is true;
	signal G8836: std_logic; attribute dont_touch of G8836: signal is true;
	signal G8837: std_logic; attribute dont_touch of G8837: signal is true;
	signal G8838: std_logic; attribute dont_touch of G8838: signal is true;
	signal G8839: std_logic; attribute dont_touch of G8839: signal is true;
	signal G8840: std_logic; attribute dont_touch of G8840: signal is true;
	signal G8841: std_logic; attribute dont_touch of G8841: signal is true;
	signal G8842: std_logic; attribute dont_touch of G8842: signal is true;
	signal G8843: std_logic; attribute dont_touch of G8843: signal is true;
	signal G8844: std_logic; attribute dont_touch of G8844: signal is true;
	signal G8845: std_logic; attribute dont_touch of G8845: signal is true;
	signal G8846: std_logic; attribute dont_touch of G8846: signal is true;
	signal G8847: std_logic; attribute dont_touch of G8847: signal is true;
	signal G8848: std_logic; attribute dont_touch of G8848: signal is true;
	signal G8849: std_logic; attribute dont_touch of G8849: signal is true;
	signal G8850: std_logic; attribute dont_touch of G8850: signal is true;
	signal G8851: std_logic; attribute dont_touch of G8851: signal is true;
	signal G8852: std_logic; attribute dont_touch of G8852: signal is true;
	signal G8853: std_logic; attribute dont_touch of G8853: signal is true;
	signal G8854: std_logic; attribute dont_touch of G8854: signal is true;
	signal G8855: std_logic; attribute dont_touch of G8855: signal is true;
	signal G8856: std_logic; attribute dont_touch of G8856: signal is true;
	signal G8857: std_logic; attribute dont_touch of G8857: signal is true;
	signal G8858: std_logic; attribute dont_touch of G8858: signal is true;
	signal G8859: std_logic; attribute dont_touch of G8859: signal is true;
	signal G8860: std_logic; attribute dont_touch of G8860: signal is true;
	signal G8861: std_logic; attribute dont_touch of G8861: signal is true;
	signal G8862: std_logic; attribute dont_touch of G8862: signal is true;
	signal G8863: std_logic; attribute dont_touch of G8863: signal is true;
	signal G8864: std_logic; attribute dont_touch of G8864: signal is true;
	signal G8865: std_logic; attribute dont_touch of G8865: signal is true;
	signal G8866: std_logic; attribute dont_touch of G8866: signal is true;
	signal G8867: std_logic; attribute dont_touch of G8867: signal is true;
	signal G8868: std_logic; attribute dont_touch of G8868: signal is true;
	signal G8869: std_logic; attribute dont_touch of G8869: signal is true;
	signal G8870: std_logic; attribute dont_touch of G8870: signal is true;
	signal G8871: std_logic; attribute dont_touch of G8871: signal is true;
	signal G8873: std_logic; attribute dont_touch of G8873: signal is true;
	signal G8874: std_logic; attribute dont_touch of G8874: signal is true;
	signal G8875: std_logic; attribute dont_touch of G8875: signal is true;
	signal G8876: std_logic; attribute dont_touch of G8876: signal is true;
	signal G8877: std_logic; attribute dont_touch of G8877: signal is true;
	signal G8878: std_logic; attribute dont_touch of G8878: signal is true;
	signal G8879: std_logic; attribute dont_touch of G8879: signal is true;
	signal G8880: std_logic; attribute dont_touch of G8880: signal is true;
	signal G8881: std_logic; attribute dont_touch of G8881: signal is true;
	signal G8882: std_logic; attribute dont_touch of G8882: signal is true;
	signal G8883: std_logic; attribute dont_touch of G8883: signal is true;
	signal G8884: std_logic; attribute dont_touch of G8884: signal is true;
	signal G8885: std_logic; attribute dont_touch of G8885: signal is true;
	signal G8886: std_logic; attribute dont_touch of G8886: signal is true;
	signal G8887: std_logic; attribute dont_touch of G8887: signal is true;
	signal G8888: std_logic; attribute dont_touch of G8888: signal is true;
	signal G8889: std_logic; attribute dont_touch of G8889: signal is true;
	signal G8890: std_logic; attribute dont_touch of G8890: signal is true;
	signal G8891: std_logic; attribute dont_touch of G8891: signal is true;
	signal G8892: std_logic; attribute dont_touch of G8892: signal is true;
	signal G8893: std_logic; attribute dont_touch of G8893: signal is true;
	signal G8894: std_logic; attribute dont_touch of G8894: signal is true;
	signal G8895: std_logic; attribute dont_touch of G8895: signal is true;
	signal G8896: std_logic; attribute dont_touch of G8896: signal is true;
	signal G8897: std_logic; attribute dont_touch of G8897: signal is true;
	signal G8898: std_logic; attribute dont_touch of G8898: signal is true;
	signal G8899: std_logic; attribute dont_touch of G8899: signal is true;
	signal G8900: std_logic; attribute dont_touch of G8900: signal is true;
	signal G8901: std_logic; attribute dont_touch of G8901: signal is true;
	signal G8902: std_logic; attribute dont_touch of G8902: signal is true;
	signal G8903: std_logic; attribute dont_touch of G8903: signal is true;
	signal G8904: std_logic; attribute dont_touch of G8904: signal is true;
	signal G8905: std_logic; attribute dont_touch of G8905: signal is true;
	signal G8906: std_logic; attribute dont_touch of G8906: signal is true;
	signal G8907: std_logic; attribute dont_touch of G8907: signal is true;
	signal G8908: std_logic; attribute dont_touch of G8908: signal is true;
	signal G8909: std_logic; attribute dont_touch of G8909: signal is true;
	signal G8910: std_logic; attribute dont_touch of G8910: signal is true;
	signal G8911: std_logic; attribute dont_touch of G8911: signal is true;
	signal G8912: std_logic; attribute dont_touch of G8912: signal is true;
	signal G8913: std_logic; attribute dont_touch of G8913: signal is true;
	signal G8914: std_logic; attribute dont_touch of G8914: signal is true;
	signal G8915: std_logic; attribute dont_touch of G8915: signal is true;
	signal G8916: std_logic; attribute dont_touch of G8916: signal is true;
	signal G8917: std_logic; attribute dont_touch of G8917: signal is true;
	signal G8918: std_logic; attribute dont_touch of G8918: signal is true;
	signal G8919: std_logic; attribute dont_touch of G8919: signal is true;
	signal G8920: std_logic; attribute dont_touch of G8920: signal is true;
	signal G8921: std_logic; attribute dont_touch of G8921: signal is true;
	signal G8922: std_logic; attribute dont_touch of G8922: signal is true;
	signal G8923: std_logic; attribute dont_touch of G8923: signal is true;
	signal G8924: std_logic; attribute dont_touch of G8924: signal is true;
	signal G8925: std_logic; attribute dont_touch of G8925: signal is true;
	signal G8926: std_logic; attribute dont_touch of G8926: signal is true;
	signal G8927: std_logic; attribute dont_touch of G8927: signal is true;
	signal G8928: std_logic; attribute dont_touch of G8928: signal is true;
	signal G8929: std_logic; attribute dont_touch of G8929: signal is true;
	signal G8930: std_logic; attribute dont_touch of G8930: signal is true;
	signal G8931: std_logic; attribute dont_touch of G8931: signal is true;
	signal G8932: std_logic; attribute dont_touch of G8932: signal is true;
	signal G8933: std_logic; attribute dont_touch of G8933: signal is true;
	signal G8934: std_logic; attribute dont_touch of G8934: signal is true;
	signal G8935: std_logic; attribute dont_touch of G8935: signal is true;
	signal G8936: std_logic; attribute dont_touch of G8936: signal is true;
	signal G8937: std_logic; attribute dont_touch of G8937: signal is true;
	signal G8938: std_logic; attribute dont_touch of G8938: signal is true;
	signal G8939: std_logic; attribute dont_touch of G8939: signal is true;
	signal G8940: std_logic; attribute dont_touch of G8940: signal is true;
	signal G8941: std_logic; attribute dont_touch of G8941: signal is true;
	signal G8942: std_logic; attribute dont_touch of G8942: signal is true;
	signal G8943: std_logic; attribute dont_touch of G8943: signal is true;
	signal G8944: std_logic; attribute dont_touch of G8944: signal is true;
	signal G8945: std_logic; attribute dont_touch of G8945: signal is true;
	signal G8946: std_logic; attribute dont_touch of G8946: signal is true;
	signal G8947: std_logic; attribute dont_touch of G8947: signal is true;
	signal G8948: std_logic; attribute dont_touch of G8948: signal is true;
	signal G8949: std_logic; attribute dont_touch of G8949: signal is true;
	signal G8950: std_logic; attribute dont_touch of G8950: signal is true;
	signal G8951: std_logic; attribute dont_touch of G8951: signal is true;
	signal G8952: std_logic; attribute dont_touch of G8952: signal is true;
	signal G8953: std_logic; attribute dont_touch of G8953: signal is true;
	signal G8954: std_logic; attribute dont_touch of G8954: signal is true;
	signal G8955: std_logic; attribute dont_touch of G8955: signal is true;
	signal G8956: std_logic; attribute dont_touch of G8956: signal is true;
	signal G8957: std_logic; attribute dont_touch of G8957: signal is true;
	signal G8959: std_logic; attribute dont_touch of G8959: signal is true;
	signal G8960: std_logic; attribute dont_touch of G8960: signal is true;
	signal G8961: std_logic; attribute dont_touch of G8961: signal is true;
	signal G8962: std_logic; attribute dont_touch of G8962: signal is true;
	signal G8963: std_logic; attribute dont_touch of G8963: signal is true;
	signal G8964: std_logic; attribute dont_touch of G8964: signal is true;
	signal G8965: std_logic; attribute dont_touch of G8965: signal is true;
	signal G8966: std_logic; attribute dont_touch of G8966: signal is true;
	signal G8967: std_logic; attribute dont_touch of G8967: signal is true;
	signal G8968: std_logic; attribute dont_touch of G8968: signal is true;
	signal G8969: std_logic; attribute dont_touch of G8969: signal is true;
	signal G8970: std_logic; attribute dont_touch of G8970: signal is true;
	signal G8971: std_logic; attribute dont_touch of G8971: signal is true;
	signal G8972: std_logic; attribute dont_touch of G8972: signal is true;
	signal G8973: std_logic; attribute dont_touch of G8973: signal is true;
	signal G8974: std_logic; attribute dont_touch of G8974: signal is true;
	signal G8975: std_logic; attribute dont_touch of G8975: signal is true;
	signal G8976: std_logic; attribute dont_touch of G8976: signal is true;
	signal G8977: std_logic; attribute dont_touch of G8977: signal is true;
	signal G8978: std_logic; attribute dont_touch of G8978: signal is true;
	signal G8979: std_logic; attribute dont_touch of G8979: signal is true;
	signal G8980: std_logic; attribute dont_touch of G8980: signal is true;
	signal G8981: std_logic; attribute dont_touch of G8981: signal is true;
	signal G8982: std_logic; attribute dont_touch of G8982: signal is true;
	signal G8983: std_logic; attribute dont_touch of G8983: signal is true;
	signal G8984: std_logic; attribute dont_touch of G8984: signal is true;
	signal G8985: std_logic; attribute dont_touch of G8985: signal is true;
	signal G8986: std_logic; attribute dont_touch of G8986: signal is true;
	signal G8987: std_logic; attribute dont_touch of G8987: signal is true;
	signal G8988: std_logic; attribute dont_touch of G8988: signal is true;
	signal G8989: std_logic; attribute dont_touch of G8989: signal is true;
	signal G8990: std_logic; attribute dont_touch of G8990: signal is true;
	signal G8991: std_logic; attribute dont_touch of G8991: signal is true;
	signal G8992: std_logic; attribute dont_touch of G8992: signal is true;
	signal G8993: std_logic; attribute dont_touch of G8993: signal is true;
	signal G8994: std_logic; attribute dont_touch of G8994: signal is true;
	signal G8995: std_logic; attribute dont_touch of G8995: signal is true;
	signal G8996: std_logic; attribute dont_touch of G8996: signal is true;
	signal G8997: std_logic; attribute dont_touch of G8997: signal is true;
	signal G8998: std_logic; attribute dont_touch of G8998: signal is true;
	signal G8999: std_logic; attribute dont_touch of G8999: signal is true;
	signal G9000: std_logic; attribute dont_touch of G9000: signal is true;
	signal G9001: std_logic; attribute dont_touch of G9001: signal is true;
	signal G9002: std_logic; attribute dont_touch of G9002: signal is true;
	signal G9003: std_logic; attribute dont_touch of G9003: signal is true;
	signal G9004: std_logic; attribute dont_touch of G9004: signal is true;
	signal G9005: std_logic; attribute dont_touch of G9005: signal is true;
	signal G9006: std_logic; attribute dont_touch of G9006: signal is true;
	signal G9007: std_logic; attribute dont_touch of G9007: signal is true;
	signal G9008: std_logic; attribute dont_touch of G9008: signal is true;
	signal G9009: std_logic; attribute dont_touch of G9009: signal is true;
	signal G9010: std_logic; attribute dont_touch of G9010: signal is true;
	signal G9011: std_logic; attribute dont_touch of G9011: signal is true;
	signal G9012: std_logic; attribute dont_touch of G9012: signal is true;
	signal G9013: std_logic; attribute dont_touch of G9013: signal is true;
	signal G9014: std_logic; attribute dont_touch of G9014: signal is true;
	signal G9015: std_logic; attribute dont_touch of G9015: signal is true;
	signal G9016: std_logic; attribute dont_touch of G9016: signal is true;
	signal G9017: std_logic; attribute dont_touch of G9017: signal is true;
	signal G9018: std_logic; attribute dont_touch of G9018: signal is true;
	signal G9019: std_logic; attribute dont_touch of G9019: signal is true;
	signal G9020: std_logic; attribute dont_touch of G9020: signal is true;
	signal G9021: std_logic; attribute dont_touch of G9021: signal is true;
	signal G9022: std_logic; attribute dont_touch of G9022: signal is true;
	signal G9023: std_logic; attribute dont_touch of G9023: signal is true;
	signal G9024: std_logic; attribute dont_touch of G9024: signal is true;
	signal G9025: std_logic; attribute dont_touch of G9025: signal is true;
	signal G9026: std_logic; attribute dont_touch of G9026: signal is true;
	signal G9027: std_logic; attribute dont_touch of G9027: signal is true;
	signal G9028: std_logic; attribute dont_touch of G9028: signal is true;
	signal G9029: std_logic; attribute dont_touch of G9029: signal is true;
	signal G9030: std_logic; attribute dont_touch of G9030: signal is true;
	signal G9031: std_logic; attribute dont_touch of G9031: signal is true;
	signal G9032: std_logic; attribute dont_touch of G9032: signal is true;
	signal G9033: std_logic; attribute dont_touch of G9033: signal is true;
	signal G9034: std_logic; attribute dont_touch of G9034: signal is true;
	signal G9035: std_logic; attribute dont_touch of G9035: signal is true;
	signal G9036: std_logic; attribute dont_touch of G9036: signal is true;
	signal G9037: std_logic; attribute dont_touch of G9037: signal is true;
	signal G9038: std_logic; attribute dont_touch of G9038: signal is true;
	signal G9039: std_logic; attribute dont_touch of G9039: signal is true;
	signal G9042: std_logic; attribute dont_touch of G9042: signal is true;
	signal G9043: std_logic; attribute dont_touch of G9043: signal is true;
	signal G9044: std_logic; attribute dont_touch of G9044: signal is true;
	signal G9045: std_logic; attribute dont_touch of G9045: signal is true;
	signal G9046: std_logic; attribute dont_touch of G9046: signal is true;
	signal G9047: std_logic; attribute dont_touch of G9047: signal is true;
	signal G9048: std_logic; attribute dont_touch of G9048: signal is true;
	signal G9049: std_logic; attribute dont_touch of G9049: signal is true;
	signal G9050: std_logic; attribute dont_touch of G9050: signal is true;
	signal G9051: std_logic; attribute dont_touch of G9051: signal is true;
	signal G9052: std_logic; attribute dont_touch of G9052: signal is true;
	signal G9053: std_logic; attribute dont_touch of G9053: signal is true;
	signal G9054: std_logic; attribute dont_touch of G9054: signal is true;
	signal G9055: std_logic; attribute dont_touch of G9055: signal is true;
	signal G9056: std_logic; attribute dont_touch of G9056: signal is true;
	signal G9057: std_logic; attribute dont_touch of G9057: signal is true;
	signal G9058: std_logic; attribute dont_touch of G9058: signal is true;
	signal G9059: std_logic; attribute dont_touch of G9059: signal is true;
	signal G9060: std_logic; attribute dont_touch of G9060: signal is true;
	signal G9061: std_logic; attribute dont_touch of G9061: signal is true;
	signal G9062: std_logic; attribute dont_touch of G9062: signal is true;
	signal G9063: std_logic; attribute dont_touch of G9063: signal is true;
	signal G9064: std_logic; attribute dont_touch of G9064: signal is true;
	signal G9065: std_logic; attribute dont_touch of G9065: signal is true;
	signal G9066: std_logic; attribute dont_touch of G9066: signal is true;
	signal G9067: std_logic; attribute dont_touch of G9067: signal is true;
	signal G9068: std_logic; attribute dont_touch of G9068: signal is true;
	signal G9069: std_logic; attribute dont_touch of G9069: signal is true;
	signal G9070: std_logic; attribute dont_touch of G9070: signal is true;
	signal G9071: std_logic; attribute dont_touch of G9071: signal is true;
	signal G9072: std_logic; attribute dont_touch of G9072: signal is true;
	signal G9073: std_logic; attribute dont_touch of G9073: signal is true;
	signal G9074: std_logic; attribute dont_touch of G9074: signal is true;
	signal G9075: std_logic; attribute dont_touch of G9075: signal is true;
	signal G9076: std_logic; attribute dont_touch of G9076: signal is true;
	signal G9077: std_logic; attribute dont_touch of G9077: signal is true;
	signal G9078: std_logic; attribute dont_touch of G9078: signal is true;
	signal G9079: std_logic; attribute dont_touch of G9079: signal is true;
	signal G9080: std_logic; attribute dont_touch of G9080: signal is true;
	signal G9081: std_logic; attribute dont_touch of G9081: signal is true;
	signal G9082: std_logic; attribute dont_touch of G9082: signal is true;
	signal G9083: std_logic; attribute dont_touch of G9083: signal is true;
	signal G9084: std_logic; attribute dont_touch of G9084: signal is true;
	signal G9085: std_logic; attribute dont_touch of G9085: signal is true;
	signal G9086: std_logic; attribute dont_touch of G9086: signal is true;
	signal G9087: std_logic; attribute dont_touch of G9087: signal is true;
	signal G9088: std_logic; attribute dont_touch of G9088: signal is true;
	signal G9089: std_logic; attribute dont_touch of G9089: signal is true;
	signal G9090: std_logic; attribute dont_touch of G9090: signal is true;
	signal G9091: std_logic; attribute dont_touch of G9091: signal is true;
	signal G9092: std_logic; attribute dont_touch of G9092: signal is true;
	signal G9093: std_logic; attribute dont_touch of G9093: signal is true;
	signal G9094: std_logic; attribute dont_touch of G9094: signal is true;
	signal G9095: std_logic; attribute dont_touch of G9095: signal is true;
	signal G9096: std_logic; attribute dont_touch of G9096: signal is true;
	signal G9097: std_logic; attribute dont_touch of G9097: signal is true;
	signal G9098: std_logic; attribute dont_touch of G9098: signal is true;
	signal G9099: std_logic; attribute dont_touch of G9099: signal is true;
	signal G9100: std_logic; attribute dont_touch of G9100: signal is true;
	signal G9101: std_logic; attribute dont_touch of G9101: signal is true;
	signal G9102: std_logic; attribute dont_touch of G9102: signal is true;
	signal G9103: std_logic; attribute dont_touch of G9103: signal is true;
	signal G9104: std_logic; attribute dont_touch of G9104: signal is true;
	signal G9105: std_logic; attribute dont_touch of G9105: signal is true;
	signal G9106: std_logic; attribute dont_touch of G9106: signal is true;
	signal G9107: std_logic; attribute dont_touch of G9107: signal is true;
	signal G9108: std_logic; attribute dont_touch of G9108: signal is true;
	signal G9109: std_logic; attribute dont_touch of G9109: signal is true;
	signal G9110: std_logic; attribute dont_touch of G9110: signal is true;
	signal G9111: std_logic; attribute dont_touch of G9111: signal is true;
	signal G9112: std_logic; attribute dont_touch of G9112: signal is true;
	signal G9113: std_logic; attribute dont_touch of G9113: signal is true;
	signal G9114: std_logic; attribute dont_touch of G9114: signal is true;
	signal G9115: std_logic; attribute dont_touch of G9115: signal is true;
	signal G9116: std_logic; attribute dont_touch of G9116: signal is true;
	signal G9117: std_logic; attribute dont_touch of G9117: signal is true;
	signal G9118: std_logic; attribute dont_touch of G9118: signal is true;
	signal G9119: std_logic; attribute dont_touch of G9119: signal is true;
	signal G9120: std_logic; attribute dont_touch of G9120: signal is true;
	signal G9121: std_logic; attribute dont_touch of G9121: signal is true;
	signal G9122: std_logic; attribute dont_touch of G9122: signal is true;
	signal G9123: std_logic; attribute dont_touch of G9123: signal is true;
	signal G9124: std_logic; attribute dont_touch of G9124: signal is true;
	signal G9125: std_logic; attribute dont_touch of G9125: signal is true;
	signal G9126: std_logic; attribute dont_touch of G9126: signal is true;
	signal G9127: std_logic; attribute dont_touch of G9127: signal is true;
	signal G9129: std_logic; attribute dont_touch of G9129: signal is true;
	signal G9130: std_logic; attribute dont_touch of G9130: signal is true;
	signal G9131: std_logic; attribute dont_touch of G9131: signal is true;
	signal G9133: std_logic; attribute dont_touch of G9133: signal is true;
	signal G9134: std_logic; attribute dont_touch of G9134: signal is true;
	signal G9135: std_logic; attribute dont_touch of G9135: signal is true;
	signal G9136: std_logic; attribute dont_touch of G9136: signal is true;
	signal G9137: std_logic; attribute dont_touch of G9137: signal is true;
	signal G9138: std_logic; attribute dont_touch of G9138: signal is true;
	signal G9139: std_logic; attribute dont_touch of G9139: signal is true;
	signal G9140: std_logic; attribute dont_touch of G9140: signal is true;
	signal G9141: std_logic; attribute dont_touch of G9141: signal is true;
	signal G9142: std_logic; attribute dont_touch of G9142: signal is true;
	signal G9143: std_logic; attribute dont_touch of G9143: signal is true;
	signal G9144: std_logic; attribute dont_touch of G9144: signal is true;
	signal G9145: std_logic; attribute dont_touch of G9145: signal is true;
	signal G9146: std_logic; attribute dont_touch of G9146: signal is true;
	signal G9147: std_logic; attribute dont_touch of G9147: signal is true;
	signal G9148: std_logic; attribute dont_touch of G9148: signal is true;
	signal G9151: std_logic; attribute dont_touch of G9151: signal is true;
	signal G9154: std_logic; attribute dont_touch of G9154: signal is true;
	signal G9157: std_logic; attribute dont_touch of G9157: signal is true;
	signal G9158: std_logic; attribute dont_touch of G9158: signal is true;
	signal G9159: std_logic; attribute dont_touch of G9159: signal is true;
	signal G9160: std_logic; attribute dont_touch of G9160: signal is true;
	signal G9161: std_logic; attribute dont_touch of G9161: signal is true;
	signal G9162: std_logic; attribute dont_touch of G9162: signal is true;
	signal G9165: std_logic; attribute dont_touch of G9165: signal is true;
	signal G9168: std_logic; attribute dont_touch of G9168: signal is true;
	signal G9171: std_logic; attribute dont_touch of G9171: signal is true;
	signal G9174: std_logic; attribute dont_touch of G9174: signal is true;
	signal G9177: std_logic; attribute dont_touch of G9177: signal is true;
	signal G9178: std_logic; attribute dont_touch of G9178: signal is true;
	signal G9179: std_logic; attribute dont_touch of G9179: signal is true;
	signal G9180: std_logic; attribute dont_touch of G9180: signal is true;
	signal G9181: std_logic; attribute dont_touch of G9181: signal is true;
	signal G9182: std_logic; attribute dont_touch of G9182: signal is true;
	signal G9183: std_logic; attribute dont_touch of G9183: signal is true;
	signal G9184: std_logic; attribute dont_touch of G9184: signal is true;
	signal G9185: std_logic; attribute dont_touch of G9185: signal is true;
	signal G9186: std_logic; attribute dont_touch of G9186: signal is true;
	signal G9187: std_logic; attribute dont_touch of G9187: signal is true;
	signal G9188: std_logic; attribute dont_touch of G9188: signal is true;
	signal G9189: std_logic; attribute dont_touch of G9189: signal is true;
	signal G9190: std_logic; attribute dont_touch of G9190: signal is true;
	signal G9191: std_logic; attribute dont_touch of G9191: signal is true;
	signal G9192: std_logic; attribute dont_touch of G9192: signal is true;
	signal G9193: std_logic; attribute dont_touch of G9193: signal is true;
	signal G9194: std_logic; attribute dont_touch of G9194: signal is true;
	signal G9195: std_logic; attribute dont_touch of G9195: signal is true;
	signal G9196: std_logic; attribute dont_touch of G9196: signal is true;
	signal G9197: std_logic; attribute dont_touch of G9197: signal is true;
	signal G9198: std_logic; attribute dont_touch of G9198: signal is true;
	signal G9199: std_logic; attribute dont_touch of G9199: signal is true;
	signal G9200: std_logic; attribute dont_touch of G9200: signal is true;
	signal G9201: std_logic; attribute dont_touch of G9201: signal is true;
	signal G9202: std_logic; attribute dont_touch of G9202: signal is true;
	signal G9203: std_logic; attribute dont_touch of G9203: signal is true;
	signal G9205: std_logic; attribute dont_touch of G9205: signal is true;
	signal G9206: std_logic; attribute dont_touch of G9206: signal is true;
	signal G9207: std_logic; attribute dont_touch of G9207: signal is true;
	signal G9208: std_logic; attribute dont_touch of G9208: signal is true;
	signal G9209: std_logic; attribute dont_touch of G9209: signal is true;
	signal G9210: std_logic; attribute dont_touch of G9210: signal is true;
	signal G9211: std_logic; attribute dont_touch of G9211: signal is true;
	signal G9212: std_logic; attribute dont_touch of G9212: signal is true;
	signal G9213: std_logic; attribute dont_touch of G9213: signal is true;
	signal G9214: std_logic; attribute dont_touch of G9214: signal is true;
	signal G9215: std_logic; attribute dont_touch of G9215: signal is true;
	signal G9216: std_logic; attribute dont_touch of G9216: signal is true;
	signal G9217: std_logic; attribute dont_touch of G9217: signal is true;
	signal G9218: std_logic; attribute dont_touch of G9218: signal is true;
	signal G9219: std_logic; attribute dont_touch of G9219: signal is true;
	signal G9220: std_logic; attribute dont_touch of G9220: signal is true;
	signal G9221: std_logic; attribute dont_touch of G9221: signal is true;
	signal G9222: std_logic; attribute dont_touch of G9222: signal is true;
	signal G9223: std_logic; attribute dont_touch of G9223: signal is true;
	signal G9226: std_logic; attribute dont_touch of G9226: signal is true;
	signal G9227: std_logic; attribute dont_touch of G9227: signal is true;
	signal G9230: std_logic; attribute dont_touch of G9230: signal is true;
	signal G9233: std_logic; attribute dont_touch of G9233: signal is true;
	signal G9234: std_logic; attribute dont_touch of G9234: signal is true;
	signal G9235: std_logic; attribute dont_touch of G9235: signal is true;
	signal G9236: std_logic; attribute dont_touch of G9236: signal is true;
	signal G9237: std_logic; attribute dont_touch of G9237: signal is true;
	signal G9238: std_logic; attribute dont_touch of G9238: signal is true;
	signal G9239: std_logic; attribute dont_touch of G9239: signal is true;
	signal G9240: std_logic; attribute dont_touch of G9240: signal is true;
	signal G9241: std_logic; attribute dont_touch of G9241: signal is true;
	signal G9244: std_logic; attribute dont_touch of G9244: signal is true;
	signal G9247: std_logic; attribute dont_touch of G9247: signal is true;
	signal G9248: std_logic; attribute dont_touch of G9248: signal is true;
	signal G9251: std_logic; attribute dont_touch of G9251: signal is true;
	signal G9252: std_logic; attribute dont_touch of G9252: signal is true;
	signal G9255: std_logic; attribute dont_touch of G9255: signal is true;
	signal G9258: std_logic; attribute dont_touch of G9258: signal is true;
	signal G9259: std_logic; attribute dont_touch of G9259: signal is true;
	signal G9260: std_logic; attribute dont_touch of G9260: signal is true;
	signal G9261: std_logic; attribute dont_touch of G9261: signal is true;
	signal G9264: std_logic; attribute dont_touch of G9264: signal is true;
	signal G9267: std_logic; attribute dont_touch of G9267: signal is true;
	signal G9270: std_logic; attribute dont_touch of G9270: signal is true;
	signal G9271: std_logic; attribute dont_touch of G9271: signal is true;
	signal G9272: std_logic; attribute dont_touch of G9272: signal is true;
	signal G9273: std_logic; attribute dont_touch of G9273: signal is true;
	signal G9274: std_logic; attribute dont_touch of G9274: signal is true;
	signal G9275: std_logic; attribute dont_touch of G9275: signal is true;
	signal G9276: std_logic; attribute dont_touch of G9276: signal is true;
	signal G9277: std_logic; attribute dont_touch of G9277: signal is true;
	signal G9278: std_logic; attribute dont_touch of G9278: signal is true;
	signal G9279: std_logic; attribute dont_touch of G9279: signal is true;
	signal G9281: std_logic; attribute dont_touch of G9281: signal is true;
	signal G9282: std_logic; attribute dont_touch of G9282: signal is true;
	signal G9285: std_logic; attribute dont_touch of G9285: signal is true;
	signal G9288: std_logic; attribute dont_touch of G9288: signal is true;
	signal G9291: std_logic; attribute dont_touch of G9291: signal is true;
	signal G9294: std_logic; attribute dont_touch of G9294: signal is true;
	signal G9298: std_logic; attribute dont_touch of G9298: signal is true;
	signal G9300: std_logic; attribute dont_touch of G9300: signal is true;
	signal G9301: std_logic; attribute dont_touch of G9301: signal is true;
	signal G9302: std_logic; attribute dont_touch of G9302: signal is true;
	signal G9303: std_logic; attribute dont_touch of G9303: signal is true;
	signal G9304: std_logic; attribute dont_touch of G9304: signal is true;
	signal G9306: std_logic; attribute dont_touch of G9306: signal is true;
	signal G9307: std_logic; attribute dont_touch of G9307: signal is true;
	signal G9309: std_logic; attribute dont_touch of G9309: signal is true;
	signal G9311: std_logic; attribute dont_touch of G9311: signal is true;
	signal G9313: std_logic; attribute dont_touch of G9313: signal is true;
	signal G9315: std_logic; attribute dont_touch of G9315: signal is true;
	signal G9316: std_logic; attribute dont_touch of G9316: signal is true;
	signal G9317: std_logic; attribute dont_touch of G9317: signal is true;
	signal G9318: std_logic; attribute dont_touch of G9318: signal is true;
	signal G9319: std_logic; attribute dont_touch of G9319: signal is true;
	signal G9320: std_logic; attribute dont_touch of G9320: signal is true;
	signal G9321: std_logic; attribute dont_touch of G9321: signal is true;
	signal G9322: std_logic; attribute dont_touch of G9322: signal is true;
	signal G9323: std_logic; attribute dont_touch of G9323: signal is true;
	signal G9324: std_logic; attribute dont_touch of G9324: signal is true;
	signal G9327: std_logic; attribute dont_touch of G9327: signal is true;
	signal G9328: std_logic; attribute dont_touch of G9328: signal is true;
	signal G9329: std_logic; attribute dont_touch of G9329: signal is true;
	signal G9330: std_logic; attribute dont_touch of G9330: signal is true;
	signal G9331: std_logic; attribute dont_touch of G9331: signal is true;
	signal G9332: std_logic; attribute dont_touch of G9332: signal is true;
	signal G9333: std_logic; attribute dont_touch of G9333: signal is true;
	signal G9334: std_logic; attribute dont_touch of G9334: signal is true;
	signal G9335: std_logic; attribute dont_touch of G9335: signal is true;
	signal G9336: std_logic; attribute dont_touch of G9336: signal is true;
	signal G9337: std_logic; attribute dont_touch of G9337: signal is true;
	signal G9338: std_logic; attribute dont_touch of G9338: signal is true;
	signal G9339: std_logic; attribute dont_touch of G9339: signal is true;
	signal G9340: std_logic; attribute dont_touch of G9340: signal is true;
	signal G9343: std_logic; attribute dont_touch of G9343: signal is true;
	signal G9344: std_logic; attribute dont_touch of G9344: signal is true;
	signal G9345: std_logic; attribute dont_touch of G9345: signal is true;
	signal G9346: std_logic; attribute dont_touch of G9346: signal is true;
	signal G9347: std_logic; attribute dont_touch of G9347: signal is true;
	signal G9348: std_logic; attribute dont_touch of G9348: signal is true;
	signal G9349: std_logic; attribute dont_touch of G9349: signal is true;
	signal G9350: std_logic; attribute dont_touch of G9350: signal is true;
	signal G9351: std_logic; attribute dont_touch of G9351: signal is true;
	signal G9352: std_logic; attribute dont_touch of G9352: signal is true;
	signal G9353: std_logic; attribute dont_touch of G9353: signal is true;
	signal G9354: std_logic; attribute dont_touch of G9354: signal is true;
	signal G9355: std_logic; attribute dont_touch of G9355: signal is true;
	signal G9356: std_logic; attribute dont_touch of G9356: signal is true;
	signal G9357: std_logic; attribute dont_touch of G9357: signal is true;
	signal G9358: std_logic; attribute dont_touch of G9358: signal is true;
	signal G9359: std_logic; attribute dont_touch of G9359: signal is true;
	signal G9360: std_logic; attribute dont_touch of G9360: signal is true;
	signal G9361: std_logic; attribute dont_touch of G9361: signal is true;
	signal G9362: std_logic; attribute dont_touch of G9362: signal is true;
	signal G9363: std_logic; attribute dont_touch of G9363: signal is true;
	signal G9366: std_logic; attribute dont_touch of G9366: signal is true;
	signal G9367: std_logic; attribute dont_touch of G9367: signal is true;
	signal G9368: std_logic; attribute dont_touch of G9368: signal is true;
	signal G9369: std_logic; attribute dont_touch of G9369: signal is true;
	signal G9370: std_logic; attribute dont_touch of G9370: signal is true;
	signal G9371: std_logic; attribute dont_touch of G9371: signal is true;
	signal G9372: std_logic; attribute dont_touch of G9372: signal is true;
	signal G9373: std_logic; attribute dont_touch of G9373: signal is true;
	signal G9374: std_logic; attribute dont_touch of G9374: signal is true;
	signal G9375: std_logic; attribute dont_touch of G9375: signal is true;
	signal G9376: std_logic; attribute dont_touch of G9376: signal is true;
	signal G9377: std_logic; attribute dont_touch of G9377: signal is true;
	signal G9379: std_logic; attribute dont_touch of G9379: signal is true;
	signal G9380: std_logic; attribute dont_touch of G9380: signal is true;
	signal G9381: std_logic; attribute dont_touch of G9381: signal is true;
	signal G9382: std_logic; attribute dont_touch of G9382: signal is true;
	signal G9383: std_logic; attribute dont_touch of G9383: signal is true;
	signal G9384: std_logic; attribute dont_touch of G9384: signal is true;
	signal G9385: std_logic; attribute dont_touch of G9385: signal is true;
	signal G9386: std_logic; attribute dont_touch of G9386: signal is true;
	signal G9387: std_logic; attribute dont_touch of G9387: signal is true;
	signal G9388: std_logic; attribute dont_touch of G9388: signal is true;
	signal G9389: std_logic; attribute dont_touch of G9389: signal is true;
	signal I5353: std_logic; attribute dont_touch of I5353: signal is true;
	signal I5356: std_logic; attribute dont_touch of I5356: signal is true;
	signal I5359: std_logic; attribute dont_touch of I5359: signal is true;
	signal I5362: std_logic; attribute dont_touch of I5362: signal is true;
	signal I5365: std_logic; attribute dont_touch of I5365: signal is true;
	signal I5368: std_logic; attribute dont_touch of I5368: signal is true;
	signal I5371: std_logic; attribute dont_touch of I5371: signal is true;
	signal I5374: std_logic; attribute dont_touch of I5374: signal is true;
	signal I5377: std_logic; attribute dont_touch of I5377: signal is true;
	signal I5380: std_logic; attribute dont_touch of I5380: signal is true;
	signal I5383: std_logic; attribute dont_touch of I5383: signal is true;
	signal I5386: std_logic; attribute dont_touch of I5386: signal is true;
	signal I5389: std_logic; attribute dont_touch of I5389: signal is true;
	signal I5392: std_logic; attribute dont_touch of I5392: signal is true;
	signal I5395: std_logic; attribute dont_touch of I5395: signal is true;
	signal I5398: std_logic; attribute dont_touch of I5398: signal is true;
	signal I5401: std_logic; attribute dont_touch of I5401: signal is true;
	signal I5404: std_logic; attribute dont_touch of I5404: signal is true;
	signal I5407: std_logic; attribute dont_touch of I5407: signal is true;
	signal I5410: std_logic; attribute dont_touch of I5410: signal is true;
	signal I5413: std_logic; attribute dont_touch of I5413: signal is true;
	signal I5416: std_logic; attribute dont_touch of I5416: signal is true;
	signal I5419: std_logic; attribute dont_touch of I5419: signal is true;
	signal I5422: std_logic; attribute dont_touch of I5422: signal is true;
	signal I5425: std_logic; attribute dont_touch of I5425: signal is true;
	signal I5428: std_logic; attribute dont_touch of I5428: signal is true;
	signal I5432: std_logic; attribute dont_touch of I5432: signal is true;
	signal I5435: std_logic; attribute dont_touch of I5435: signal is true;
	signal I5466: std_logic; attribute dont_touch of I5466: signal is true;
	signal I5471: std_logic; attribute dont_touch of I5471: signal is true;
	signal I5475: std_logic; attribute dont_touch of I5475: signal is true;
	signal I5478: std_logic; attribute dont_touch of I5478: signal is true;
	signal I5505: std_logic; attribute dont_touch of I5505: signal is true;
	signal I5506: std_logic; attribute dont_touch of I5506: signal is true;
	signal I5507: std_logic; attribute dont_touch of I5507: signal is true;
	signal I5512: std_logic; attribute dont_touch of I5512: signal is true;
	signal I5515: std_logic; attribute dont_touch of I5515: signal is true;
	signal I5519: std_logic; attribute dont_touch of I5519: signal is true;
	signal I5520: std_logic; attribute dont_touch of I5520: signal is true;
	signal I5521: std_logic; attribute dont_touch of I5521: signal is true;
	signal I5528: std_logic; attribute dont_touch of I5528: signal is true;
	signal I5531: std_logic; attribute dont_touch of I5531: signal is true;
	signal I5535: std_logic; attribute dont_touch of I5535: signal is true;
	signal I5542: std_logic; attribute dont_touch of I5542: signal is true;
	signal I5545: std_logic; attribute dont_touch of I5545: signal is true;
	signal I5548: std_logic; attribute dont_touch of I5548: signal is true;
	signal I5552: std_logic; attribute dont_touch of I5552: signal is true;
	signal I5555: std_logic; attribute dont_touch of I5555: signal is true;
	signal I5559: std_logic; attribute dont_touch of I5559: signal is true;
	signal I5562: std_logic; attribute dont_touch of I5562: signal is true;
	signal I5565: std_logic; attribute dont_touch of I5565: signal is true;
	signal I5568: std_logic; attribute dont_touch of I5568: signal is true;
	signal I5577: std_logic; attribute dont_touch of I5577: signal is true;
	signal I5598: std_logic; attribute dont_touch of I5598: signal is true;
	signal I5599: std_logic; attribute dont_touch of I5599: signal is true;
	signal I5600: std_logic; attribute dont_touch of I5600: signal is true;
	signal I5605: std_logic; attribute dont_touch of I5605: signal is true;
	signal I5609: std_logic; attribute dont_touch of I5609: signal is true;
	signal I5616: std_logic; attribute dont_touch of I5616: signal is true;
	signal I5619: std_logic; attribute dont_touch of I5619: signal is true;
	signal I5620: std_logic; attribute dont_touch of I5620: signal is true;
	signal I5621: std_logic; attribute dont_touch of I5621: signal is true;
	signal I5633: std_logic; attribute dont_touch of I5633: signal is true;
	signal I5636: std_logic; attribute dont_touch of I5636: signal is true;
	signal I5646: std_logic; attribute dont_touch of I5646: signal is true;
	signal I5649: std_logic; attribute dont_touch of I5649: signal is true;
	signal I5654: std_logic; attribute dont_touch of I5654: signal is true;
	signal I5657: std_logic; attribute dont_touch of I5657: signal is true;
	signal I5664: std_logic; attribute dont_touch of I5664: signal is true;
	signal I5667: std_logic; attribute dont_touch of I5667: signal is true;
	signal I5670: std_logic; attribute dont_touch of I5670: signal is true;
	signal I5676: std_logic; attribute dont_touch of I5676: signal is true;
	signal I5679: std_logic; attribute dont_touch of I5679: signal is true;
	signal I5682: std_logic; attribute dont_touch of I5682: signal is true;
	signal I5689: std_logic; attribute dont_touch of I5689: signal is true;
	signal I5692: std_logic; attribute dont_touch of I5692: signal is true;
	signal I5695: std_logic; attribute dont_touch of I5695: signal is true;
	signal I5696: std_logic; attribute dont_touch of I5696: signal is true;
	signal I5697: std_logic; attribute dont_touch of I5697: signal is true;
	signal I5706: std_logic; attribute dont_touch of I5706: signal is true;
	signal I5709: std_logic; attribute dont_touch of I5709: signal is true;
	signal I5715: std_logic; attribute dont_touch of I5715: signal is true;
	signal I5718: std_logic; attribute dont_touch of I5718: signal is true;
	signal I5732: std_logic; attribute dont_touch of I5732: signal is true;
	signal I5747: std_logic; attribute dont_touch of I5747: signal is true;
	signal I5751: std_logic; attribute dont_touch of I5751: signal is true;
	signal I5754: std_logic; attribute dont_touch of I5754: signal is true;
	signal I5757: std_logic; attribute dont_touch of I5757: signal is true;
	signal I5763: std_logic; attribute dont_touch of I5763: signal is true;
	signal I5766: std_logic; attribute dont_touch of I5766: signal is true;
	signal I5772: std_logic; attribute dont_touch of I5772: signal is true;
	signal I5775: std_logic; attribute dont_touch of I5775: signal is true;
	signal I5781: std_logic; attribute dont_touch of I5781: signal is true;
	signal I5789: std_logic; attribute dont_touch of I5789: signal is true;
	signal I5795: std_logic; attribute dont_touch of I5795: signal is true;
	signal I5801: std_logic; attribute dont_touch of I5801: signal is true;
	signal I5812: std_logic; attribute dont_touch of I5812: signal is true;
	signal I5817: std_logic; attribute dont_touch of I5817: signal is true;
	signal I5831: std_logic; attribute dont_touch of I5831: signal is true;
	signal I5839: std_logic; attribute dont_touch of I5839: signal is true;
	signal I5842: std_logic; attribute dont_touch of I5842: signal is true;
	signal I5847: std_logic; attribute dont_touch of I5847: signal is true;
	signal I5852: std_logic; attribute dont_touch of I5852: signal is true;
	signal I5855: std_logic; attribute dont_touch of I5855: signal is true;
	signal I5861: std_logic; attribute dont_touch of I5861: signal is true;
	signal I5865: std_logic; attribute dont_touch of I5865: signal is true;
	signal I5868: std_logic; attribute dont_touch of I5868: signal is true;
	signal I5872: std_logic; attribute dont_touch of I5872: signal is true;
	signal I5879: std_logic; attribute dont_touch of I5879: signal is true;
	signal I5883: std_logic; attribute dont_touch of I5883: signal is true;
	signal I5889: std_logic; attribute dont_touch of I5889: signal is true;
	signal I5894: std_logic; attribute dont_touch of I5894: signal is true;
	signal I5897: std_logic; attribute dont_touch of I5897: signal is true;
	signal I5901: std_logic; attribute dont_touch of I5901: signal is true;
	signal I5908: std_logic; attribute dont_touch of I5908: signal is true;
	signal I5911: std_logic; attribute dont_touch of I5911: signal is true;
	signal I5914: std_logic; attribute dont_touch of I5914: signal is true;
	signal I5920: std_logic; attribute dont_touch of I5920: signal is true;
	signal I5923: std_logic; attribute dont_touch of I5923: signal is true;
	signal I5926: std_logic; attribute dont_touch of I5926: signal is true;
	signal I5933: std_logic; attribute dont_touch of I5933: signal is true;
	signal I5936: std_logic; attribute dont_touch of I5936: signal is true;
	signal I5939: std_logic; attribute dont_touch of I5939: signal is true;
	signal I5942: std_logic; attribute dont_touch of I5942: signal is true;
	signal I5945: std_logic; attribute dont_touch of I5945: signal is true;
	signal I5948: std_logic; attribute dont_touch of I5948: signal is true;
	signal I5954: std_logic; attribute dont_touch of I5954: signal is true;
	signal I5957: std_logic; attribute dont_touch of I5957: signal is true;
	signal I5960: std_logic; attribute dont_touch of I5960: signal is true;
	signal I5963: std_logic; attribute dont_touch of I5963: signal is true;
	signal I5966: std_logic; attribute dont_touch of I5966: signal is true;
	signal I5969: std_logic; attribute dont_touch of I5969: signal is true;
	signal I5972: std_logic; attribute dont_touch of I5972: signal is true;
	signal I5975: std_logic; attribute dont_touch of I5975: signal is true;
	signal I5978: std_logic; attribute dont_touch of I5978: signal is true;
	signal I5981: std_logic; attribute dont_touch of I5981: signal is true;
	signal I5984: std_logic; attribute dont_touch of I5984: signal is true;
	signal I5989: std_logic; attribute dont_touch of I5989: signal is true;
	signal I5997: std_logic; attribute dont_touch of I5997: signal is true;
	signal I6000: std_logic; attribute dont_touch of I6000: signal is true;
	signal I6003: std_logic; attribute dont_touch of I6003: signal is true;
	signal I6006: std_logic; attribute dont_touch of I6006: signal is true;
	signal I6009: std_logic; attribute dont_touch of I6009: signal is true;
	signal I6012: std_logic; attribute dont_touch of I6012: signal is true;
	signal I6015: std_logic; attribute dont_touch of I6015: signal is true;
	signal I6018: std_logic; attribute dont_touch of I6018: signal is true;
	signal I6021: std_logic; attribute dont_touch of I6021: signal is true;
	signal I6024: std_logic; attribute dont_touch of I6024: signal is true;
	signal I6029: std_logic; attribute dont_touch of I6029: signal is true;
	signal I6033: std_logic; attribute dont_touch of I6033: signal is true;
	signal I6036: std_logic; attribute dont_touch of I6036: signal is true;
	signal I6039: std_logic; attribute dont_touch of I6039: signal is true;
	signal I6042: std_logic; attribute dont_touch of I6042: signal is true;
	signal I6045: std_logic; attribute dont_touch of I6045: signal is true;
	signal I6048: std_logic; attribute dont_touch of I6048: signal is true;
	signal I6051: std_logic; attribute dont_touch of I6051: signal is true;
	signal I6054: std_logic; attribute dont_touch of I6054: signal is true;
	signal I6057: std_logic; attribute dont_touch of I6057: signal is true;
	signal I6060: std_logic; attribute dont_touch of I6060: signal is true;
	signal I6064: std_logic; attribute dont_touch of I6064: signal is true;
	signal I6065: std_logic; attribute dont_touch of I6065: signal is true;
	signal I6066: std_logic; attribute dont_touch of I6066: signal is true;
	signal I6072: std_logic; attribute dont_touch of I6072: signal is true;
	signal I6075: std_logic; attribute dont_touch of I6075: signal is true;
	signal I6078: std_logic; attribute dont_touch of I6078: signal is true;
	signal I6081: std_logic; attribute dont_touch of I6081: signal is true;
	signal I6084: std_logic; attribute dont_touch of I6084: signal is true;
	signal I6087: std_logic; attribute dont_touch of I6087: signal is true;
	signal I6090: std_logic; attribute dont_touch of I6090: signal is true;
	signal I6093: std_logic; attribute dont_touch of I6093: signal is true;
	signal I6096: std_logic; attribute dont_touch of I6096: signal is true;
	signal I6099: std_logic; attribute dont_touch of I6099: signal is true;
	signal I6102: std_logic; attribute dont_touch of I6102: signal is true;
	signal I6103: std_logic; attribute dont_touch of I6103: signal is true;
	signal I6104: std_logic; attribute dont_touch of I6104: signal is true;
	signal I6109: std_logic; attribute dont_touch of I6109: signal is true;
	signal I6112: std_logic; attribute dont_touch of I6112: signal is true;
	signal I6115: std_logic; attribute dont_touch of I6115: signal is true;
	signal I6118: std_logic; attribute dont_touch of I6118: signal is true;
	signal I6121: std_logic; attribute dont_touch of I6121: signal is true;
	signal I6124: std_logic; attribute dont_touch of I6124: signal is true;
	signal I6127: std_logic; attribute dont_touch of I6127: signal is true;
	signal I6130: std_logic; attribute dont_touch of I6130: signal is true;
	signal I6133: std_logic; attribute dont_touch of I6133: signal is true;
	signal I6134: std_logic; attribute dont_touch of I6134: signal is true;
	signal I6135: std_logic; attribute dont_touch of I6135: signal is true;
	signal I6143: std_logic; attribute dont_touch of I6143: signal is true;
	signal I6148: std_logic; attribute dont_touch of I6148: signal is true;
	signal I6151: std_logic; attribute dont_touch of I6151: signal is true;
	signal I6154: std_logic; attribute dont_touch of I6154: signal is true;
	signal I6157: std_logic; attribute dont_touch of I6157: signal is true;
	signal I6160: std_logic; attribute dont_touch of I6160: signal is true;
	signal I6163: std_logic; attribute dont_touch of I6163: signal is true;
	signal I6166: std_logic; attribute dont_touch of I6166: signal is true;
	signal I6170: std_logic; attribute dont_touch of I6170: signal is true;
	signal I6171: std_logic; attribute dont_touch of I6171: signal is true;
	signal I6172: std_logic; attribute dont_touch of I6172: signal is true;
	signal I6178: std_logic; attribute dont_touch of I6178: signal is true;
	signal I6183: std_logic; attribute dont_touch of I6183: signal is true;
	signal I6186: std_logic; attribute dont_touch of I6186: signal is true;
	signal I6189: std_logic; attribute dont_touch of I6189: signal is true;
	signal I6192: std_logic; attribute dont_touch of I6192: signal is true;
	signal I6195: std_logic; attribute dont_touch of I6195: signal is true;
	signal I6198: std_logic; attribute dont_touch of I6198: signal is true;
	signal I6201: std_logic; attribute dont_touch of I6201: signal is true;
	signal I6202: std_logic; attribute dont_touch of I6202: signal is true;
	signal I6203: std_logic; attribute dont_touch of I6203: signal is true;
	signal I6208: std_logic; attribute dont_touch of I6208: signal is true;
	signal I6209: std_logic; attribute dont_touch of I6209: signal is true;
	signal I6214: std_logic; attribute dont_touch of I6214: signal is true;
	signal I6217: std_logic; attribute dont_touch of I6217: signal is true;
	signal I6220: std_logic; attribute dont_touch of I6220: signal is true;
	signal I6223: std_logic; attribute dont_touch of I6223: signal is true;
	signal I6226: std_logic; attribute dont_touch of I6226: signal is true;
	signal I6229: std_logic; attribute dont_touch of I6229: signal is true;
	signal I6232: std_logic; attribute dont_touch of I6232: signal is true;
	signal I6233: std_logic; attribute dont_touch of I6233: signal is true;
	signal I6234: std_logic; attribute dont_touch of I6234: signal is true;
	signal I6239: std_logic; attribute dont_touch of I6239: signal is true;
	signal I6242: std_logic; attribute dont_touch of I6242: signal is true;
	signal I6245: std_logic; attribute dont_touch of I6245: signal is true;
	signal I6248: std_logic; attribute dont_touch of I6248: signal is true;
	signal I6251: std_logic; attribute dont_touch of I6251: signal is true;
	signal I6254: std_logic; attribute dont_touch of I6254: signal is true;
	signal I6257: std_logic; attribute dont_touch of I6257: signal is true;
	signal I6258: std_logic; attribute dont_touch of I6258: signal is true;
	signal I6259: std_logic; attribute dont_touch of I6259: signal is true;
	signal I6267: std_logic; attribute dont_touch of I6267: signal is true;
	signal I6270: std_logic; attribute dont_touch of I6270: signal is true;
	signal I6273: std_logic; attribute dont_touch of I6273: signal is true;
	signal I6274: std_logic; attribute dont_touch of I6274: signal is true;
	signal I6275: std_logic; attribute dont_touch of I6275: signal is true;
	signal I6286: std_logic; attribute dont_touch of I6286: signal is true;
	signal I6291: std_logic; attribute dont_touch of I6291: signal is true;
	signal I6294: std_logic; attribute dont_touch of I6294: signal is true;
	signal I6299: std_logic; attribute dont_touch of I6299: signal is true;
	signal I6302: std_logic; attribute dont_touch of I6302: signal is true;
	signal I6305: std_logic; attribute dont_touch of I6305: signal is true;
	signal I6309: std_logic; attribute dont_touch of I6309: signal is true;
	signal I6317: std_logic; attribute dont_touch of I6317: signal is true;
	signal I6323: std_logic; attribute dont_touch of I6323: signal is true;
	signal I6326: std_logic; attribute dont_touch of I6326: signal is true;
	signal I6333: std_logic; attribute dont_touch of I6333: signal is true;
	signal I6337: std_logic; attribute dont_touch of I6337: signal is true;
	signal I6341: std_logic; attribute dont_touch of I6341: signal is true;
	signal I6348: std_logic; attribute dont_touch of I6348: signal is true;
	signal I6354: std_logic; attribute dont_touch of I6354: signal is true;
	signal I6358: std_logic; attribute dont_touch of I6358: signal is true;
	signal I6363: std_logic; attribute dont_touch of I6363: signal is true;
	signal I6368: std_logic; attribute dont_touch of I6368: signal is true;
	signal I6371: std_logic; attribute dont_touch of I6371: signal is true;
	signal I6376: std_logic; attribute dont_touch of I6376: signal is true;
	signal I6416: std_logic; attribute dont_touch of I6416: signal is true;
	signal I6419: std_logic; attribute dont_touch of I6419: signal is true;
	signal I6422: std_logic; attribute dont_touch of I6422: signal is true;
	signal I6425: std_logic; attribute dont_touch of I6425: signal is true;
	signal I6428: std_logic; attribute dont_touch of I6428: signal is true;
	signal I6431: std_logic; attribute dont_touch of I6431: signal is true;
	signal I6434: std_logic; attribute dont_touch of I6434: signal is true;
	signal I6437: std_logic; attribute dont_touch of I6437: signal is true;
	signal I6440: std_logic; attribute dont_touch of I6440: signal is true;
	signal I6443: std_logic; attribute dont_touch of I6443: signal is true;
	signal I6446: std_logic; attribute dont_touch of I6446: signal is true;
	signal I6451: std_logic; attribute dont_touch of I6451: signal is true;
	signal I6454: std_logic; attribute dont_touch of I6454: signal is true;
	signal I6457: std_logic; attribute dont_touch of I6457: signal is true;
	signal I6460: std_logic; attribute dont_touch of I6460: signal is true;
	signal I6463: std_logic; attribute dont_touch of I6463: signal is true;
	signal I6468: std_logic; attribute dont_touch of I6468: signal is true;
	signal I6471: std_logic; attribute dont_touch of I6471: signal is true;
	signal I6474: std_logic; attribute dont_touch of I6474: signal is true;
	signal I6499: std_logic; attribute dont_touch of I6499: signal is true;
	signal I6500: std_logic; attribute dont_touch of I6500: signal is true;
	signal I6501: std_logic; attribute dont_touch of I6501: signal is true;
	signal I6509: std_logic; attribute dont_touch of I6509: signal is true;
	signal I6517: std_logic; attribute dont_touch of I6517: signal is true;
	signal I6522: std_logic; attribute dont_touch of I6522: signal is true;
	signal I6523: std_logic; attribute dont_touch of I6523: signal is true;
	signal I6524: std_logic; attribute dont_touch of I6524: signal is true;
	signal I6532: std_logic; attribute dont_touch of I6532: signal is true;
	signal I6538: std_logic; attribute dont_touch of I6538: signal is true;
	signal I6539: std_logic; attribute dont_touch of I6539: signal is true;
	signal I6540: std_logic; attribute dont_touch of I6540: signal is true;
	signal I6553: std_logic; attribute dont_touch of I6553: signal is true;
	signal I6561: std_logic; attribute dont_touch of I6561: signal is true;
	signal I6564: std_logic; attribute dont_touch of I6564: signal is true;
	signal I6571: std_logic; attribute dont_touch of I6571: signal is true;
	signal I6574: std_logic; attribute dont_touch of I6574: signal is true;
	signal I6578: std_logic; attribute dont_touch of I6578: signal is true;
	signal I6587: std_logic; attribute dont_touch of I6587: signal is true;
	signal I6590: std_logic; attribute dont_touch of I6590: signal is true;
	signal I6597: std_logic; attribute dont_touch of I6597: signal is true;
	signal I6608: std_logic; attribute dont_touch of I6608: signal is true;
	signal I6615: std_logic; attribute dont_touch of I6615: signal is true;
	signal I6629: std_logic; attribute dont_touch of I6629: signal is true;
	signal I6636: std_logic; attribute dont_touch of I6636: signal is true;
	signal I6643: std_logic; attribute dont_touch of I6643: signal is true;
	signal I6646: std_logic; attribute dont_touch of I6646: signal is true;
	signal I6652: std_logic; attribute dont_touch of I6652: signal is true;
	signal I6657: std_logic; attribute dont_touch of I6657: signal is true;
	signal I6663: std_logic; attribute dont_touch of I6663: signal is true;
	signal I6669: std_logic; attribute dont_touch of I6669: signal is true;
	signal I6673: std_logic; attribute dont_touch of I6673: signal is true;
	signal I6676: std_logic; attribute dont_touch of I6676: signal is true;
	signal I6680: std_logic; attribute dont_touch of I6680: signal is true;
	signal I6686: std_logic; attribute dont_touch of I6686: signal is true;
	signal I6695: std_logic; attribute dont_touch of I6695: signal is true;
	signal I6703: std_logic; attribute dont_touch of I6703: signal is true;
	signal I6711: std_logic; attribute dont_touch of I6711: signal is true;
	signal I6716: std_logic; attribute dont_touch of I6716: signal is true;
	signal I6723: std_logic; attribute dont_touch of I6723: signal is true;
	signal I6728: std_logic; attribute dont_touch of I6728: signal is true;
	signal I6733: std_logic; attribute dont_touch of I6733: signal is true;
	signal I6739: std_logic; attribute dont_touch of I6739: signal is true;
	signal I6740: std_logic; attribute dont_touch of I6740: signal is true;
	signal I6741: std_logic; attribute dont_touch of I6741: signal is true;
	signal I6750: std_logic; attribute dont_touch of I6750: signal is true;
	signal I6751: std_logic; attribute dont_touch of I6751: signal is true;
	signal I6752: std_logic; attribute dont_touch of I6752: signal is true;
	signal I6757: std_logic; attribute dont_touch of I6757: signal is true;
	signal I6758: std_logic; attribute dont_touch of I6758: signal is true;
	signal I6759: std_logic; attribute dont_touch of I6759: signal is true;
	signal I6764: std_logic; attribute dont_touch of I6764: signal is true;
	signal I6767: std_logic; attribute dont_touch of I6767: signal is true;
	signal I6770: std_logic; attribute dont_touch of I6770: signal is true;
	signal I6774: std_logic; attribute dont_touch of I6774: signal is true;
	signal I6775: std_logic; attribute dont_touch of I6775: signal is true;
	signal I6776: std_logic; attribute dont_touch of I6776: signal is true;
	signal I6784: std_logic; attribute dont_touch of I6784: signal is true;
	signal I6788: std_logic; attribute dont_touch of I6788: signal is true;
	signal I6791: std_logic; attribute dont_touch of I6791: signal is true;
	signal I6795: std_logic; attribute dont_touch of I6795: signal is true;
	signal I6800: std_logic; attribute dont_touch of I6800: signal is true;
	signal I6805: std_logic; attribute dont_touch of I6805: signal is true;
	signal I6813: std_logic; attribute dont_touch of I6813: signal is true;
	signal I6814: std_logic; attribute dont_touch of I6814: signal is true;
	signal I6815: std_logic; attribute dont_touch of I6815: signal is true;
	signal I6820: std_logic; attribute dont_touch of I6820: signal is true;
	signal I6826: std_logic; attribute dont_touch of I6826: signal is true;
	signal I6831: std_logic; attribute dont_touch of I6831: signal is true;
	signal I6834: std_logic; attribute dont_touch of I6834: signal is true;
	signal I6839: std_logic; attribute dont_touch of I6839: signal is true;
	signal I6842: std_logic; attribute dont_touch of I6842: signal is true;
	signal I6843: std_logic; attribute dont_touch of I6843: signal is true;
	signal I6844: std_logic; attribute dont_touch of I6844: signal is true;
	signal I6849: std_logic; attribute dont_touch of I6849: signal is true;
	signal I6853: std_logic; attribute dont_touch of I6853: signal is true;
	signal I6856: std_logic; attribute dont_touch of I6856: signal is true;
	signal I6860: std_logic; attribute dont_touch of I6860: signal is true;
	signal I6864: std_logic; attribute dont_touch of I6864: signal is true;
	signal I6868: std_logic; attribute dont_touch of I6868: signal is true;
	signal I6872: std_logic; attribute dont_touch of I6872: signal is true;
	signal I6876: std_logic; attribute dont_touch of I6876: signal is true;
	signal I6877: std_logic; attribute dont_touch of I6877: signal is true;
	signal I6878: std_logic; attribute dont_touch of I6878: signal is true;
	signal I6887: std_logic; attribute dont_touch of I6887: signal is true;
	signal I6894: std_logic; attribute dont_touch of I6894: signal is true;
	signal I6900: std_logic; attribute dont_touch of I6900: signal is true;
	signal I6904: std_logic; attribute dont_touch of I6904: signal is true;
	signal I6905: std_logic; attribute dont_touch of I6905: signal is true;
	signal I6906: std_logic; attribute dont_touch of I6906: signal is true;
	signal I6911: std_logic; attribute dont_touch of I6911: signal is true;
	signal I6916: std_logic; attribute dont_touch of I6916: signal is true;
	signal I6917: std_logic; attribute dont_touch of I6917: signal is true;
	signal I6918: std_logic; attribute dont_touch of I6918: signal is true;
	signal I6923: std_logic; attribute dont_touch of I6923: signal is true;
	signal I6924: std_logic; attribute dont_touch of I6924: signal is true;
	signal I6925: std_logic; attribute dont_touch of I6925: signal is true;
	signal I6930: std_logic; attribute dont_touch of I6930: signal is true;
	signal I6936: std_logic; attribute dont_touch of I6936: signal is true;
	signal I6939: std_logic; attribute dont_touch of I6939: signal is true;
	signal I6940: std_logic; attribute dont_touch of I6940: signal is true;
	signal I6941: std_logic; attribute dont_touch of I6941: signal is true;
	signal I6946: std_logic; attribute dont_touch of I6946: signal is true;
	signal I6949: std_logic; attribute dont_touch of I6949: signal is true;
	signal I6952: std_logic; attribute dont_touch of I6952: signal is true;
	signal I6956: std_logic; attribute dont_touch of I6956: signal is true;
	signal I6959: std_logic; attribute dont_touch of I6959: signal is true;
	signal I6963: std_logic; attribute dont_touch of I6963: signal is true;
	signal I6970: std_logic; attribute dont_touch of I6970: signal is true;
	signal I6974: std_logic; attribute dont_touch of I6974: signal is true;
	signal I6996: std_logic; attribute dont_touch of I6996: signal is true;
	signal I6997: std_logic; attribute dont_touch of I6997: signal is true;
	signal I6998: std_logic; attribute dont_touch of I6998: signal is true;
	signal I7009: std_logic; attribute dont_touch of I7009: signal is true;
	signal I7010: std_logic; attribute dont_touch of I7010: signal is true;
	signal I7011: std_logic; attribute dont_touch of I7011: signal is true;
	signal I7029: std_logic; attribute dont_touch of I7029: signal is true;
	signal I7036: std_logic; attribute dont_touch of I7036: signal is true;
	signal I7041: std_logic; attribute dont_touch of I7041: signal is true;
	signal I7044: std_logic; attribute dont_touch of I7044: signal is true;
	signal I7053: std_logic; attribute dont_touch of I7053: signal is true;
	signal I7061: std_logic; attribute dont_touch of I7061: signal is true;
	signal I7064: std_logic; attribute dont_touch of I7064: signal is true;
	signal I7068: std_logic; attribute dont_touch of I7068: signal is true;
	signal I7069: std_logic; attribute dont_touch of I7069: signal is true;
	signal I7070: std_logic; attribute dont_touch of I7070: signal is true;
	signal I7079: std_logic; attribute dont_touch of I7079: signal is true;
	signal I7082: std_logic; attribute dont_touch of I7082: signal is true;
	signal I7085: std_logic; attribute dont_touch of I7085: signal is true;
	signal I7086: std_logic; attribute dont_touch of I7086: signal is true;
	signal I7087: std_logic; attribute dont_touch of I7087: signal is true;
	signal I7095: std_logic; attribute dont_touch of I7095: signal is true;
	signal I7098: std_logic; attribute dont_touch of I7098: signal is true;
	signal I7101: std_logic; attribute dont_touch of I7101: signal is true;
	signal I7104: std_logic; attribute dont_touch of I7104: signal is true;
	signal I7107: std_logic; attribute dont_touch of I7107: signal is true;
	signal I7112: std_logic; attribute dont_touch of I7112: signal is true;
	signal I7115: std_logic; attribute dont_touch of I7115: signal is true;
	signal I7118: std_logic; attribute dont_touch of I7118: signal is true;
	signal I7126: std_logic; attribute dont_touch of I7126: signal is true;
	signal I7129: std_logic; attribute dont_touch of I7129: signal is true;
	signal I7132: std_logic; attribute dont_touch of I7132: signal is true;
	signal I7138: std_logic; attribute dont_touch of I7138: signal is true;
	signal I7139: std_logic; attribute dont_touch of I7139: signal is true;
	signal I7140: std_logic; attribute dont_touch of I7140: signal is true;
	signal I7145: std_logic; attribute dont_touch of I7145: signal is true;
	signal I7148: std_logic; attribute dont_touch of I7148: signal is true;
	signal I7149: std_logic; attribute dont_touch of I7149: signal is true;
	signal I7150: std_logic; attribute dont_touch of I7150: signal is true;
	signal I7156: std_logic; attribute dont_touch of I7156: signal is true;
	signal I7157: std_logic; attribute dont_touch of I7157: signal is true;
	signal I7158: std_logic; attribute dont_touch of I7158: signal is true;
	signal I7164: std_logic; attribute dont_touch of I7164: signal is true;
	signal I7167: std_logic; attribute dont_touch of I7167: signal is true;
	signal I7172: std_logic; attribute dont_touch of I7172: signal is true;
	signal I7173: std_logic; attribute dont_touch of I7173: signal is true;
	signal I7174: std_logic; attribute dont_touch of I7174: signal is true;
	signal I7179: std_logic; attribute dont_touch of I7179: signal is true;
	signal I7180: std_logic; attribute dont_touch of I7180: signal is true;
	signal I7181: std_logic; attribute dont_touch of I7181: signal is true;
	signal I7186: std_logic; attribute dont_touch of I7186: signal is true;
	signal I7187: std_logic; attribute dont_touch of I7187: signal is true;
	signal I7188: std_logic; attribute dont_touch of I7188: signal is true;
	signal I7195: std_logic; attribute dont_touch of I7195: signal is true;
	signal I7198: std_logic; attribute dont_touch of I7198: signal is true;
	signal I7204: std_logic; attribute dont_touch of I7204: signal is true;
	signal I7211: std_logic; attribute dont_touch of I7211: signal is true;
	signal I7214: std_logic; attribute dont_touch of I7214: signal is true;
	signal I7215: std_logic; attribute dont_touch of I7215: signal is true;
	signal I7216: std_logic; attribute dont_touch of I7216: signal is true;
	signal I7232: std_logic; attribute dont_touch of I7232: signal is true;
	signal I7233: std_logic; attribute dont_touch of I7233: signal is true;
	signal I7239: std_logic; attribute dont_touch of I7239: signal is true;
	signal I7240: std_logic; attribute dont_touch of I7240: signal is true;
	signal I7241: std_logic; attribute dont_touch of I7241: signal is true;
	signal I7255: std_logic; attribute dont_touch of I7255: signal is true;
	signal I7262: std_logic; attribute dont_touch of I7262: signal is true;
	signal I7268: std_logic; attribute dont_touch of I7268: signal is true;
	signal I7269: std_logic; attribute dont_touch of I7269: signal is true;
	signal I7270: std_logic; attribute dont_touch of I7270: signal is true;
	signal I7277: std_logic; attribute dont_touch of I7277: signal is true;
	signal I7278: std_logic; attribute dont_touch of I7278: signal is true;
	signal I7279: std_logic; attribute dont_touch of I7279: signal is true;
	signal I7287: std_logic; attribute dont_touch of I7287: signal is true;
	signal I7290: std_logic; attribute dont_touch of I7290: signal is true;
	signal I7293: std_logic; attribute dont_touch of I7293: signal is true;
	signal I7296: std_logic; attribute dont_touch of I7296: signal is true;
	signal I7299: std_logic; attribute dont_touch of I7299: signal is true;
	signal I7302: std_logic; attribute dont_touch of I7302: signal is true;
	signal I7305: std_logic; attribute dont_touch of I7305: signal is true;
	signal I7308: std_logic; attribute dont_touch of I7308: signal is true;
	signal I7311: std_logic; attribute dont_touch of I7311: signal is true;
	signal I7314: std_logic; attribute dont_touch of I7314: signal is true;
	signal I7317: std_logic; attribute dont_touch of I7317: signal is true;
	signal I7320: std_logic; attribute dont_touch of I7320: signal is true;
	signal I7323: std_logic; attribute dont_touch of I7323: signal is true;
	signal I7326: std_logic; attribute dont_touch of I7326: signal is true;
	signal I7329: std_logic; attribute dont_touch of I7329: signal is true;
	signal I7332: std_logic; attribute dont_touch of I7332: signal is true;
	signal I7335: std_logic; attribute dont_touch of I7335: signal is true;
	signal I7338: std_logic; attribute dont_touch of I7338: signal is true;
	signal I7341: std_logic; attribute dont_touch of I7341: signal is true;
	signal I7344: std_logic; attribute dont_touch of I7344: signal is true;
	signal I7347: std_logic; attribute dont_touch of I7347: signal is true;
	signal I7350: std_logic; attribute dont_touch of I7350: signal is true;
	signal I7353: std_logic; attribute dont_touch of I7353: signal is true;
	signal I7356: std_logic; attribute dont_touch of I7356: signal is true;
	signal I7359: std_logic; attribute dont_touch of I7359: signal is true;
	signal I7362: std_logic; attribute dont_touch of I7362: signal is true;
	signal I7365: std_logic; attribute dont_touch of I7365: signal is true;
	signal I7368: std_logic; attribute dont_touch of I7368: signal is true;
	signal I7371: std_logic; attribute dont_touch of I7371: signal is true;
	signal I7374: std_logic; attribute dont_touch of I7374: signal is true;
	signal I7377: std_logic; attribute dont_touch of I7377: signal is true;
	signal I7380: std_logic; attribute dont_touch of I7380: signal is true;
	signal I7383: std_logic; attribute dont_touch of I7383: signal is true;
	signal I7386: std_logic; attribute dont_touch of I7386: signal is true;
	signal I7389: std_logic; attribute dont_touch of I7389: signal is true;
	signal I7392: std_logic; attribute dont_touch of I7392: signal is true;
	signal I7400: std_logic; attribute dont_touch of I7400: signal is true;
	signal I7417: std_logic; attribute dont_touch of I7417: signal is true;
	signal I7421: std_logic; attribute dont_touch of I7421: signal is true;
	signal I7422: std_logic; attribute dont_touch of I7422: signal is true;
	signal I7423: std_logic; attribute dont_touch of I7423: signal is true;
	signal I7428: std_logic; attribute dont_touch of I7428: signal is true;
	signal I7429: std_logic; attribute dont_touch of I7429: signal is true;
	signal I7430: std_logic; attribute dont_touch of I7430: signal is true;
	signal I7436: std_logic; attribute dont_touch of I7436: signal is true;
	signal I7437: std_logic; attribute dont_touch of I7437: signal is true;
	signal I7438: std_logic; attribute dont_touch of I7438: signal is true;
	signal I7443: std_logic; attribute dont_touch of I7443: signal is true;
	signal I7444: std_logic; attribute dont_touch of I7444: signal is true;
	signal I7445: std_logic; attribute dont_touch of I7445: signal is true;
	signal I7452: std_logic; attribute dont_touch of I7452: signal is true;
	signal I7453: std_logic; attribute dont_touch of I7453: signal is true;
	signal I7454: std_logic; attribute dont_touch of I7454: signal is true;
	signal I7459: std_logic; attribute dont_touch of I7459: signal is true;
	signal I7460: std_logic; attribute dont_touch of I7460: signal is true;
	signal I7461: std_logic; attribute dont_touch of I7461: signal is true;
	signal I7466: std_logic; attribute dont_touch of I7466: signal is true;
	signal I7467: std_logic; attribute dont_touch of I7467: signal is true;
	signal I7468: std_logic; attribute dont_touch of I7468: signal is true;
	signal I7473: std_logic; attribute dont_touch of I7473: signal is true;
	signal I7478: std_logic; attribute dont_touch of I7478: signal is true;
	signal I7479: std_logic; attribute dont_touch of I7479: signal is true;
	signal I7480: std_logic; attribute dont_touch of I7480: signal is true;
	signal I7485: std_logic; attribute dont_touch of I7485: signal is true;
	signal I7486: std_logic; attribute dont_touch of I7486: signal is true;
	signal I7487: std_logic; attribute dont_touch of I7487: signal is true;
	signal I7492: std_logic; attribute dont_touch of I7492: signal is true;
	signal I7495: std_logic; attribute dont_touch of I7495: signal is true;
	signal I7498: std_logic; attribute dont_touch of I7498: signal is true;
	signal I7503: std_logic; attribute dont_touch of I7503: signal is true;
	signal I7504: std_logic; attribute dont_touch of I7504: signal is true;
	signal I7505: std_logic; attribute dont_touch of I7505: signal is true;
	signal I7510: std_logic; attribute dont_touch of I7510: signal is true;
	signal I7511: std_logic; attribute dont_touch of I7511: signal is true;
	signal I7512: std_logic; attribute dont_touch of I7512: signal is true;
	signal I7517: std_logic; attribute dont_touch of I7517: signal is true;
	signal I7520: std_logic; attribute dont_touch of I7520: signal is true;
	signal I7523: std_logic; attribute dont_touch of I7523: signal is true;
	signal I7526: std_logic; attribute dont_touch of I7526: signal is true;
	signal I7531: std_logic; attribute dont_touch of I7531: signal is true;
	signal I7532: std_logic; attribute dont_touch of I7532: signal is true;
	signal I7533: std_logic; attribute dont_touch of I7533: signal is true;
	signal I7538: std_logic; attribute dont_touch of I7538: signal is true;
	signal I7539: std_logic; attribute dont_touch of I7539: signal is true;
	signal I7540: std_logic; attribute dont_touch of I7540: signal is true;
	signal I7545: std_logic; attribute dont_touch of I7545: signal is true;
	signal I7548: std_logic; attribute dont_touch of I7548: signal is true;
	signal I7551: std_logic; attribute dont_touch of I7551: signal is true;
	signal I7554: std_logic; attribute dont_touch of I7554: signal is true;
	signal I7558: std_logic; attribute dont_touch of I7558: signal is true;
	signal I7561: std_logic; attribute dont_touch of I7561: signal is true;
	signal I7564: std_logic; attribute dont_touch of I7564: signal is true;
	signal I7567: std_logic; attribute dont_touch of I7567: signal is true;
	signal I7568: std_logic; attribute dont_touch of I7568: signal is true;
	signal I7569: std_logic; attribute dont_touch of I7569: signal is true;
	signal I7574: std_logic; attribute dont_touch of I7574: signal is true;
	signal I7575: std_logic; attribute dont_touch of I7575: signal is true;
	signal I7576: std_logic; attribute dont_touch of I7576: signal is true;
	signal I7581: std_logic; attribute dont_touch of I7581: signal is true;
	signal I7584: std_logic; attribute dont_touch of I7584: signal is true;
	signal I7588: std_logic; attribute dont_touch of I7588: signal is true;
	signal I7592: std_logic; attribute dont_touch of I7592: signal is true;
	signal I7595: std_logic; attribute dont_touch of I7595: signal is true;
	signal I7599: std_logic; attribute dont_touch of I7599: signal is true;
	signal I7602: std_logic; attribute dont_touch of I7602: signal is true;
	signal I7605: std_logic; attribute dont_touch of I7605: signal is true;
	signal I7609: std_logic; attribute dont_touch of I7609: signal is true;
	signal I7610: std_logic; attribute dont_touch of I7610: signal is true;
	signal I7611: std_logic; attribute dont_touch of I7611: signal is true;
	signal I7616: std_logic; attribute dont_touch of I7616: signal is true;
	signal I7617: std_logic; attribute dont_touch of I7617: signal is true;
	signal I7618: std_logic; attribute dont_touch of I7618: signal is true;
	signal I7623: std_logic; attribute dont_touch of I7623: signal is true;
	signal I7626: std_logic; attribute dont_touch of I7626: signal is true;
	signal I7629: std_logic; attribute dont_touch of I7629: signal is true;
	signal I7632: std_logic; attribute dont_touch of I7632: signal is true;
	signal I7635: std_logic; attribute dont_touch of I7635: signal is true;
	signal I7640: std_logic; attribute dont_touch of I7640: signal is true;
	signal I7644: std_logic; attribute dont_touch of I7644: signal is true;
	signal I7648: std_logic; attribute dont_touch of I7648: signal is true;
	signal I7651: std_logic; attribute dont_touch of I7651: signal is true;
	signal I7655: std_logic; attribute dont_touch of I7655: signal is true;
	signal I7658: std_logic; attribute dont_touch of I7658: signal is true;
	signal I7662: std_logic; attribute dont_touch of I7662: signal is true;
	signal I7667: std_logic; attribute dont_touch of I7667: signal is true;
	signal I7672: std_logic; attribute dont_touch of I7672: signal is true;
	signal I7676: std_logic; attribute dont_touch of I7676: signal is true;
	signal I7680: std_logic; attribute dont_touch of I7680: signal is true;
	signal I7683: std_logic; attribute dont_touch of I7683: signal is true;
	signal I7688: std_logic; attribute dont_touch of I7688: signal is true;
	signal I7691: std_logic; attribute dont_touch of I7691: signal is true;
	signal I7697: std_logic; attribute dont_touch of I7697: signal is true;
	signal I7702: std_logic; attribute dont_touch of I7702: signal is true;
	signal I7706: std_logic; attribute dont_touch of I7706: signal is true;
	signal I7712: std_logic; attribute dont_touch of I7712: signal is true;
	signal I7716: std_logic; attribute dont_touch of I7716: signal is true;
	signal I7723: std_logic; attribute dont_touch of I7723: signal is true;
	signal I7728: std_logic; attribute dont_touch of I7728: signal is true;
	signal I7731: std_logic; attribute dont_touch of I7731: signal is true;
	signal I7734: std_logic; attribute dont_touch of I7734: signal is true;
	signal I7738: std_logic; attribute dont_touch of I7738: signal is true;
	signal I7746: std_logic; attribute dont_touch of I7746: signal is true;
	signal I7749: std_logic; attribute dont_touch of I7749: signal is true;
	signal I7752: std_logic; attribute dont_touch of I7752: signal is true;
	signal I7755: std_logic; attribute dont_touch of I7755: signal is true;
	signal I7758: std_logic; attribute dont_touch of I7758: signal is true;
	signal I7762: std_logic; attribute dont_touch of I7762: signal is true;
	signal I7765: std_logic; attribute dont_touch of I7765: signal is true;
	signal I7769: std_logic; attribute dont_touch of I7769: signal is true;
	signal I7775: std_logic; attribute dont_touch of I7775: signal is true;
	signal I7778: std_logic; attribute dont_touch of I7778: signal is true;
	signal I7781: std_logic; attribute dont_touch of I7781: signal is true;
	signal I7785: std_logic; attribute dont_touch of I7785: signal is true;
	signal I7788: std_logic; attribute dont_touch of I7788: signal is true;
	signal I7792: std_logic; attribute dont_touch of I7792: signal is true;
	signal I7797: std_logic; attribute dont_touch of I7797: signal is true;
	signal I7800: std_logic; attribute dont_touch of I7800: signal is true;
	signal I7804: std_logic; attribute dont_touch of I7804: signal is true;
	signal I7807: std_logic; attribute dont_touch of I7807: signal is true;
	signal I7811: std_logic; attribute dont_touch of I7811: signal is true;
	signal I7814: std_logic; attribute dont_touch of I7814: signal is true;
	signal I7832: std_logic; attribute dont_touch of I7832: signal is true;
	signal I7838: std_logic; attribute dont_touch of I7838: signal is true;
	signal I7844: std_logic; attribute dont_touch of I7844: signal is true;
	signal I7847: std_logic; attribute dont_touch of I7847: signal is true;
	signal I7850: std_logic; attribute dont_touch of I7850: signal is true;
	signal I7856: std_logic; attribute dont_touch of I7856: signal is true;
	signal I7859: std_logic; attribute dont_touch of I7859: signal is true;
	signal I7864: std_logic; attribute dont_touch of I7864: signal is true;
	signal I7867: std_logic; attribute dont_touch of I7867: signal is true;
	signal I7870: std_logic; attribute dont_touch of I7870: signal is true;
	signal I7875: std_logic; attribute dont_touch of I7875: signal is true;
	signal I7878: std_logic; attribute dont_touch of I7878: signal is true;
	signal I7882: std_logic; attribute dont_touch of I7882: signal is true;
	signal I7885: std_logic; attribute dont_touch of I7885: signal is true;
	signal I7888: std_logic; attribute dont_touch of I7888: signal is true;
	signal I7891: std_logic; attribute dont_touch of I7891: signal is true;
	signal I7892: std_logic; attribute dont_touch of I7892: signal is true;
	signal I7893: std_logic; attribute dont_touch of I7893: signal is true;
	signal I7899: std_logic; attribute dont_touch of I7899: signal is true;
	signal I7902: std_logic; attribute dont_touch of I7902: signal is true;
	signal I7905: std_logic; attribute dont_touch of I7905: signal is true;
	signal I7908: std_logic; attribute dont_touch of I7908: signal is true;
	signal I7911: std_logic; attribute dont_touch of I7911: signal is true;
	signal I7919: std_logic; attribute dont_touch of I7919: signal is true;
	signal I7922: std_logic; attribute dont_touch of I7922: signal is true;
	signal I7925: std_logic; attribute dont_touch of I7925: signal is true;
	signal I7928: std_logic; attribute dont_touch of I7928: signal is true;
	signal I7931: std_logic; attribute dont_touch of I7931: signal is true;
	signal I7937: std_logic; attribute dont_touch of I7937: signal is true;
	signal I7938: std_logic; attribute dont_touch of I7938: signal is true;
	signal I7939: std_logic; attribute dont_touch of I7939: signal is true;
	signal I7944: std_logic; attribute dont_touch of I7944: signal is true;
	signal I7947: std_logic; attribute dont_touch of I7947: signal is true;
	signal I7950: std_logic; attribute dont_touch of I7950: signal is true;
	signal I7953: std_logic; attribute dont_touch of I7953: signal is true;
	signal I7956: std_logic; attribute dont_touch of I7956: signal is true;
	signal I7959: std_logic; attribute dont_touch of I7959: signal is true;
	signal I7964: std_logic; attribute dont_touch of I7964: signal is true;
	signal I7967: std_logic; attribute dont_touch of I7967: signal is true;
	signal I7970: std_logic; attribute dont_touch of I7970: signal is true;
	signal I7973: std_logic; attribute dont_touch of I7973: signal is true;
	signal I7978: std_logic; attribute dont_touch of I7978: signal is true;
	signal I7981: std_logic; attribute dont_touch of I7981: signal is true;
	signal I7987: std_logic; attribute dont_touch of I7987: signal is true;
	signal I7994: std_logic; attribute dont_touch of I7994: signal is true;
	signal I7995: std_logic; attribute dont_touch of I7995: signal is true;
	signal I8000: std_logic; attribute dont_touch of I8000: signal is true;
	signal I8001: std_logic; attribute dont_touch of I8001: signal is true;
	signal I8005: std_logic; attribute dont_touch of I8005: signal is true;
	signal I8006: std_logic; attribute dont_touch of I8006: signal is true;
	signal I8011: std_logic; attribute dont_touch of I8011: signal is true;
	signal I8014: std_logic; attribute dont_touch of I8014: signal is true;
	signal I8015: std_logic; attribute dont_touch of I8015: signal is true;
	signal I8019: std_logic; attribute dont_touch of I8019: signal is true;
	signal I8020: std_logic; attribute dont_touch of I8020: signal is true;
	signal I8024: std_logic; attribute dont_touch of I8024: signal is true;
	signal I8028: std_logic; attribute dont_touch of I8028: signal is true;
	signal I8029: std_logic; attribute dont_touch of I8029: signal is true;
	signal I8033: std_logic; attribute dont_touch of I8033: signal is true;
	signal I8034: std_logic; attribute dont_touch of I8034: signal is true;
	signal I8040: std_logic; attribute dont_touch of I8040: signal is true;
	signal I8041: std_logic; attribute dont_touch of I8041: signal is true;
	signal I8045: std_logic; attribute dont_touch of I8045: signal is true;
	signal I8046: std_logic; attribute dont_touch of I8046: signal is true;
	signal I8052: std_logic; attribute dont_touch of I8052: signal is true;
	signal I8053: std_logic; attribute dont_touch of I8053: signal is true;
	signal I8057: std_logic; attribute dont_touch of I8057: signal is true;
	signal I8058: std_logic; attribute dont_touch of I8058: signal is true;
	signal I8063: std_logic; attribute dont_touch of I8063: signal is true;
	signal I8064: std_logic; attribute dont_touch of I8064: signal is true;
	signal I8071: std_logic; attribute dont_touch of I8071: signal is true;
	signal I8072: std_logic; attribute dont_touch of I8072: signal is true;
	signal I8078: std_logic; attribute dont_touch of I8078: signal is true;
	signal I8079: std_logic; attribute dont_touch of I8079: signal is true;
	signal I8084: std_logic; attribute dont_touch of I8084: signal is true;
	signal I8089: std_logic; attribute dont_touch of I8089: signal is true;
	signal I8090: std_logic; attribute dont_touch of I8090: signal is true;
	signal I8094: std_logic; attribute dont_touch of I8094: signal is true;
	signal I8097: std_logic; attribute dont_touch of I8097: signal is true;
	signal I8101: std_logic; attribute dont_touch of I8101: signal is true;
	signal I8105: std_logic; attribute dont_touch of I8105: signal is true;
	signal I8108: std_logic; attribute dont_touch of I8108: signal is true;
	signal I8109: std_logic; attribute dont_touch of I8109: signal is true;
	signal I8114: std_logic; attribute dont_touch of I8114: signal is true;
	signal I8115: std_logic; attribute dont_touch of I8115: signal is true;
	signal I8119: std_logic; attribute dont_touch of I8119: signal is true;
	signal I8120: std_logic; attribute dont_touch of I8120: signal is true;
	signal I8121: std_logic; attribute dont_touch of I8121: signal is true;
	signal I8127: std_logic; attribute dont_touch of I8127: signal is true;
	signal I8132: std_logic; attribute dont_touch of I8132: signal is true;
	signal I8133: std_logic; attribute dont_touch of I8133: signal is true;
	signal I8134: std_logic; attribute dont_touch of I8134: signal is true;
	signal I8140: std_logic; attribute dont_touch of I8140: signal is true;
	signal I8143: std_logic; attribute dont_touch of I8143: signal is true;
	signal I8150: std_logic; attribute dont_touch of I8150: signal is true;
	signal I8151: std_logic; attribute dont_touch of I8151: signal is true;
	signal I8152: std_logic; attribute dont_touch of I8152: signal is true;
	signal I8157: std_logic; attribute dont_touch of I8157: signal is true;
	signal I8161: std_logic; attribute dont_touch of I8161: signal is true;
	signal I8164: std_logic; attribute dont_touch of I8164: signal is true;
	signal I8165: std_logic; attribute dont_touch of I8165: signal is true;
	signal I8166: std_logic; attribute dont_touch of I8166: signal is true;
	signal I8172: std_logic; attribute dont_touch of I8172: signal is true;
	signal I8177: std_logic; attribute dont_touch of I8177: signal is true;
	signal I8180: std_logic; attribute dont_touch of I8180: signal is true;
	signal I8186: std_logic; attribute dont_touch of I8186: signal is true;
	signal I8190: std_logic; attribute dont_touch of I8190: signal is true;
	signal I8193: std_logic; attribute dont_touch of I8193: signal is true;
	signal I8196: std_logic; attribute dont_touch of I8196: signal is true;
	signal I8202: std_logic; attribute dont_touch of I8202: signal is true;
	signal I8205: std_logic; attribute dont_touch of I8205: signal is true;
	signal I8209: std_logic; attribute dont_touch of I8209: signal is true;
	signal I8215: std_logic; attribute dont_touch of I8215: signal is true;
	signal I8218: std_logic; attribute dont_touch of I8218: signal is true;
	signal I8224: std_logic; attribute dont_touch of I8224: signal is true;
	signal I8225: std_logic; attribute dont_touch of I8225: signal is true;
	signal I8233: std_logic; attribute dont_touch of I8233: signal is true;
	signal I8237: std_logic; attribute dont_touch of I8237: signal is true;
	signal I8240: std_logic; attribute dont_touch of I8240: signal is true;
	signal I8243: std_logic; attribute dont_touch of I8243: signal is true;
	signal I8244: std_logic; attribute dont_touch of I8244: signal is true;
	signal I8245: std_logic; attribute dont_touch of I8245: signal is true;
	signal I8253: std_logic; attribute dont_touch of I8253: signal is true;
	signal I8254: std_logic; attribute dont_touch of I8254: signal is true;
	signal I8255: std_logic; attribute dont_touch of I8255: signal is true;
	signal I8261: std_logic; attribute dont_touch of I8261: signal is true;
	signal I8264: std_logic; attribute dont_touch of I8264: signal is true;
	signal I8268: std_logic; attribute dont_touch of I8268: signal is true;
	signal I8273: std_logic; attribute dont_touch of I8273: signal is true;
	signal I8277: std_logic; attribute dont_touch of I8277: signal is true;
	signal I8282: std_logic; attribute dont_touch of I8282: signal is true;
	signal I8288: std_logic; attribute dont_touch of I8288: signal is true;
	signal I8291: std_logic; attribute dont_touch of I8291: signal is true;
	signal I8296: std_logic; attribute dont_touch of I8296: signal is true;
	signal I8299: std_logic; attribute dont_touch of I8299: signal is true;
	signal I8308: std_logic; attribute dont_touch of I8308: signal is true;
	signal I8315: std_logic; attribute dont_touch of I8315: signal is true;
	signal I8326: std_logic; attribute dont_touch of I8326: signal is true;
	signal I8327: std_logic; attribute dont_touch of I8327: signal is true;
	signal I8328: std_logic; attribute dont_touch of I8328: signal is true;
	signal I8333: std_logic; attribute dont_touch of I8333: signal is true;
	signal I8338: std_logic; attribute dont_touch of I8338: signal is true;
	signal I8339: std_logic; attribute dont_touch of I8339: signal is true;
	signal I8340: std_logic; attribute dont_touch of I8340: signal is true;
	signal I8351: std_logic; attribute dont_touch of I8351: signal is true;
	signal I8354: std_logic; attribute dont_touch of I8354: signal is true;
	signal I8357: std_logic; attribute dont_touch of I8357: signal is true;
	signal I8360: std_logic; attribute dont_touch of I8360: signal is true;
	signal I8363: std_logic; attribute dont_touch of I8363: signal is true;
	signal I8373: std_logic; attribute dont_touch of I8373: signal is true;
	signal I8392: std_logic; attribute dont_touch of I8392: signal is true;
	signal I8393: std_logic; attribute dont_touch of I8393: signal is true;
	signal I8394: std_logic; attribute dont_touch of I8394: signal is true;
	signal I8400: std_logic; attribute dont_touch of I8400: signal is true;
	signal I8401: std_logic; attribute dont_touch of I8401: signal is true;
	signal I8412: std_logic; attribute dont_touch of I8412: signal is true;
	signal I8413: std_logic; attribute dont_touch of I8413: signal is true;
	signal I8417: std_logic; attribute dont_touch of I8417: signal is true;
	signal I8418: std_logic; attribute dont_touch of I8418: signal is true;
	signal I8428: std_logic; attribute dont_touch of I8428: signal is true;
	signal I8431: std_logic; attribute dont_touch of I8431: signal is true;
	signal I8432: std_logic; attribute dont_touch of I8432: signal is true;
	signal I8436: std_logic; attribute dont_touch of I8436: signal is true;
	signal I8437: std_logic; attribute dont_touch of I8437: signal is true;
	signal I8446: std_logic; attribute dont_touch of I8446: signal is true;
	signal I8449: std_logic; attribute dont_touch of I8449: signal is true;
	signal I8452: std_logic; attribute dont_touch of I8452: signal is true;
	signal I8455: std_logic; attribute dont_touch of I8455: signal is true;
	signal I8456: std_logic; attribute dont_touch of I8456: signal is true;
	signal I8460: std_logic; attribute dont_touch of I8460: signal is true;
	signal I8461: std_logic; attribute dont_touch of I8461: signal is true;
	signal I8470: std_logic; attribute dont_touch of I8470: signal is true;
	signal I8471: std_logic; attribute dont_touch of I8471: signal is true;
	signal I8472: std_logic; attribute dont_touch of I8472: signal is true;
	signal I8477: std_logic; attribute dont_touch of I8477: signal is true;
	signal I8480: std_logic; attribute dont_touch of I8480: signal is true;
	signal I8483: std_logic; attribute dont_touch of I8483: signal is true;
	signal I8486: std_logic; attribute dont_touch of I8486: signal is true;
	signal I8490: std_logic; attribute dont_touch of I8490: signal is true;
	signal I8491: std_logic; attribute dont_touch of I8491: signal is true;
	signal I8495: std_logic; attribute dont_touch of I8495: signal is true;
	signal I8496: std_logic; attribute dont_touch of I8496: signal is true;
	signal I8502: std_logic; attribute dont_touch of I8502: signal is true;
	signal I8503: std_logic; attribute dont_touch of I8503: signal is true;
	signal I8504: std_logic; attribute dont_touch of I8504: signal is true;
	signal I8510: std_logic; attribute dont_touch of I8510: signal is true;
	signal I8511: std_logic; attribute dont_touch of I8511: signal is true;
	signal I8512: std_logic; attribute dont_touch of I8512: signal is true;
	signal I8517: std_logic; attribute dont_touch of I8517: signal is true;
	signal I8520: std_logic; attribute dont_touch of I8520: signal is true;
	signal I8523: std_logic; attribute dont_touch of I8523: signal is true;
	signal I8524: std_logic; attribute dont_touch of I8524: signal is true;
	signal I8528: std_logic; attribute dont_touch of I8528: signal is true;
	signal I8529: std_logic; attribute dont_touch of I8529: signal is true;
	signal I8536: std_logic; attribute dont_touch of I8536: signal is true;
	signal I8537: std_logic; attribute dont_touch of I8537: signal is true;
	signal I8538: std_logic; attribute dont_touch of I8538: signal is true;
	signal I8543: std_logic; attribute dont_touch of I8543: signal is true;
	signal I8546: std_logic; attribute dont_touch of I8546: signal is true;
	signal I8547: std_logic; attribute dont_touch of I8547: signal is true;
	signal I8551: std_logic; attribute dont_touch of I8551: signal is true;
	signal I8552: std_logic; attribute dont_touch of I8552: signal is true;
	signal I8558: std_logic; attribute dont_touch of I8558: signal is true;
	signal I8559: std_logic; attribute dont_touch of I8559: signal is true;
	signal I8560: std_logic; attribute dont_touch of I8560: signal is true;
	signal I8565: std_logic; attribute dont_touch of I8565: signal is true;
	signal I8568: std_logic; attribute dont_touch of I8568: signal is true;
	signal I8569: std_logic; attribute dont_touch of I8569: signal is true;
	signal I8573: std_logic; attribute dont_touch of I8573: signal is true;
	signal I8574: std_logic; attribute dont_touch of I8574: signal is true;
	signal I8581: std_logic; attribute dont_touch of I8581: signal is true;
	signal I8582: std_logic; attribute dont_touch of I8582: signal is true;
	signal I8583: std_logic; attribute dont_touch of I8583: signal is true;
	signal I8588: std_logic; attribute dont_touch of I8588: signal is true;
	signal I8589: std_logic; attribute dont_touch of I8589: signal is true;
	signal I8593: std_logic; attribute dont_touch of I8593: signal is true;
	signal I8594: std_logic; attribute dont_touch of I8594: signal is true;
	signal I8605: std_logic; attribute dont_touch of I8605: signal is true;
	signal I8606: std_logic; attribute dont_touch of I8606: signal is true;
	signal I8607: std_logic; attribute dont_touch of I8607: signal is true;
	signal I8612: std_logic; attribute dont_touch of I8612: signal is true;
	signal I8613: std_logic; attribute dont_touch of I8613: signal is true;
	signal I8617: std_logic; attribute dont_touch of I8617: signal is true;
	signal I8618: std_logic; attribute dont_touch of I8618: signal is true;
	signal I8635: std_logic; attribute dont_touch of I8635: signal is true;
	signal I8636: std_logic; attribute dont_touch of I8636: signal is true;
	signal I8637: std_logic; attribute dont_touch of I8637: signal is true;
	signal I8642: std_logic; attribute dont_touch of I8642: signal is true;
	signal I8643: std_logic; attribute dont_touch of I8643: signal is true;
	signal I8658: std_logic; attribute dont_touch of I8658: signal is true;
	signal I8659: std_logic; attribute dont_touch of I8659: signal is true;
	signal I8660: std_logic; attribute dont_touch of I8660: signal is true;
	signal I8665: std_logic; attribute dont_touch of I8665: signal is true;
	signal I8678: std_logic; attribute dont_touch of I8678: signal is true;
	signal I8679: std_logic; attribute dont_touch of I8679: signal is true;
	signal I8680: std_logic; attribute dont_touch of I8680: signal is true;
	signal I8706: std_logic; attribute dont_touch of I8706: signal is true;
	signal I8709: std_logic; attribute dont_touch of I8709: signal is true;
	signal I8712: std_logic; attribute dont_touch of I8712: signal is true;
	signal I8715: std_logic; attribute dont_touch of I8715: signal is true;
	signal I8718: std_logic; attribute dont_touch of I8718: signal is true;
	signal I8721: std_logic; attribute dont_touch of I8721: signal is true;
	signal I8724: std_logic; attribute dont_touch of I8724: signal is true;
	signal I8727: std_logic; attribute dont_touch of I8727: signal is true;
	signal I8730: std_logic; attribute dont_touch of I8730: signal is true;
	signal I8733: std_logic; attribute dont_touch of I8733: signal is true;
	signal I8736: std_logic; attribute dont_touch of I8736: signal is true;
	signal I8739: std_logic; attribute dont_touch of I8739: signal is true;
	signal I8742: std_logic; attribute dont_touch of I8742: signal is true;
	signal I8745: std_logic; attribute dont_touch of I8745: signal is true;
	signal I8748: std_logic; attribute dont_touch of I8748: signal is true;
	signal I8751: std_logic; attribute dont_touch of I8751: signal is true;
	signal I8754: std_logic; attribute dont_touch of I8754: signal is true;
	signal I8757: std_logic; attribute dont_touch of I8757: signal is true;
	signal I8760: std_logic; attribute dont_touch of I8760: signal is true;
	signal I8763: std_logic; attribute dont_touch of I8763: signal is true;
	signal I8766: std_logic; attribute dont_touch of I8766: signal is true;
	signal I8769: std_logic; attribute dont_touch of I8769: signal is true;
	signal I8772: std_logic; attribute dont_touch of I8772: signal is true;
	signal I8775: std_logic; attribute dont_touch of I8775: signal is true;
	signal I8778: std_logic; attribute dont_touch of I8778: signal is true;
	signal I8781: std_logic; attribute dont_touch of I8781: signal is true;
	signal I8784: std_logic; attribute dont_touch of I8784: signal is true;
	signal I8787: std_logic; attribute dont_touch of I8787: signal is true;
	signal I8790: std_logic; attribute dont_touch of I8790: signal is true;
	signal I8793: std_logic; attribute dont_touch of I8793: signal is true;
	signal I8796: std_logic; attribute dont_touch of I8796: signal is true;
	signal I8799: std_logic; attribute dont_touch of I8799: signal is true;
	signal I8802: std_logic; attribute dont_touch of I8802: signal is true;
	signal I8805: std_logic; attribute dont_touch of I8805: signal is true;
	signal I8808: std_logic; attribute dont_touch of I8808: signal is true;
	signal I8811: std_logic; attribute dont_touch of I8811: signal is true;
	signal I8814: std_logic; attribute dont_touch of I8814: signal is true;
	signal I8817: std_logic; attribute dont_touch of I8817: signal is true;
	signal I8820: std_logic; attribute dont_touch of I8820: signal is true;
	signal I8823: std_logic; attribute dont_touch of I8823: signal is true;
	signal I8826: std_logic; attribute dont_touch of I8826: signal is true;
	signal I8829: std_logic; attribute dont_touch of I8829: signal is true;
	signal I8832: std_logic; attribute dont_touch of I8832: signal is true;
	signal I8835: std_logic; attribute dont_touch of I8835: signal is true;
	signal I8838: std_logic; attribute dont_touch of I8838: signal is true;
	signal I8841: std_logic; attribute dont_touch of I8841: signal is true;
	signal I8844: std_logic; attribute dont_touch of I8844: signal is true;
	signal I8847: std_logic; attribute dont_touch of I8847: signal is true;
	signal I8850: std_logic; attribute dont_touch of I8850: signal is true;
	signal I8853: std_logic; attribute dont_touch of I8853: signal is true;
	signal I8856: std_logic; attribute dont_touch of I8856: signal is true;
	signal I8859: std_logic; attribute dont_touch of I8859: signal is true;
	signal I8862: std_logic; attribute dont_touch of I8862: signal is true;
	signal I8865: std_logic; attribute dont_touch of I8865: signal is true;
	signal I8868: std_logic; attribute dont_touch of I8868: signal is true;
	signal I8871: std_logic; attribute dont_touch of I8871: signal is true;
	signal I8874: std_logic; attribute dont_touch of I8874: signal is true;
	signal I8877: std_logic; attribute dont_touch of I8877: signal is true;
	signal I8880: std_logic; attribute dont_touch of I8880: signal is true;
	signal I8883: std_logic; attribute dont_touch of I8883: signal is true;
	signal I8886: std_logic; attribute dont_touch of I8886: signal is true;
	signal I8889: std_logic; attribute dont_touch of I8889: signal is true;
	signal I8892: std_logic; attribute dont_touch of I8892: signal is true;
	signal I8895: std_logic; attribute dont_touch of I8895: signal is true;
	signal I8898: std_logic; attribute dont_touch of I8898: signal is true;
	signal I8901: std_logic; attribute dont_touch of I8901: signal is true;
	signal I8904: std_logic; attribute dont_touch of I8904: signal is true;
	signal I8907: std_logic; attribute dont_touch of I8907: signal is true;
	signal I8910: std_logic; attribute dont_touch of I8910: signal is true;
	signal I8913: std_logic; attribute dont_touch of I8913: signal is true;
	signal I8916: std_logic; attribute dont_touch of I8916: signal is true;
	signal I8919: std_logic; attribute dont_touch of I8919: signal is true;
	signal I8922: std_logic; attribute dont_touch of I8922: signal is true;
	signal I8925: std_logic; attribute dont_touch of I8925: signal is true;
	signal I8928: std_logic; attribute dont_touch of I8928: signal is true;
	signal I8932: std_logic; attribute dont_touch of I8932: signal is true;
	signal I8935: std_logic; attribute dont_touch of I8935: signal is true;
	signal I8938: std_logic; attribute dont_touch of I8938: signal is true;
	signal I8939: std_logic; attribute dont_touch of I8939: signal is true;
	signal I8940: std_logic; attribute dont_touch of I8940: signal is true;
	signal I8945: std_logic; attribute dont_touch of I8945: signal is true;
	signal I8949: std_logic; attribute dont_touch of I8949: signal is true;
	signal I8952: std_logic; attribute dont_touch of I8952: signal is true;
	signal I8955: std_logic; attribute dont_touch of I8955: signal is true;
	signal I8956: std_logic; attribute dont_touch of I8956: signal is true;
	signal I8957: std_logic; attribute dont_touch of I8957: signal is true;
	signal I8962: std_logic; attribute dont_touch of I8962: signal is true;
	signal I8966: std_logic; attribute dont_touch of I8966: signal is true;
	signal I8971: std_logic; attribute dont_touch of I8971: signal is true;
	signal I8974: std_logic; attribute dont_touch of I8974: signal is true;
	signal I8977: std_logic; attribute dont_touch of I8977: signal is true;
	signal I8980: std_logic; attribute dont_touch of I8980: signal is true;
	signal I8983: std_logic; attribute dont_touch of I8983: signal is true;
	signal I8986: std_logic; attribute dont_touch of I8986: signal is true;
	signal I8989: std_logic; attribute dont_touch of I8989: signal is true;
	signal I8994: std_logic; attribute dont_touch of I8994: signal is true;
	signal I8998: std_logic; attribute dont_touch of I8998: signal is true;
	signal I9001: std_logic; attribute dont_touch of I9001: signal is true;
	signal I9005: std_logic; attribute dont_touch of I9005: signal is true;
	signal I9009: std_logic; attribute dont_touch of I9009: signal is true;
	signal I9014: std_logic; attribute dont_touch of I9014: signal is true;
	signal I9018: std_logic; attribute dont_touch of I9018: signal is true;
	signal I9021: std_logic; attribute dont_touch of I9021: signal is true;
	signal I9025: std_logic; attribute dont_touch of I9025: signal is true;
	signal I9029: std_logic; attribute dont_touch of I9029: signal is true;
	signal I9034: std_logic; attribute dont_touch of I9034: signal is true;
	signal I9038: std_logic; attribute dont_touch of I9038: signal is true;
	signal I9041: std_logic; attribute dont_touch of I9041: signal is true;
	signal I9044: std_logic; attribute dont_touch of I9044: signal is true;
	signal I9047: std_logic; attribute dont_touch of I9047: signal is true;
	signal I9050: std_logic; attribute dont_touch of I9050: signal is true;
	signal I9053: std_logic; attribute dont_touch of I9053: signal is true;
	signal I9057: std_logic; attribute dont_touch of I9057: signal is true;
	signal I9058: std_logic; attribute dont_touch of I9058: signal is true;
	signal I9059: std_logic; attribute dont_touch of I9059: signal is true;
	signal I9064: std_logic; attribute dont_touch of I9064: signal is true;
	signal I9069: std_logic; attribute dont_touch of I9069: signal is true;
	signal I9070: std_logic; attribute dont_touch of I9070: signal is true;
	signal I9071: std_logic; attribute dont_touch of I9071: signal is true;
	signal I9076: std_logic; attribute dont_touch of I9076: signal is true;
	signal I9081: std_logic; attribute dont_touch of I9081: signal is true;
	signal I9084: std_logic; attribute dont_touch of I9084: signal is true;
	signal I9089: std_logic; attribute dont_touch of I9089: signal is true;
	signal I9095: std_logic; attribute dont_touch of I9095: signal is true;
	signal I9099: std_logic; attribute dont_touch of I9099: signal is true;
	signal I9103: std_logic; attribute dont_touch of I9103: signal is true;
	signal I9107: std_logic; attribute dont_touch of I9107: signal is true;
	signal I9111: std_logic; attribute dont_touch of I9111: signal is true;
	signal I9116: std_logic; attribute dont_touch of I9116: signal is true;
	signal I9123: std_logic; attribute dont_touch of I9123: signal is true;
	signal I9126: std_logic; attribute dont_touch of I9126: signal is true;
	signal I9129: std_logic; attribute dont_touch of I9129: signal is true;
	signal I9132: std_logic; attribute dont_touch of I9132: signal is true;
	signal I9136: std_logic; attribute dont_touch of I9136: signal is true;
	signal I9139: std_logic; attribute dont_touch of I9139: signal is true;
	signal I9142: std_logic; attribute dont_touch of I9142: signal is true;
	signal I9145: std_logic; attribute dont_touch of I9145: signal is true;
	signal I9148: std_logic; attribute dont_touch of I9148: signal is true;
	signal I9151: std_logic; attribute dont_touch of I9151: signal is true;
	signal I9152: std_logic; attribute dont_touch of I9152: signal is true;
	signal I9153: std_logic; attribute dont_touch of I9153: signal is true;
	signal I9158: std_logic; attribute dont_touch of I9158: signal is true;
	signal I9162: std_logic; attribute dont_touch of I9162: signal is true;
	signal I9166: std_logic; attribute dont_touch of I9166: signal is true;
	signal I9169: std_logic; attribute dont_touch of I9169: signal is true;
	signal I9170: std_logic; attribute dont_touch of I9170: signal is true;
	signal I9171: std_logic; attribute dont_touch of I9171: signal is true;
	signal I9177: std_logic; attribute dont_touch of I9177: signal is true;
	signal I9181: std_logic; attribute dont_touch of I9181: signal is true;
	signal I9182: std_logic; attribute dont_touch of I9182: signal is true;
	signal I9183: std_logic; attribute dont_touch of I9183: signal is true;
	signal I9194: std_logic; attribute dont_touch of I9194: signal is true;
	signal I9195: std_logic; attribute dont_touch of I9195: signal is true;
	signal I9196: std_logic; attribute dont_touch of I9196: signal is true;
	signal I9202: std_logic; attribute dont_touch of I9202: signal is true;
	signal I9209: std_logic; attribute dont_touch of I9209: signal is true;
	signal I9217: std_logic; attribute dont_touch of I9217: signal is true;
	signal I9222: std_logic; attribute dont_touch of I9222: signal is true;
	signal I9233: std_logic; attribute dont_touch of I9233: signal is true;
	signal I9234: std_logic; attribute dont_touch of I9234: signal is true;
	signal I9235: std_logic; attribute dont_touch of I9235: signal is true;
	signal I9241: std_logic; attribute dont_touch of I9241: signal is true;
	signal I9242: std_logic; attribute dont_touch of I9242: signal is true;
	signal I9243: std_logic; attribute dont_touch of I9243: signal is true;
	signal I9250: std_logic; attribute dont_touch of I9250: signal is true;
	signal I9258: std_logic; attribute dont_touch of I9258: signal is true;
	signal I9261: std_logic; attribute dont_touch of I9261: signal is true;
	signal I9271: std_logic; attribute dont_touch of I9271: signal is true;
	signal I9276: std_logic; attribute dont_touch of I9276: signal is true;
	signal I9277: std_logic; attribute dont_touch of I9277: signal is true;
	signal I9278: std_logic; attribute dont_touch of I9278: signal is true;
	signal I9301: std_logic; attribute dont_touch of I9301: signal is true;
	signal I9310: std_logic; attribute dont_touch of I9310: signal is true;
	signal I9325: std_logic; attribute dont_touch of I9325: signal is true;
	signal I9330: std_logic; attribute dont_touch of I9330: signal is true;
	signal I9333: std_logic; attribute dont_touch of I9333: signal is true;
	signal I9336: std_logic; attribute dont_touch of I9336: signal is true;
	signal I9341: std_logic; attribute dont_touch of I9341: signal is true;
	signal I9344: std_logic; attribute dont_touch of I9344: signal is true;
	signal I9347: std_logic; attribute dont_touch of I9347: signal is true;
	signal I9350: std_logic; attribute dont_touch of I9350: signal is true;
	signal I9360: std_logic; attribute dont_touch of I9360: signal is true;
	signal I9363: std_logic; attribute dont_touch of I9363: signal is true;
	signal I9366: std_logic; attribute dont_touch of I9366: signal is true;
	signal I9369: std_logic; attribute dont_touch of I9369: signal is true;
	signal I9372: std_logic; attribute dont_touch of I9372: signal is true;
	signal I9381: std_logic; attribute dont_touch of I9381: signal is true;
	signal I9382: std_logic; attribute dont_touch of I9382: signal is true;
	signal I9383: std_logic; attribute dont_touch of I9383: signal is true;
	signal I9393: std_logic; attribute dont_touch of I9393: signal is true;
	signal I9396: std_logic; attribute dont_touch of I9396: signal is true;
	signal I9407: std_logic; attribute dont_touch of I9407: signal is true;
	signal I9416: std_logic; attribute dont_touch of I9416: signal is true;
	signal I9419: std_logic; attribute dont_touch of I9419: signal is true;
	signal I9422: std_logic; attribute dont_touch of I9422: signal is true;
	signal I9425: std_logic; attribute dont_touch of I9425: signal is true;
	signal I9440: std_logic; attribute dont_touch of I9440: signal is true;
	signal I9443: std_logic; attribute dont_touch of I9443: signal is true;
	signal I9446: std_logic; attribute dont_touch of I9446: signal is true;
	signal I9457: std_logic; attribute dont_touch of I9457: signal is true;
	signal I9460: std_logic; attribute dont_touch of I9460: signal is true;
	signal I9463: std_logic; attribute dont_touch of I9463: signal is true;
	signal I9466: std_logic; attribute dont_touch of I9466: signal is true;
	signal I9475: std_logic; attribute dont_touch of I9475: signal is true;
	signal I9476: std_logic; attribute dont_touch of I9476: signal is true;
	signal I9477: std_logic; attribute dont_touch of I9477: signal is true;
	signal I9484: std_logic; attribute dont_touch of I9484: signal is true;
	signal I9493: std_logic; attribute dont_touch of I9493: signal is true;
	signal I9496: std_logic; attribute dont_touch of I9496: signal is true;
	signal I9499: std_logic; attribute dont_touch of I9499: signal is true;
	signal I9502: std_logic; attribute dont_touch of I9502: signal is true;
	signal I9505: std_logic; attribute dont_touch of I9505: signal is true;
	signal I9512: std_logic; attribute dont_touch of I9512: signal is true;
	signal I9515: std_logic; attribute dont_touch of I9515: signal is true;
	signal I9520: std_logic; attribute dont_touch of I9520: signal is true;
	signal I9525: std_logic; attribute dont_touch of I9525: signal is true;
	signal I9528: std_logic; attribute dont_touch of I9528: signal is true;
	signal I9531: std_logic; attribute dont_touch of I9531: signal is true;
	signal I9534: std_logic; attribute dont_touch of I9534: signal is true;
	signal I9535: std_logic; attribute dont_touch of I9535: signal is true;
	signal I9539: std_logic; attribute dont_touch of I9539: signal is true;
	signal I9543: std_logic; attribute dont_touch of I9543: signal is true;
	signal I9547: std_logic; attribute dont_touch of I9547: signal is true;
	signal I9548: std_logic; attribute dont_touch of I9548: signal is true;
	signal I9549: std_logic; attribute dont_touch of I9549: signal is true;
	signal I9555: std_logic; attribute dont_touch of I9555: signal is true;
	signal I9558: std_logic; attribute dont_touch of I9558: signal is true;
	signal I9561: std_logic; attribute dont_touch of I9561: signal is true;
	signal I9564: std_logic; attribute dont_touch of I9564: signal is true;
	signal I9567: std_logic; attribute dont_touch of I9567: signal is true;
	signal I9570: std_logic; attribute dont_touch of I9570: signal is true;
	signal I9573: std_logic; attribute dont_touch of I9573: signal is true;
	signal I9576: std_logic; attribute dont_touch of I9576: signal is true;
	signal I9579: std_logic; attribute dont_touch of I9579: signal is true;
	signal I9582: std_logic; attribute dont_touch of I9582: signal is true;
	signal I9585: std_logic; attribute dont_touch of I9585: signal is true;
	signal I9588: std_logic; attribute dont_touch of I9588: signal is true;
	signal I9591: std_logic; attribute dont_touch of I9591: signal is true;
	signal I9594: std_logic; attribute dont_touch of I9594: signal is true;
	signal I9597: std_logic; attribute dont_touch of I9597: signal is true;
	signal I9600: std_logic; attribute dont_touch of I9600: signal is true;
	signal I9603: std_logic; attribute dont_touch of I9603: signal is true;
	signal I9606: std_logic; attribute dont_touch of I9606: signal is true;
	signal I9609: std_logic; attribute dont_touch of I9609: signal is true;
	signal I9612: std_logic; attribute dont_touch of I9612: signal is true;
	signal I9615: std_logic; attribute dont_touch of I9615: signal is true;
	signal I9618: std_logic; attribute dont_touch of I9618: signal is true;
	signal I9621: std_logic; attribute dont_touch of I9621: signal is true;
	signal I9624: std_logic; attribute dont_touch of I9624: signal is true;
	signal I9627: std_logic; attribute dont_touch of I9627: signal is true;
	signal I9630: std_logic; attribute dont_touch of I9630: signal is true;
	signal I9633: std_logic; attribute dont_touch of I9633: signal is true;
	signal I9636: std_logic; attribute dont_touch of I9636: signal is true;
	signal I9639: std_logic; attribute dont_touch of I9639: signal is true;
	signal I9642: std_logic; attribute dont_touch of I9642: signal is true;
	signal I9645: std_logic; attribute dont_touch of I9645: signal is true;
	signal I9648: std_logic; attribute dont_touch of I9648: signal is true;
	signal I9651: std_logic; attribute dont_touch of I9651: signal is true;
	signal I9654: std_logic; attribute dont_touch of I9654: signal is true;
	signal I9657: std_logic; attribute dont_touch of I9657: signal is true;
	signal I9660: std_logic; attribute dont_touch of I9660: signal is true;
	signal I9663: std_logic; attribute dont_touch of I9663: signal is true;
	signal I9666: std_logic; attribute dont_touch of I9666: signal is true;
	signal I9669: std_logic; attribute dont_touch of I9669: signal is true;
	signal I9672: std_logic; attribute dont_touch of I9672: signal is true;
	signal I9675: std_logic; attribute dont_touch of I9675: signal is true;
	signal I9678: std_logic; attribute dont_touch of I9678: signal is true;
	signal I9681: std_logic; attribute dont_touch of I9681: signal is true;
	signal I9684: std_logic; attribute dont_touch of I9684: signal is true;
	signal I9687: std_logic; attribute dont_touch of I9687: signal is true;
	signal I9691: std_logic; attribute dont_touch of I9691: signal is true;
	signal I9692: std_logic; attribute dont_touch of I9692: signal is true;
	signal I9693: std_logic; attribute dont_touch of I9693: signal is true;
	signal I9745: std_logic; attribute dont_touch of I9745: signal is true;
	signal I9746: std_logic; attribute dont_touch of I9746: signal is true;
	signal I9747: std_logic; attribute dont_touch of I9747: signal is true;
	signal I9752: std_logic; attribute dont_touch of I9752: signal is true;
	signal I9760: std_logic; attribute dont_touch of I9760: signal is true;
	signal I9767: std_logic; attribute dont_touch of I9767: signal is true;
	signal I9768: std_logic; attribute dont_touch of I9768: signal is true;
	signal I9769: std_logic; attribute dont_touch of I9769: signal is true;
	signal I9774: std_logic; attribute dont_touch of I9774: signal is true;
	signal I9782: std_logic; attribute dont_touch of I9782: signal is true;
	signal I9785: std_logic; attribute dont_touch of I9785: signal is true;
	signal I9788: std_logic; attribute dont_touch of I9788: signal is true;
	signal I9791: std_logic; attribute dont_touch of I9791: signal is true;
	signal I9794: std_logic; attribute dont_touch of I9794: signal is true;
	signal I9804: std_logic; attribute dont_touch of I9804: signal is true;
	signal I9819: std_logic; attribute dont_touch of I9819: signal is true;
	signal I9823: std_logic; attribute dont_touch of I9823: signal is true;
	signal I9826: std_logic; attribute dont_touch of I9826: signal is true;
	signal I9827: std_logic; attribute dont_touch of I9827: signal is true;
	signal I9828: std_logic; attribute dont_touch of I9828: signal is true;
	signal I9834: std_logic; attribute dont_touch of I9834: signal is true;
	signal I9837: std_logic; attribute dont_touch of I9837: signal is true;
	signal I9840: std_logic; attribute dont_touch of I9840: signal is true;
	signal I9845: std_logic; attribute dont_touch of I9845: signal is true;
	signal I9850: std_logic; attribute dont_touch of I9850: signal is true;
	signal I9884: std_logic; attribute dont_touch of I9884: signal is true;
	signal I9889: std_logic; attribute dont_touch of I9889: signal is true;
	signal I9892: std_logic; attribute dont_touch of I9892: signal is true;
	signal I9907: std_logic; attribute dont_touch of I9907: signal is true;
	signal I9910: std_logic; attribute dont_touch of I9910: signal is true;
	signal I9918: std_logic; attribute dont_touch of I9918: signal is true;
	signal I9929: std_logic; attribute dont_touch of I9929: signal is true;
	signal I9935: std_logic; attribute dont_touch of I9935: signal is true;
	signal I9938: std_logic; attribute dont_touch of I9938: signal is true;
	signal I9946: std_logic; attribute dont_touch of I9946: signal is true;
	signal I9947: std_logic; attribute dont_touch of I9947: signal is true;
	signal I9948: std_logic; attribute dont_touch of I9948: signal is true;
	signal I9953: std_logic; attribute dont_touch of I9953: signal is true;
	signal I9954: std_logic; attribute dont_touch of I9954: signal is true;
	signal I9955: std_logic; attribute dont_touch of I9955: signal is true;
	signal I9963: std_logic; attribute dont_touch of I9963: signal is true;
	signal I9964: std_logic; attribute dont_touch of I9964: signal is true;
	signal I9965: std_logic; attribute dont_touch of I9965: signal is true;
	signal I9974: std_logic; attribute dont_touch of I9974: signal is true;
	signal I9978: std_logic; attribute dont_touch of I9978: signal is true;
	signal I9979: std_logic; attribute dont_touch of I9979: signal is true;
	signal I9980: std_logic; attribute dont_touch of I9980: signal is true;
	signal I9985: std_logic; attribute dont_touch of I9985: signal is true;
	signal I9986: std_logic; attribute dont_touch of I9986: signal is true;
	signal I9987: std_logic; attribute dont_touch of I9987: signal is true;
	signal I9992: std_logic; attribute dont_touch of I9992: signal is true;
	signal I9993: std_logic; attribute dont_touch of I9993: signal is true;
	signal I9994: std_logic; attribute dont_touch of I9994: signal is true;
	signal I9999: std_logic; attribute dont_touch of I9999: signal is true;
	signal I10000: std_logic; attribute dont_touch of I10000: signal is true;
	signal I10001: std_logic; attribute dont_touch of I10001: signal is true;
	signal I10009: std_logic; attribute dont_touch of I10009: signal is true;
	signal I10010: std_logic; attribute dont_touch of I10010: signal is true;
	signal I10011: std_logic; attribute dont_touch of I10011: signal is true;
	signal I10017: std_logic; attribute dont_touch of I10017: signal is true;
	signal I10018: std_logic; attribute dont_touch of I10018: signal is true;
	signal I10019: std_logic; attribute dont_touch of I10019: signal is true;
	signal I10028: std_logic; attribute dont_touch of I10028: signal is true;
	signal I10032: std_logic; attribute dont_touch of I10032: signal is true;
	signal I10038: std_logic; attribute dont_touch of I10038: signal is true;
	signal I10039: std_logic; attribute dont_touch of I10039: signal is true;
	signal I10040: std_logic; attribute dont_touch of I10040: signal is true;
	signal I10046: std_logic; attribute dont_touch of I10046: signal is true;
	signal I10060: std_logic; attribute dont_touch of I10060: signal is true;
	signal I10061: std_logic; attribute dont_touch of I10061: signal is true;
	signal I10062: std_logic; attribute dont_touch of I10062: signal is true;
	signal I10071: std_logic; attribute dont_touch of I10071: signal is true;
	signal I10072: std_logic; attribute dont_touch of I10072: signal is true;
	signal I10073: std_logic; attribute dont_touch of I10073: signal is true;
	signal I10078: std_logic; attribute dont_touch of I10078: signal is true;
	signal I10079: std_logic; attribute dont_touch of I10079: signal is true;
	signal I10080: std_logic; attribute dont_touch of I10080: signal is true;
	signal I10092: std_logic; attribute dont_touch of I10092: signal is true;
	signal I10093: std_logic; attribute dont_touch of I10093: signal is true;
	signal I10094: std_logic; attribute dont_touch of I10094: signal is true;
	signal I10125: std_logic; attribute dont_touch of I10125: signal is true;
	signal I10128: std_logic; attribute dont_touch of I10128: signal is true;
	signal I10135: std_logic; attribute dont_touch of I10135: signal is true;
	signal I10142: std_logic; attribute dont_touch of I10142: signal is true;
	signal I10143: std_logic; attribute dont_touch of I10143: signal is true;
	signal I10144: std_logic; attribute dont_touch of I10144: signal is true;
	signal I10151: std_logic; attribute dont_touch of I10151: signal is true;
	signal I10154: std_logic; attribute dont_touch of I10154: signal is true;
	signal I10157: std_logic; attribute dont_touch of I10157: signal is true;
	signal I10160: std_logic; attribute dont_touch of I10160: signal is true;
	signal I10166: std_logic; attribute dont_touch of I10166: signal is true;
	signal I10169: std_logic; attribute dont_touch of I10169: signal is true;
	signal I10172: std_logic; attribute dont_touch of I10172: signal is true;
	signal I10177: std_logic; attribute dont_touch of I10177: signal is true;
	signal I10180: std_logic; attribute dont_touch of I10180: signal is true;
	signal I10183: std_logic; attribute dont_touch of I10183: signal is true;
	signal I10186: std_logic; attribute dont_touch of I10186: signal is true;
	signal I10190: std_logic; attribute dont_touch of I10190: signal is true;
	signal I10193: std_logic; attribute dont_touch of I10193: signal is true;
	signal I10196: std_logic; attribute dont_touch of I10196: signal is true;
	signal I10197: std_logic; attribute dont_touch of I10197: signal is true;
	signal I10198: std_logic; attribute dont_touch of I10198: signal is true;
	signal I10204: std_logic; attribute dont_touch of I10204: signal is true;
	signal I10207: std_logic; attribute dont_touch of I10207: signal is true;
	signal I10223: std_logic; attribute dont_touch of I10223: signal is true;
	signal I10224: std_logic; attribute dont_touch of I10224: signal is true;
	signal I10225: std_logic; attribute dont_touch of I10225: signal is true;
	signal I10236: std_logic; attribute dont_touch of I10236: signal is true;
	signal I10243: std_logic; attribute dont_touch of I10243: signal is true;
	signal I10247: std_logic; attribute dont_touch of I10247: signal is true;
	signal I10250: std_logic; attribute dont_touch of I10250: signal is true;
	signal I10253: std_logic; attribute dont_touch of I10253: signal is true;
	signal I10256: std_logic; attribute dont_touch of I10256: signal is true;
	signal I10259: std_logic; attribute dont_touch of I10259: signal is true;
	signal I10262: std_logic; attribute dont_touch of I10262: signal is true;
	signal I10265: std_logic; attribute dont_touch of I10265: signal is true;
	signal I10268: std_logic; attribute dont_touch of I10268: signal is true;
	signal I10271: std_logic; attribute dont_touch of I10271: signal is true;
	signal I10274: std_logic; attribute dont_touch of I10274: signal is true;
	signal I10277: std_logic; attribute dont_touch of I10277: signal is true;
	signal I10280: std_logic; attribute dont_touch of I10280: signal is true;
	signal I10283: std_logic; attribute dont_touch of I10283: signal is true;
	signal I10286: std_logic; attribute dont_touch of I10286: signal is true;
	signal I10289: std_logic; attribute dont_touch of I10289: signal is true;
	signal I10292: std_logic; attribute dont_touch of I10292: signal is true;
	signal I10295: std_logic; attribute dont_touch of I10295: signal is true;
	signal I10298: std_logic; attribute dont_touch of I10298: signal is true;
	signal I10299: std_logic; attribute dont_touch of I10299: signal is true;
	signal I10300: std_logic; attribute dont_touch of I10300: signal is true;
	signal I10305: std_logic; attribute dont_touch of I10305: signal is true;
	signal I10306: std_logic; attribute dont_touch of I10306: signal is true;
	signal I10307: std_logic; attribute dont_touch of I10307: signal is true;
	signal I10313: std_logic; attribute dont_touch of I10313: signal is true;
	signal I10314: std_logic; attribute dont_touch of I10314: signal is true;
	signal I10315: std_logic; attribute dont_touch of I10315: signal is true;
	signal I10320: std_logic; attribute dont_touch of I10320: signal is true;
	signal I10321: std_logic; attribute dont_touch of I10321: signal is true;
	signal I10322: std_logic; attribute dont_touch of I10322: signal is true;
	signal I10327: std_logic; attribute dont_touch of I10327: signal is true;
	signal I10328: std_logic; attribute dont_touch of I10328: signal is true;
	signal I10329: std_logic; attribute dont_touch of I10329: signal is true;
	signal I10334: std_logic; attribute dont_touch of I10334: signal is true;
	signal I10335: std_logic; attribute dont_touch of I10335: signal is true;
	signal I10336: std_logic; attribute dont_touch of I10336: signal is true;
	signal I10343: std_logic; attribute dont_touch of I10343: signal is true;
	signal I10347: std_logic; attribute dont_touch of I10347: signal is true;
	signal I10350: std_logic; attribute dont_touch of I10350: signal is true;
	signal I10353: std_logic; attribute dont_touch of I10353: signal is true;
	signal I10356: std_logic; attribute dont_touch of I10356: signal is true;
	signal I10359: std_logic; attribute dont_touch of I10359: signal is true;
	signal I10360: std_logic; attribute dont_touch of I10360: signal is true;
	signal I10361: std_logic; attribute dont_touch of I10361: signal is true;
	signal I10366: std_logic; attribute dont_touch of I10366: signal is true;
	signal I10369: std_logic; attribute dont_touch of I10369: signal is true;
	signal I10373: std_logic; attribute dont_touch of I10373: signal is true;
	signal I10377: std_logic; attribute dont_touch of I10377: signal is true;
	signal I10380: std_logic; attribute dont_touch of I10380: signal is true;
	signal I10384: std_logic; attribute dont_touch of I10384: signal is true;
	signal I10387: std_logic; attribute dont_touch of I10387: signal is true;
	signal I10390: std_logic; attribute dont_touch of I10390: signal is true;
	signal I10393: std_logic; attribute dont_touch of I10393: signal is true;
	signal I10397: std_logic; attribute dont_touch of I10397: signal is true;
	signal I10400: std_logic; attribute dont_touch of I10400: signal is true;
	signal I10403: std_logic; attribute dont_touch of I10403: signal is true;
	signal I10406: std_logic; attribute dont_touch of I10406: signal is true;
	signal I10409: std_logic; attribute dont_touch of I10409: signal is true;
	signal I10412: std_logic; attribute dont_touch of I10412: signal is true;
	signal I10415: std_logic; attribute dont_touch of I10415: signal is true;
	signal I10418: std_logic; attribute dont_touch of I10418: signal is true;
	signal I10421: std_logic; attribute dont_touch of I10421: signal is true;
	signal I10424: std_logic; attribute dont_touch of I10424: signal is true;
	signal I10427: std_logic; attribute dont_touch of I10427: signal is true;
	signal I10430: std_logic; attribute dont_touch of I10430: signal is true;
	signal I10433: std_logic; attribute dont_touch of I10433: signal is true;
	signal I10436: std_logic; attribute dont_touch of I10436: signal is true;
	signal I10439: std_logic; attribute dont_touch of I10439: signal is true;
	signal I10442: std_logic; attribute dont_touch of I10442: signal is true;
	signal I10445: std_logic; attribute dont_touch of I10445: signal is true;
	signal I10448: std_logic; attribute dont_touch of I10448: signal is true;
	signal I10451: std_logic; attribute dont_touch of I10451: signal is true;
	signal I10454: std_logic; attribute dont_touch of I10454: signal is true;
	signal I10457: std_logic; attribute dont_touch of I10457: signal is true;
	signal I10460: std_logic; attribute dont_touch of I10460: signal is true;
	signal I10463: std_logic; attribute dont_touch of I10463: signal is true;
	signal I10466: std_logic; attribute dont_touch of I10466: signal is true;
	signal I10469: std_logic; attribute dont_touch of I10469: signal is true;
	signal I10472: std_logic; attribute dont_touch of I10472: signal is true;
	signal I10475: std_logic; attribute dont_touch of I10475: signal is true;
	signal I10479: std_logic; attribute dont_touch of I10479: signal is true;
	signal I10482: std_logic; attribute dont_touch of I10482: signal is true;
	signal I10485: std_logic; attribute dont_touch of I10485: signal is true;
	signal I10488: std_logic; attribute dont_touch of I10488: signal is true;
	signal I10491: std_logic; attribute dont_touch of I10491: signal is true;
	signal I10494: std_logic; attribute dont_touch of I10494: signal is true;
	signal I10497: std_logic; attribute dont_touch of I10497: signal is true;
	signal I10500: std_logic; attribute dont_touch of I10500: signal is true;
	signal I10503: std_logic; attribute dont_touch of I10503: signal is true;
	signal I10506: std_logic; attribute dont_touch of I10506: signal is true;
	signal I10509: std_logic; attribute dont_touch of I10509: signal is true;
	signal I10512: std_logic; attribute dont_touch of I10512: signal is true;
	signal I10516: std_logic; attribute dont_touch of I10516: signal is true;
	signal I10519: std_logic; attribute dont_touch of I10519: signal is true;
	signal I10522: std_logic; attribute dont_touch of I10522: signal is true;
	signal I10525: std_logic; attribute dont_touch of I10525: signal is true;
	signal I10528: std_logic; attribute dont_touch of I10528: signal is true;
	signal I10532: std_logic; attribute dont_touch of I10532: signal is true;
	signal I10535: std_logic; attribute dont_touch of I10535: signal is true;
	signal I10538: std_logic; attribute dont_touch of I10538: signal is true;
	signal I10541: std_logic; attribute dont_touch of I10541: signal is true;
	signal I10545: std_logic; attribute dont_touch of I10545: signal is true;
	signal I10548: std_logic; attribute dont_touch of I10548: signal is true;
	signal I10552: std_logic; attribute dont_touch of I10552: signal is true;
	signal I10555: std_logic; attribute dont_touch of I10555: signal is true;
	signal I10558: std_logic; attribute dont_touch of I10558: signal is true;
	signal I10561: std_logic; attribute dont_touch of I10561: signal is true;
	signal I10565: std_logic; attribute dont_touch of I10565: signal is true;
	signal I10569: std_logic; attribute dont_touch of I10569: signal is true;
	signal I10574: std_logic; attribute dont_touch of I10574: signal is true;
	signal I10579: std_logic; attribute dont_touch of I10579: signal is true;
	signal I10582: std_logic; attribute dont_touch of I10582: signal is true;
	signal I10587: std_logic; attribute dont_touch of I10587: signal is true;
	signal I10592: std_logic; attribute dont_touch of I10592: signal is true;
	signal I10597: std_logic; attribute dont_touch of I10597: signal is true;
	signal I10605: std_logic; attribute dont_touch of I10605: signal is true;
	signal I10608: std_logic; attribute dont_touch of I10608: signal is true;
	signal I10614: std_logic; attribute dont_touch of I10614: signal is true;
	signal I10617: std_logic; attribute dont_touch of I10617: signal is true;
	signal I10625: std_logic; attribute dont_touch of I10625: signal is true;
	signal I10626: std_logic; attribute dont_touch of I10626: signal is true;
	signal I10627: std_logic; attribute dont_touch of I10627: signal is true;
	signal I10639: std_logic; attribute dont_touch of I10639: signal is true;
	signal I10643: std_logic; attribute dont_touch of I10643: signal is true;
	signal I10646: std_logic; attribute dont_touch of I10646: signal is true;
	signal I10649: std_logic; attribute dont_touch of I10649: signal is true;
	signal I10675: std_logic; attribute dont_touch of I10675: signal is true;
	signal I10678: std_logic; attribute dont_touch of I10678: signal is true;
	signal I10681: std_logic; attribute dont_touch of I10681: signal is true;
	signal I10684: std_logic; attribute dont_touch of I10684: signal is true;
	signal I10687: std_logic; attribute dont_touch of I10687: signal is true;
	signal I10690: std_logic; attribute dont_touch of I10690: signal is true;
	signal I10694: std_logic; attribute dont_touch of I10694: signal is true;
	signal I10702: std_logic; attribute dont_touch of I10702: signal is true;
	signal I10705: std_logic; attribute dont_touch of I10705: signal is true;
	signal I10708: std_logic; attribute dont_touch of I10708: signal is true;
	signal I10716: std_logic; attribute dont_touch of I10716: signal is true;
	signal I10719: std_logic; attribute dont_touch of I10719: signal is true;
	signal I10739: std_logic; attribute dont_touch of I10739: signal is true;
	signal I10743: std_logic; attribute dont_touch of I10743: signal is true;
	signal I10744: std_logic; attribute dont_touch of I10744: signal is true;
	signal I10745: std_logic; attribute dont_touch of I10745: signal is true;
	signal I10752: std_logic; attribute dont_touch of I10752: signal is true;
	signal I10758: std_logic; attribute dont_touch of I10758: signal is true;
	signal I10761: std_logic; attribute dont_touch of I10761: signal is true;
	signal I10766: std_logic; attribute dont_touch of I10766: signal is true;
	signal I10770: std_logic; attribute dont_touch of I10770: signal is true;
	signal I10773: std_logic; attribute dont_touch of I10773: signal is true;
	signal I10776: std_logic; attribute dont_touch of I10776: signal is true;
	signal I10780: std_logic; attribute dont_touch of I10780: signal is true;
	signal I10783: std_logic; attribute dont_touch of I10783: signal is true;
	signal I10786: std_logic; attribute dont_touch of I10786: signal is true;
	signal I10789: std_logic; attribute dont_touch of I10789: signal is true;
	signal I10790: std_logic; attribute dont_touch of I10790: signal is true;
	signal I10791: std_logic; attribute dont_touch of I10791: signal is true;
	signal I10796: std_logic; attribute dont_touch of I10796: signal is true;
	signal I10801: std_logic; attribute dont_touch of I10801: signal is true;
	signal I10804: std_logic; attribute dont_touch of I10804: signal is true;
	signal I10807: std_logic; attribute dont_touch of I10807: signal is true;
	signal I10810: std_logic; attribute dont_touch of I10810: signal is true;
	signal I10815: std_logic; attribute dont_touch of I10815: signal is true;
	signal I10818: std_logic; attribute dont_touch of I10818: signal is true;
	signal I10819: std_logic; attribute dont_touch of I10819: signal is true;
	signal I10820: std_logic; attribute dont_touch of I10820: signal is true;
	signal I10826: std_logic; attribute dont_touch of I10826: signal is true;
	signal I10829: std_logic; attribute dont_touch of I10829: signal is true;
	signal I10834: std_logic; attribute dont_touch of I10834: signal is true;
	signal I10835: std_logic; attribute dont_touch of I10835: signal is true;
	signal I10836: std_logic; attribute dont_touch of I10836: signal is true;
	signal I10842: std_logic; attribute dont_touch of I10842: signal is true;
	signal I10847: std_logic; attribute dont_touch of I10847: signal is true;
	signal I10848: std_logic; attribute dont_touch of I10848: signal is true;
	signal I10849: std_logic; attribute dont_touch of I10849: signal is true;
	signal I10854: std_logic; attribute dont_touch of I10854: signal is true;
	signal I10855: std_logic; attribute dont_touch of I10855: signal is true;
	signal I10856: std_logic; attribute dont_touch of I10856: signal is true;
	signal I10862: std_logic; attribute dont_touch of I10862: signal is true;
	signal I10866: std_logic; attribute dont_touch of I10866: signal is true;
	signal I10867: std_logic; attribute dont_touch of I10867: signal is true;
	signal I10868: std_logic; attribute dont_touch of I10868: signal is true;
	signal I10873: std_logic; attribute dont_touch of I10873: signal is true;
	signal I10874: std_logic; attribute dont_touch of I10874: signal is true;
	signal I10875: std_logic; attribute dont_touch of I10875: signal is true;
	signal I10882: std_logic; attribute dont_touch of I10882: signal is true;
	signal I10888: std_logic; attribute dont_touch of I10888: signal is true;
	signal I10889: std_logic; attribute dont_touch of I10889: signal is true;
	signal I10890: std_logic; attribute dont_touch of I10890: signal is true;
	signal I10896: std_logic; attribute dont_touch of I10896: signal is true;
	signal I10899: std_logic; attribute dont_touch of I10899: signal is true;
	signal I10900: std_logic; attribute dont_touch of I10900: signal is true;
	signal I10901: std_logic; attribute dont_touch of I10901: signal is true;
	signal I10906: std_logic; attribute dont_touch of I10906: signal is true;
	signal I10907: std_logic; attribute dont_touch of I10907: signal is true;
	signal I10908: std_logic; attribute dont_touch of I10908: signal is true;
	signal I10914: std_logic; attribute dont_touch of I10914: signal is true;
	signal I10919: std_logic; attribute dont_touch of I10919: signal is true;
	signal I10923: std_logic; attribute dont_touch of I10923: signal is true;
	signal I10924: std_logic; attribute dont_touch of I10924: signal is true;
	signal I10925: std_logic; attribute dont_touch of I10925: signal is true;
	signal I10930: std_logic; attribute dont_touch of I10930: signal is true;
	signal I10933: std_logic; attribute dont_touch of I10933: signal is true;
	signal I10937: std_logic; attribute dont_touch of I10937: signal is true;
	signal I10940: std_logic; attribute dont_touch of I10940: signal is true;
	signal I10946: std_logic; attribute dont_touch of I10946: signal is true;
	signal I10949: std_logic; attribute dont_touch of I10949: signal is true;
	signal I10952: std_logic; attribute dont_touch of I10952: signal is true;
	signal I10953: std_logic; attribute dont_touch of I10953: signal is true;
	signal I10954: std_logic; attribute dont_touch of I10954: signal is true;
	signal I10962: std_logic; attribute dont_touch of I10962: signal is true;
	signal I10965: std_logic; attribute dont_touch of I10965: signal is true;
	signal I10969: std_logic; attribute dont_touch of I10969: signal is true;
	signal I10973: std_logic; attribute dont_touch of I10973: signal is true;
	signal I10976: std_logic; attribute dont_touch of I10976: signal is true;
	signal I10980: std_logic; attribute dont_touch of I10980: signal is true;
	signal I10981: std_logic; attribute dont_touch of I10981: signal is true;
	signal I10982: std_logic; attribute dont_touch of I10982: signal is true;
	signal I10987: std_logic; attribute dont_touch of I10987: signal is true;
	signal I10991: std_logic; attribute dont_touch of I10991: signal is true;
	signal I10992: std_logic; attribute dont_touch of I10992: signal is true;
	signal I10993: std_logic; attribute dont_touch of I10993: signal is true;
	signal I10998: std_logic; attribute dont_touch of I10998: signal is true;
	signal I11001: std_logic; attribute dont_touch of I11001: signal is true;
	signal I11004: std_logic; attribute dont_touch of I11004: signal is true;
	signal I11008: std_logic; attribute dont_touch of I11008: signal is true;
	signal I11011: std_logic; attribute dont_touch of I11011: signal is true;
	signal I11014: std_logic; attribute dont_touch of I11014: signal is true;
	signal I11018: std_logic; attribute dont_touch of I11018: signal is true;
	signal I11021: std_logic; attribute dont_touch of I11021: signal is true;
	signal I11025: std_logic; attribute dont_touch of I11025: signal is true;
	signal I11028: std_logic; attribute dont_touch of I11028: signal is true;
	signal I11031: std_logic; attribute dont_touch of I11031: signal is true;
	signal I11034: std_logic; attribute dont_touch of I11034: signal is true;
	signal I11037: std_logic; attribute dont_touch of I11037: signal is true;
	signal I11040: std_logic; attribute dont_touch of I11040: signal is true;
	signal I11043: std_logic; attribute dont_touch of I11043: signal is true;
	signal I11047: std_logic; attribute dont_touch of I11047: signal is true;
	signal I11050: std_logic; attribute dont_touch of I11050: signal is true;
	signal I11055: std_logic; attribute dont_touch of I11055: signal is true;
	signal I11060: std_logic; attribute dont_touch of I11060: signal is true;
	signal I11066: std_logic; attribute dont_touch of I11066: signal is true;
	signal I11069: std_logic; attribute dont_touch of I11069: signal is true;
	signal I11078: std_logic; attribute dont_touch of I11078: signal is true;
	signal I11079: std_logic; attribute dont_touch of I11079: signal is true;
	signal I11080: std_logic; attribute dont_touch of I11080: signal is true;
	signal I11086: std_logic; attribute dont_touch of I11086: signal is true;
	signal I11090: std_logic; attribute dont_touch of I11090: signal is true;
	signal I11094: std_logic; attribute dont_touch of I11094: signal is true;
	signal I11095: std_logic; attribute dont_touch of I11095: signal is true;
	signal I11096: std_logic; attribute dont_touch of I11096: signal is true;
	signal I11101: std_logic; attribute dont_touch of I11101: signal is true;
	signal I11102: std_logic; attribute dont_touch of I11102: signal is true;
	signal I11103: std_logic; attribute dont_touch of I11103: signal is true;
	signal I11108: std_logic; attribute dont_touch of I11108: signal is true;
	signal I11109: std_logic; attribute dont_touch of I11109: signal is true;
	signal I11110: std_logic; attribute dont_touch of I11110: signal is true;
	signal I11115: std_logic; attribute dont_touch of I11115: signal is true;
	signal I11116: std_logic; attribute dont_touch of I11116: signal is true;
	signal I11117: std_logic; attribute dont_touch of I11117: signal is true;
	signal I11122: std_logic; attribute dont_touch of I11122: signal is true;
	signal I11123: std_logic; attribute dont_touch of I11123: signal is true;
	signal I11124: std_logic; attribute dont_touch of I11124: signal is true;
	signal I11129: std_logic; attribute dont_touch of I11129: signal is true;
	signal I11132: std_logic; attribute dont_touch of I11132: signal is true;
	signal I11135: std_logic; attribute dont_touch of I11135: signal is true;
	signal I11136: std_logic; attribute dont_touch of I11136: signal is true;
	signal I11137: std_logic; attribute dont_touch of I11137: signal is true;
	signal I11142: std_logic; attribute dont_touch of I11142: signal is true;
	signal I11143: std_logic; attribute dont_touch of I11143: signal is true;
	signal I11144: std_logic; attribute dont_touch of I11144: signal is true;
	signal I11149: std_logic; attribute dont_touch of I11149: signal is true;
	signal I11150: std_logic; attribute dont_touch of I11150: signal is true;
	signal I11151: std_logic; attribute dont_touch of I11151: signal is true;
	signal I11156: std_logic; attribute dont_touch of I11156: signal is true;
	signal I11157: std_logic; attribute dont_touch of I11157: signal is true;
	signal I11158: std_logic; attribute dont_touch of I11158: signal is true;
	signal I11163: std_logic; attribute dont_touch of I11163: signal is true;
	signal I11164: std_logic; attribute dont_touch of I11164: signal is true;
	signal I11165: std_logic; attribute dont_touch of I11165: signal is true;
	signal I11170: std_logic; attribute dont_touch of I11170: signal is true;
	signal I11171: std_logic; attribute dont_touch of I11171: signal is true;
	signal I11172: std_logic; attribute dont_touch of I11172: signal is true;
	signal I11177: std_logic; attribute dont_touch of I11177: signal is true;
	signal I11178: std_logic; attribute dont_touch of I11178: signal is true;
	signal I11179: std_logic; attribute dont_touch of I11179: signal is true;
	signal I11184: std_logic; attribute dont_touch of I11184: signal is true;
	signal I11185: std_logic; attribute dont_touch of I11185: signal is true;
	signal I11186: std_logic; attribute dont_touch of I11186: signal is true;
	signal I11191: std_logic; attribute dont_touch of I11191: signal is true;
	signal I11194: std_logic; attribute dont_touch of I11194: signal is true;
	signal I11197: std_logic; attribute dont_touch of I11197: signal is true;
	signal I11200: std_logic; attribute dont_touch of I11200: signal is true;
	signal I11203: std_logic; attribute dont_touch of I11203: signal is true;
	signal I11206: std_logic; attribute dont_touch of I11206: signal is true;
	signal I11209: std_logic; attribute dont_touch of I11209: signal is true;
	signal I11212: std_logic; attribute dont_touch of I11212: signal is true;
	signal I11215: std_logic; attribute dont_touch of I11215: signal is true;
	signal I11218: std_logic; attribute dont_touch of I11218: signal is true;
	signal I11221: std_logic; attribute dont_touch of I11221: signal is true;
	signal I11224: std_logic; attribute dont_touch of I11224: signal is true;
	signal I11227: std_logic; attribute dont_touch of I11227: signal is true;
	signal I11230: std_logic; attribute dont_touch of I11230: signal is true;
	signal I11233: std_logic; attribute dont_touch of I11233: signal is true;
	signal I11236: std_logic; attribute dont_touch of I11236: signal is true;
	signal I11239: std_logic; attribute dont_touch of I11239: signal is true;
	signal I11242: std_logic; attribute dont_touch of I11242: signal is true;
	signal I11245: std_logic; attribute dont_touch of I11245: signal is true;
	signal I11248: std_logic; attribute dont_touch of I11248: signal is true;
	signal I11251: std_logic; attribute dont_touch of I11251: signal is true;
	signal I11254: std_logic; attribute dont_touch of I11254: signal is true;
	signal I11257: std_logic; attribute dont_touch of I11257: signal is true;
	signal I11260: std_logic; attribute dont_touch of I11260: signal is true;
	signal I11263: std_logic; attribute dont_touch of I11263: signal is true;
	signal I11266: std_logic; attribute dont_touch of I11266: signal is true;
	signal I11269: std_logic; attribute dont_touch of I11269: signal is true;
	signal I11272: std_logic; attribute dont_touch of I11272: signal is true;
	signal I11275: std_logic; attribute dont_touch of I11275: signal is true;
	signal I11278: std_logic; attribute dont_touch of I11278: signal is true;
	signal I11281: std_logic; attribute dont_touch of I11281: signal is true;
	signal I11284: std_logic; attribute dont_touch of I11284: signal is true;
	signal I11287: std_logic; attribute dont_touch of I11287: signal is true;
	signal I11290: std_logic; attribute dont_touch of I11290: signal is true;
	signal I11293: std_logic; attribute dont_touch of I11293: signal is true;
	signal I11296: std_logic; attribute dont_touch of I11296: signal is true;
	signal I11299: std_logic; attribute dont_touch of I11299: signal is true;
	signal I11302: std_logic; attribute dont_touch of I11302: signal is true;
	signal I11305: std_logic; attribute dont_touch of I11305: signal is true;
	signal I11308: std_logic; attribute dont_touch of I11308: signal is true;
	signal I11311: std_logic; attribute dont_touch of I11311: signal is true;
	signal I11314: std_logic; attribute dont_touch of I11314: signal is true;
	signal I11317: std_logic; attribute dont_touch of I11317: signal is true;
	signal I11320: std_logic; attribute dont_touch of I11320: signal is true;
	signal I11323: std_logic; attribute dont_touch of I11323: signal is true;
	signal I11326: std_logic; attribute dont_touch of I11326: signal is true;
	signal I11329: std_logic; attribute dont_touch of I11329: signal is true;
	signal I11332: std_logic; attribute dont_touch of I11332: signal is true;
	signal I11335: std_logic; attribute dont_touch of I11335: signal is true;
	signal I11338: std_logic; attribute dont_touch of I11338: signal is true;
	signal I11341: std_logic; attribute dont_touch of I11341: signal is true;
	signal I11344: std_logic; attribute dont_touch of I11344: signal is true;
	signal I11347: std_logic; attribute dont_touch of I11347: signal is true;
	signal I11350: std_logic; attribute dont_touch of I11350: signal is true;
	signal I11353: std_logic; attribute dont_touch of I11353: signal is true;
	signal I11356: std_logic; attribute dont_touch of I11356: signal is true;
	signal I11359: std_logic; attribute dont_touch of I11359: signal is true;
	signal I11362: std_logic; attribute dont_touch of I11362: signal is true;
	signal I11365: std_logic; attribute dont_touch of I11365: signal is true;
	signal I11368: std_logic; attribute dont_touch of I11368: signal is true;
	signal I11371: std_logic; attribute dont_touch of I11371: signal is true;
	signal I11374: std_logic; attribute dont_touch of I11374: signal is true;
	signal I11377: std_logic; attribute dont_touch of I11377: signal is true;
	signal I11380: std_logic; attribute dont_touch of I11380: signal is true;
	signal I11383: std_logic; attribute dont_touch of I11383: signal is true;
	signal I11386: std_logic; attribute dont_touch of I11386: signal is true;
	signal I11389: std_logic; attribute dont_touch of I11389: signal is true;
	signal I11392: std_logic; attribute dont_touch of I11392: signal is true;
	signal I11395: std_logic; attribute dont_touch of I11395: signal is true;
	signal I11398: std_logic; attribute dont_touch of I11398: signal is true;
	signal I11401: std_logic; attribute dont_touch of I11401: signal is true;
	signal I11404: std_logic; attribute dont_touch of I11404: signal is true;
	signal I11407: std_logic; attribute dont_touch of I11407: signal is true;
	signal I11410: std_logic; attribute dont_touch of I11410: signal is true;
	signal I11413: std_logic; attribute dont_touch of I11413: signal is true;
	signal I11416: std_logic; attribute dont_touch of I11416: signal is true;
	signal I11419: std_logic; attribute dont_touch of I11419: signal is true;
	signal I11422: std_logic; attribute dont_touch of I11422: signal is true;
	signal I11425: std_logic; attribute dont_touch of I11425: signal is true;
	signal I11428: std_logic; attribute dont_touch of I11428: signal is true;
	signal I11431: std_logic; attribute dont_touch of I11431: signal is true;
	signal I11434: std_logic; attribute dont_touch of I11434: signal is true;
	signal I11437: std_logic; attribute dont_touch of I11437: signal is true;
	signal I11440: std_logic; attribute dont_touch of I11440: signal is true;
	signal I11443: std_logic; attribute dont_touch of I11443: signal is true;
	signal I11446: std_logic; attribute dont_touch of I11446: signal is true;
	signal I11449: std_logic; attribute dont_touch of I11449: signal is true;
	signal I11452: std_logic; attribute dont_touch of I11452: signal is true;
	signal I11455: std_logic; attribute dont_touch of I11455: signal is true;
	signal I11458: std_logic; attribute dont_touch of I11458: signal is true;
	signal I11461: std_logic; attribute dont_touch of I11461: signal is true;
	signal I11464: std_logic; attribute dont_touch of I11464: signal is true;
	signal I11467: std_logic; attribute dont_touch of I11467: signal is true;
	signal I11470: std_logic; attribute dont_touch of I11470: signal is true;
	signal I11473: std_logic; attribute dont_touch of I11473: signal is true;
	signal I11476: std_logic; attribute dont_touch of I11476: signal is true;
	signal I11479: std_logic; attribute dont_touch of I11479: signal is true;
	signal I11482: std_logic; attribute dont_touch of I11482: signal is true;
	signal I11485: std_logic; attribute dont_touch of I11485: signal is true;
	signal I11488: std_logic; attribute dont_touch of I11488: signal is true;
	signal I11491: std_logic; attribute dont_touch of I11491: signal is true;
	signal I11494: std_logic; attribute dont_touch of I11494: signal is true;
	signal I11497: std_logic; attribute dont_touch of I11497: signal is true;
	signal I11500: std_logic; attribute dont_touch of I11500: signal is true;
	signal I11503: std_logic; attribute dont_touch of I11503: signal is true;
	signal I11506: std_logic; attribute dont_touch of I11506: signal is true;
	signal I11512: std_logic; attribute dont_touch of I11512: signal is true;
	signal I11515: std_logic; attribute dont_touch of I11515: signal is true;
	signal I11522: std_logic; attribute dont_touch of I11522: signal is true;
	signal I11525: std_logic; attribute dont_touch of I11525: signal is true;
	signal I11533: std_logic; attribute dont_touch of I11533: signal is true;
	signal I11549: std_logic; attribute dont_touch of I11549: signal is true;
	signal I11550: std_logic; attribute dont_touch of I11550: signal is true;
	signal I11551: std_logic; attribute dont_touch of I11551: signal is true;
	signal I11556: std_logic; attribute dont_touch of I11556: signal is true;
	signal I11559: std_logic; attribute dont_touch of I11559: signal is true;
	signal I11562: std_logic; attribute dont_touch of I11562: signal is true;
	signal I11569: std_logic; attribute dont_touch of I11569: signal is true;
	signal I11574: std_logic; attribute dont_touch of I11574: signal is true;
	signal I11575: std_logic; attribute dont_touch of I11575: signal is true;
	signal I11576: std_logic; attribute dont_touch of I11576: signal is true;
	signal I11586: std_logic; attribute dont_touch of I11586: signal is true;
	signal I11591: std_logic; attribute dont_touch of I11591: signal is true;
	signal I11596: std_logic; attribute dont_touch of I11596: signal is true;
	signal I11603: std_logic; attribute dont_touch of I11603: signal is true;
	signal I11607: std_logic; attribute dont_touch of I11607: signal is true;
	signal I11614: std_logic; attribute dont_touch of I11614: signal is true;
	signal I11615: std_logic; attribute dont_touch of I11615: signal is true;
	signal I11616: std_logic; attribute dont_touch of I11616: signal is true;
	signal I11622: std_logic; attribute dont_touch of I11622: signal is true;
	signal I11627: std_logic; attribute dont_touch of I11627: signal is true;
	signal I11633: std_logic; attribute dont_touch of I11633: signal is true;
	signal I11638: std_logic; attribute dont_touch of I11638: signal is true;
	signal I11641: std_logic; attribute dont_touch of I11641: signal is true;
	signal I11645: std_logic; attribute dont_touch of I11645: signal is true;
	signal I11648: std_logic; attribute dont_touch of I11648: signal is true;
	signal I11652: std_logic; attribute dont_touch of I11652: signal is true;
	signal I11656: std_logic; attribute dont_touch of I11656: signal is true;
	signal I11659: std_logic; attribute dont_touch of I11659: signal is true;
	signal I11662: std_logic; attribute dont_touch of I11662: signal is true;
	signal I11666: std_logic; attribute dont_touch of I11666: signal is true;
	signal I11669: std_logic; attribute dont_touch of I11669: signal is true;
	signal I11672: std_logic; attribute dont_touch of I11672: signal is true;
	signal I11677: std_logic; attribute dont_touch of I11677: signal is true;
	signal I11680: std_logic; attribute dont_touch of I11680: signal is true;
	signal I11683: std_logic; attribute dont_touch of I11683: signal is true;
	signal I11686: std_logic; attribute dont_touch of I11686: signal is true;
	signal I11689: std_logic; attribute dont_touch of I11689: signal is true;
	signal I11693: std_logic; attribute dont_touch of I11693: signal is true;
	signal I11696: std_logic; attribute dont_touch of I11696: signal is true;
	signal I11701: std_logic; attribute dont_touch of I11701: signal is true;
	signal I11704: std_logic; attribute dont_touch of I11704: signal is true;
	signal I11707: std_logic; attribute dont_touch of I11707: signal is true;
	signal I11710: std_logic; attribute dont_touch of I11710: signal is true;
	signal I11714: std_logic; attribute dont_touch of I11714: signal is true;
	signal I11718: std_logic; attribute dont_touch of I11718: signal is true;
	signal I11722: std_logic; attribute dont_touch of I11722: signal is true;
	signal I11725: std_logic; attribute dont_touch of I11725: signal is true;
	signal I11729: std_logic; attribute dont_touch of I11729: signal is true;
	signal I11732: std_logic; attribute dont_touch of I11732: signal is true;
	signal I11736: std_logic; attribute dont_touch of I11736: signal is true;
	signal I11740: std_logic; attribute dont_touch of I11740: signal is true;
	signal I11744: std_logic; attribute dont_touch of I11744: signal is true;
	signal I11747: std_logic; attribute dont_touch of I11747: signal is true;
	signal I11750: std_logic; attribute dont_touch of I11750: signal is true;
	signal I11751: std_logic; attribute dont_touch of I11751: signal is true;
	signal I11752: std_logic; attribute dont_touch of I11752: signal is true;
	signal I11757: std_logic; attribute dont_touch of I11757: signal is true;
	signal I11758: std_logic; attribute dont_touch of I11758: signal is true;
	signal I11759: std_logic; attribute dont_touch of I11759: signal is true;
	signal I11764: std_logic; attribute dont_touch of I11764: signal is true;
	signal I11773: std_logic; attribute dont_touch of I11773: signal is true;
	signal I11778: std_logic; attribute dont_touch of I11778: signal is true;
	signal I11781: std_logic; attribute dont_touch of I11781: signal is true;
	signal I11787: std_logic; attribute dont_touch of I11787: signal is true;
	signal I11790: std_logic; attribute dont_touch of I11790: signal is true;
	signal I11793: std_logic; attribute dont_touch of I11793: signal is true;
	signal I11796: std_logic; attribute dont_touch of I11796: signal is true;
	signal I11800: std_logic; attribute dont_touch of I11800: signal is true;
	signal I11803: std_logic; attribute dont_touch of I11803: signal is true;
	signal I11806: std_logic; attribute dont_touch of I11806: signal is true;
	signal I11809: std_logic; attribute dont_touch of I11809: signal is true;
	signal I11815: std_logic; attribute dont_touch of I11815: signal is true;
	signal I11818: std_logic; attribute dont_touch of I11818: signal is true;
	signal I11821: std_logic; attribute dont_touch of I11821: signal is true;
	signal I11824: std_logic; attribute dont_touch of I11824: signal is true;
	signal I11827: std_logic; attribute dont_touch of I11827: signal is true;
	signal I11832: std_logic; attribute dont_touch of I11832: signal is true;
	signal I11835: std_logic; attribute dont_touch of I11835: signal is true;
	signal I11838: std_logic; attribute dont_touch of I11838: signal is true;
	signal I11841: std_logic; attribute dont_touch of I11841: signal is true;
	signal I11842: std_logic; attribute dont_touch of I11842: signal is true;
	signal I11843: std_logic; attribute dont_touch of I11843: signal is true;
	signal I11848: std_logic; attribute dont_touch of I11848: signal is true;
	signal I11851: std_logic; attribute dont_touch of I11851: signal is true;
	signal I11855: std_logic; attribute dont_touch of I11855: signal is true;
	signal I11858: std_logic; attribute dont_touch of I11858: signal is true;
	signal I11861: std_logic; attribute dont_touch of I11861: signal is true;
	signal I11864: std_logic; attribute dont_touch of I11864: signal is true;
	signal I11867: std_logic; attribute dont_touch of I11867: signal is true;
	signal I11870: std_logic; attribute dont_touch of I11870: signal is true;
	signal I11873: std_logic; attribute dont_touch of I11873: signal is true;
	signal I11874: std_logic; attribute dont_touch of I11874: signal is true;
	signal I11875: std_logic; attribute dont_touch of I11875: signal is true;
	signal I11880: std_logic; attribute dont_touch of I11880: signal is true;
	signal I11884: std_logic; attribute dont_touch of I11884: signal is true;
	signal I11887: std_logic; attribute dont_touch of I11887: signal is true;
	signal I11890: std_logic; attribute dont_touch of I11890: signal is true;
	signal I11894: std_logic; attribute dont_touch of I11894: signal is true;
	signal I11897: std_logic; attribute dont_touch of I11897: signal is true;
	signal I11900: std_logic; attribute dont_touch of I11900: signal is true;
	signal I11903: std_logic; attribute dont_touch of I11903: signal is true;
	signal I11908: std_logic; attribute dont_touch of I11908: signal is true;
	signal I11912: std_logic; attribute dont_touch of I11912: signal is true;
	signal I11917: std_logic; attribute dont_touch of I11917: signal is true;
	signal I11920: std_logic; attribute dont_touch of I11920: signal is true;
	signal I11923: std_logic; attribute dont_touch of I11923: signal is true;
	signal I11926: std_logic; attribute dont_touch of I11926: signal is true;
	signal I11929: std_logic; attribute dont_touch of I11929: signal is true;
	signal I11933: std_logic; attribute dont_touch of I11933: signal is true;
	signal I11936: std_logic; attribute dont_touch of I11936: signal is true;
	signal I11939: std_logic; attribute dont_touch of I11939: signal is true;
	signal I11942: std_logic; attribute dont_touch of I11942: signal is true;
	signal I11945: std_logic; attribute dont_touch of I11945: signal is true;
	signal I11948: std_logic; attribute dont_touch of I11948: signal is true;
	signal I11951: std_logic; attribute dont_touch of I11951: signal is true;
	signal I11955: std_logic; attribute dont_touch of I11955: signal is true;
	signal I11958: std_logic; attribute dont_touch of I11958: signal is true;
	signal I11961: std_logic; attribute dont_touch of I11961: signal is true;
	signal I11964: std_logic; attribute dont_touch of I11964: signal is true;
	signal I11967: std_logic; attribute dont_touch of I11967: signal is true;
	signal I11971: std_logic; attribute dont_touch of I11971: signal is true;
	signal I11974: std_logic; attribute dont_touch of I11974: signal is true;
	signal I11978: std_logic; attribute dont_touch of I11978: signal is true;
	signal I11981: std_logic; attribute dont_touch of I11981: signal is true;
	signal I11984: std_logic; attribute dont_touch of I11984: signal is true;
	signal I11987: std_logic; attribute dont_touch of I11987: signal is true;
	signal I11991: std_logic; attribute dont_touch of I11991: signal is true;
	signal I11994: std_logic; attribute dont_touch of I11994: signal is true;
	signal I11998: std_logic; attribute dont_touch of I11998: signal is true;
	signal I12003: std_logic; attribute dont_touch of I12003: signal is true;
	signal I12008: std_logic; attribute dont_touch of I12008: signal is true;
	signal I12011: std_logic; attribute dont_touch of I12011: signal is true;
	signal I12015: std_logic; attribute dont_touch of I12015: signal is true;
	signal I12016: std_logic; attribute dont_touch of I12016: signal is true;
	signal I12017: std_logic; attribute dont_touch of I12017: signal is true;
	signal I12022: std_logic; attribute dont_touch of I12022: signal is true;
	signal I12025: std_logic; attribute dont_touch of I12025: signal is true;
	signal I12031: std_logic; attribute dont_touch of I12031: signal is true;
	signal I12032: std_logic; attribute dont_touch of I12032: signal is true;
	signal I12033: std_logic; attribute dont_touch of I12033: signal is true;
	signal I12038: std_logic; attribute dont_touch of I12038: signal is true;
	signal I12041: std_logic; attribute dont_touch of I12041: signal is true;
	signal I12044: std_logic; attribute dont_touch of I12044: signal is true;
	signal I12051: std_logic; attribute dont_touch of I12051: signal is true;
	signal I12052: std_logic; attribute dont_touch of I12052: signal is true;
	signal I12053: std_logic; attribute dont_touch of I12053: signal is true;
	signal I12059: std_logic; attribute dont_touch of I12059: signal is true;
	signal I12062: std_logic; attribute dont_touch of I12062: signal is true;
	signal I12065: std_logic; attribute dont_touch of I12065: signal is true;
	signal I12068: std_logic; attribute dont_touch of I12068: signal is true;
	signal I12078: std_logic; attribute dont_touch of I12078: signal is true;
	signal I12079: std_logic; attribute dont_touch of I12079: signal is true;
	signal I12080: std_logic; attribute dont_touch of I12080: signal is true;
	signal I12085: std_logic; attribute dont_touch of I12085: signal is true;
	signal I12088: std_logic; attribute dont_touch of I12088: signal is true;
	signal I12091: std_logic; attribute dont_touch of I12091: signal is true;
	signal I12098: std_logic; attribute dont_touch of I12098: signal is true;
	signal I12101: std_logic; attribute dont_touch of I12101: signal is true;
	signal I12108: std_logic; attribute dont_touch of I12108: signal is true;
	signal I12111: std_logic; attribute dont_touch of I12111: signal is true;
	signal I12117: std_logic; attribute dont_touch of I12117: signal is true;
	signal I12120: std_logic; attribute dont_touch of I12120: signal is true;
	signal I12124: std_logic; attribute dont_touch of I12124: signal is true;
	signal I12128: std_logic; attribute dont_touch of I12128: signal is true;
	signal I12131: std_logic; attribute dont_touch of I12131: signal is true;
	signal I12135: std_logic; attribute dont_touch of I12135: signal is true;
	signal I12138: std_logic; attribute dont_touch of I12138: signal is true;
	signal I12141: std_logic; attribute dont_touch of I12141: signal is true;
	signal I12145: std_logic; attribute dont_touch of I12145: signal is true;
	signal I12148: std_logic; attribute dont_touch of I12148: signal is true;
	signal I12151: std_logic; attribute dont_touch of I12151: signal is true;
	signal I12154: std_logic; attribute dont_touch of I12154: signal is true;
	signal I12158: std_logic; attribute dont_touch of I12158: signal is true;
	signal I12161: std_logic; attribute dont_touch of I12161: signal is true;
	signal I12164: std_logic; attribute dont_touch of I12164: signal is true;
	signal I12167: std_logic; attribute dont_touch of I12167: signal is true;
	signal I12170: std_logic; attribute dont_touch of I12170: signal is true;
	signal I12173: std_logic; attribute dont_touch of I12173: signal is true;
	signal I12176: std_logic; attribute dont_touch of I12176: signal is true;
	signal I12179: std_logic; attribute dont_touch of I12179: signal is true;
	signal I12180: std_logic; attribute dont_touch of I12180: signal is true;
	signal I12181: std_logic; attribute dont_touch of I12181: signal is true;
	signal I12187: std_logic; attribute dont_touch of I12187: signal is true;
	signal I12190: std_logic; attribute dont_touch of I12190: signal is true;
	signal I12193: std_logic; attribute dont_touch of I12193: signal is true;
	signal I12196: std_logic; attribute dont_touch of I12196: signal is true;
	signal I12199: std_logic; attribute dont_touch of I12199: signal is true;
	signal I12202: std_logic; attribute dont_touch of I12202: signal is true;
	signal I12205: std_logic; attribute dont_touch of I12205: signal is true;
	signal I12208: std_logic; attribute dont_touch of I12208: signal is true;
	signal I12211: std_logic; attribute dont_touch of I12211: signal is true;
	signal I12214: std_logic; attribute dont_touch of I12214: signal is true;
	signal I12217: std_logic; attribute dont_touch of I12217: signal is true;
	signal I12220: std_logic; attribute dont_touch of I12220: signal is true;
	signal I12223: std_logic; attribute dont_touch of I12223: signal is true;
	signal I12226: std_logic; attribute dont_touch of I12226: signal is true;
	signal I12229: std_logic; attribute dont_touch of I12229: signal is true;
	signal I12232: std_logic; attribute dont_touch of I12232: signal is true;
	signal I12235: std_logic; attribute dont_touch of I12235: signal is true;
	signal I12238: std_logic; attribute dont_touch of I12238: signal is true;
	signal I12241: std_logic; attribute dont_touch of I12241: signal is true;
	signal I12244: std_logic; attribute dont_touch of I12244: signal is true;
	signal I12247: std_logic; attribute dont_touch of I12247: signal is true;
	signal I12250: std_logic; attribute dont_touch of I12250: signal is true;
	signal I12253: std_logic; attribute dont_touch of I12253: signal is true;
	signal I12256: std_logic; attribute dont_touch of I12256: signal is true;
	signal I12259: std_logic; attribute dont_touch of I12259: signal is true;
	signal I12262: std_logic; attribute dont_touch of I12262: signal is true;
	signal I12265: std_logic; attribute dont_touch of I12265: signal is true;
	signal I12268: std_logic; attribute dont_touch of I12268: signal is true;
	signal I12271: std_logic; attribute dont_touch of I12271: signal is true;
	signal I12274: std_logic; attribute dont_touch of I12274: signal is true;
	signal I12277: std_logic; attribute dont_touch of I12277: signal is true;
	signal I12280: std_logic; attribute dont_touch of I12280: signal is true;
	signal I12283: std_logic; attribute dont_touch of I12283: signal is true;
	signal I12286: std_logic; attribute dont_touch of I12286: signal is true;
	signal I12289: std_logic; attribute dont_touch of I12289: signal is true;
	signal I12292: std_logic; attribute dont_touch of I12292: signal is true;
	signal I12295: std_logic; attribute dont_touch of I12295: signal is true;
	signal I12298: std_logic; attribute dont_touch of I12298: signal is true;
	signal I12301: std_logic; attribute dont_touch of I12301: signal is true;
	signal I12304: std_logic; attribute dont_touch of I12304: signal is true;
	signal I12307: std_logic; attribute dont_touch of I12307: signal is true;
	signal I12310: std_logic; attribute dont_touch of I12310: signal is true;
	signal I12313: std_logic; attribute dont_touch of I12313: signal is true;
	signal I12316: std_logic; attribute dont_touch of I12316: signal is true;
	signal I12319: std_logic; attribute dont_touch of I12319: signal is true;
	signal I12322: std_logic; attribute dont_touch of I12322: signal is true;
	signal I12325: std_logic; attribute dont_touch of I12325: signal is true;
	signal I12328: std_logic; attribute dont_touch of I12328: signal is true;
	signal I12331: std_logic; attribute dont_touch of I12331: signal is true;
	signal I12334: std_logic; attribute dont_touch of I12334: signal is true;
	signal I12337: std_logic; attribute dont_touch of I12337: signal is true;
	signal I12340: std_logic; attribute dont_touch of I12340: signal is true;
	signal I12343: std_logic; attribute dont_touch of I12343: signal is true;
	signal I12346: std_logic; attribute dont_touch of I12346: signal is true;
	signal I12349: std_logic; attribute dont_touch of I12349: signal is true;
	signal I12352: std_logic; attribute dont_touch of I12352: signal is true;
	signal I12355: std_logic; attribute dont_touch of I12355: signal is true;
	signal I12358: std_logic; attribute dont_touch of I12358: signal is true;
	signal I12361: std_logic; attribute dont_touch of I12361: signal is true;
	signal I12364: std_logic; attribute dont_touch of I12364: signal is true;
	signal I12367: std_logic; attribute dont_touch of I12367: signal is true;
	signal I12370: std_logic; attribute dont_touch of I12370: signal is true;
	signal I12373: std_logic; attribute dont_touch of I12373: signal is true;
	signal I12376: std_logic; attribute dont_touch of I12376: signal is true;
	signal I12379: std_logic; attribute dont_touch of I12379: signal is true;
	signal I12382: std_logic; attribute dont_touch of I12382: signal is true;
	signal I12385: std_logic; attribute dont_touch of I12385: signal is true;
	signal I12388: std_logic; attribute dont_touch of I12388: signal is true;
	signal I12391: std_logic; attribute dont_touch of I12391: signal is true;
	signal I12394: std_logic; attribute dont_touch of I12394: signal is true;
	signal I12397: std_logic; attribute dont_touch of I12397: signal is true;
	signal I12400: std_logic; attribute dont_touch of I12400: signal is true;
	signal I12403: std_logic; attribute dont_touch of I12403: signal is true;
	signal I12406: std_logic; attribute dont_touch of I12406: signal is true;
	signal I12409: std_logic; attribute dont_touch of I12409: signal is true;
	signal I12412: std_logic; attribute dont_touch of I12412: signal is true;
	signal I12415: std_logic; attribute dont_touch of I12415: signal is true;
	signal I12418: std_logic; attribute dont_touch of I12418: signal is true;
	signal I12421: std_logic; attribute dont_touch of I12421: signal is true;
	signal I12424: std_logic; attribute dont_touch of I12424: signal is true;
	signal I12427: std_logic; attribute dont_touch of I12427: signal is true;
	signal I12430: std_logic; attribute dont_touch of I12430: signal is true;
	signal I12433: std_logic; attribute dont_touch of I12433: signal is true;
	signal I12436: std_logic; attribute dont_touch of I12436: signal is true;
	signal I12439: std_logic; attribute dont_touch of I12439: signal is true;
	signal I12442: std_logic; attribute dont_touch of I12442: signal is true;
	signal I12445: std_logic; attribute dont_touch of I12445: signal is true;
	signal I12448: std_logic; attribute dont_touch of I12448: signal is true;
	signal I12451: std_logic; attribute dont_touch of I12451: signal is true;
	signal I12454: std_logic; attribute dont_touch of I12454: signal is true;
	signal I12457: std_logic; attribute dont_touch of I12457: signal is true;
	signal I12460: std_logic; attribute dont_touch of I12460: signal is true;
	signal I12463: std_logic; attribute dont_touch of I12463: signal is true;
	signal I12466: std_logic; attribute dont_touch of I12466: signal is true;
	signal I12469: std_logic; attribute dont_touch of I12469: signal is true;
	signal I12472: std_logic; attribute dont_touch of I12472: signal is true;
	signal I12475: std_logic; attribute dont_touch of I12475: signal is true;
	signal I12478: std_logic; attribute dont_touch of I12478: signal is true;
	signal I12481: std_logic; attribute dont_touch of I12481: signal is true;
	signal I12484: std_logic; attribute dont_touch of I12484: signal is true;
	signal I12487: std_logic; attribute dont_touch of I12487: signal is true;
	signal I12490: std_logic; attribute dont_touch of I12490: signal is true;
	signal I12493: std_logic; attribute dont_touch of I12493: signal is true;
	signal I12496: std_logic; attribute dont_touch of I12496: signal is true;
	signal I12499: std_logic; attribute dont_touch of I12499: signal is true;
	signal I12502: std_logic; attribute dont_touch of I12502: signal is true;
	signal I12505: std_logic; attribute dont_touch of I12505: signal is true;
	signal I12508: std_logic; attribute dont_touch of I12508: signal is true;
	signal I12511: std_logic; attribute dont_touch of I12511: signal is true;
	signal I12514: std_logic; attribute dont_touch of I12514: signal is true;
	signal I12517: std_logic; attribute dont_touch of I12517: signal is true;
	signal I12520: std_logic; attribute dont_touch of I12520: signal is true;
	signal I12523: std_logic; attribute dont_touch of I12523: signal is true;
	signal I12526: std_logic; attribute dont_touch of I12526: signal is true;
	signal I12529: std_logic; attribute dont_touch of I12529: signal is true;
	signal I12532: std_logic; attribute dont_touch of I12532: signal is true;
	signal I12535: std_logic; attribute dont_touch of I12535: signal is true;
	signal I12538: std_logic; attribute dont_touch of I12538: signal is true;
	signal I12541: std_logic; attribute dont_touch of I12541: signal is true;
	signal I12544: std_logic; attribute dont_touch of I12544: signal is true;
	signal I12547: std_logic; attribute dont_touch of I12547: signal is true;
	signal I12550: std_logic; attribute dont_touch of I12550: signal is true;
	signal I12551: std_logic; attribute dont_touch of I12551: signal is true;
	signal I12552: std_logic; attribute dont_touch of I12552: signal is true;
	signal I12558: std_logic; attribute dont_touch of I12558: signal is true;
	signal I12561: std_logic; attribute dont_touch of I12561: signal is true;
	signal I12564: std_logic; attribute dont_touch of I12564: signal is true;
	signal I12567: std_logic; attribute dont_touch of I12567: signal is true;
	signal I12571: std_logic; attribute dont_touch of I12571: signal is true;
	signal I12575: std_logic; attribute dont_touch of I12575: signal is true;
	signal I12576: std_logic; attribute dont_touch of I12576: signal is true;
	signal I12577: std_logic; attribute dont_touch of I12577: signal is true;
	signal I12582: std_logic; attribute dont_touch of I12582: signal is true;
	signal I12586: std_logic; attribute dont_touch of I12586: signal is true;
	signal I12592: std_logic; attribute dont_touch of I12592: signal is true;
	signal I12596: std_logic; attribute dont_touch of I12596: signal is true;
	signal I12597: std_logic; attribute dont_touch of I12597: signal is true;
	signal I12598: std_logic; attribute dont_touch of I12598: signal is true;
	signal I12609: std_logic; attribute dont_touch of I12609: signal is true;
	signal I12629: std_logic; attribute dont_touch of I12629: signal is true;
	signal I12632: std_logic; attribute dont_touch of I12632: signal is true;
	signal I12635: std_logic; attribute dont_touch of I12635: signal is true;
	signal I12639: std_logic; attribute dont_touch of I12639: signal is true;
	signal I12643: std_logic; attribute dont_touch of I12643: signal is true;
	signal I12646: std_logic; attribute dont_touch of I12646: signal is true;
	signal I12649: std_logic; attribute dont_touch of I12649: signal is true;
	signal I12652: std_logic; attribute dont_touch of I12652: signal is true;
	signal I12655: std_logic; attribute dont_touch of I12655: signal is true;
	signal I12659: std_logic; attribute dont_touch of I12659: signal is true;
	signal I12666: std_logic; attribute dont_touch of I12666: signal is true;
	signal I12669: std_logic; attribute dont_touch of I12669: signal is true;
	signal I12672: std_logic; attribute dont_touch of I12672: signal is true;
	signal I12675: std_logic; attribute dont_touch of I12675: signal is true;
	signal I12678: std_logic; attribute dont_touch of I12678: signal is true;
	signal I12681: std_logic; attribute dont_touch of I12681: signal is true;
	signal I12684: std_logic; attribute dont_touch of I12684: signal is true;
	signal I12687: std_logic; attribute dont_touch of I12687: signal is true;
	signal I12690: std_logic; attribute dont_touch of I12690: signal is true;
	signal I12696: std_logic; attribute dont_touch of I12696: signal is true;
	signal I12699: std_logic; attribute dont_touch of I12699: signal is true;
	signal I12702: std_logic; attribute dont_touch of I12702: signal is true;
	signal I12708: std_logic; attribute dont_touch of I12708: signal is true;
	signal I12712: std_logic; attribute dont_touch of I12712: signal is true;
	signal I12717: std_logic; attribute dont_touch of I12717: signal is true;
	signal I12722: std_logic; attribute dont_touch of I12722: signal is true;
	signal I12725: std_logic; attribute dont_touch of I12725: signal is true;
	signal I12731: std_logic; attribute dont_touch of I12731: signal is true;
	signal I12737: std_logic; attribute dont_touch of I12737: signal is true;
	signal I12742: std_logic; attribute dont_touch of I12742: signal is true;
	signal I12748: std_logic; attribute dont_touch of I12748: signal is true;
	signal I12753: std_logic; attribute dont_touch of I12753: signal is true;
	signal I12757: std_logic; attribute dont_touch of I12757: signal is true;
	signal I12760: std_logic; attribute dont_touch of I12760: signal is true;
	signal I12763: std_logic; attribute dont_touch of I12763: signal is true;
	signal I12768: std_logic; attribute dont_touch of I12768: signal is true;
	signal I12771: std_logic; attribute dont_touch of I12771: signal is true;
	signal I12776: std_logic; attribute dont_touch of I12776: signal is true;
	signal I12779: std_logic; attribute dont_touch of I12779: signal is true;
	signal I12782: std_logic; attribute dont_touch of I12782: signal is true;
	signal I12806: std_logic; attribute dont_touch of I12806: signal is true;
	signal I12810: std_logic; attribute dont_touch of I12810: signal is true;
	signal I12813: std_logic; attribute dont_touch of I12813: signal is true;
	signal I12826: std_logic; attribute dont_touch of I12826: signal is true;
	signal I12829: std_logic; attribute dont_touch of I12829: signal is true;
	signal I12832: std_logic; attribute dont_touch of I12832: signal is true;
	signal I12833: std_logic; attribute dont_touch of I12833: signal is true;
	signal I12834: std_logic; attribute dont_touch of I12834: signal is true;
	signal I12839: std_logic; attribute dont_touch of I12839: signal is true;
	signal I12852: std_logic; attribute dont_touch of I12852: signal is true;
	signal I12853: std_logic; attribute dont_touch of I12853: signal is true;
	signal I12854: std_logic; attribute dont_touch of I12854: signal is true;
	signal I12866: std_logic; attribute dont_touch of I12866: signal is true;
	signal I12869: std_logic; attribute dont_touch of I12869: signal is true;
	signal I12870: std_logic; attribute dont_touch of I12870: signal is true;
	signal I12871: std_logic; attribute dont_touch of I12871: signal is true;
	signal I12877: std_logic; attribute dont_touch of I12877: signal is true;
	signal I12881: std_logic; attribute dont_touch of I12881: signal is true;
	signal I12885: std_logic; attribute dont_touch of I12885: signal is true;
	signal I12888: std_logic; attribute dont_touch of I12888: signal is true;
	signal I12891: std_logic; attribute dont_touch of I12891: signal is true;
	signal I12894: std_logic; attribute dont_touch of I12894: signal is true;
	signal I12897: std_logic; attribute dont_touch of I12897: signal is true;
	signal I12900: std_logic; attribute dont_touch of I12900: signal is true;
	signal I12903: std_logic; attribute dont_touch of I12903: signal is true;
	signal I12906: std_logic; attribute dont_touch of I12906: signal is true;
	signal I12909: std_logic; attribute dont_touch of I12909: signal is true;
	signal I12912: std_logic; attribute dont_touch of I12912: signal is true;
	signal I12915: std_logic; attribute dont_touch of I12915: signal is true;
	signal I12918: std_logic; attribute dont_touch of I12918: signal is true;
	signal I12921: std_logic; attribute dont_touch of I12921: signal is true;
	signal I12924: std_logic; attribute dont_touch of I12924: signal is true;
	signal I12927: std_logic; attribute dont_touch of I12927: signal is true;
	signal I12930: std_logic; attribute dont_touch of I12930: signal is true;
	signal I12933: std_logic; attribute dont_touch of I12933: signal is true;
	signal I12936: std_logic; attribute dont_touch of I12936: signal is true;
	signal I12939: std_logic; attribute dont_touch of I12939: signal is true;
	signal I12942: std_logic; attribute dont_touch of I12942: signal is true;
	signal I12945: std_logic; attribute dont_touch of I12945: signal is true;
	signal I12948: std_logic; attribute dont_touch of I12948: signal is true;
	signal I12951: std_logic; attribute dont_touch of I12951: signal is true;
	signal I12952: std_logic; attribute dont_touch of I12952: signal is true;
	signal I12953: std_logic; attribute dont_touch of I12953: signal is true;
	signal I12958: std_logic; attribute dont_touch of I12958: signal is true;
	signal I12961: std_logic; attribute dont_touch of I12961: signal is true;
	signal I12965: std_logic; attribute dont_touch of I12965: signal is true;
	signal I12968: std_logic; attribute dont_touch of I12968: signal is true;
	signal I12973: std_logic; attribute dont_touch of I12973: signal is true;
	signal I12976: std_logic; attribute dont_touch of I12976: signal is true;
	signal I12980: std_logic; attribute dont_touch of I12980: signal is true;
	signal I12983: std_logic; attribute dont_touch of I12983: signal is true;
	signal I12986: std_logic; attribute dont_touch of I12986: signal is true;
	signal I12989: std_logic; attribute dont_touch of I12989: signal is true;
	signal I12993: std_logic; attribute dont_touch of I12993: signal is true;
	signal I12996: std_logic; attribute dont_touch of I12996: signal is true;
	signal I12999: std_logic; attribute dont_touch of I12999: signal is true;
	signal I13002: std_logic; attribute dont_touch of I13002: signal is true;
	signal I13003: std_logic; attribute dont_touch of I13003: signal is true;
	signal I13004: std_logic; attribute dont_touch of I13004: signal is true;
	signal I13009: std_logic; attribute dont_touch of I13009: signal is true;
	signal I13012: std_logic; attribute dont_touch of I13012: signal is true;
	signal I13016: std_logic; attribute dont_touch of I13016: signal is true;
	signal I13017: std_logic; attribute dont_touch of I13017: signal is true;
	signal I13018: std_logic; attribute dont_touch of I13018: signal is true;
	signal I13023: std_logic; attribute dont_touch of I13023: signal is true;
	signal I13028: std_logic; attribute dont_touch of I13028: signal is true;
	signal I13031: std_logic; attribute dont_touch of I13031: signal is true;
	signal I13035: std_logic; attribute dont_touch of I13035: signal is true;
	signal I13039: std_logic; attribute dont_touch of I13039: signal is true;
	signal I13042: std_logic; attribute dont_touch of I13042: signal is true;
	signal I13045: std_logic; attribute dont_touch of I13045: signal is true;
	signal I13048: std_logic; attribute dont_touch of I13048: signal is true;
	signal I13051: std_logic; attribute dont_touch of I13051: signal is true;
	signal I13054: std_logic; attribute dont_touch of I13054: signal is true;
	signal I13057: std_logic; attribute dont_touch of I13057: signal is true;
	signal I13060: std_logic; attribute dont_touch of I13060: signal is true;
	signal I13063: std_logic; attribute dont_touch of I13063: signal is true;
	signal I13066: std_logic; attribute dont_touch of I13066: signal is true;
	signal I13072: std_logic; attribute dont_touch of I13072: signal is true;
	signal I13075: std_logic; attribute dont_touch of I13075: signal is true;
	signal I13084: std_logic; attribute dont_touch of I13084: signal is true;
	signal I13088: std_logic; attribute dont_touch of I13088: signal is true;
	signal I13092: std_logic; attribute dont_touch of I13092: signal is true;
	signal I13099: std_logic; attribute dont_touch of I13099: signal is true;
	signal I13103: std_logic; attribute dont_touch of I13103: signal is true;
	signal I13106: std_logic; attribute dont_touch of I13106: signal is true;
	signal I13109: std_logic; attribute dont_touch of I13109: signal is true;
	signal I13112: std_logic; attribute dont_touch of I13112: signal is true;
	signal I13118: std_logic; attribute dont_touch of I13118: signal is true;
	signal I13122: std_logic; attribute dont_touch of I13122: signal is true;
	signal I13126: std_logic; attribute dont_touch of I13126: signal is true;
	signal I13131: std_logic; attribute dont_touch of I13131: signal is true;
	signal I13134: std_logic; attribute dont_touch of I13134: signal is true;
	signal I13137: std_logic; attribute dont_touch of I13137: signal is true;
	signal I13140: std_logic; attribute dont_touch of I13140: signal is true;
	signal I13144: std_logic; attribute dont_touch of I13144: signal is true;
	signal I13147: std_logic; attribute dont_touch of I13147: signal is true;
	signal I13152: std_logic; attribute dont_touch of I13152: signal is true;
	signal I13157: std_logic; attribute dont_touch of I13157: signal is true;
	signal I13161: std_logic; attribute dont_touch of I13161: signal is true;
	signal I13164: std_logic; attribute dont_touch of I13164: signal is true;
	signal I13173: std_logic; attribute dont_touch of I13173: signal is true;
	signal I13185: std_logic; attribute dont_touch of I13185: signal is true;
	signal I13189: std_logic; attribute dont_touch of I13189: signal is true;
	signal I13193: std_logic; attribute dont_touch of I13193: signal is true;
	signal I13196: std_logic; attribute dont_touch of I13196: signal is true;
	signal I13199: std_logic; attribute dont_touch of I13199: signal is true;
	signal I13203: std_logic; attribute dont_touch of I13203: signal is true;
	signal I13209: std_logic; attribute dont_touch of I13209: signal is true;
	signal I13213: std_logic; attribute dont_touch of I13213: signal is true;
	signal I13214: std_logic; attribute dont_touch of I13214: signal is true;
	signal I13215: std_logic; attribute dont_touch of I13215: signal is true;
	signal I13220: std_logic; attribute dont_touch of I13220: signal is true;
	signal I13225: std_logic; attribute dont_touch of I13225: signal is true;
	signal I13228: std_logic; attribute dont_touch of I13228: signal is true;
	signal I13231: std_logic; attribute dont_touch of I13231: signal is true;
	signal I13234: std_logic; attribute dont_touch of I13234: signal is true;
	signal I13238: std_logic; attribute dont_touch of I13238: signal is true;
	signal I13241: std_logic; attribute dont_touch of I13241: signal is true;
	signal I13244: std_logic; attribute dont_touch of I13244: signal is true;
	signal I13247: std_logic; attribute dont_touch of I13247: signal is true;
	signal I13250: std_logic; attribute dont_touch of I13250: signal is true;
	signal I13255: std_logic; attribute dont_touch of I13255: signal is true;
	signal I13258: std_logic; attribute dont_touch of I13258: signal is true;
	signal I13261: std_logic; attribute dont_touch of I13261: signal is true;
	signal I13264: std_logic; attribute dont_touch of I13264: signal is true;
	signal I13267: std_logic; attribute dont_touch of I13267: signal is true;
	signal I13271: std_logic; attribute dont_touch of I13271: signal is true;
	signal I13274: std_logic; attribute dont_touch of I13274: signal is true;
	signal I13277: std_logic; attribute dont_touch of I13277: signal is true;
	signal I13281: std_logic; attribute dont_touch of I13281: signal is true;
	signal I13284: std_logic; attribute dont_touch of I13284: signal is true;
	signal I13287: std_logic; attribute dont_touch of I13287: signal is true;
	signal I13290: std_logic; attribute dont_touch of I13290: signal is true;
	signal I13293: std_logic; attribute dont_touch of I13293: signal is true;
	signal I13296: std_logic; attribute dont_touch of I13296: signal is true;
	signal I13299: std_logic; attribute dont_touch of I13299: signal is true;
	signal I13302: std_logic; attribute dont_touch of I13302: signal is true;
	signal I13305: std_logic; attribute dont_touch of I13305: signal is true;
	signal I13308: std_logic; attribute dont_touch of I13308: signal is true;
	signal I13311: std_logic; attribute dont_touch of I13311: signal is true;
	signal I13314: std_logic; attribute dont_touch of I13314: signal is true;
	signal I13317: std_logic; attribute dont_touch of I13317: signal is true;
	signal I13320: std_logic; attribute dont_touch of I13320: signal is true;
	signal I13323: std_logic; attribute dont_touch of I13323: signal is true;
	signal I13326: std_logic; attribute dont_touch of I13326: signal is true;
	signal I13329: std_logic; attribute dont_touch of I13329: signal is true;
	signal I13332: std_logic; attribute dont_touch of I13332: signal is true;
	signal I13335: std_logic; attribute dont_touch of I13335: signal is true;
	signal I13338: std_logic; attribute dont_touch of I13338: signal is true;
	signal I13341: std_logic; attribute dont_touch of I13341: signal is true;
	signal I13344: std_logic; attribute dont_touch of I13344: signal is true;
	signal I13347: std_logic; attribute dont_touch of I13347: signal is true;
	signal I13350: std_logic; attribute dont_touch of I13350: signal is true;
	signal I13353: std_logic; attribute dont_touch of I13353: signal is true;
	signal I13356: std_logic; attribute dont_touch of I13356: signal is true;
	signal I13359: std_logic; attribute dont_touch of I13359: signal is true;
	signal I13362: std_logic; attribute dont_touch of I13362: signal is true;
	signal I13365: std_logic; attribute dont_touch of I13365: signal is true;
	signal I13369: std_logic; attribute dont_touch of I13369: signal is true;
	signal I13373: std_logic; attribute dont_touch of I13373: signal is true;
	signal I13376: std_logic; attribute dont_touch of I13376: signal is true;
	signal I13377: std_logic; attribute dont_touch of I13377: signal is true;
	signal I13378: std_logic; attribute dont_touch of I13378: signal is true;
	signal I13383: std_logic; attribute dont_touch of I13383: signal is true;
	signal I13388: std_logic; attribute dont_touch of I13388: signal is true;
	signal I13395: std_logic; attribute dont_touch of I13395: signal is true;
	signal I13396: std_logic; attribute dont_touch of I13396: signal is true;
	signal I13397: std_logic; attribute dont_touch of I13397: signal is true;
	signal I13403: std_logic; attribute dont_touch of I13403: signal is true;
	signal I13407: std_logic; attribute dont_touch of I13407: signal is true;
	signal I13410: std_logic; attribute dont_touch of I13410: signal is true;
	signal I13413: std_logic; attribute dont_touch of I13413: signal is true;
	signal I13416: std_logic; attribute dont_touch of I13416: signal is true;
	signal I13419: std_logic; attribute dont_touch of I13419: signal is true;
	signal I13422: std_logic; attribute dont_touch of I13422: signal is true;
	signal I13425: std_logic; attribute dont_touch of I13425: signal is true;
	signal I13428: std_logic; attribute dont_touch of I13428: signal is true;
	signal I13432: std_logic; attribute dont_touch of I13432: signal is true;
	signal I13435: std_logic; attribute dont_touch of I13435: signal is true;
	signal I13438: std_logic; attribute dont_touch of I13438: signal is true;
	signal I13441: std_logic; attribute dont_touch of I13441: signal is true;
	signal I13444: std_logic; attribute dont_touch of I13444: signal is true;
	signal I13447: std_logic; attribute dont_touch of I13447: signal is true;
	signal I13451: std_logic; attribute dont_touch of I13451: signal is true;
	signal I13454: std_logic; attribute dont_touch of I13454: signal is true;
	signal I13457: std_logic; attribute dont_touch of I13457: signal is true;
	signal I13460: std_logic; attribute dont_touch of I13460: signal is true;
	signal I13463: std_logic; attribute dont_touch of I13463: signal is true;
	signal I13466: std_logic; attribute dont_touch of I13466: signal is true;
	signal I13469: std_logic; attribute dont_touch of I13469: signal is true;
	signal I13472: std_logic; attribute dont_touch of I13472: signal is true;
	signal I13475: std_logic; attribute dont_touch of I13475: signal is true;
	signal I13478: std_logic; attribute dont_touch of I13478: signal is true;
	signal I13481: std_logic; attribute dont_touch of I13481: signal is true;
	signal I13484: std_logic; attribute dont_touch of I13484: signal is true;
	signal I13487: std_logic; attribute dont_touch of I13487: signal is true;
	signal I13490: std_logic; attribute dont_touch of I13490: signal is true;
	signal I13493: std_logic; attribute dont_touch of I13493: signal is true;
	signal I13496: std_logic; attribute dont_touch of I13496: signal is true;
	signal I13499: std_logic; attribute dont_touch of I13499: signal is true;
	signal I13502: std_logic; attribute dont_touch of I13502: signal is true;
	signal I13506: std_logic; attribute dont_touch of I13506: signal is true;
	signal I13509: std_logic; attribute dont_touch of I13509: signal is true;
	signal I13512: std_logic; attribute dont_touch of I13512: signal is true;
	signal I13515: std_logic; attribute dont_touch of I13515: signal is true;
	signal I13518: std_logic; attribute dont_touch of I13518: signal is true;
	signal I13524: std_logic; attribute dont_touch of I13524: signal is true;
	signal I13527: std_logic; attribute dont_touch of I13527: signal is true;
	signal I13533: std_logic; attribute dont_touch of I13533: signal is true;
	signal I13537: std_logic; attribute dont_touch of I13537: signal is true;
	signal I13541: std_logic; attribute dont_touch of I13541: signal is true;
	signal I13544: std_logic; attribute dont_touch of I13544: signal is true;
	signal I13547: std_logic; attribute dont_touch of I13547: signal is true;
	signal I13550: std_logic; attribute dont_touch of I13550: signal is true;
	signal I13553: std_logic; attribute dont_touch of I13553: signal is true;
	signal I13559: std_logic; attribute dont_touch of I13559: signal is true;
	signal I13562: std_logic; attribute dont_touch of I13562: signal is true;
	signal I13565: std_logic; attribute dont_touch of I13565: signal is true;
	signal I13570: std_logic; attribute dont_touch of I13570: signal is true;
	signal I13574: std_logic; attribute dont_touch of I13574: signal is true;
	signal I13577: std_logic; attribute dont_touch of I13577: signal is true;
	signal I13580: std_logic; attribute dont_touch of I13580: signal is true;
	signal I13583: std_logic; attribute dont_touch of I13583: signal is true;
	signal I13587: std_logic; attribute dont_touch of I13587: signal is true;
	signal I13588: std_logic; attribute dont_touch of I13588: signal is true;
	signal I13589: std_logic; attribute dont_touch of I13589: signal is true;
	signal I13595: std_logic; attribute dont_touch of I13595: signal is true;
	signal I13598: std_logic; attribute dont_touch of I13598: signal is true;
	signal I13599: std_logic; attribute dont_touch of I13599: signal is true;
	signal I13600: std_logic; attribute dont_touch of I13600: signal is true;
	signal I13605: std_logic; attribute dont_touch of I13605: signal is true;
	signal I13610: std_logic; attribute dont_touch of I13610: signal is true;
	signal I13613: std_logic; attribute dont_touch of I13613: signal is true;
	signal I13617: std_logic; attribute dont_touch of I13617: signal is true;
	signal I13622: std_logic; attribute dont_touch of I13622: signal is true;
	signal I13628: std_logic; attribute dont_touch of I13628: signal is true;
	signal I13631: std_logic; attribute dont_touch of I13631: signal is true;
	signal I13635: std_logic; attribute dont_touch of I13635: signal is true;
	signal I13638: std_logic; attribute dont_touch of I13638: signal is true;
	signal I13639: std_logic; attribute dont_touch of I13639: signal is true;
	signal I13640: std_logic; attribute dont_touch of I13640: signal is true;
	signal I13646: std_logic; attribute dont_touch of I13646: signal is true;
	signal I13649: std_logic; attribute dont_touch of I13649: signal is true;
	signal I13653: std_logic; attribute dont_touch of I13653: signal is true;
	signal I13656: std_logic; attribute dont_touch of I13656: signal is true;
	signal I13659: std_logic; attribute dont_touch of I13659: signal is true;
	signal I13663: std_logic; attribute dont_touch of I13663: signal is true;
	signal I13666: std_logic; attribute dont_touch of I13666: signal is true;
	signal I13669: std_logic; attribute dont_touch of I13669: signal is true;
	signal I13672: std_logic; attribute dont_touch of I13672: signal is true;
	signal I13676: std_logic; attribute dont_touch of I13676: signal is true;
	signal I13679: std_logic; attribute dont_touch of I13679: signal is true;
	signal I13682: std_logic; attribute dont_touch of I13682: signal is true;
	signal I13685: std_logic; attribute dont_touch of I13685: signal is true;
	signal I13686: std_logic; attribute dont_touch of I13686: signal is true;
	signal I13687: std_logic; attribute dont_touch of I13687: signal is true;
	signal I13692: std_logic; attribute dont_touch of I13692: signal is true;
	signal I13695: std_logic; attribute dont_touch of I13695: signal is true;
	signal I13698: std_logic; attribute dont_touch of I13698: signal is true;
	signal I13701: std_logic; attribute dont_touch of I13701: signal is true;
	signal I13704: std_logic; attribute dont_touch of I13704: signal is true;
	signal I13707: std_logic; attribute dont_touch of I13707: signal is true;
	signal I13710: std_logic; attribute dont_touch of I13710: signal is true;
	signal I13713: std_logic; attribute dont_touch of I13713: signal is true;
	signal I13716: std_logic; attribute dont_touch of I13716: signal is true;
	signal I13719: std_logic; attribute dont_touch of I13719: signal is true;
	signal I13722: std_logic; attribute dont_touch of I13722: signal is true;
	signal I13725: std_logic; attribute dont_touch of I13725: signal is true;
	signal I13728: std_logic; attribute dont_touch of I13728: signal is true;
	signal I13731: std_logic; attribute dont_touch of I13731: signal is true;
	signal I13734: std_logic; attribute dont_touch of I13734: signal is true;
	signal I13737: std_logic; attribute dont_touch of I13737: signal is true;
	signal I13740: std_logic; attribute dont_touch of I13740: signal is true;
	signal I13743: std_logic; attribute dont_touch of I13743: signal is true;
	signal I13746: std_logic; attribute dont_touch of I13746: signal is true;
	signal I13749: std_logic; attribute dont_touch of I13749: signal is true;
	signal I13752: std_logic; attribute dont_touch of I13752: signal is true;
	signal I13755: std_logic; attribute dont_touch of I13755: signal is true;
	signal I13758: std_logic; attribute dont_touch of I13758: signal is true;
	signal I13761: std_logic; attribute dont_touch of I13761: signal is true;
	signal I13764: std_logic; attribute dont_touch of I13764: signal is true;
	signal I13767: std_logic; attribute dont_touch of I13767: signal is true;
	signal I13770: std_logic; attribute dont_touch of I13770: signal is true;
	signal I13773: std_logic; attribute dont_touch of I13773: signal is true;
	signal I13776: std_logic; attribute dont_touch of I13776: signal is true;
	signal I13779: std_logic; attribute dont_touch of I13779: signal is true;
	signal I13782: std_logic; attribute dont_touch of I13782: signal is true;
	signal I13785: std_logic; attribute dont_touch of I13785: signal is true;
	signal I13786: std_logic; attribute dont_touch of I13786: signal is true;
	signal I13787: std_logic; attribute dont_touch of I13787: signal is true;
	signal I13794: std_logic; attribute dont_touch of I13794: signal is true;
	signal I13797: std_logic; attribute dont_touch of I13797: signal is true;
	signal I13800: std_logic; attribute dont_touch of I13800: signal is true;
	signal I13801: std_logic; attribute dont_touch of I13801: signal is true;
	signal I13802: std_logic; attribute dont_touch of I13802: signal is true;
	signal I13807: std_logic; attribute dont_touch of I13807: signal is true;
	signal I13810: std_logic; attribute dont_touch of I13810: signal is true;
	signal I13813: std_logic; attribute dont_touch of I13813: signal is true;
	signal I13816: std_logic; attribute dont_touch of I13816: signal is true;
	signal I13819: std_logic; attribute dont_touch of I13819: signal is true;
	signal I13822: std_logic; attribute dont_touch of I13822: signal is true;
	signal I13825: std_logic; attribute dont_touch of I13825: signal is true;
	signal I13828: std_logic; attribute dont_touch of I13828: signal is true;
	signal I13831: std_logic; attribute dont_touch of I13831: signal is true;
	signal I13834: std_logic; attribute dont_touch of I13834: signal is true;
	signal I13837: std_logic; attribute dont_touch of I13837: signal is true;
	signal I13843: std_logic; attribute dont_touch of I13843: signal is true;
	signal I13846: std_logic; attribute dont_touch of I13846: signal is true;
	signal I13850: std_logic; attribute dont_touch of I13850: signal is true;
	signal I13854: std_logic; attribute dont_touch of I13854: signal is true;
	signal I13858: std_logic; attribute dont_touch of I13858: signal is true;
	signal I13861: std_logic; attribute dont_touch of I13861: signal is true;
	signal I13865: std_logic; attribute dont_touch of I13865: signal is true;
	signal I13869: std_logic; attribute dont_touch of I13869: signal is true;
	signal I13873: std_logic; attribute dont_touch of I13873: signal is true;
	signal I13876: std_logic; attribute dont_touch of I13876: signal is true;
	signal I13879: std_logic; attribute dont_touch of I13879: signal is true;
	signal I13882: std_logic; attribute dont_touch of I13882: signal is true;
	signal I13885: std_logic; attribute dont_touch of I13885: signal is true;
	signal I13888: std_logic; attribute dont_touch of I13888: signal is true;
	signal I13891: std_logic; attribute dont_touch of I13891: signal is true;
	signal I13894: std_logic; attribute dont_touch of I13894: signal is true;
	signal I13897: std_logic; attribute dont_touch of I13897: signal is true;
	signal I13900: std_logic; attribute dont_touch of I13900: signal is true;
	signal I13903: std_logic; attribute dont_touch of I13903: signal is true;
	signal I13906: std_logic; attribute dont_touch of I13906: signal is true;
	signal I13909: std_logic; attribute dont_touch of I13909: signal is true;
	signal I13912: std_logic; attribute dont_touch of I13912: signal is true;
	signal I13915: std_logic; attribute dont_touch of I13915: signal is true;
	signal I13918: std_logic; attribute dont_touch of I13918: signal is true;
	signal I13921: std_logic; attribute dont_touch of I13921: signal is true;
	signal I13924: std_logic; attribute dont_touch of I13924: signal is true;
	signal I13927: std_logic; attribute dont_touch of I13927: signal is true;
	signal I13930: std_logic; attribute dont_touch of I13930: signal is true;
	signal I13940: std_logic; attribute dont_touch of I13940: signal is true;
	signal I13956: std_logic; attribute dont_touch of I13956: signal is true;
	signal I13962: std_logic; attribute dont_touch of I13962: signal is true;
	signal I13979: std_logic; attribute dont_touch of I13979: signal is true;
	signal I13997: std_logic; attribute dont_touch of I13997: signal is true;
	signal I14001: std_logic; attribute dont_touch of I14001: signal is true;
	signal I14005: std_logic; attribute dont_touch of I14005: signal is true;
	signal I14009: std_logic; attribute dont_touch of I14009: signal is true;
	signal I14012: std_logic; attribute dont_touch of I14012: signal is true;
	signal I14015: std_logic; attribute dont_touch of I14015: signal is true;
	signal I14019: std_logic; attribute dont_touch of I14019: signal is true;
	signal I14022: std_logic; attribute dont_touch of I14022: signal is true;
	signal I14025: std_logic; attribute dont_touch of I14025: signal is true;
	signal I14028: std_logic; attribute dont_touch of I14028: signal is true;
	signal I14031: std_logic; attribute dont_touch of I14031: signal is true;
	signal I14035: std_logic; attribute dont_touch of I14035: signal is true;
	signal I14039: std_logic; attribute dont_touch of I14039: signal is true;
	signal I14042: std_logic; attribute dont_touch of I14042: signal is true;
	signal I14046: std_logic; attribute dont_touch of I14046: signal is true;
	signal I14049: std_logic; attribute dont_touch of I14049: signal is true;
	signal I14052: std_logic; attribute dont_touch of I14052: signal is true;
	signal I14055: std_logic; attribute dont_touch of I14055: signal is true;
	signal I14058: std_logic; attribute dont_touch of I14058: signal is true;
	signal I14061: std_logic; attribute dont_touch of I14061: signal is true;
	signal I14064: std_logic; attribute dont_touch of I14064: signal is true;
	signal I14067: std_logic; attribute dont_touch of I14067: signal is true;
	signal I14070: std_logic; attribute dont_touch of I14070: signal is true;
	signal I14073: std_logic; attribute dont_touch of I14073: signal is true;
	signal I14076: std_logic; attribute dont_touch of I14076: signal is true;
	signal I14079: std_logic; attribute dont_touch of I14079: signal is true;
	signal I14082: std_logic; attribute dont_touch of I14082: signal is true;
	signal I14085: std_logic; attribute dont_touch of I14085: signal is true;
	signal I14088: std_logic; attribute dont_touch of I14088: signal is true;
	signal I14091: std_logic; attribute dont_touch of I14091: signal is true;
	signal I14094: std_logic; attribute dont_touch of I14094: signal is true;
	signal I14097: std_logic; attribute dont_touch of I14097: signal is true;
	signal I14100: std_logic; attribute dont_touch of I14100: signal is true;
	signal I14103: std_logic; attribute dont_touch of I14103: signal is true;
	signal I14106: std_logic; attribute dont_touch of I14106: signal is true;
	signal I14109: std_logic; attribute dont_touch of I14109: signal is true;
	signal I14112: std_logic; attribute dont_touch of I14112: signal is true;
	signal I14115: std_logic; attribute dont_touch of I14115: signal is true;
	signal I14118: std_logic; attribute dont_touch of I14118: signal is true;
	signal I14121: std_logic; attribute dont_touch of I14121: signal is true;
	signal I14124: std_logic; attribute dont_touch of I14124: signal is true;
	signal I14127: std_logic; attribute dont_touch of I14127: signal is true;
	signal I14130: std_logic; attribute dont_touch of I14130: signal is true;
	signal I14133: std_logic; attribute dont_touch of I14133: signal is true;
	signal I14136: std_logic; attribute dont_touch of I14136: signal is true;
	signal I14139: std_logic; attribute dont_touch of I14139: signal is true;
	signal I14142: std_logic; attribute dont_touch of I14142: signal is true;
	signal I14145: std_logic; attribute dont_touch of I14145: signal is true;
	signal I14148: std_logic; attribute dont_touch of I14148: signal is true;
	signal I14151: std_logic; attribute dont_touch of I14151: signal is true;
	signal I14154: std_logic; attribute dont_touch of I14154: signal is true;
	signal I14157: std_logic; attribute dont_touch of I14157: signal is true;
	signal I14160: std_logic; attribute dont_touch of I14160: signal is true;
	signal I14163: std_logic; attribute dont_touch of I14163: signal is true;
	signal I14166: std_logic; attribute dont_touch of I14166: signal is true;
	signal I14169: std_logic; attribute dont_touch of I14169: signal is true;
	signal I14172: std_logic; attribute dont_touch of I14172: signal is true;
	signal I14175: std_logic; attribute dont_touch of I14175: signal is true;
	signal I14178: std_logic; attribute dont_touch of I14178: signal is true;
	signal I14181: std_logic; attribute dont_touch of I14181: signal is true;
	signal I14184: std_logic; attribute dont_touch of I14184: signal is true;
	signal I14187: std_logic; attribute dont_touch of I14187: signal is true;
	signal I14190: std_logic; attribute dont_touch of I14190: signal is true;
	signal I14193: std_logic; attribute dont_touch of I14193: signal is true;
	signal I14196: std_logic; attribute dont_touch of I14196: signal is true;
	signal I14199: std_logic; attribute dont_touch of I14199: signal is true;
	signal I14202: std_logic; attribute dont_touch of I14202: signal is true;
	signal I14205: std_logic; attribute dont_touch of I14205: signal is true;
	signal I14208: std_logic; attribute dont_touch of I14208: signal is true;
	signal I14211: std_logic; attribute dont_touch of I14211: signal is true;
	signal I14214: std_logic; attribute dont_touch of I14214: signal is true;
	signal I14219: std_logic; attribute dont_touch of I14219: signal is true;
	signal I14224: std_logic; attribute dont_touch of I14224: signal is true;
	signal I14227: std_logic; attribute dont_touch of I14227: signal is true;
	signal I14231: std_logic; attribute dont_touch of I14231: signal is true;
	signal I14234: std_logic; attribute dont_touch of I14234: signal is true;
	signal I14238: std_logic; attribute dont_touch of I14238: signal is true;
	signal I14244: std_logic; attribute dont_touch of I14244: signal is true;
	signal I14245: std_logic; attribute dont_touch of I14245: signal is true;
	signal I14246: std_logic; attribute dont_touch of I14246: signal is true;
	signal I14251: std_logic; attribute dont_touch of I14251: signal is true;
	signal I14257: std_logic; attribute dont_touch of I14257: signal is true;
	signal I14260: std_logic; attribute dont_touch of I14260: signal is true;
	signal I14264: std_logic; attribute dont_touch of I14264: signal is true;
	signal I14267: std_logic; attribute dont_touch of I14267: signal is true;
	signal I14270: std_logic; attribute dont_touch of I14270: signal is true;
	signal I14273: std_logic; attribute dont_touch of I14273: signal is true;
	signal I14276: std_logic; attribute dont_touch of I14276: signal is true;
	signal I14279: std_logic; attribute dont_touch of I14279: signal is true;
	signal I14282: std_logic; attribute dont_touch of I14282: signal is true;
	signal I14285: std_logic; attribute dont_touch of I14285: signal is true;
	signal I14288: std_logic; attribute dont_touch of I14288: signal is true;
	signal I14291: std_logic; attribute dont_touch of I14291: signal is true;
	signal I14294: std_logic; attribute dont_touch of I14294: signal is true;
	signal I14298: std_logic; attribute dont_touch of I14298: signal is true;
	signal I14302: std_logic; attribute dont_touch of I14302: signal is true;
	signal I14305: std_logic; attribute dont_touch of I14305: signal is true;
	signal I14311: std_logic; attribute dont_touch of I14311: signal is true;
	signal I14315: std_logic; attribute dont_touch of I14315: signal is true;
	signal I14318: std_logic; attribute dont_touch of I14318: signal is true;
	signal I14325: std_logic; attribute dont_touch of I14325: signal is true;
	signal I14330: std_logic; attribute dont_touch of I14330: signal is true;
	signal I14334: std_logic; attribute dont_touch of I14334: signal is true;
	signal I14338: std_logic; attribute dont_touch of I14338: signal is true;
	signal I14342: std_logic; attribute dont_touch of I14342: signal is true;
	signal I14349: std_logic; attribute dont_touch of I14349: signal is true;
	signal I14366: std_logic; attribute dont_touch of I14366: signal is true;
	signal I14370: std_logic; attribute dont_touch of I14370: signal is true;
	signal I14374: std_logic; attribute dont_touch of I14374: signal is true;
	signal I14378: std_logic; attribute dont_touch of I14378: signal is true;
	signal I14381: std_logic; attribute dont_touch of I14381: signal is true;
	signal I14388: std_logic; attribute dont_touch of I14388: signal is true;
	signal I14394: std_logic; attribute dont_touch of I14394: signal is true;
	signal I14397: std_logic; attribute dont_touch of I14397: signal is true;
	signal I14400: std_logic; attribute dont_touch of I14400: signal is true;
	signal I14403: std_logic; attribute dont_touch of I14403: signal is true;
	signal I14406: std_logic; attribute dont_touch of I14406: signal is true;
	signal I14410: std_logic; attribute dont_touch of I14410: signal is true;
	signal I14413: std_logic; attribute dont_touch of I14413: signal is true;
	signal I14416: std_logic; attribute dont_touch of I14416: signal is true;
	signal I14420: std_logic; attribute dont_touch of I14420: signal is true;
	signal I14424: std_logic; attribute dont_touch of I14424: signal is true;
	signal I14427: std_logic; attribute dont_touch of I14427: signal is true;
	signal I14430: std_logic; attribute dont_touch of I14430: signal is true;
	signal I14433: std_logic; attribute dont_touch of I14433: signal is true;
	signal I14436: std_logic; attribute dont_touch of I14436: signal is true;
	signal I14439: std_logic; attribute dont_touch of I14439: signal is true;
	signal I14442: std_logic; attribute dont_touch of I14442: signal is true;
	signal I14445: std_logic; attribute dont_touch of I14445: signal is true;
	signal I14448: std_logic; attribute dont_touch of I14448: signal is true;
	signal I14451: std_logic; attribute dont_touch of I14451: signal is true;
	signal I14454: std_logic; attribute dont_touch of I14454: signal is true;
	signal I14457: std_logic; attribute dont_touch of I14457: signal is true;
	signal I14460: std_logic; attribute dont_touch of I14460: signal is true;
	signal I14463: std_logic; attribute dont_touch of I14463: signal is true;
	signal I14467: std_logic; attribute dont_touch of I14467: signal is true;
	signal I14468: std_logic; attribute dont_touch of I14468: signal is true;
	signal I14472: std_logic; attribute dont_touch of I14472: signal is true;
	signal I14473: std_logic; attribute dont_touch of I14473: signal is true;
	signal I14474: std_logic; attribute dont_touch of I14474: signal is true;
	signal I14479: std_logic; attribute dont_touch of I14479: signal is true;
	signal I14480: std_logic; attribute dont_touch of I14480: signal is true;
	signal I14484: std_logic; attribute dont_touch of I14484: signal is true;
	signal I14485: std_logic; attribute dont_touch of I14485: signal is true;
	signal I14489: std_logic; attribute dont_touch of I14489: signal is true;
	signal I14492: std_logic; attribute dont_touch of I14492: signal is true;
	signal I14495: std_logic; attribute dont_touch of I14495: signal is true;
	signal I14496: std_logic; attribute dont_touch of I14496: signal is true;
	signal I14531: std_logic; attribute dont_touch of I14531: signal is true;
	signal I14573: std_logic; attribute dont_touch of I14573: signal is true;
	signal I14603: std_logic; attribute dont_touch of I14603: signal is true;
	signal I14614: std_logic; attribute dont_touch of I14614: signal is true;
	signal I14623: std_logic; attribute dont_touch of I14623: signal is true;
	signal I14637: std_logic; attribute dont_touch of I14637: signal is true;
	signal I14643: std_logic; attribute dont_touch of I14643: signal is true;
	signal I14646: std_logic; attribute dont_touch of I14646: signal is true;
	signal I14657: std_logic; attribute dont_touch of I14657: signal is true;
	signal I14662: std_logic; attribute dont_touch of I14662: signal is true;
	signal I14668: std_logic; attribute dont_touch of I14668: signal is true;
	signal I14674: std_logic; attribute dont_touch of I14674: signal is true;
	signal I14677: std_logic; attribute dont_touch of I14677: signal is true;
	signal I14680: std_logic; attribute dont_touch of I14680: signal is true;
	signal I14683: std_logic; attribute dont_touch of I14683: signal is true;
	signal I14687: std_logic; attribute dont_touch of I14687: signal is true;
	signal I14695: std_logic; attribute dont_touch of I14695: signal is true;
	signal I14709: std_logic; attribute dont_touch of I14709: signal is true;
	signal I14712: std_logic; attribute dont_touch of I14712: signal is true;
	signal I14718: std_logic; attribute dont_touch of I14718: signal is true;
	signal I14722: std_logic; attribute dont_touch of I14722: signal is true;
	signal I14725: std_logic; attribute dont_touch of I14725: signal is true;
	signal I14728: std_logic; attribute dont_touch of I14728: signal is true;
	signal I14732: std_logic; attribute dont_touch of I14732: signal is true;
	signal I14739: std_logic; attribute dont_touch of I14739: signal is true;
	signal I14743: std_logic; attribute dont_touch of I14743: signal is true;
	signal I14747: std_logic; attribute dont_touch of I14747: signal is true;
	signal I14753: std_logic; attribute dont_touch of I14753: signal is true;
	signal I14754: std_logic; attribute dont_touch of I14754: signal is true;
	signal I14758: std_logic; attribute dont_touch of I14758: signal is true;
	signal I14759: std_logic; attribute dont_touch of I14759: signal is true;
	signal I14763: std_logic; attribute dont_touch of I14763: signal is true;
	signal I14766: std_logic; attribute dont_touch of I14766: signal is true;
	signal I14767: std_logic; attribute dont_touch of I14767: signal is true;
	signal I14771: std_logic; attribute dont_touch of I14771: signal is true;
	signal I14772: std_logic; attribute dont_touch of I14772: signal is true;
	signal I14777: std_logic; attribute dont_touch of I14777: signal is true;
	signal I14780: std_logic; attribute dont_touch of I14780: signal is true;
	signal I14783: std_logic; attribute dont_touch of I14783: signal is true;
	signal I14786: std_logic; attribute dont_touch of I14786: signal is true;
	signal I14789: std_logic; attribute dont_touch of I14789: signal is true;
	signal I14792: std_logic; attribute dont_touch of I14792: signal is true;
	signal I14795: std_logic; attribute dont_touch of I14795: signal is true;
	signal I14798: std_logic; attribute dont_touch of I14798: signal is true;
	signal I14801: std_logic; attribute dont_touch of I14801: signal is true;
	signal I14804: std_logic; attribute dont_touch of I14804: signal is true;
	signal I14807: std_logic; attribute dont_touch of I14807: signal is true;
	signal I14810: std_logic; attribute dont_touch of I14810: signal is true;
	signal I14813: std_logic; attribute dont_touch of I14813: signal is true;
	signal I14816: std_logic; attribute dont_touch of I14816: signal is true;
	signal I14819: std_logic; attribute dont_touch of I14819: signal is true;
	signal I14822: std_logic; attribute dont_touch of I14822: signal is true;
	signal I14825: std_logic; attribute dont_touch of I14825: signal is true;
	signal I14828: std_logic; attribute dont_touch of I14828: signal is true;
	signal I14831: std_logic; attribute dont_touch of I14831: signal is true;
	signal I14834: std_logic; attribute dont_touch of I14834: signal is true;
	signal I14837: std_logic; attribute dont_touch of I14837: signal is true;
	signal I14838: std_logic; attribute dont_touch of I14838: signal is true;
	signal I14839: std_logic; attribute dont_touch of I14839: signal is true;
	signal I14844: std_logic; attribute dont_touch of I14844: signal is true;
	signal I14848: std_logic; attribute dont_touch of I14848: signal is true;
	signal I14851: std_logic; attribute dont_touch of I14851: signal is true;
	signal I14857: std_logic; attribute dont_touch of I14857: signal is true;
	signal I14904: std_logic; attribute dont_touch of I14904: signal is true;
	signal I14925: std_logic; attribute dont_touch of I14925: signal is true;
	signal I14932: std_logic; attribute dont_touch of I14932: signal is true;
	signal I14933: std_logic; attribute dont_touch of I14933: signal is true;
	signal I14941: std_logic; attribute dont_touch of I14941: signal is true;
	signal I14942: std_logic; attribute dont_touch of I14942: signal is true;
	signal I14951: std_logic; attribute dont_touch of I14951: signal is true;
	signal I14952: std_logic; attribute dont_touch of I14952: signal is true;
	signal I14959: std_logic; attribute dont_touch of I14959: signal is true;
	signal I14960: std_logic; attribute dont_touch of I14960: signal is true;
	signal I14964: std_logic; attribute dont_touch of I14964: signal is true;
	signal I14969: std_logic; attribute dont_touch of I14969: signal is true;
	signal I14970: std_logic; attribute dont_touch of I14970: signal is true;
	signal I14974: std_logic; attribute dont_touch of I14974: signal is true;
	signal I14980: std_logic; attribute dont_touch of I14980: signal is true;
	signal I14985: std_logic; attribute dont_touch of I14985: signal is true;
	signal I14990: std_logic; attribute dont_touch of I14990: signal is true;
	signal I14996: std_logic; attribute dont_touch of I14996: signal is true;
	signal I15003: std_logic; attribute dont_touch of I15003: signal is true;
	signal I15007: std_logic; attribute dont_touch of I15007: signal is true;
	signal I15010: std_logic; attribute dont_touch of I15010: signal is true;
	signal I15014: std_logic; attribute dont_touch of I15014: signal is true;
	signal I15017: std_logic; attribute dont_touch of I15017: signal is true;
	signal I15018: std_logic; attribute dont_touch of I15018: signal is true;
	signal I15019: std_logic; attribute dont_touch of I15019: signal is true;
	signal I15020: std_logic; attribute dont_touch of I15020: signal is true;
	signal I15021: std_logic; attribute dont_touch of I15021: signal is true;
	signal I15029: std_logic; attribute dont_touch of I15029: signal is true;
	signal I15030: std_logic; attribute dont_touch of I15030: signal is true;
	signal I15031: std_logic; attribute dont_touch of I15031: signal is true;
	signal I15032: std_logic; attribute dont_touch of I15032: signal is true;
	signal I15033: std_logic; attribute dont_touch of I15033: signal is true;
	signal I15040: std_logic; attribute dont_touch of I15040: signal is true;
	signal I15041: std_logic; attribute dont_touch of I15041: signal is true;
	signal I15042: std_logic; attribute dont_touch of I15042: signal is true;
	signal I15043: std_logic; attribute dont_touch of I15043: signal is true;
	signal I15044: std_logic; attribute dont_touch of I15044: signal is true;
	signal I15051: std_logic; attribute dont_touch of I15051: signal is true;
	signal I15052: std_logic; attribute dont_touch of I15052: signal is true;
	signal I15053: std_logic; attribute dont_touch of I15053: signal is true;
	signal I15054: std_logic; attribute dont_touch of I15054: signal is true;
	signal I15055: std_logic; attribute dont_touch of I15055: signal is true;
	signal I15062: std_logic; attribute dont_touch of I15062: signal is true;
	signal I15065: std_logic; attribute dont_touch of I15065: signal is true;
	signal I15068: std_logic; attribute dont_touch of I15068: signal is true;
	signal I15071: std_logic; attribute dont_touch of I15071: signal is true;
	signal I15072: std_logic; attribute dont_touch of I15072: signal is true;
	signal I15073: std_logic; attribute dont_touch of I15073: signal is true;
	signal I15074: std_logic; attribute dont_touch of I15074: signal is true;
	signal I15075: std_logic; attribute dont_touch of I15075: signal is true;
	signal I15082: std_logic; attribute dont_touch of I15082: signal is true;
	signal I15083: std_logic; attribute dont_touch of I15083: signal is true;
	signal I15084: std_logic; attribute dont_touch of I15084: signal is true;
	signal I15085: std_logic; attribute dont_touch of I15085: signal is true;
	signal I15086: std_logic; attribute dont_touch of I15086: signal is true;
	signal I15098: std_logic; attribute dont_touch of I15098: signal is true;
	signal I15099: std_logic; attribute dont_touch of I15099: signal is true;
	signal I15100: std_logic; attribute dont_touch of I15100: signal is true;
	signal I15101: std_logic; attribute dont_touch of I15101: signal is true;
	signal I15102: std_logic; attribute dont_touch of I15102: signal is true;
	signal I15109: std_logic; attribute dont_touch of I15109: signal is true;
	signal I15110: std_logic; attribute dont_touch of I15110: signal is true;
	signal I15111: std_logic; attribute dont_touch of I15111: signal is true;
	signal I15112: std_logic; attribute dont_touch of I15112: signal is true;
	signal I15113: std_logic; attribute dont_touch of I15113: signal is true;
	signal I15147: std_logic; attribute dont_touch of I15147: signal is true;
	signal I15152: std_logic; attribute dont_touch of I15152: signal is true;
	signal I15160: std_logic; attribute dont_touch of I15160: signal is true;
	signal I15165: std_logic; attribute dont_touch of I15165: signal is true;
	signal I15169: std_logic; attribute dont_touch of I15169: signal is true;
	signal I15172: std_logic; attribute dont_touch of I15172: signal is true;
	signal I15175: std_logic; attribute dont_touch of I15175: signal is true;
	signal I15178: std_logic; attribute dont_touch of I15178: signal is true;
	signal I15181: std_logic; attribute dont_touch of I15181: signal is true;
	signal I15184: std_logic; attribute dont_touch of I15184: signal is true;
	signal I15187: std_logic; attribute dont_touch of I15187: signal is true;
	signal I15190: std_logic; attribute dont_touch of I15190: signal is true;
	signal I15193: std_logic; attribute dont_touch of I15193: signal is true;
	signal I15196: std_logic; attribute dont_touch of I15196: signal is true;
	signal I15199: std_logic; attribute dont_touch of I15199: signal is true;
	signal I15202: std_logic; attribute dont_touch of I15202: signal is true;
	signal I15205: std_logic; attribute dont_touch of I15205: signal is true;
	signal I15208: std_logic; attribute dont_touch of I15208: signal is true;
	signal I15211: std_logic; attribute dont_touch of I15211: signal is true;
	signal I15218: std_logic; attribute dont_touch of I15218: signal is true;
	signal I15222: std_logic; attribute dont_touch of I15222: signal is true;
	signal I15225: std_logic; attribute dont_touch of I15225: signal is true;
	signal I15228: std_logic; attribute dont_touch of I15228: signal is true;
	signal I15229: std_logic; attribute dont_touch of I15229: signal is true;
	signal I15230: std_logic; attribute dont_touch of I15230: signal is true;
	signal I15231: std_logic; attribute dont_touch of I15231: signal is true;
	signal I15232: std_logic; attribute dont_touch of I15232: signal is true;
	signal I15239: std_logic; attribute dont_touch of I15239: signal is true;
	signal I15240: std_logic; attribute dont_touch of I15240: signal is true;
	signal I15241: std_logic; attribute dont_touch of I15241: signal is true;
	signal I15242: std_logic; attribute dont_touch of I15242: signal is true;
	signal I15243: std_logic; attribute dont_touch of I15243: signal is true;
	signal I15250: std_logic; attribute dont_touch of I15250: signal is true;
	signal I15251: std_logic; attribute dont_touch of I15251: signal is true;
	signal I15252: std_logic; attribute dont_touch of I15252: signal is true;
	signal I15253: std_logic; attribute dont_touch of I15253: signal is true;
	signal I15254: std_logic; attribute dont_touch of I15254: signal is true;
	signal I15261: std_logic; attribute dont_touch of I15261: signal is true;
	signal I15262: std_logic; attribute dont_touch of I15262: signal is true;
	signal I15263: std_logic; attribute dont_touch of I15263: signal is true;
	signal I15264: std_logic; attribute dont_touch of I15264: signal is true;
	signal I15265: std_logic; attribute dont_touch of I15265: signal is true;
	signal I15272: std_logic; attribute dont_touch of I15272: signal is true;
	signal I15273: std_logic; attribute dont_touch of I15273: signal is true;
	signal I15274: std_logic; attribute dont_touch of I15274: signal is true;
	signal I15275: std_logic; attribute dont_touch of I15275: signal is true;
	signal I15276: std_logic; attribute dont_touch of I15276: signal is true;
	signal I15283: std_logic; attribute dont_touch of I15283: signal is true;
	signal I15284: std_logic; attribute dont_touch of I15284: signal is true;
	signal I15285: std_logic; attribute dont_touch of I15285: signal is true;
	signal I15290: std_logic; attribute dont_touch of I15290: signal is true;
	signal I15291: std_logic; attribute dont_touch of I15291: signal is true;
	signal I15292: std_logic; attribute dont_touch of I15292: signal is true;
	signal I15297: std_logic; attribute dont_touch of I15297: signal is true;
	signal I15298: std_logic; attribute dont_touch of I15298: signal is true;
	signal I15308: std_logic; attribute dont_touch of I15308: signal is true;
	signal I15315: std_logic; attribute dont_touch of I15315: signal is true;
	signal I15324: std_logic; attribute dont_touch of I15324: signal is true;
	signal I15329: std_logic; attribute dont_touch of I15329: signal is true;
	signal I15334: std_logic; attribute dont_touch of I15334: signal is true;
	signal I15337: std_logic; attribute dont_touch of I15337: signal is true;
	signal I15340: std_logic; attribute dont_touch of I15340: signal is true;
	signal I15379: std_logic; attribute dont_touch of I15379: signal is true;
	signal I15382: std_logic; attribute dont_touch of I15382: signal is true;
	signal I15385: std_logic; attribute dont_touch of I15385: signal is true;
	signal I15388: std_logic; attribute dont_touch of I15388: signal is true;
	signal I15391: std_logic; attribute dont_touch of I15391: signal is true;
	signal I15394: std_logic; attribute dont_touch of I15394: signal is true;
	signal I15400: std_logic; attribute dont_touch of I15400: signal is true;
	signal I15405: std_logic; attribute dont_touch of I15405: signal is true;
	signal I15408: std_logic; attribute dont_touch of I15408: signal is true;
	signal I15411: std_logic; attribute dont_touch of I15411: signal is true;
	signal I15414: std_logic; attribute dont_touch of I15414: signal is true;
	signal I15417: std_logic; attribute dont_touch of I15417: signal is true;
	signal I15420: std_logic; attribute dont_touch of I15420: signal is true;
	signal I15423: std_logic; attribute dont_touch of I15423: signal is true;
	signal I15426: std_logic; attribute dont_touch of I15426: signal is true;
	signal I15429: std_logic; attribute dont_touch of I15429: signal is true;
	signal I15433: std_logic; attribute dont_touch of I15433: signal is true;
	signal I15475: std_logic; attribute dont_touch of I15475: signal is true;
	signal I15478: std_logic; attribute dont_touch of I15478: signal is true;
	signal I15481: std_logic; attribute dont_touch of I15481: signal is true;
	signal I15484: std_logic; attribute dont_touch of I15484: signal is true;
	signal I15492: std_logic; attribute dont_touch of I15492: signal is true;
	signal I15495: std_logic; attribute dont_touch of I15495: signal is true;
	signal I15498: std_logic; attribute dont_touch of I15498: signal is true;
	signal I15501: std_logic; attribute dont_touch of I15501: signal is true;
	signal I15504: std_logic; attribute dont_touch of I15504: signal is true;
	signal I15507: std_logic; attribute dont_touch of I15507: signal is true;
	signal I15510: std_logic; attribute dont_touch of I15510: signal is true;
	signal I15513: std_logic; attribute dont_touch of I15513: signal is true;
	signal I15516: std_logic; attribute dont_touch of I15516: signal is true;
	signal I15519: std_logic; attribute dont_touch of I15519: signal is true;
	signal I15522: std_logic; attribute dont_touch of I15522: signal is true;
	signal I15527: std_logic; attribute dont_touch of I15527: signal is true;
	signal I15530: std_logic; attribute dont_touch of I15530: signal is true;
	signal I15533: std_logic; attribute dont_touch of I15533: signal is true;
	signal I15536: std_logic; attribute dont_touch of I15536: signal is true;
	signal I15539: std_logic; attribute dont_touch of I15539: signal is true;
	signal I15543: std_logic; attribute dont_touch of I15543: signal is true;
	signal I15546: std_logic; attribute dont_touch of I15546: signal is true;
	signal I15550: std_logic; attribute dont_touch of I15550: signal is true;
	signal I15553: std_logic; attribute dont_touch of I15553: signal is true;
	signal I15557: std_logic; attribute dont_touch of I15557: signal is true;
	signal I15562: std_logic; attribute dont_touch of I15562: signal is true;
	signal I15565: std_logic; attribute dont_touch of I15565: signal is true;
	signal I15568: std_logic; attribute dont_touch of I15568: signal is true;
	signal I15571: std_logic; attribute dont_touch of I15571: signal is true;
	signal I15574: std_logic; attribute dont_touch of I15574: signal is true;
	signal I15577: std_logic; attribute dont_touch of I15577: signal is true;
	signal I15580: std_logic; attribute dont_touch of I15580: signal is true;
	signal I15583: std_logic; attribute dont_touch of I15583: signal is true;
	signal I15586: std_logic; attribute dont_touch of I15586: signal is true;
	signal I15589: std_logic; attribute dont_touch of I15589: signal is true;
	signal I15592: std_logic; attribute dont_touch of I15592: signal is true;
	signal I15595: std_logic; attribute dont_touch of I15595: signal is true;
	signal I15598: std_logic; attribute dont_touch of I15598: signal is true;
	signal I15601: std_logic; attribute dont_touch of I15601: signal is true;
	signal I15604: std_logic; attribute dont_touch of I15604: signal is true;
	signal I15607: std_logic; attribute dont_touch of I15607: signal is true;
	signal I15610: std_logic; attribute dont_touch of I15610: signal is true;
	signal I15613: std_logic; attribute dont_touch of I15613: signal is true;
	signal I15616: std_logic; attribute dont_touch of I15616: signal is true;
	signal I15619: std_logic; attribute dont_touch of I15619: signal is true;
	signal I15622: std_logic; attribute dont_touch of I15622: signal is true;
	signal I15625: std_logic; attribute dont_touch of I15625: signal is true;
	signal I15628: std_logic; attribute dont_touch of I15628: signal is true;
	signal I15631: std_logic; attribute dont_touch of I15631: signal is true;
	signal I15635: std_logic; attribute dont_touch of I15635: signal is true;
	signal I15638: std_logic; attribute dont_touch of I15638: signal is true;
	signal I15641: std_logic; attribute dont_touch of I15641: signal is true;
	signal I15645: std_logic; attribute dont_touch of I15645: signal is true;
	signal I15648: std_logic; attribute dont_touch of I15648: signal is true;
	signal I15651: std_logic; attribute dont_touch of I15651: signal is true;
	signal I15654: std_logic; attribute dont_touch of I15654: signal is true;
	signal I15657: std_logic; attribute dont_touch of I15657: signal is true;
	signal I15660: std_logic; attribute dont_touch of I15660: signal is true;
	signal I15663: std_logic; attribute dont_touch of I15663: signal is true;
	signal I15666: std_logic; attribute dont_touch of I15666: signal is true;
	signal I15669: std_logic; attribute dont_touch of I15669: signal is true;
	signal I15672: std_logic; attribute dont_touch of I15672: signal is true;
	signal I15675: std_logic; attribute dont_touch of I15675: signal is true;
	signal I15678: std_logic; attribute dont_touch of I15678: signal is true;
	signal I15681: std_logic; attribute dont_touch of I15681: signal is true;
	signal I15684: std_logic; attribute dont_touch of I15684: signal is true;
	signal I15687: std_logic; attribute dont_touch of I15687: signal is true;
	signal I15690: std_logic; attribute dont_touch of I15690: signal is true;
	signal I15693: std_logic; attribute dont_touch of I15693: signal is true;
	signal I15696: std_logic; attribute dont_touch of I15696: signal is true;
	signal I15699: std_logic; attribute dont_touch of I15699: signal is true;
	signal I15702: std_logic; attribute dont_touch of I15702: signal is true;
	signal I15705: std_logic; attribute dont_touch of I15705: signal is true;
	signal I15708: std_logic; attribute dont_touch of I15708: signal is true;
	signal I15711: std_logic; attribute dont_touch of I15711: signal is true;
	signal I15714: std_logic; attribute dont_touch of I15714: signal is true;
	signal I15717: std_logic; attribute dont_touch of I15717: signal is true;
	signal I15720: std_logic; attribute dont_touch of I15720: signal is true;
	signal I15723: std_logic; attribute dont_touch of I15723: signal is true;
	signal I15726: std_logic; attribute dont_touch of I15726: signal is true;
	signal I15729: std_logic; attribute dont_touch of I15729: signal is true;
	signal I15732: std_logic; attribute dont_touch of I15732: signal is true;
	signal I15735: std_logic; attribute dont_touch of I15735: signal is true;
	signal I15738: std_logic; attribute dont_touch of I15738: signal is true;
	signal I15741: std_logic; attribute dont_touch of I15741: signal is true;
	signal I15747: std_logic; attribute dont_touch of I15747: signal is true;
	signal I15753: std_logic; attribute dont_touch of I15753: signal is true;
	signal I15756: std_logic; attribute dont_touch of I15756: signal is true;
	signal I15759: std_logic; attribute dont_touch of I15759: signal is true;
	signal I15762: std_logic; attribute dont_touch of I15762: signal is true;
	signal I15765: std_logic; attribute dont_touch of I15765: signal is true;
	signal I15770: std_logic; attribute dont_touch of I15770: signal is true;
	signal I15773: std_logic; attribute dont_touch of I15773: signal is true;
	signal I15776: std_logic; attribute dont_touch of I15776: signal is true;
	signal I15784: std_logic; attribute dont_touch of I15784: signal is true;
	signal I15791: std_logic; attribute dont_touch of I15791: signal is true;
	signal I15803: std_logic; attribute dont_touch of I15803: signal is true;
	signal I15811: std_logic; attribute dont_touch of I15811: signal is true;
	signal I15814: std_logic; attribute dont_touch of I15814: signal is true;
	signal I15817: std_logic; attribute dont_touch of I15817: signal is true;
	signal I15818: std_logic; attribute dont_touch of I15818: signal is true;
	signal I15819: std_logic; attribute dont_touch of I15819: signal is true;
	signal I15824: std_logic; attribute dont_touch of I15824: signal is true;
	signal I15830: std_logic; attribute dont_touch of I15830: signal is true;
	signal I15833: std_logic; attribute dont_touch of I15833: signal is true;
	signal I15836: std_logic; attribute dont_touch of I15836: signal is true;
	signal I15839: std_logic; attribute dont_touch of I15839: signal is true;
	signal I15842: std_logic; attribute dont_touch of I15842: signal is true;
	signal I15845: std_logic; attribute dont_touch of I15845: signal is true;
	signal I15848: std_logic; attribute dont_touch of I15848: signal is true;
	signal I15849: std_logic; attribute dont_touch of I15849: signal is true;
	signal I15850: std_logic; attribute dont_touch of I15850: signal is true;
	signal I15855: std_logic; attribute dont_touch of I15855: signal is true;
	signal I15856: std_logic; attribute dont_touch of I15856: signal is true;
	signal I15857: std_logic; attribute dont_touch of I15857: signal is true;
	signal I15862: std_logic; attribute dont_touch of I15862: signal is true;
	signal I15863: std_logic; attribute dont_touch of I15863: signal is true;
	signal I15864: std_logic; attribute dont_touch of I15864: signal is true;
	signal I15871: std_logic; attribute dont_touch of I15871: signal is true;
	signal I15880: std_logic; attribute dont_touch of I15880: signal is true;
	signal I15881: std_logic; attribute dont_touch of I15881: signal is true;
	signal I15882: std_logic; attribute dont_touch of I15882: signal is true;
	signal I15887: std_logic; attribute dont_touch of I15887: signal is true;
	signal I15888: std_logic; attribute dont_touch of I15888: signal is true;
	signal I15889: std_logic; attribute dont_touch of I15889: signal is true;
	signal I15894: std_logic; attribute dont_touch of I15894: signal is true;
	signal I15897: std_logic; attribute dont_touch of I15897: signal is true;
	signal I15898: std_logic; attribute dont_touch of I15898: signal is true;
	signal I15899: std_logic; attribute dont_touch of I15899: signal is true;
	signal I15909: std_logic; attribute dont_touch of I15909: signal is true;
	signal I15912: std_logic; attribute dont_touch of I15912: signal is true;
	signal I15915: std_logic; attribute dont_touch of I15915: signal is true;
	signal I15918: std_logic; attribute dont_touch of I15918: signal is true;
	signal I15921: std_logic; attribute dont_touch of I15921: signal is true;
	signal I15924: std_logic; attribute dont_touch of I15924: signal is true;
	signal I15927: std_logic; attribute dont_touch of I15927: signal is true;
	signal I15930: std_logic; attribute dont_touch of I15930: signal is true;
	signal I15933: std_logic; attribute dont_touch of I15933: signal is true;
	signal I15937: std_logic; attribute dont_touch of I15937: signal is true;
	signal I15940: std_logic; attribute dont_touch of I15940: signal is true;
	signal I15943: std_logic; attribute dont_touch of I15943: signal is true;
	signal I15947: std_logic; attribute dont_touch of I15947: signal is true;
	signal I15950: std_logic; attribute dont_touch of I15950: signal is true;
	signal I15953: std_logic; attribute dont_touch of I15953: signal is true;
	signal I15956: std_logic; attribute dont_touch of I15956: signal is true;
	signal I15959: std_logic; attribute dont_touch of I15959: signal is true;
	signal I15962: std_logic; attribute dont_touch of I15962: signal is true;
	signal I15965: std_logic; attribute dont_touch of I15965: signal is true;
	signal I15971: std_logic; attribute dont_touch of I15971: signal is true;
	signal I15974: std_logic; attribute dont_touch of I15974: signal is true;
	signal I15978: std_logic; attribute dont_touch of I15978: signal is true;
	signal I15982: std_logic; attribute dont_touch of I15982: signal is true;
	signal I15985: std_logic; attribute dont_touch of I15985: signal is true;
	signal I15990: std_logic; attribute dont_touch of I15990: signal is true;
	signal I16006: std_logic; attribute dont_touch of I16006: signal is true;
	signal I16009: std_logic; attribute dont_touch of I16009: signal is true;
	signal I16017: std_logic; attribute dont_touch of I16017: signal is true;
	signal I16020: std_logic; attribute dont_touch of I16020: signal is true;
	signal I16023: std_logic; attribute dont_touch of I16023: signal is true;
	signal I16026: std_logic; attribute dont_touch of I16026: signal is true;
	signal I16033: std_logic; attribute dont_touch of I16033: signal is true;
	signal I16036: std_logic; attribute dont_touch of I16036: signal is true;
	signal I16040: std_logic; attribute dont_touch of I16040: signal is true;
	signal I16043: std_logic; attribute dont_touch of I16043: signal is true;
	signal I16046: std_logic; attribute dont_touch of I16046: signal is true;
	signal I16049: std_logic; attribute dont_touch of I16049: signal is true;
	signal I16052: std_logic; attribute dont_touch of I16052: signal is true;
	signal I16055: std_logic; attribute dont_touch of I16055: signal is true;
	signal I16058: std_logic; attribute dont_touch of I16058: signal is true;
	signal I16061: std_logic; attribute dont_touch of I16061: signal is true;
	signal I16072: std_logic; attribute dont_touch of I16072: signal is true;
	signal I16084: std_logic; attribute dont_touch of I16084: signal is true;
	signal I16090: std_logic; attribute dont_touch of I16090: signal is true;
	signal I16100: std_logic; attribute dont_touch of I16100: signal is true;
	signal I16103: std_logic; attribute dont_touch of I16103: signal is true;
	signal I16107: std_logic; attribute dont_touch of I16107: signal is true;
	signal I16116: std_logic; attribute dont_touch of I16116: signal is true;
	signal I16119: std_logic; attribute dont_touch of I16119: signal is true;
	signal I16122: std_logic; attribute dont_touch of I16122: signal is true;
	signal I16126: std_logic; attribute dont_touch of I16126: signal is true;
	signal I16129: std_logic; attribute dont_touch of I16129: signal is true;
	signal I16132: std_logic; attribute dont_touch of I16132: signal is true;
	signal I16135: std_logic; attribute dont_touch of I16135: signal is true;
	signal I16138: std_logic; attribute dont_touch of I16138: signal is true;
	signal I16142: std_logic; attribute dont_touch of I16142: signal is true;
	signal I16145: std_logic; attribute dont_touch of I16145: signal is true;
	signal I16148: std_logic; attribute dont_touch of I16148: signal is true;
	signal I16151: std_logic; attribute dont_touch of I16151: signal is true;
	signal I16154: std_logic; attribute dont_touch of I16154: signal is true;
	signal I16158: std_logic; attribute dont_touch of I16158: signal is true;
	signal I16161: std_logic; attribute dont_touch of I16161: signal is true;
	signal I16165: std_logic; attribute dont_touch of I16165: signal is true;
	signal I16168: std_logic; attribute dont_touch of I16168: signal is true;
	signal I16173: std_logic; attribute dont_touch of I16173: signal is true;
	signal I16176: std_logic; attribute dont_touch of I16176: signal is true;
	signal I16180: std_logic; attribute dont_touch of I16180: signal is true;
	signal I16183: std_logic; attribute dont_touch of I16183: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			G2<=G9361;
			G3<=G9360;
			G4<=G9372;
			G5<=G9373;
			G6<=G9374;
			G7<=G9375;
			G8<=G9376;
			G12<=G8662;
			G13<=G7308;
			G16<=G1404;
			G20<=G6386;
			G33<=G5184;
			G38<=G5746;
			G46<=G8955;
			G47<=G9389;
			G48<=G9362;
			G52<=G6781;
			G55<=G7733;
			G58<=G7734;
			G62<=G7509;
			G65<=G4598;
			G68<=G6774;
			G71<=G6775;
			G74<=G6776;
			G77<=G6777;
			G80<=G6778;
			G83<=G6779;
			G86<=G6780;
			G89<=G92;
			G92<=G6794;
			G93<=G5145;
			G94<=G6782;
			G95<=G94;
			G98<=G5146;
			G99<=G6783;
			G100<=G99;
			G103<=G5157;
			G104<=G6784;
			G105<=G104;
			G108<=G5147;
			G109<=G6785;
			G110<=G109;
			G113<=G5148;
			G114<=G6786;
			G117<=G5153;
			G118<=G6787;
			G121<=G5154;
			G122<=G6788;
			G125<=G5155;
			G126<=G6789;
			G129<=G5156;
			G130<=G6790;
			G133<=G5149;
			G134<=G6791;
			G137<=G5150;
			G138<=G6792;
			G141<=G5151;
			G142<=G6793;
			G145<=G5152;
			G146<=G7735;
			G150<=G7738;
			G154<=G7739;
			G158<=G7740;
			G162<=G7741;
			G168<=G7742;
			G172<=G1270;
			G173<=G7736;
			G174<=G7737;
			G179<=G5159;
			G180<=G5158;
			G181<=G5160;
			G182<=G5161;
			G183<=G6309;
			G184<=G6310;
			G185<=G4599;
			G186<=G3830;
			G187<=G5730;
			G190<=G201;
			G195<=G3831;
			G196<=G5731;
			G199<=G3832;
			G200<=G199;
			G201<=G200;
			G202<=G5732;
			G205<=G3835;
			G207<=G5733;
			G210<=G3834;
			G211<=G4600;
			G212<=G4601;
			G213<=G4602;
			G214<=G4603;
			G215<=G4604;
			G216<=G6311;
			G219<=G6312;
			G222<=G6313;
			G225<=G6314;
			G228<=G6315;
			G231<=G4605;
			G232<=G4606;
			G233<=G4607;
			G234<=G4608;
			G235<=G4609;
			G236<=G4610;
			G237<=G6316;
			G240<=G6317;
			G243<=G6318;
			G246<=G6319;
			G249<=G6320;
			G252<=G6321;
			G255<=G9087;
			G258<=G9088;
			G261<=G9089;
			G264<=G9090;
			G267<=G9091;
			G270<=G9092;
			G273<=G4611;
			G274<=G4612;
			G275<=G6322;
			G278<=G6323;
			G281<=G9085;
			G284<=G9086;
			G287<=G3836;
			G290<=G287;
			G292<=G4613;
			G293<=G4614;
			G294<=G4615;
			G295<=G4616;
			G296<=G4617;
			G297<=G6324;
			G300<=G6325;
			G303<=G6326;
			G306<=G6327;
			G309<=G6328;
			G312<=G4618;
			G313<=G4619;
			G314<=G4620;
			G315<=G4621;
			G316<=G4622;
			G317<=G4623;
			G318<=G6329;
			G321<=G6330;
			G324<=G6331;
			G327<=G6332;
			G330<=G6333;
			G333<=G6334;
			G336<=G9095;
			G339<=G9096;
			G342<=G9097;
			G345<=G9098;
			G348<=G9099;
			G351<=G9100;
			G354<=G4624;
			G355<=G4625;
			G356<=G6335;
			G359<=G6336;
			G362<=G9093;
			G365<=G9094;
			G368<=G3838;
			G371<=G368;
			G373<=G4626;
			G374<=G4627;
			G375<=G4628;
			G376<=G4629;
			G377<=G4630;
			G378<=G6337;
			G381<=G6338;
			G384<=G6339;
			G387<=G6340;
			G390<=G6341;
			G393<=G4631;
			G394<=G4632;
			G395<=G4633;
			G396<=G4634;
			G397<=G4635;
			G398<=G4636;
			G399<=G6342;
			G402<=G6343;
			G405<=G6344;
			G408<=G6345;
			G411<=G6346;
			G414<=G6347;
			G417<=G9103;
			G420<=G9104;
			G423<=G9105;
			G426<=G9106;
			G429<=G9107;
			G432<=G9108;
			G435<=G4637;
			G436<=G4638;
			G437<=G6348;
			G440<=G6349;
			G443<=G9101;
			G446<=G9102;
			G449<=G3840;
			G452<=G449;
			G454<=G4639;
			G455<=G4640;
			G456<=G4641;
			G457<=G4642;
			G458<=G4643;
			G459<=G6350;
			G462<=G6351;
			G465<=G6352;
			G468<=G6353;
			G471<=G6354;
			G474<=G4644;
			G475<=G4645;
			G476<=G4646;
			G477<=G4647;
			G478<=G4648;
			G479<=G4649;
			G480<=G6355;
			G483<=G6356;
			G486<=G6357;
			G489<=G6358;
			G492<=G6359;
			G495<=G6360;
			G498<=G9111;
			G501<=G9112;
			G504<=G9113;
			G507<=G9114;
			G510<=G9115;
			G513<=G9116;
			G516<=G4650;
			G517<=G4651;
			G518<=G6361;
			G521<=G6362;
			G524<=G9109;
			G527<=G9110;
			G530<=G3842;
			G533<=G530;
			G535<=G3844;
			G536<=G6363;
			G539<=G3845;
			G540<=G6364;
			G543<=G3846;
			G544<=G6365;
			G547<=G9026;
			G550<=G9027;
			G553<=G9028;
			G556<=G3847;
			G557<=G6366;
			G560<=G6370;
			G563<=G9029;
			G566<=G3848;
			G567<=G6367;
			G570<=G9030;
			G573<=G9033;
			G576<=G3849;
			G579<=G3850;
			G580<=G6368;
			G583<=G3851;
			G584<=G6369;
			G587<=G3852;
			G588<=G9031;
			G591<=G9032;
			G595<=G576;
			G596<=G6795;
			G597<=G6796;
			G598<=G6797;
			G599<=G6798;
			G600<=G6807;
			G601<=G6799;
			G602<=G6800;
			G603<=G6801;
			G604<=G6802;
			G605<=G6803;
			G606<=G6804;
			G607<=G6805;
			G608<=G6806;
			G609<=G6808;
			G610<=G6809;
			G611<=G6810;
			G612<=G6811;
			G613<=G6820;
			G614<=G6812;
			G615<=G6813;
			G616<=G6814;
			G617<=G6815;
			G618<=G6816;
			G619<=G6817;
			G620<=G6818;
			G621<=G6819;
			G622<=G6821;
			G623<=G6822;
			G624<=G6831;
			G625<=G6823;
			G626<=G6824;
			G627<=G6825;
			G628<=G6826;
			G629<=G6827;
			G630<=G6828;
			G631<=G6829;
			G632<=G6830;
			G646<=G4652;
			G652<=G646;
			G661<=G7743;
			G665<=G7744;
			G669<=G7745;
			G673<=G7746;
			G677<=G7747;
			G681<=G7748;
			G685<=G7749;
			G689<=G6371;
			G706<=G7750;
			G710<=G7751;
			G714<=G7752;
			G718<=G7753;
			G727<=G8228;
			G730<=G7754;
			G734<=G7755;
			G741<=G9386;
			G746<=G8956;
			G758<=G6840;
			G759<=G6832;
			G760<=G6833;
			G761<=G6834;
			G762<=G6835;
			G763<=G6836;
			G764<=G6837;
			G765<=G6838;
			G766<=G6839;
			G767<=G6841;
			G768<=G6842;
			G769<=G6843;
			G770<=G6844;
			G771<=G6845;
			G772<=G6846;
			G773<=G6847;
			G774<=G6848;
			G775<=G7759;
			G778<=G7296;
			G782<=G5734;
			G789<=G7297;
			G792<=G5162;
			G799<=G7756;
			G803<=G7757;
			G806<=G7510;
			G809<=G7511;
			G812<=G7758;
			G815<=G7760;
			G819<=G7761;
			G822<=G7512;
			G825<=G7513;
			G828<=G7762;
			G831<=G2651;
			G834<=G2650;
			G837<=G2649;
			G840<=G2648;
			G843<=G2647;
			G846<=G2646;
			G849<=G2645;
			G852<=G2644;
			G855<=G8220;
			G859<=G8221;
			G863<=G8222;
			G866<=G5163;
			G871<=G5167;
			G874<=G4654;
			G875<=G5165;
			G878<=G890;
			G883<=G921;
			G887<=G7099;
			G888<=G7100;
			G889<=G7101;
			G890<=G7102;
			G891<=G3855;
			G896<=G891;
			G901<=G896;
			G906<=G901;
			G911<=G906;
			G916<=G911;
			G921<=G916;
			G926<=G878;
			G933<=G5166;
			G936<=G5168;
			G940<=G5735;
			G942<=G2652;
			G943<=G8671;
			G944<=G6372;
			G945<=G5170;
			G948<=G8664;
			G949<=G8665;
			G950<=G8666;
			G951<=G8667;
			G952<=G8668;
			G953<=G8669;
			G954<=G8670;
			G959<=G5169;
			G963<=G7764;
			G966<=G8223;
			G969<=G966;
			G970<=G963;
			G971<=G5171;
			G972<=G2653;
			G973<=G8672;
			G976<=G8864;
			G979<=G7104;
			G984<=G9133;
			G985<=G7515;
			G990<=G7516;
			G995<=G7517;
			G998<=G1005;
			G999<=G8865;
			G1004<=G7105;
			G1005<=G1004;
			G1007<=G8867;
			G1012<=G6851;
			G1013<=G1014;
			G1014<=G1012;
			G1018<=G8869;
			G1021<=G8870;
			G1025<=G8871;
			G1029<=G2654;
			G1030<=G7518;
			G1033<=G9034;
			G1034<=G8957;
			G1037<=G7519;
			G1041<=G7765;
			G1045<=G8224;
			G1049<=G8673;
			G1053<=G8873;
			G1057<=G8959;
			G1061<=G9035;
			G1065<=G9117;
			G1069<=G9134;
			G1073<=G9145;
			G1077<=G7767;
			G1081<=G6852;
			G1084<=G7106;
			G1087<=G6853;
			G1092<=G7520;
			G1097<=G1185;
			G1098<=G6854;
			G1102<=G6855;
			G1106<=G7107;
			G1110<=G7299;
			G1114<=G7521;
			G1118<=G7766;
			G1122<=G8225;
			G1126<=G8674;
			G1130<=G7522;
			G1134<=G7523;
			G1138<=G7524;
			G1142<=G8874;
			G1146<=G1612;
			G1147<=G1146;
			G1148<=G1147;
			G1149<=G7525;
			G1153<=G6856;
			G1154<=G1153;
			G1155<=G1154;
			G1156<=G1081;
			G1157<=G1156;
			G1158<=G1159;
			G1159<=G1157;
			G1160<=G1163;
			G1163<=G2655;
			G1166<=G1167;
			G1167<=G1170;
			G1170<=G1173;
			G1173<=G7526;
			G1176<=G5172;
			G1179<=G1186;
			G1182<=G1160;
			G1185<=G1155;
			G1186<=G1182;
			G1189<=G6392;
			G1190<=G8677;
			G1191<=G6373;
			G1192<=G1191;
			G1193<=G1192;
			G1195<=G6374;
			G1197<=G1196;
			G1199<=G6375;
			G1200<=G1199;
			G1201<=G1200;
			G1204<=G1203;
			G1205<=G1204;
			G1207<=G5173;
			G1211<=G5174;
			G1214<=G5736;
			G1217<=G6377;
			G1220<=G6378;
			G1223<=G6379;
			G1224<=G6857;
			G1225<=G6858;
			G1226<=G6859;
			G1227<=G7108;
			G1228<=G7109;
			G1229<=G7110;
			G1230<=G7300;
			G1231<=G1236;
			G1236<=G1240;
			G1240<=G1235;
			G1243<=G2660;
			G1244<=G2659;
			G1245<=G1244;
			G1247<=G6380;
			G1250<=G7111;
			G1251<=G6860;
			G1252<=G2661;
			G1253<=G5741;
			G1254<=G6381;
			G1257<=G5738;
			G1260<=G6382;
			G1263<=G5737;
			G1266<=G5739;
			G1267<=G4656;
			G1268<=G5175;
			G1269<=G5740;
			G1270<=G1271;
			G1271<=G5176;
			G1272<=G6383;
			G1276<=G6384;
			G1280<=G7112;
			G1284<=G7301;
			G1288<=G7527;
			G1292<=G7302;
			G1296<=G7304;
			G1300<=G7303;
			G1304<=G1312;
			G1307<=G3858;
			G1308<=G6385;
			G1309<=G1308;
			G1310<=G1309;
			G1311<=G1310;
			G1312<=G1311;
			G1313<=G5742;
			G1317<=G5743;
			G1318<=G6861;
			G1319<=G7113;
			G1320<=G7114;
			G1321<=G7115;
			G1322<=G7116;
			G1323<=G7117;
			G1324<=G7118;
			G1325<=G7305;
			G1326<=G7306;
			G1327<=G7307;
			G1328<=G7309;
			G1329<=G2663;
			G1330<=G6862;
			G1333<=G6863;
			G1336<=G6864;
			G1339<=G6865;
			G1342<=G7119;
			G1345<=G7528;
			G1348<=G7529;
			G1351<=G7530;
			G1354<=G7768;
			G1357<=G8675;
			G1360<=G8676;
			G1363<=G6877;
			G1364<=G6878;
			G1365<=G6867;
			G1366<=G6866;
			G1367<=G6873;
			G1368<=G6874;
			G1369<=G6875;
			G1370<=G6876;
			G1371<=G6868;
			G1372<=G6870;
			G1373<=G6871;
			G1374<=G6872;
			G1375<=G6869;
			G1376<=G6890;
			G1377<=G6891;
			G1378<=G6880;
			G1379<=G6879;
			G1380<=G6886;
			G1381<=G6887;
			G1382<=G6888;
			G1383<=G6889;
			G1384<=G6881;
			G1385<=G6883;
			G1386<=G6884;
			G1387<=G6885;
			G1388<=G6882;
			G1389<=G4658;
			G1390<=G4659;
			G1391<=G1390;
			G1392<=G6387;
			G1393<=G2664;
			G1394<=G6388;
			G1395<=G1393;
			G1396<=G4662;
			G1397<=G6389;
			G1398<=G1396;
			G1399<=G3861;
			G1400<=G6390;
			G1401<=G1399;
			G1402<=G6391;
			G1403<=G1402;
			G1404<=G1403;
			G1405<=G5744;
			G1408<=G5177;
			G1409<=G5178;
			G1412<=G5745;
			G1415<=G5180;
			G1416<=G4665;
			G1421<=G5179;
			G1424<=G3862;
			G1428<=G2672;
			G1429<=G2671;
			G1430<=G4666;
			G1431<=G2673;
			G1432<=G5183;
			G1435<=G5181;
			G1439<=G5182;
			G1443<=G4667;
			G1444<=G5185;
			G1450<=G5186;
			G1454<=G5187;
			G1459<=G3863;
			G1460<=G4668;
			G1461<=G4669;
			G1462<=G8678;
			G1467<=G8875;
			G1472<=G8960;
			G1477<=G9036;
			G1481<=G7769;
			G1486<=G8226;
			G1489<=G7770;
			G1494<=G7771;
			G1499<=G7772;
			G1504<=G7773;
			G1509<=G7774;
			G1513<=G1524;
			G1514<=G7775;
			G1519<=G8227;
			G1524<=G6393;
			G1528<=G7776;
			G1532<=G7781;
			G1537<=G7777;
			G1541<=G7778;
			G1545<=G7779;
			G1549<=G7780;
		end if;
	end process;
	G206<= not I5353;
	G291<= not I5356;
	G372<= not I5359;
	G453<= not I5362;
	G534<= not I5365;
	G594<= not I5368;
	G636<= not I5371;
	G639<= not I5374;
	G642<= not I5377;
	G649<= not I5380;
	G655<= not I5383;
	G658<= not I5386;
	G691<= not I5389;
	G695<= not I5392;
	G699<= not I5395;
	G703<= not I5398;
	G724<= not I5401;
	G738<= not I5404;
	G785<= not I5407;
	G1006<= not I5410;
	G1011<= not I5413;
	G1015<= not I5416;
	G1017<= not I5419;
	G1235<= not I5422;
	G1246<= not I5425;
	G1555<= not I5428;
	G1556<= not G65;
	G1557<= not I5432;
	G1558<= not I5435;
	G1562<= not G636;
	G1563<= not G639;
	G1564<= not G642;
	G1565<= not G649;
	G1566<= not G652;
	G1567<= not G655;
	G1568<= not G658;
	G1569<= not G661;
	G1570<= not G665;
	G1571<= not G669;
	G1572<= not G673;
	G1573<= not G677;
	G1574<= not G681;
	G1575<= not G685;
	G1576<= not G691;
	G1577<= not G695;
	G1578<= not G699;
	G1579<= not G703;
	G1580<= not G706;
	G1581<= not G710;
	G1582<= not G714;
	G1583<= not G718;
	G1584<= not G738;
	G1585<= not G724;
	G1586<= not G730;
	G1587<= not G734;
	G1588<= not G741;
	G1589<= not G746;
	G1590<= not I5466;
	G1597<= not G973;
	G1600<= not G976;
	G1603<= not I5471;
	G1611<= not G1073;
	G1612<= not I5475;
	G1616<= not I5478;
	G1637<= not G1087;
	G1638<= not G1092;
	G1639<= not G1207;
	G1643<= not G1211;
	G1646<= not G1214;
	G1649<= not G1217;
	G1652<= not G1220;
	G1655<= not G1231;
	G1658<= not G1313;
	G1661<= not G1405;
	G1662<= not G1412;
	G1663<= not G1416;
	G1664<= not G1462;
	G1665<= not G1467;
	G1666<= not G1472;
	G1667<= not G1481;
	G1670<= not G1489;
	G1671<= not G1494;
	G1672<= not G1499;
	G1673<= not G1504;
	G1674<= not G1514;
	G1675<= not G1519;
	G1676<= not G727;
	G1677<= not G1532;
	G1679<= not I5512;
	G1680<= not I5515;
	G1681<= not G929;
	G1683<= not G795;
	G1684<= not G1;
	G1685<= not I5528;
	G1686<= not I5531;
	G1687<= not G10;
	G1688<= not I5535;
	G1689<= not G855;
	G1694<= not G21;
	G1695<= not G778;
	G1698<= not I5542;
	G1701<= not I5545;
	G1704<= not I5548;
	G1707<= not G955;
	G1708<= not I5552;
	G1711<= not I5555;
	G1715<= not I5559;
	G1718<= not I5562;
	G1721<= not I5565;
	G1724<= not I5568;
	G1726<= not G158;
	G1727<= not G596;
	G1732<= not G1439;
	G1736<= not I5577;
	G1737<= not G597;
	G1738<= not G741;
	G1742<= not G1486;
	G1743<= not G598;
	G1744<= not G600;
	G1745<= not G746;
	G1746<= not G290;
	G1747<= not G599;
	G1748<= not G601;
	G1749<= not G371;
	G1750<= not G602;
	G1751<= not G452;
	G1752<= not G603;
	G1756<= not G533;
	G1757<= not G604;
	G1758<= not G1084;
	G1760<= not I5605;
	G1768<= not G605;
	G1769<= not I5609;
	G1770<= not G606;
	G1771<= not G609;
	G1772<= not G607;
	G1773<= not G610;
	G1774<= not I5616;
	G1776<= not G608;
	G1777<= not G611;
	G1778<= not G613;
	G1779<= not G612;
	G1780<= not G614;
	G1781<= not G622;
	G1782<= not G624;
	G1783<= not I5633;
	G1784<= not I5636;
	G1785<= not G615;
	G1786<= not G623;
	G1787<= not G625;
	G1788<= not G984;
	G1789<= not G1034;
	G1792<= not G616;
	G1793<= not G626;
	G1794<= not I5646;
	G1795<= not I5649;
	G1796<= not G617;
	G1797<= not G627;
	G1798<= not I5654;
	G1799<= not I5657;
	G1800<= not G1477;
	G1801<= not G618;
	G1802<= not G628;
	G1803<= not G758;
	G1804<= not I5664;
	G1805<= not I5667;
	G1806<= not I5670;
	G1807<= not G619;
	G1808<= not G629;
	G1809<= not G759;
	G1810<= not I5676;
	G1811<= not I5679;
	G1812<= not I5682;
	G1813<= not G620;
	G1814<= not G630;
	G1815<= not G760;
	G1816<= not G767;
	G1817<= not I5689;
	G1818<= not I5692;
	G1820<= not G621;
	G1821<= not G631;
	G1822<= not G761;
	G1823<= not G768;
	G1824<= not I5706;
	G1825<= not I5709;
	G1826<= not G632;
	G1827<= not G762;
	G1828<= not G769;
	G1829<= not I5715;
	G1830<= not I5718;
	G1831<= not G689;
	G1832<= not G763;
	G1833<= not G770;
	G1837<= not G1007;
	G1838<= not G1450;
	G1842<= not G764;
	G1843<= not G771;
	G1847<= not G765;
	G1848<= not G772;
	G1849<= not I5732;
	G1852<= not G887;
	G1853<= not G766;
	G1854<= not G773;
	G1855<= not G866;
	G1856<= not G774;
	G1857<= not G889;
	G1860<= not G162;
	G1863<= not G68;
	G1864<= not G162;
	G1865<= not G1013;
	G1866<= not G71;
	G1867<= not G878;
	G1868<= not I5747;
	G1869<= not G74;
	G1870<= not I5751;
	G1871<= not I5754;
	G1876<= not G77;
	G1877<= not G595;
	G1878<= not G80;
	G1879<= not I5763;
	G1886<= not I5766;
	G1887<= not G83;
	G1888<= not G781;
	G1889<= not G1018;
	G1894<= not I5772;
	G1895<= not I5775;
	G1896<= not G86;
	G1897<= not G789;
	G1901<= not I5781;
	G1904<= not G1021;
	G1907<= not G52;
	G1908<= not G812;
	G1909<= not G998;
	G1911<= not I5789;
	G1912<= not G1524;
	G1916<= not G775;
	G1917<= not I5795;
	G1918<= not G822;
	G1922<= not G1251;
	G1923<= not I5801;
	G1924<= not G174;
	G1925<= not G825;
	G1926<= not G874;
	G1929<= not G1224;
	G1933<= not G1247;
	G1934<= not G154;
	G1935<= not G1280;
	G1938<= not G1288;
	G1941<= not I5812;
	G1942<= not G828;
	G1943<= not G1025;
	G1944<= not I5817;
	G1945<= not G1081;
	G1948<= not G1250;
	G1949<= not G1292;
	G1952<= not G1333;
	G1958<= not G786;
	G1959<= not G1252;
	G1960<= not G1268;
	G1961<= not G1345;
	G1967<= not G1432;
	G1970<= not I5831;
	G1974<= not G803;
	G1975<= not G1253;
	G1976<= not G1269;
	G1977<= not G1357;
	G1983<= not I5839;
	G1987<= not I5842;
	G2006<= not G806;
	G2007<= not G1223;
	G2011<= not I5847;
	G2015<= not G33;
	G2016<= not I5852;
	G2020<= not I5855;
	G2038<= not G809;
	G2039<= not G1228;
	G2044<= not I5861;
	G2052<= not I5865;
	G2057<= not I5868;
	G2073<= not G1254;
	G2074<= not I5872;
	G2091<= not G819;
	G2092<= not G1225;
	G2096<= not G1226;
	G2100<= not G1227;
	G2104<= not I5879;
	G2105<= not G1444;
	G2106<= not I5883;
	G2128<= not G1284;
	G2131<= not G1300;
	G2134<= not G1317;
	G2137<= not I5889;
	G2145<= not G1296;
	G2148<= not G1304;
	G2149<= not I5894;
	G2157<= not I5897;
	G2161<= not G1454;
	G2162<= not I5901;
	G2170<= not G1229;
	G2174<= not G1319;
	G2177<= not G1322;
	G2180<= not G1318;
	G2183<= not I5908;
	G2184<= not I5911;
	G2185<= not I5914;
	G2202<= not G1321;
	G2205<= not G13;
	G2207<= not I5920;
	G2208<= not I5923;
	G2209<= not I5926;
	G2210<= not G1326;
	G2215<= not G1416;
	G2216<= not I5933;
	G2221<= not I5936;
	G2222<= not I5939;
	G2223<= not I5942;
	G2224<= not I5945;
	G2225<= not I5948;
	G2226<= not G1320;
	G2231<= not I5954;
	G2232<= not I5957;
	G2233<= not I5960;
	G2234<= not I5963;
	G2235<= not I5966;
	G2236<= not I5969;
	G2237<= not I5972;
	G2238<= not I5975;
	G2239<= not I5978;
	G2240<= not I5981;
	G2241<= not I5984;
	G2242<= not G985;
	G2245<= not G999;
	G2246<= not I5989;
	G2253<= not G1323;
	G2256<= not G1324;
	G2259<= not G1325;
	G2263<= not G1394;
	G2264<= not I5997;
	G2265<= not I6000;
	G2266<= not I6003;
	G2267<= not I6006;
	G2268<= not I6009;
	G2269<= not I6012;
	G2270<= not I6015;
	G2271<= not I6018;
	G2272<= not I6021;
	G2273<= not I6024;
	G2274<= not G782;
	G2275<= not G990;
	G2276<= not I6029;
	G2282<= not G1400;
	G2283<= not I6033;
	G2284<= not I6036;
	G2285<= not I6039;
	G2286<= not I6042;
	G2287<= not I6045;
	G2288<= not I6048;
	G2289<= not I6051;
	G2290<= not I6054;
	G2291<= not I6057;
	G2292<= not I6060;
	G2293<= not G888;
	G2295<= not G995;
	G2298<= not I6072;
	G2306<= not I6075;
	G2307<= not I6078;
	G2308<= not I6081;
	G2309<= not I6084;
	G2310<= not I6087;
	G2311<= not I6090;
	G2312<= not I6093;
	G2313<= not I6096;
	G2314<= not I6099;
	G2316<= not I6109;
	G2323<= not I6112;
	G2324<= not I6115;
	G2325<= not I6118;
	G2326<= not I6121;
	G2327<= not I6124;
	G2328<= not I6127;
	G2329<= not I6130;
	G2331<= not G933;
	G2332<= not G926;
	G2334<= not I6143;
	G2340<= not G1327;
	G2343<= not G1392;
	G2344<= not I6148;
	G2345<= not I6151;
	G2346<= not I6154;
	G2347<= not I6157;
	G2348<= not I6160;
	G2349<= not I6163;
	G2350<= not I6166;
	G2351<= not G792;
	G2353<= not G871;
	G2354<= not I6178;
	G2359<= not G1397;
	G2360<= not G1435;
	G2361<= not I6183;
	G2362<= not I6186;
	G2363<= not I6189;
	G2364<= not I6192;
	G2365<= not I6195;
	G2366<= not I6198;
	G2371<= not G944;
	G2372<= not I6214;
	G2373<= not I6217;
	G2374<= not I6220;
	G2375<= not I6223;
	G2376<= not I6226;
	G2377<= not I6229;
	G2379<= not I6239;
	G2380<= not I6242;
	G2381<= not I6245;
	G2382<= not I6248;
	G2383<= not I6251;
	G2384<= not I6254;
	G2389<= not G1230;
	G2392<= not G11;
	G2393<= not I6267;
	G2394<= not I6270;
	G2396<= not G1033;
	G2397<= not G1272;
	G2401<= not G22;
	G2402<= not G29;
	G2403<= not G1176;
	G2404<= not G1276;
	G2407<= not I6286;
	G2424<= not G1329;
	G2452<= not G23;
	G2453<= not I6291;
	G2454<= not I6294;
	G2457<= not G24;
	G2458<= not G30;
	G2459<= not I6299;
	G2460<= not I6302;
	G2467<= not I6305;
	G2470<= not G42;
	G2471<= not I6309;
	G2477<= not G25;
	G2478<= not G31;
	G2479<= not G32;
	G2480<= not G44;
	G2481<= not I6317;
	G2484<= not G45;
	G2485<= not G62;
	G2486<= not G959;
	G2487<= not I6323;
	G2490<= not I6326;
	G2494<= not G9;
	G2495<= not G26;
	G2496<= not G942;
	G2497<= not G945;
	G2498<= not I6333;
	G2501<= not G27;
	G2502<= not I6337;
	G2505<= not G28;
	G2506<= not I6341;
	G2509<= not G37;
	G2510<= not G58;
	G2511<= not G1328;
	G2514<= not G1330;
	G2517<= not I6348;
	G2520<= not G41;
	G2522<= not G1342;
	G2525<= not I6354;
	G2528<= not G1260;
	G2532<= not I6358;
	G2533<= not G1336;
	G2536<= not G1354;
	G2539<= not I6363;
	G2540<= not G1339;
	G2543<= not G1348;
	G2546<= not I6368;
	G2547<= not I6371;
	G2548<= not G1351;
	G2551<= not G1360;
	G2554<= not I6376;
	G2555<= not G936;
	G2556<= not G1190;
	G2557<= not G940;
	G2561<= not G1555;
	G2562<= not G1652;
	G2573<= not G1649;
	G2584<= not G1646;
	G2595<= not G1643;
	G2605<= not G1639;
	G2614<= not G1562;
	G2615<= not G1563;
	G2616<= not G1564;
	G2617<= not G1565;
	G2618<= not G1566;
	G2621<= not G1567;
	G2622<= not G1568;
	G2623<= not G1585;
	G2624<= not G1569;
	G2625<= not G1570;
	G2626<= not G1571;
	G2627<= not G1572;
	G2628<= not G1573;
	G2629<= not G1574;
	G2630<= not G1575;
	G2631<= not G1586;
	G2632<= not G1576;
	G2633<= not G1577;
	G2634<= not G1578;
	G2635<= not G1579;
	G2636<= not G1580;
	G2637<= not G1581;
	G2638<= not G1582;
	G2639<= not G1583;
	G2640<= not G1584;
	G2641<= not G1587;
	G2642<= not G1588;
	G2643<= not G1589;
	G2644<= not I6416;
	G2645<= not I6419;
	G2646<= not I6422;
	G2647<= not I6425;
	G2648<= not I6428;
	G2649<= not I6431;
	G2650<= not I6434;
	G2651<= not I6437;
	G2652<= not I6440;
	G2653<= not I6443;
	G2654<= not I6446;
	G2655<= not G1611;
	G2659<= not G1655;
	G2660<= not I6451;
	G2661<= not I6454;
	G2662<= not I6457;
	G2663<= not I6460;
	G2664<= not I6463;
	G2665<= not G1661;
	G2668<= not G1662;
	G2671<= not I6468;
	G2672<= not I6471;
	G2673<= not I6474;
	G2674<= not G1675;
	G2677<= not G1664;
	G2680<= not G1665;
	G2683<= not G1666;
	G2686<= not G1667;
	G2689<= not G1670;
	G2692<= not G1671;
	G2695<= not G1672;
	G2698<= not G1673;
	G2699<= not G1674;
	G2700<= not G1744;
	G2703<= not G1809;
	G2706<= not G1821;
	G2709<= not G1747;
	G2712<= not G2039;
	G2721<= not G1803;
	G2724<= not G1814;
	G2727<= not G2424;
	G2728<= not G2256;
	G2734<= not G2170;
	G2743<= not G1808;
	G2746<= not G2259;
	G2752<= not G2389;
	G2761<= not G1820;
	G2764<= not G1802;
	G2767<= not I6509;
	G2769<= not G2424;
	G2770<= not G2210;
	G2774<= not G1813;
	G2777<= not G1797;
	G2780<= not I6517;
	G2782<= not G1616;
	G2784<= not G2340;
	G2787<= not G1807;
	G2790<= not G1793;
	G2793<= not I6532;
	G2794<= not G2185;
	G2795<= not G1801;
	G2798<= not G1787;
	G2804<= not G1796;
	G2807<= not G1782;
	G2810<= not G1922;
	G2816<= not G1685;
	G2817<= not G1849;
	G2818<= not G1792;
	G2821<= not G1786;
	G2824<= not G1688;
	G2825<= not I6553;
	G2826<= not G2183;
	G2828<= not G1980;
	G2829<= not G1785;
	G2832<= not G2184;
	G2833<= not I6561;
	G2834<= not I6564;
	G2837<= not G1780;
	G2840<= not G2207;
	G2841<= not G2208;
	G2842<= not G2209;
	G2843<= not I6571;
	G2844<= not I6574;
	G2862<= not I6578;
	G2863<= not G1778;
	G2866<= not G2221;
	G2867<= not G2222;
	G2868<= not G2223;
	G2869<= not G2224;
	G2870<= not G2225;
	G2871<= not I6587;
	G2872<= not I6590;
	G2873<= not G1779;
	G2876<= not G2231;
	G2877<= not G2232;
	G2878<= not G2233;
	G2879<= not I6597;
	G2880<= not G2234;
	G2881<= not G2235;
	G2882<= not G2236;
	G2883<= not G2237;
	G2884<= not G2238;
	G2885<= not G2239;
	G2886<= not G2240;
	G2887<= not G2241;
	G2888<= not I6608;
	G2890<= not G2264;
	G2891<= not G2265;
	G2892<= not G2266;
	G2893<= not I6615;
	G2894<= not G2267;
	G2895<= not G2268;
	G2896<= not G2269;
	G2897<= not G2270;
	G2898<= not G2271;
	G2899<= not G2272;
	G2900<= not G2273;
	G2901<= not G2284;
	G2902<= not G2285;
	G2903<= not G2286;
	G2904<= not G2287;
	G2905<= not I6629;
	G2906<= not G2288;
	G2907<= not G2289;
	G2908<= not G2290;
	G2909<= not G2291;
	G2910<= not I6636;
	G2911<= not G2292;
	G2913<= not G2307;
	G2914<= not G2308;
	G2915<= not I6643;
	G2916<= not I6646;
	G2917<= not G2309;
	G2918<= not G2310;
	G2919<= not G2311;
	G2920<= not I6652;
	G2921<= not G2312;
	G2922<= not G2313;
	G2923<= not I6657;
	G2924<= not G2314;
	G2925<= not G2324;
	G2926<= not G2325;
	G2927<= not I6663;
	G2928<= not G2326;
	G2929<= not G2327;
	G2930<= not G2328;
	G2931<= not I6669;
	G2932<= not G2329;
	G2933<= not I6673;
	G2934<= not I6676;
	G2936<= not I6680;
	G2937<= not G2346;
	G2938<= not G2347;
	G2939<= not G2348;
	G2940<= not I6686;
	G2941<= not G2349;
	G2942<= not G2350;
	G2943<= not G2362;
	G2944<= not G2363;
	G2945<= not G2364;
	G2946<= not G2365;
	G2947<= not I6695;
	G2948<= not G2366;
	G2953<= not G2373;
	G2954<= not G2374;
	G2955<= not I6703;
	G2956<= not G2375;
	G2957<= not G2376;
	G2958<= not G2377;
	G2959<= not G1926;
	G2960<= not G2381;
	G2961<= not I6711;
	G2962<= not G2382;
	G2963<= not G2383;
	G2964<= not I6716;
	G2965<= not G2384;
	G2966<= not G1856;
	G2969<= not G2393;
	G2970<= not G2394;
	G2971<= not I6723;
	G2973<= not G1854;
	G2976<= not I6728;
	G2982<= not G1848;
	G2985<= not I6733;
	G2989<= not G1843;
	G2992<= not G1833;
	G2996<= not G1828;
	G2999<= not G1823;
	G3008<= not G1816;
	G3013<= not I6764;
	G3014<= not I6767;
	G3018<= not I6770;
	G3019<= not G2007;
	G3029<= not G1929;
	G3038<= not G2092;
	G3047<= not G1736;
	G3048<= not I6784;
	G3050<= not I6788;
	G3051<= not I6791;
	G3052<= not G2096;
	G3061<= not I6795;
	G3062<= not G2100;
	G3071<= not G1948;
	G3074<= not I6800;
	G3075<= not G2216;
	G3076<= not G1831;
	G3077<= not I6805;
	G3078<= not G1603;
	G3079<= not G1603;
	G3080<= not G1679;
	G3082<= not G1680;
	G3084<= not I6820;
	G3085<= not G1945;
	G3086<= not G1852;
	G3091<= not G1603;
	G3092<= not I6826;
	G3093<= not G1686;
	G3095<= not I6831;
	G3096<= not I6834;
	G3124<= not G1857;
	G3128<= not I6839;
	G3130<= not I6849;
	G3158<= not I6853;
	G3159<= not I6856;
	G3187<= not I6860;
	G3189<= not I6864;
	G3191<= not I6868;
	G3219<= not I6872;
	G3220<= not G1889;
	G3230<= not I6887;
	G3238<= not I6894;
	G3264<= not I6900;
	G3285<= not G1689;
	G3287<= not I6911;
	G3316<= not I6930;
	G3338<= not G1901;
	G3340<= not G2474;
	G3341<= not I6936;
	G3359<= not I6946;
	G3390<= not I6949;
	G3398<= not I6952;
	G3430<= not I6956;
	G3461<= not I6959;
	G3462<= not G1743;
	G3465<= not I6963;
	G3485<= not G1737;
	G3488<= not G1727;
	G3491<= not G1800;
	G3492<= not I6970;
	G3495<= not G1616;
	G3496<= not I6974;
	G3497<= not G2185;
	G3498<= not G1616;
	G3499<= not G2185;
	G3500<= not G1616;
	G3501<= not G2185;
	G3502<= not G1616;
	G3503<= not G2407;
	G3506<= not G1781;
	G3510<= not G2185;
	G3511<= not G1616;
	G3512<= not G1616;
	G3513<= not G2407;
	G3514<= not G2424;
	G3517<= not G2283;
	G3519<= not G2185;
	G3520<= not G1616;
	G3521<= not G2185;
	G3522<= not G2407;
	G3523<= not G2407;
	G3524<= not G2306;
	G3526<= not G2185;
	G3527<= not G1616;
	G3529<= not G2323;
	G3530<= not G2185;
	G3531<= not G1616;
	G3532<= not G2407;
	G3533<= not G2397;
	G3539<= not G2424;
	G3540<= not G2424;
	G3542<= not G1777;
	G3545<= not G2344;
	G3546<= not I7029;
	G3547<= not G2345;
	G3548<= not G2185;
	G3549<= not G2404;
	G3556<= not I7036;
	G3557<= not G1773;
	G3560<= not G2361;
	G3561<= not I7041;
	G3562<= not I7044;
	G3563<= not G2007;
	G3567<= not G2407;
	G3568<= not G1935;
	G3573<= not G2424;
	G3574<= not G1771;
	G3577<= not G2372;
	G3578<= not I7053;
	G3579<= not G1929;
	G3582<= not G2407;
	G3583<= not G2128;
	G3587<= not G1964;
	G3588<= not G2379;
	G3589<= not I7061;
	G3590<= not I7064;
	G3591<= not G1789;
	G3603<= not G2092;
	G3604<= not G2407;
	G3605<= not G1938;
	G3610<= not G2424;
	G3611<= not I7079;
	G3612<= not I7082;
	G3617<= not G1655;
	G3629<= not G2424;
	G3630<= not I7095;
	G3631<= not I7098;
	G3632<= not I7101;
	G3633<= not I7104;
	G3634<= not I7107;
	G3635<= not G1949;
	G3639<= not G2424;
	G3640<= not I7112;
	G3641<= not I7115;
	G3642<= not I7118;
	G3643<= not G2453;
	G3644<= not G2131;
	G3647<= not G2424;
	G3648<= not G2424;
	G3649<= not G2424;
	G3650<= not I7126;
	G3651<= not I7129;
	G3652<= not I7132;
	G3653<= not G2459;
	G3654<= not G2521;
	G3655<= not G1844;
	G3657<= not I7145;
	G3659<= not G2293;
	G3666<= not G2134;
	G3674<= not I7164;
	G3675<= not I7167;
	G3676<= not G2380;
	G3677<= not G2485;
	G3684<= not G2180;
	G3691<= not I7195;
	G3692<= not I7198;
	G3693<= not G2424;
	G3694<= not G2174;
	G3700<= not G2514;
	G3705<= not I7204;
	G3707<= not G2226;
	G3712<= not G1952;
	G3716<= not G2522;
	G3721<= not I7211;
	G3723<= not G2096;
	G3728<= not G2202;
	G3732<= not G2533;
	G3735<= not G1961;
	G3739<= not G2536;
	G3743<= not G1776;
	G3746<= not G2100;
	G3750<= not G2177;
	G3753<= not G2540;
	G3754<= not G2543;
	G3757<= not G1977;
	G3761<= not G1772;
	G3764<= not G2039;
	G3768<= not G2253;
	G3769<= not G2548;
	G3770<= not G2551;
	G3771<= not G1853;
	G3774<= not G1770;
	G3777<= not G2170;
	G3778<= not G2145;
	G3779<= not G2511;
	G3780<= not G1847;
	G3783<= not I7255;
	G3784<= not G1768;
	G3787<= not G1842;
	G3798<= not G1757;
	G3801<= not I7262;
	G3802<= not G1832;
	G3805<= not G1752;
	G3808<= not G1827;
	G3812<= not G1750;
	G3815<= not G1822;
	G3819<= not G1748;
	G3822<= not G1815;
	G3825<= not G1826;
	G3828<= not I7287;
	G3829<= not I7290;
	G3830<= not I7293;
	G3831<= not I7296;
	G3832<= not I7299;
	G3833<= not I7302;
	G3834<= not I7305;
	G3835<= not I7308;
	G3836<= not I7311;
	G3837<= not I7314;
	G3838<= not I7317;
	G3839<= not I7320;
	G3840<= not I7323;
	G3841<= not I7326;
	G3842<= not I7329;
	G3843<= not I7332;
	G3844<= not I7335;
	G3845<= not I7338;
	G3846<= not I7341;
	G3847<= not I7344;
	G3848<= not I7347;
	G3849<= not I7350;
	G3850<= not I7353;
	G3851<= not I7356;
	G3852<= not I7359;
	G3853<= not I7362;
	G3854<= not I7365;
	G3855<= not I7368;
	G3856<= not I7371;
	G3857<= not I7374;
	G3858<= not I7377;
	G3859<= not I7380;
	G3860<= not I7383;
	G3861<= not I7386;
	G3862<= not I7389;
	G3863<= not I7392;
	G3864<= not G2943;
	G3865<= not G2944;
	G3866<= not G2945;
	G3867<= not G2946;
	G3868<= not G2948;
	G3869<= not I7400;
	G3870<= not G3466;
	G3871<= not G2953;
	G3872<= not G2954;
	G3873<= not G2956;
	G3874<= not G2957;
	G3875<= not G2958;
	G3876<= not G3466;
	G3877<= not G2960;
	G3878<= not G2962;
	G3879<= not G2963;
	G3880<= not G2965;
	G3881<= not G2969;
	G3882<= not G2970;
	G3884<= not I7417;
	G3888<= not G3097;
	G3891<= not G3097;
	G3892<= not G3131;
	G3896<= not I7473;
	G3897<= not G3131;
	G3898<= not G3160;
	G3901<= not I7492;
	G3902<= not I7495;
	G3903<= not I7498;
	G3904<= not G3160;
	G3905<= not G3192;
	G3908<= not I7517;
	G3909<= not I7520;
	G3910<= not I7523;
	G3911<= not I7526;
	G3912<= not G3192;
	G3913<= not G2834;
	G3916<= not I7545;
	G3917<= not I7548;
	G3918<= not I7551;
	G3919<= not I7554;
	G3920<= not G3097;
	G3921<= not I7558;
	G3922<= not I7561;
	G3923<= not I7564;
	G3926<= not I7581;
	G3927<= not I7584;
	G3928<= not G3097;
	G3929<= not I7588;
	G3930<= not G3097;
	G3931<= not I7592;
	G3932<= not I7595;
	G3933<= not G3131;
	G3934<= not I7599;
	G3935<= not I7602;
	G3936<= not I7605;
	G3937<= not G2845;
	G3940<= not I7623;
	G3941<= not I7626;
	G3942<= not I7629;
	G3943<= not I7632;
	G3944<= not I7635;
	G3945<= not G3097;
	G3946<= not G3097;
	G3947<= not I7640;
	G3948<= not G3131;
	G3949<= not I7644;
	G3950<= not G3131;
	G3951<= not I7648;
	G3952<= not I7651;
	G3953<= not G3160;
	G3954<= not I7655;
	G3955<= not I7658;
	G3956<= not G2845;
	G3957<= not I7662;
	G3958<= not G3097;
	G3959<= not G3097;
	G3960<= not I7667;
	G3961<= not G3131;
	G3962<= not G3131;
	G3963<= not I7672;
	G3964<= not G3160;
	G3965<= not I7676;
	G3966<= not G3160;
	G3967<= not I7680;
	G3968<= not I7683;
	G3969<= not G3192;
	G3970<= not G2845;
	G3971<= not I7688;
	G3972<= not I7691;
	G3973<= not G3097;
	G3974<= not G3131;
	G3975<= not G3131;
	G3976<= not I7697;
	G3977<= not G3160;
	G3978<= not G3160;
	G3979<= not I7702;
	G3980<= not G3192;
	G3981<= not I7706;
	G3982<= not G3192;
	G3983<= not G2845;
	G3985<= not I7712;
	G3987<= not I7716;
	G3988<= not G3097;
	G3989<= not G3131;
	G3990<= not G3160;
	G3991<= not G3160;
	G3992<= not I7723;
	G3993<= not G3192;
	G3994<= not G3192;
	G3995<= not I7728;
	G3996<= not I7731;
	G3997<= not I7734;
	G3998<= not G3097;
	G3999<= not I7738;
	G4000<= not G3131;
	G4001<= not G3160;
	G4002<= not G3192;
	G4003<= not G3192;
	G4004<= not G2845;
	G4005<= not I7746;
	G4006<= not I7749;
	G4007<= not I7752;
	G4008<= not I7755;
	G4009<= not I7758;
	G4010<= not G3097;
	G4011<= not I7762;
	G4012<= not I7765;
	G4013<= not G3131;
	G4014<= not I7769;
	G4015<= not G3160;
	G4016<= not G3192;
	G4017<= not G2845;
	G4018<= not I7775;
	G4019<= not I7778;
	G4020<= not I7781;
	G4021<= not G3131;
	G4022<= not I7785;
	G4023<= not I7788;
	G4024<= not G3160;
	G4025<= not I7792;
	G4026<= not G3192;
	G4027<= not G2845;
	G4028<= not I7797;
	G4029<= not I7800;
	G4030<= not G3160;
	G4031<= not I7804;
	G4032<= not I7807;
	G4033<= not G3192;
	G4034<= not I7811;
	G4035<= not I7814;
	G4036<= not G3192;
	G4037<= not G2845;
	G4041<= not G2605;
	G4044<= not G2595;
	G4050<= not G3080;
	G4051<= not G3093;
	G4056<= not G3082;
	G4057<= not I7832;
	G4065<= not I7838;
	G4069<= not I7844;
	G4070<= not I7847;
	G4071<= not I7850;
	G4075<= not I7856;
	G4076<= not I7859;
	G4079<= not I7864;
	G4080<= not I7867;
	G4081<= not I7870;
	G4084<= not I7875;
	G4085<= not I7878;
	G4087<= not I7882;
	G4088<= not I7885;
	G4089<= not I7888;
	G4092<= not I7899;
	G4093<= not I7902;
	G4094<= not I7905;
	G4095<= not I7908;
	G4096<= not I7911;
	G4102<= not I7919;
	G4103<= not I7922;
	G4104<= not I7925;
	G4105<= not I7928;
	G4106<= not I7931;
	G4111<= not I7944;
	G4112<= not I7947;
	G4113<= not I7950;
	G4114<= not I7953;
	G4115<= not I7956;
	G4116<= not I7959;
	G4119<= not I7964;
	G4120<= not I7967;
	G4121<= not I7970;
	G4122<= not I7973;
	G4125<= not I7978;
	G4126<= not I7981;
	G4130<= not I7987;
	G4134<= not G3676;
	G4146<= not I8011;
	G4153<= not I8024;
	G4191<= not I8084;
	G4195<= not I8094;
	G4196<= not I8097;
	G4197<= not G3591;
	G4198<= not I8101;
	G4200<= not I8105;
	G4202<= not G2810;
	G4226<= not G3591;
	G4229<= not I8140;
	G4242<= not I8161;
	G4245<= not I8172;
	G4250<= not I8177;
	G4251<= not I8180;
	G4253<= not G2734;
	G4257<= not I8190;
	G4258<= not I8193;
	G4259<= not I8196;
	G4265<= not G3591;
	G4266<= not I8202;
	G4267<= not I8205;
	G4270<= not G2573;
	G4273<= not I8215;
	G4274<= not I8218;
	G4275<= not G3790;
	G4279<= not G3340;
	G4281<= not G2562;
	G4285<= not I8233;
	G4286<= not G3790;
	G4296<= not G3790;
	G4300<= not I8261;
	G4301<= not I8264;
	G4303<= not I8268;
	G4306<= not I8273;
	G4307<= not G3700;
	G4308<= not I8277;
	G4311<= not I8282;
	G4316<= not I8291;
	G4328<= not G3086;
	G4335<= not G3659;
	G4341<= not I8308;
	G4344<= not G3124;
	G4350<= not I8315;
	G4353<= not G3665;
	G4357<= not G3679;
	G4358<= not G3680;
	G4360<= not I8333;
	G4362<= not G2810;
	G4370<= not I8351;
	G4371<= not I8354;
	G4372<= not I8357;
	G4373<= not I8360;
	G4381<= not G3466;
	G4382<= not I8373;
	G4426<= not I8428;
	G4438<= not I8446;
	G4443<= not I8449;
	G4444<= not I8452;
	G4455<= not G3811;
	G4457<= not I8477;
	G4462<= not I8480;
	G4463<= not I8483;
	G4464<= not I8486;
	G4465<= not G3677;
	G4475<= not G3818;
	G4477<= not I8517;
	G4482<= not I8520;
	G4489<= not G2826;
	G4493<= not I8543;
	G4500<= not G2832;
	G4501<= not G2801;
	G4503<= not I8565;
	G4510<= not G2840;
	G4511<= not G2841;
	G4512<= not G2842;
	G4521<= not G2866;
	G4522<= not G2867;
	G4523<= not G2868;
	G4524<= not G2869;
	G4525<= not G2870;
	G4527<= not G3466;
	G4535<= not G2876;
	G4536<= not G2877;
	G4537<= not G2878;
	G4538<= not G2880;
	G4539<= not G2881;
	G4540<= not G2882;
	G4541<= not G2883;
	G4542<= not G2884;
	G4543<= not G2885;
	G4544<= not G2886;
	G4545<= not G2887;
	G4547<= not G3466;
	G4552<= not G2890;
	G4553<= not G2891;
	G4554<= not G2892;
	G4555<= not G2894;
	G4556<= not G2895;
	G4557<= not G2896;
	G4558<= not G2897;
	G4559<= not G2898;
	G4560<= not G2899;
	G4561<= not G2900;
	G4562<= not G3466;
	G4564<= not I8665;
	G4565<= not G2901;
	G4566<= not G2902;
	G4567<= not G2903;
	G4568<= not G2904;
	G4569<= not G2906;
	G4570<= not G2907;
	G4571<= not G2908;
	G4572<= not G2909;
	G4573<= not G2911;
	G4574<= not G3466;
	G4576<= not G2913;
	G4577<= not G2914;
	G4578<= not G2917;
	G4579<= not G2918;
	G4580<= not G2919;
	G4581<= not G2921;
	G4582<= not G2922;
	G4583<= not G2924;
	G4584<= not G3466;
	G4585<= not G2925;
	G4586<= not G2926;
	G4587<= not G2928;
	G4588<= not G2929;
	G4589<= not G2930;
	G4590<= not G2932;
	G4591<= not G2937;
	G4592<= not G2938;
	G4593<= not G2939;
	G4594<= not G2941;
	G4595<= not G2942;
	G4596<= not G3466;
	G4597<= not I8706;
	G4598<= not I8709;
	G4599<= not I8712;
	G4600<= not I8715;
	G4601<= not I8718;
	G4602<= not I8721;
	G4603<= not I8724;
	G4604<= not I8727;
	G4605<= not I8730;
	G4606<= not I8733;
	G4607<= not I8736;
	G4608<= not I8739;
	G4609<= not I8742;
	G4610<= not I8745;
	G4611<= not I8748;
	G4612<= not I8751;
	G4613<= not I8754;
	G4614<= not I8757;
	G4615<= not I8760;
	G4616<= not I8763;
	G4617<= not I8766;
	G4618<= not I8769;
	G4619<= not I8772;
	G4620<= not I8775;
	G4621<= not I8778;
	G4622<= not I8781;
	G4623<= not I8784;
	G4624<= not I8787;
	G4625<= not I8790;
	G4626<= not I8793;
	G4627<= not I8796;
	G4628<= not I8799;
	G4629<= not I8802;
	G4630<= not I8805;
	G4631<= not I8808;
	G4632<= not I8811;
	G4633<= not I8814;
	G4634<= not I8817;
	G4635<= not I8820;
	G4636<= not I8823;
	G4637<= not I8826;
	G4638<= not I8829;
	G4639<= not I8832;
	G4640<= not I8835;
	G4641<= not I8838;
	G4642<= not I8841;
	G4643<= not I8844;
	G4644<= not I8847;
	G4645<= not I8850;
	G4646<= not I8853;
	G4647<= not I8856;
	G4648<= not I8859;
	G4649<= not I8862;
	G4650<= not I8865;
	G4651<= not I8868;
	G4652<= not I8871;
	G4653<= not I8874;
	G4654<= not I8877;
	G4655<= not I8880;
	G4656<= not I8883;
	G4657<= not I8886;
	G4658<= not I8889;
	G4659<= not I8892;
	G4660<= not I8895;
	G4661<= not I8898;
	G4662<= not I8901;
	G4663<= not I8904;
	G4664<= not I8907;
	G4665<= not I8910;
	G4666<= not I8913;
	G4667<= not I8916;
	G4668<= not I8919;
	G4669<= not I8922;
	G4670<= not I8925;
	G4673<= not I8928;
	G4677<= not I8932;
	G4678<= not I8935;
	G4680<= not I8945;
	G4684<= not I8949;
	G4685<= not I8952;
	G4687<= not I8962;
	G4689<= not I8966;
	G4692<= not I8971;
	G4693<= not I8974;
	G4694<= not I8977;
	G4695<= not I8980;
	G4696<= not I8983;
	G4697<= not I8986;
	G4698<= not I8989;
	G4701<= not I8994;
	G4703<= not I8998;
	G4704<= not I9001;
	G4706<= not I9005;
	G4710<= not I9009;
	G4713<= not I9014;
	G4718<= not I9018;
	G4719<= not I9021;
	G4721<= not I9025;
	G4732<= not I9034;
	G4733<= not G4202;
	G4738<= not I9050;
	G4739<= not I9053;
	G4742<= not I9064;
	G4746<= not I9076;
	G4748<= not G4465;
	G4776<= not I9081;
	G4777<= not I9084;
	G4780<= not I9089;
	G4784<= not I9095;
	G4788<= not I9103;
	G4792<= not I9111;
	G4795<= not I9116;
	G4800<= not I9123;
	G4801<= not I9126;
	G4802<= not I9129;
	G4803<= not I9132;
	G4805<= not I9136;
	G4806<= not I9139;
	G4807<= not I9142;
	G4808<= not I9145;
	G4809<= not I9148;
	G4811<= not I9158;
	G4813<= not I9162;
	G4822<= not I9177;
	G4841<= not G4250;
	G4867<= not I9209;
	G4873<= not I9217;
	G4882<= not G4069;
	G4885<= not G4070;
	G4886<= not G4071;
	G4890<= not G4075;
	G4891<= not G4076;
	G4892<= not I9250;
	G4895<= not G4078;
	G4898<= not G4079;
	G4899<= not G4080;
	G4900<= not I9258;
	G4903<= not G4084;
	G4904<= not G4085;
	G4907<= not G4087;
	G4908<= not G4088;
	G4909<= not I9271;
	G4913<= not G4092;
	G4914<= not G4093;
	G4915<= not G4094;
	G4916<= not G4202;
	G4917<= not G4102;
	G4918<= not G4103;
	G4919<= not G4104;
	G4920<= not G4105;
	G4921<= not G4202;
	G4922<= not G4111;
	G4923<= not G4112;
	G4924<= not G4113;
	G4925<= not G4114;
	G4926<= not G4202;
	G4928<= not G4119;
	G4929<= not G4120;
	G4930<= not G4121;
	G4931<= not I9301;
	G4932<= not G4202;
	G4934<= not G4125;
	G4935<= not G4202;
	G4938<= not I9310;
	G4960<= not G4259;
	G4963<= not G4328;
	G5000<= not I9325;
	G5002<= not G4335;
	G5006<= not I9333;
	G5007<= not I9336;
	G5009<= not G4344;
	G5013<= not I9341;
	G5014<= not I9344;
	G5015<= not I9347;
	G5016<= not I9350;
	G5022<= not G4438;
	G5024<= not I9360;
	G5025<= not I9363;
	G5026<= not I9366;
	G5027<= not I9369;
	G5028<= not I9372;
	G5037<= not G4438;
	G5038<= not G4457;
	G5041<= not I9393;
	G5042<= not I9396;
	G5051<= not I9407;
	G5053<= not G4438;
	G5054<= not G4457;
	G5055<= not G4477;
	G5058<= not I9416;
	G5059<= not I9419;
	G5060<= not I9422;
	G5061<= not I9425;
	G5071<= not G4438;
	G5072<= not G4457;
	G5073<= not G4477;
	G5074<= not I9440;
	G5075<= not I9443;
	G5076<= not I9446;
	G5083<= not G4457;
	G5084<= not G4477;
	G5085<= not I9457;
	G5086<= not I9460;
	G5087<= not I9463;
	G5088<= not I9466;
	G5099<= not G4477;
	G5100<= not I9484;
	G5101<= not G4259;
	G5109<= not I9493;
	G5112<= not I9496;
	G5113<= not I9499;
	G5114<= not I9502;
	G5115<= not I9505;
	G5120<= not I9512;
	G5121<= not I9515;
	G5124<= not I9520;
	G5127<= not I9525;
	G5128<= not I9528;
	G5129<= not I9531;
	G5137<= not I9539;
	G5139<= not I9543;
	G5143<= not I9555;
	G5144<= not I9558;
	G5145<= not I9561;
	G5146<= not I9564;
	G5147<= not I9567;
	G5148<= not I9570;
	G5149<= not I9573;
	G5150<= not I9576;
	G5151<= not I9579;
	G5152<= not I9582;
	G5153<= not I9585;
	G5154<= not I9588;
	G5155<= not I9591;
	G5156<= not I9594;
	G5157<= not I9597;
	G5158<= not I9600;
	G5159<= not I9603;
	G5160<= not I9606;
	G5161<= not I9609;
	G5162<= not I9612;
	G5163<= not I9615;
	G5164<= not I9618;
	G5165<= not I9621;
	G5166<= not I9624;
	G5167<= not I9627;
	G5168<= not I9630;
	G5169<= not I9633;
	G5170<= not I9636;
	G5171<= not I9639;
	G5172<= not I9642;
	G5173<= not I9645;
	G5174<= not I9648;
	G5175<= not I9651;
	G5176<= not I9654;
	G5177<= not I9657;
	G5178<= not I9660;
	G5179<= not I9663;
	G5180<= not I9666;
	G5181<= not I9669;
	G5182<= not I9672;
	G5183<= not I9675;
	G5184<= not I9678;
	G5185<= not I9681;
	G5186<= not I9684;
	G5187<= not I9687;
	G5190<= not G4938;
	G5191<= not G4969;
	G5192<= not G4841;
	G5197<= not G4938;
	G5198<= not G4969;
	G5199<= not G4841;
	G5206<= not G4938;
	G5207<= not G4673;
	G5224<= not G5114;
	G5240<= not I9752;
	G5246<= not I9760;
	G5258<= not I9774;
	G5261<= not G4748;
	G5266<= not I9782;
	G5267<= not I9785;
	G5268<= not I9788;
	G5269<= not I9791;
	G5278<= not I9794;
	G5285<= not G4841;
	G5286<= not G4714;
	G5294<= not G5087;
	G5299<= not I9804;
	G5302<= not G5028;
	G5309<= not G4969;
	G5311<= not G4938;
	G5335<= not G4677;
	G5344<= not I9819;
	G5362<= not I9823;
	G5364<= not G5124;
	G5367<= not I9834;
	G5384<= not I9837;
	G5395<= not I9840;
	G5396<= not G4692;
	G5397<= not G5076;
	G5401<= not I9845;
	G5402<= not G5000;
	G5403<= not G5088;
	G5412<= not I9850;
	G5417<= not G5006;
	G5418<= not G5100;
	G5426<= not G5013;
	G5427<= not G5115;
	G5433<= not G5024;
	G5434<= not G5112;
	G5435<= not G5121;
	G5437<= not G5041;
	G5439<= not G5058;
	G5444<= not G5074;
	G5445<= not G5059;
	G5448<= not G5137;
	G5453<= not G4680;
	G5459<= not G4882;
	G5460<= not G4684;
	G5461<= not G4885;
	G5462<= not G4886;
	G5463<= not G5085;
	G5466<= not G4890;
	G5467<= not G4891;
	G5468<= not I9884;
	G5469<= not G4898;
	G5470<= not G4899;
	G5471<= not I9889;
	G5472<= not I9892;
	G5473<= not G4903;
	G5474<= not G4904;
	G5476<= not G4907;
	G5477<= not G4908;
	G5478<= not G5025;
	G5480<= not G4913;
	G5481<= not G4914;
	G5482<= not G4915;
	G5487<= not I9907;
	G5488<= not I9910;
	G5490<= not G4917;
	G5491<= not G4918;
	G5492<= not G4919;
	G5493<= not G4920;
	G5494<= not I9918;
	G5514<= not G4922;
	G5515<= not G4923;
	G5516<= not G4924;
	G5517<= not G4925;
	G5519<= not I9929;
	G5520<= not G4928;
	G5521<= not G4929;
	G5522<= not G4930;
	G5523<= not I9935;
	G5524<= not I9938;
	G5525<= not G4934;
	G5526<= not G5086;
	G5529<= not G4689;
	G5541<= not G4814;
	G5542<= not G5061;
	G5551<= not I9974;
	G5569<= not I10028;
	G5571<= not I10032;
	G5574<= not G4969;
	G5577<= not I10046;
	G5578<= not G4841;
	G5580<= not G4938;
	G5581<= not G4969;
	G5582<= not G4969;
	G5584<= not G4841;
	G5586<= not G4938;
	G5587<= not G4938;
	G5591<= not G4841;
	G5592<= not G4969;
	G5596<= not G4841;
	G5597<= not G4969;
	G5598<= not G4938;
	G5600<= not G5128;
	G5603<= not G4938;
	G5604<= not G4969;
	G5606<= not G4748;
	G5607<= not G4938;
	G5608<= not G4969;
	G5609<= not G4748;
	G5610<= not G4938;
	G5611<= not G4969;
	G5612<= not G4814;
	G5613<= not G4748;
	G5616<= not G4938;
	G5617<= not G4969;
	G5618<= not G5015;
	G5621<= not G4748;
	G5622<= not G4938;
	G5623<= not G4969;
	G5626<= not G4748;
	G5627<= not G4673;
	G5628<= not G4748;
	G5631<= not G4938;
	G5633<= not G4895;
	G5638<= not G4748;
	G5639<= not G4748;
	G5642<= not I10125;
	G5643<= not I10128;
	G5644<= not G4748;
	G5645<= not G4748;
	G5648<= not G4748;
	G5649<= not G4748;
	G5652<= not I10135;
	G5653<= not G4748;
	G5654<= not G4748;
	G5658<= not G4748;
	G5662<= not G5027;
	G5665<= not G4748;
	G5668<= not I10151;
	G5669<= not I10154;
	G5670<= not I10157;
	G5671<= not I10160;
	G5674<= not G5042;
	G5677<= not I10166;
	G5678<= not I10169;
	G5679<= not I10172;
	G5680<= not G5101;
	G5682<= not I10177;
	G5683<= not I10180;
	G5684<= not I10183;
	G5685<= not I10186;
	G5687<= not I10190;
	G5688<= not I10193;
	G5690<= not G4748;
	G5693<= not I10204;
	G5696<= not I10207;
	G5701<= not G5120;
	G5705<= not G4841;
	G5709<= not G4841;
	G5713<= not G4841;
	G5717<= not G4969;
	G5718<= not G4841;
	G5719<= not I10236;
	G5723<= not G4938;
	G5724<= not G4969;
	G5725<= not G4841;
	G5726<= not I10243;
	G5729<= not G5144;
	G5730<= not I10247;
	G5731<= not I10250;
	G5732<= not I10253;
	G5733<= not I10256;
	G5734<= not I10259;
	G5735<= not I10262;
	G5736<= not I10265;
	G5737<= not I10268;
	G5738<= not I10271;
	G5739<= not I10274;
	G5740<= not I10277;
	G5741<= not I10280;
	G5742<= not I10283;
	G5743<= not I10286;
	G5744<= not I10289;
	G5745<= not I10292;
	G5746<= not I10295;
	G5749<= not G5207;
	G5754<= not G5403;
	G5755<= not G5494;
	G5756<= not I10343;
	G5757<= not G5261;
	G5758<= not I10347;
	G5759<= not I10350;
	G5760<= not I10353;
	G5761<= not I10356;
	G5763<= not I10366;
	G5764<= not I10369;
	G5766<= not I10373;
	G5768<= not I10377;
	G5769<= not I10380;
	G5779<= not I10384;
	G5780<= not I10387;
	G5781<= not I10390;
	G5782<= not I10393;
	G5784<= not I10397;
	G5785<= not I10400;
	G5786<= not I10403;
	G5787<= not I10406;
	G5788<= not I10409;
	G5789<= not I10412;
	G5790<= not I10415;
	G5793<= not I10418;
	G5794<= not I10421;
	G5795<= not I10424;
	G5796<= not I10427;
	G5797<= not I10430;
	G5798<= not I10433;
	G5799<= not I10436;
	G5800<= not I10439;
	G5801<= not I10442;
	G5802<= not I10445;
	G5805<= not I10448;
	G5806<= not I10451;
	G5807<= not I10454;
	G5808<= not I10457;
	G5809<= not I10460;
	G5810<= not I10463;
	G5811<= not I10466;
	G5812<= not I10469;
	G5813<= not I10472;
	G5814<= not I10475;
	G5818<= not I10479;
	G5819<= not I10482;
	G5820<= not I10485;
	G5821<= not I10488;
	G5822<= not I10491;
	G5823<= not I10494;
	G5824<= not I10497;
	G5825<= not I10500;
	G5826<= not I10503;
	G5827<= not I10506;
	G5828<= not I10509;
	G5829<= not I10512;
	G5831<= not I10516;
	G5832<= not I10519;
	G5833<= not I10522;
	G5834<= not I10525;
	G5835<= not I10528;
	G5836<= not G5529;
	G5839<= not I10532;
	G5840<= not I10535;
	G5841<= not I10538;
	G5842<= not I10541;
	G5843<= not G5367;
	G5844<= not I10545;
	G5845<= not I10548;
	G5846<= not G5367;
	G5847<= not I10552;
	G5868<= not I10555;
	G5871<= not I10558;
	G5872<= not I10561;
	G5873<= not G5367;
	G5874<= not I10565;
	G5897<= not I10569;
	G5916<= not G5384;
	G5917<= not G5412;
	G5918<= not I10574;
	G5938<= not G5412;
	G5939<= not I10579;
	G5956<= not I10582;
	G5971<= not I10587;
	G5987<= not G5294;
	G5988<= not I10592;
	G6004<= not G5494;
	G6007<= not G5494;
	G6008<= not G5367;
	G6009<= not I10605;
	G6010<= not I10608;
	G6011<= not G5494;
	G6012<= not G5367;
	G6014<= not I10614;
	G6015<= not I10617;
	G6018<= not G5494;
	G6019<= not G5367;
	G6020<= not G5367;
	G6024<= not G5494;
	G6025<= not G5367;
	G6026<= not G5384;
	G6027<= not G5384;
	G6028<= not G5529;
	G6032<= not G5494;
	G6033<= not G5384;
	G6034<= not I10639;
	G6035<= not G5494;
	G6036<= not I10643;
	G6037<= not I10646;
	G6038<= not I10649;
	G6048<= not G5246;
	G6050<= not G5246;
	G6051<= not G5246;
	G6059<= not G5317;
	G6062<= not I10675;
	G6063<= not I10678;
	G6064<= not I10681;
	G6065<= not I10684;
	G6068<= not I10687;
	G6069<= not I10690;
	G6070<= not G5317;
	G6071<= not I10694;
	G6072<= not G5345;
	G6073<= not G5384;
	G6074<= not G5317;
	G6075<= not G5345;
	G6076<= not G5287;
	G6083<= not I10702;
	G6087<= not I10705;
	G6088<= not I10708;
	G6089<= not G5317;
	G6090<= not G5529;
	G6092<= not G5317;
	G6093<= not G5345;
	G6094<= not I10716;
	G6095<= not I10719;
	G6096<= not G5317;
	G6097<= not G5345;
	G6101<= not G5317;
	G6102<= not G5345;
	G6103<= not G5317;
	G6104<= not G5345;
	G6106<= not G5345;
	G6108<= not G5345;
	G6110<= not G5335;
	G6111<= not G5453;
	G6117<= not I10739;
	G6118<= not G5549;
	G6122<= not I10752;
	G6129<= not I10758;
	G6130<= not I10761;
	G6131<= not G5529;
	G6133<= not I10766;
	G6134<= not G5428;
	G6135<= not I10770;
	G6136<= not I10773;
	G6137<= not I10776;
	G6139<= not I10780;
	G6140<= not I10783;
	G6141<= not I10786;
	G6143<= not I10796;
	G6146<= not I10801;
	G6147<= not I10804;
	G6148<= not I10807;
	G6149<= not I10810;
	G6150<= not G5287;
	G6152<= not I10815;
	G6155<= not I10826;
	G6156<= not I10829;
	G6161<= not I10842;
	G6167<= not I10862;
	G6173<= not I10882;
	G6179<= not I10896;
	G6183<= not I10914;
	G6186<= not I10919;
	G6189<= not I10930;
	G6190<= not I10933;
	G6194<= not I10937;
	G6195<= not I10940;
	G6198<= not G5335;
	G6201<= not I10946;
	G6202<= not I10949;
	G6205<= not G5628;
	G6206<= not G5639;
	G6207<= not I10962;
	G6208<= not I10965;
	G6210<= not I10969;
	G6211<= not G5645;
	G6212<= not I10973;
	G6213<= not I10976;
	G6216<= not I10987;
	G6217<= not G5649;
	G6219<= not I10998;
	G6220<= not I11001;
	G6221<= not I11004;
	G6222<= not G5654;
	G6223<= not I11008;
	G6224<= not I11011;
	G6225<= not I11014;
	G6226<= not G5658;
	G6227<= not I11018;
	G6228<= not I11021;
	G6229<= not G5665;
	G6230<= not I11025;
	G6231<= not I11028;
	G6232<= not I11031;
	G6235<= not I11034;
	G6236<= not I11037;
	G6237<= not I11040;
	G6238<= not I11043;
	G6242<= not I11047;
	G6243<= not I11050;
	G6244<= not G5670;
	G6245<= not G5690;
	G6246<= not I11055;
	G6250<= not G5679;
	G6251<= not I11060;
	G6252<= not G5418;
	G6253<= not G5403;
	G6254<= not G5683;
	G6255<= not I11066;
	G6256<= not I11069;
	G6257<= not G5685;
	G6258<= not G5427;
	G6263<= not G5688;
	G6264<= not G5403;
	G6267<= not I11086;
	G6269<= not I11090;
	G6278<= not I11129;
	G6279<= not I11132;
	G6288<= not I11191;
	G6289<= not I11194;
	G6290<= not I11197;
	G6291<= not I11200;
	G6292<= not I11203;
	G6293<= not I11206;
	G6294<= not I11209;
	G6295<= not I11212;
	G6296<= not I11215;
	G6297<= not I11218;
	G6298<= not I11221;
	G6299<= not I11224;
	G6300<= not I11227;
	G6301<= not I11230;
	G6302<= not I11233;
	G6303<= not I11236;
	G6304<= not I11239;
	G6305<= not I11242;
	G6306<= not I11245;
	G6307<= not I11248;
	G6308<= not I11251;
	G6309<= not I11254;
	G6310<= not I11257;
	G6311<= not I11260;
	G6312<= not I11263;
	G6313<= not I11266;
	G6314<= not I11269;
	G6315<= not I11272;
	G6316<= not I11275;
	G6317<= not I11278;
	G6318<= not I11281;
	G6319<= not I11284;
	G6320<= not I11287;
	G6321<= not I11290;
	G6322<= not I11293;
	G6323<= not I11296;
	G6324<= not I11299;
	G6325<= not I11302;
	G6326<= not I11305;
	G6327<= not I11308;
	G6328<= not I11311;
	G6329<= not I11314;
	G6330<= not I11317;
	G6331<= not I11320;
	G6332<= not I11323;
	G6333<= not I11326;
	G6334<= not I11329;
	G6335<= not I11332;
	G6336<= not I11335;
	G6337<= not I11338;
	G6338<= not I11341;
	G6339<= not I11344;
	G6340<= not I11347;
	G6341<= not I11350;
	G6342<= not I11353;
	G6343<= not I11356;
	G6344<= not I11359;
	G6345<= not I11362;
	G6346<= not I11365;
	G6347<= not I11368;
	G6348<= not I11371;
	G6349<= not I11374;
	G6350<= not I11377;
	G6351<= not I11380;
	G6352<= not I11383;
	G6353<= not I11386;
	G6354<= not I11389;
	G6355<= not I11392;
	G6356<= not I11395;
	G6357<= not I11398;
	G6358<= not I11401;
	G6359<= not I11404;
	G6360<= not I11407;
	G6361<= not I11410;
	G6362<= not I11413;
	G6363<= not I11416;
	G6364<= not I11419;
	G6365<= not I11422;
	G6366<= not I11425;
	G6367<= not I11428;
	G6368<= not I11431;
	G6369<= not I11434;
	G6370<= not I11437;
	G6371<= not I11440;
	G6372<= not I11443;
	G6373<= not I11446;
	G6374<= not I11449;
	G6375<= not I11452;
	G6376<= not I11455;
	G6377<= not I11458;
	G6378<= not I11461;
	G6379<= not I11464;
	G6380<= not I11467;
	G6381<= not I11470;
	G6382<= not I11473;
	G6383<= not I11476;
	G6384<= not I11479;
	G6385<= not I11482;
	G6386<= not I11485;
	G6387<= not I11488;
	G6388<= not I11491;
	G6389<= not I11494;
	G6390<= not I11497;
	G6391<= not I11500;
	G6392<= not I11503;
	G6393<= not I11506;
	G6397<= not I11512;
	G6398<= not I11515;
	G6403<= not I11522;
	G6404<= not I11525;
	G6410<= not I11533;
	G6425<= not I11556;
	G6426<= not I11559;
	G6427<= not I11562;
	G6432<= not I11569;
	G6441<= not I11586;
	G6446<= not I11591;
	G6449<= not I11596;
	G6461<= not I11607;
	G6468<= not I11622;
	G6471<= not I11627;
	G6475<= not I11633;
	G6478<= not I11638;
	G6481<= not I11641;
	G6483<= not I11645;
	G6486<= not I11648;
	G6488<= not I11652;
	G6490<= not I11656;
	G6493<= not I11659;
	G6496<= not I11662;
	G6498<= not I11666;
	G6501<= not I11669;
	G6502<= not I11672;
	G6505<= not I11677;
	G6506<= not I11680;
	G6507<= not I11683;
	G6508<= not I11686;
	G6509<= not I11689;
	G6511<= not I11693;
	G6514<= not I11696;
	G6515<= not G6125;
	G6517<= not I11701;
	G6520<= not I11704;
	G6523<= not I11707;
	G6524<= not I11710;
	G6538<= not I11714;
	G6542<= not I11718;
	G6552<= not I11722;
	G6553<= not I11725;
	G6555<= not I11729;
	G6556<= not I11732;
	G6562<= not I11736;
	G6566<= not I11740;
	G6568<= not I11744;
	G6569<= not I11747;
	G6572<= not I11764;
	G6573<= not G5868;
	G6581<= not I11773;
	G6586<= not I11778;
	G6587<= not I11781;
	G6588<= not G5836;
	G6589<= not G6083;
	G6591<= not I11787;
	G6592<= not I11790;
	G6593<= not I11793;
	G6594<= not I11796;
	G6595<= not G6083;
	G6596<= not I11800;
	G6597<= not I11803;
	G6598<= not I11806;
	G6599<= not I11809;
	G6601<= not G6083;
	G6603<= not I11815;
	G6604<= not I11818;
	G6605<= not I11821;
	G6606<= not I11824;
	G6607<= not I11827;
	G6612<= not I11832;
	G6613<= not I11835;
	G6614<= not I11838;
	G6616<= not I11848;
	G6617<= not I11851;
	G6618<= not G6003;
	G6621<= not I11855;
	G6622<= not I11858;
	G6623<= not I11861;
	G6624<= not I11864;
	G6625<= not I11867;
	G6626<= not I11870;
	G6628<= not I11880;
	G6630<= not I11884;
	G6631<= not I11887;
	G6632<= not I11890;
	G6634<= not I11894;
	G6635<= not I11897;
	G6636<= not I11900;
	G6637<= not I11903;
	G6639<= not G6198;
	G6640<= not I11908;
	G6642<= not I11912;
	G6644<= not G6208;
	G6645<= not I11917;
	G6646<= not I11920;
	G6647<= not I11923;
	G6648<= not I11926;
	G6649<= not I11929;
	G6650<= not G6213;
	G6651<= not I11933;
	G6652<= not I11936;
	G6653<= not I11939;
	G6654<= not I11942;
	G6655<= not I11945;
	G6656<= not I11948;
	G6657<= not I11951;
	G6658<= not G6224;
	G6659<= not I11955;
	G6660<= not I11958;
	G6661<= not I11961;
	G6662<= not I11964;
	G6663<= not I11967;
	G6671<= not I11971;
	G6672<= not I11974;
	G6674<= not I11978;
	G6675<= not I11981;
	G6676<= not I11984;
	G6677<= not I11987;
	G6681<= not I11991;
	G6682<= not I11994;
	G6683<= not G6237;
	G6684<= not I11998;
	G6687<= not I12003;
	G6692<= not I12008;
	G6693<= not I12011;
	G6696<= not I12022;
	G6697<= not I12025;
	G6700<= not G6244;
	G6702<= not I12038;
	G6703<= not I12041;
	G6704<= not I12044;
	G6708<= not G6250;
	G6711<= not I12059;
	G6712<= not I12062;
	G6713<= not I12065;
	G6714<= not I12068;
	G6720<= not G6254;
	G6721<= not G6257;
	G6723<= not I12085;
	G6724<= not I12088;
	G6725<= not I12091;
	G6729<= not G6263;
	G6730<= not I12098;
	G6731<= not I12101;
	G6736<= not I12108;
	G6737<= not I12111;
	G6741<= not I12117;
	G6742<= not I12120;
	G6744<= not I12124;
	G6751<= not I12128;
	G6752<= not I12131;
	G6754<= not I12135;
	G6755<= not I12138;
	G6756<= not I12141;
	G6758<= not I12145;
	G6759<= not I12148;
	G6760<= not I12151;
	G6761<= not I12154;
	G6763<= not I12158;
	G6764<= not I12161;
	G6765<= not I12164;
	G6766<= not I12167;
	G6767<= not I12170;
	G6768<= not I12173;
	G6769<= not I12176;
	G6772<= not I12187;
	G6773<= not I12190;
	G6774<= not I12193;
	G6775<= not I12196;
	G6776<= not I12199;
	G6777<= not I12202;
	G6778<= not I12205;
	G6779<= not I12208;
	G6780<= not I12211;
	G6781<= not I12214;
	G6782<= not I12217;
	G6783<= not I12220;
	G6784<= not I12223;
	G6785<= not I12226;
	G6786<= not I12229;
	G6787<= not I12232;
	G6788<= not I12235;
	G6789<= not I12238;
	G6790<= not I12241;
	G6791<= not I12244;
	G6792<= not I12247;
	G6793<= not I12250;
	G6794<= not I12253;
	G6795<= not I12256;
	G6796<= not I12259;
	G6797<= not I12262;
	G6798<= not I12265;
	G6799<= not I12268;
	G6800<= not I12271;
	G6801<= not I12274;
	G6802<= not I12277;
	G6803<= not I12280;
	G6804<= not I12283;
	G6805<= not I12286;
	G6806<= not I12289;
	G6807<= not I12292;
	G6808<= not I12295;
	G6809<= not I12298;
	G6810<= not I12301;
	G6811<= not I12304;
	G6812<= not I12307;
	G6813<= not I12310;
	G6814<= not I12313;
	G6815<= not I12316;
	G6816<= not I12319;
	G6817<= not I12322;
	G6818<= not I12325;
	G6819<= not I12328;
	G6820<= not I12331;
	G6821<= not I12334;
	G6822<= not I12337;
	G6823<= not I12340;
	G6824<= not I12343;
	G6825<= not I12346;
	G6826<= not I12349;
	G6827<= not I12352;
	G6828<= not I12355;
	G6829<= not I12358;
	G6830<= not I12361;
	G6831<= not I12364;
	G6832<= not I12367;
	G6833<= not I12370;
	G6834<= not I12373;
	G6835<= not I12376;
	G6836<= not I12379;
	G6837<= not I12382;
	G6838<= not I12385;
	G6839<= not I12388;
	G6840<= not I12391;
	G6841<= not I12394;
	G6842<= not I12397;
	G6843<= not I12400;
	G6844<= not I12403;
	G6845<= not I12406;
	G6846<= not I12409;
	G6847<= not I12412;
	G6848<= not I12415;
	G6849<= not I12418;
	G6850<= not I12421;
	G6851<= not I12424;
	G6852<= not I12427;
	G6853<= not I12430;
	G6854<= not I12433;
	G6855<= not I12436;
	G6856<= not I12439;
	G6857<= not I12442;
	G6858<= not I12445;
	G6859<= not I12448;
	G6860<= not I12451;
	G6861<= not I12454;
	G6862<= not I12457;
	G6863<= not I12460;
	G6864<= not I12463;
	G6865<= not I12466;
	G6866<= not I12469;
	G6867<= not I12472;
	G6868<= not I12475;
	G6869<= not I12478;
	G6870<= not I12481;
	G6871<= not I12484;
	G6872<= not I12487;
	G6873<= not I12490;
	G6874<= not I12493;
	G6875<= not I12496;
	G6876<= not I12499;
	G6877<= not I12502;
	G6878<= not I12505;
	G6879<= not I12508;
	G6880<= not I12511;
	G6881<= not I12514;
	G6882<= not I12517;
	G6883<= not I12520;
	G6884<= not I12523;
	G6885<= not I12526;
	G6886<= not I12529;
	G6887<= not I12532;
	G6888<= not I12535;
	G6889<= not I12538;
	G6890<= not I12541;
	G6891<= not I12544;
	G6892<= not I12547;
	G6894<= not G6525;
	G6895<= not I12558;
	G6896<= not I12561;
	G6897<= not I12564;
	G6898<= not I12567;
	G6899<= not G6525;
	G6900<= not I12571;
	G6901<= not G6525;
	G6903<= not I12582;
	G6904<= not G6426;
	G6905<= not I12586;
	G6909<= not I12592;
	G6918<= not I12609;
	G6922<= not G6525;
	G6936<= not I12629;
	G6937<= not I12632;
	G6938<= not I12635;
	G6939<= not G6543;
	G6940<= not I12639;
	G6944<= not I12643;
	G6945<= not I12646;
	G6946<= not I12649;
	G6947<= not I12652;
	G6948<= not I12655;
	G6950<= not I12659;
	G6953<= not G6745;
	G6955<= not I12666;
	G6956<= not I12669;
	G6957<= not I12672;
	G6958<= not I12675;
	G6959<= not I12678;
	G6960<= not I12681;
	G6961<= not I12684;
	G6962<= not I12687;
	G6963<= not I12690;
	G6967<= not I12696;
	G6968<= not I12699;
	G6969<= not I12702;
	G6973<= not I12708;
	G6975<= not I12712;
	G6977<= not G6664;
	G6978<= not I12717;
	G6983<= not I12722;
	G6984<= not I12725;
	G6993<= not I12731;
	G6997<= not I12737;
	G7000<= not I12742;
	G7006<= not I12748;
	G7009<= not I12753;
	G7013<= not I12757;
	G7014<= not I12760;
	G7015<= not I12763;
	G7018<= not I12768;
	G7019<= not I12771;
	G7022<= not I12776;
	G7023<= not I12779;
	G7024<= not I12782;
	G7028<= not G6525;
	G7032<= not G6525;
	G7034<= not G6525;
	G7035<= not G6543;
	G7037<= not G6525;
	G7039<= not G6543;
	G7042<= not G6543;
	G7043<= not G6543;
	G7044<= not G6543;
	G7045<= not G6490;
	G7046<= not I12806;
	G7047<= not G6498;
	G7048<= not I12810;
	G7049<= not I12813;
	G7050<= not G6618;
	G7054<= not G6511;
	G7055<= not G6517;
	G7056<= not G6520;
	G7057<= not G6644;
	G7058<= not G6649;
	G7059<= not G6538;
	G7060<= not G6654;
	G7061<= not G6650;
	G7063<= not I12826;
	G7064<= not I12829;
	G7066<= not I12839;
	G7067<= not G6658;
	G7068<= not G6556;
	G7070<= not G6562;
	G7077<= not G6676;
	G7078<= not G6683;
	G7090<= not G6525;
	G7091<= not G6525;
	G7092<= not I12866;
	G7094<= not G6525;
	G7095<= not I12877;
	G7097<= not I12881;
	G7098<= not G6525;
	G7099<= not I12885;
	G7100<= not I12888;
	G7101<= not I12891;
	G7102<= not I12894;
	G7103<= not I12897;
	G7104<= not I12900;
	G7105<= not I12903;
	G7106<= not I12906;
	G7107<= not I12909;
	G7108<= not I12912;
	G7109<= not I12915;
	G7110<= not I12918;
	G7111<= not I12921;
	G7112<= not I12924;
	G7113<= not I12927;
	G7114<= not I12930;
	G7115<= not I12933;
	G7116<= not I12936;
	G7117<= not I12939;
	G7118<= not I12942;
	G7119<= not I12945;
	G7120<= not I12948;
	G7122<= not I12958;
	G7123<= not I12961;
	G7124<= not G6896;
	G7125<= not I12965;
	G7126<= not I12968;
	G7127<= not G6974;
	G7129<= not I12973;
	G7130<= not I12976;
	G7131<= not G6976;
	G7132<= not I12980;
	G7133<= not I12983;
	G7134<= not I12986;
	G7135<= not I12989;
	G7137<= not I12993;
	G7138<= not I12996;
	G7139<= not I12999;
	G7141<= not I13009;
	G7142<= not I13012;
	G7143<= not G6996;
	G7145<= not I13023;
	G7146<= not G6998;
	G7147<= not G6904;
	G7148<= not I13028;
	G7149<= not I13031;
	G7150<= not G6952;
	G7151<= not I13035;
	G7155<= not I13039;
	G7156<= not I13042;
	G7157<= not I13045;
	G7158<= not I13048;
	G7159<= not I13051;
	G7160<= not I13054;
	G7161<= not I13057;
	G7162<= not I13060;
	G7163<= not I13063;
	G7164<= not I13066;
	G7168<= not I13072;
	G7169<= not I13075;
	G7171<= not G7071;
	G7172<= not G7092;
	G7173<= not G6980;
	G7174<= not G7097;
	G7176<= not I13084;
	G7178<= not I13088;
	G7180<= not I13092;
	G7185<= not I13099;
	G7187<= not I13103;
	G7188<= not I13106;
	G7189<= not I13109;
	G7190<= not I13112;
	G7194<= not I13118;
	G7196<= not I13122;
	G7198<= not I13126;
	G7205<= not I13131;
	G7206<= not I13134;
	G7207<= not I13137;
	G7208<= not I13140;
	G7210<= not I13144;
	G7211<= not I13147;
	G7216<= not I13152;
	G7221<= not I13157;
	G7223<= not I13161;
	G7224<= not I13164;
	G7225<= not G6936;
	G7226<= not G6937;
	G7229<= not G6938;
	G7231<= not I13173;
	G7233<= not G6940;
	G7236<= not G6944;
	G7239<= not G6945;
	G7241<= not I13185;
	G7243<= not I13189;
	G7245<= not I13193;
	G7246<= not I13196;
	G7247<= not I13199;
	G7251<= not I13203;
	G7253<= not G7049;
	G7255<= not I13209;
	G7256<= not G7058;
	G7259<= not G7060;
	G7260<= not G7064;
	G7261<= not I13225;
	G7262<= not I13228;
	G7263<= not I13231;
	G7264<= not I13234;
	G7265<= not G7077;
	G7266<= not I13238;
	G7267<= not I13241;
	G7268<= not I13244;
	G7269<= not I13247;
	G7270<= not I13250;
	G7273<= not I13255;
	G7274<= not I13258;
	G7275<= not I13261;
	G7276<= not I13264;
	G7277<= not I13267;
	G7279<= not I13271;
	G7280<= not I13274;
	G7281<= not I13277;
	G7283<= not I13281;
	G7284<= not I13284;
	G7285<= not I13287;
	G7286<= not I13290;
	G7287<= not I13293;
	G7288<= not I13296;
	G7289<= not I13299;
	G7290<= not I13302;
	G7291<= not I13305;
	G7292<= not I13308;
	G7293<= not I13311;
	G7294<= not I13314;
	G7295<= not I13317;
	G7296<= not I13320;
	G7297<= not I13323;
	G7298<= not I13326;
	G7299<= not I13329;
	G7300<= not I13332;
	G7301<= not I13335;
	G7302<= not I13338;
	G7303<= not I13341;
	G7304<= not I13344;
	G7305<= not I13347;
	G7306<= not I13350;
	G7307<= not I13353;
	G7308<= not I13356;
	G7309<= not I13359;
	G7310<= not I13362;
	G7311<= not I13365;
	G7313<= not I13369;
	G7315<= not I13373;
	G7317<= not I13383;
	G7319<= not G7124;
	G7320<= not I13388;
	G7327<= not I13403;
	G7329<= not I13407;
	G7330<= not I13410;
	G7331<= not I13413;
	G7332<= not I13416;
	G7333<= not I13419;
	G7334<= not I13422;
	G7335<= not I13425;
	G7336<= not I13428;
	G7338<= not I13432;
	G7339<= not I13435;
	G7340<= not I13438;
	G7341<= not I13441;
	G7342<= not I13444;
	G7343<= not I13447;
	G7344<= not G7150;
	G7345<= not I13451;
	G7346<= not I13454;
	G7347<= not I13457;
	G7348<= not I13460;
	G7349<= not I13463;
	G7350<= not I13466;
	G7351<= not I13469;
	G7352<= not I13472;
	G7353<= not I13475;
	G7354<= not I13478;
	G7355<= not I13481;
	G7356<= not I13484;
	G7357<= not I13487;
	G7358<= not I13490;
	G7359<= not I13493;
	G7360<= not I13496;
	G7361<= not I13499;
	G7362<= not I13502;
	G7364<= not I13506;
	G7365<= not I13509;
	G7366<= not I13512;
	G7367<= not I13515;
	G7405<= not I13518;
	G7411<= not G7202;
	G7413<= not I13524;
	G7414<= not I13527;
	G7418<= not I13533;
	G7420<= not I13537;
	G7422<= not I13541;
	G7423<= not I13544;
	G7424<= not I13547;
	G7425<= not I13550;
	G7432<= not I13559;
	G7433<= not I13562;
	G7434<= not I13565;
	G7437<= not I13570;
	G7439<= not I13574;
	G7440<= not I13577;
	G7441<= not I13580;
	G7442<= not I13583;
	G7446<= not I13595;
	G7448<= not I13605;
	G7454<= not I13610;
	G7455<= not I13613;
	G7456<= not G7174;
	G7459<= not I13617;
	G7460<= not G7172;
	G7463<= not G7239;
	G7466<= not I13622;
	G7467<= not G7236;
	G7470<= not G7253;
	G7471<= not G7233;
	G7474<= not I13628;
	G7475<= not I13631;
	G7476<= not G7229;
	G7479<= not I13635;
	G7483<= not G7226;
	G7486<= not I13646;
	G7487<= not I13649;
	G7488<= not G7225;
	G7491<= not I13653;
	G7492<= not I13656;
	G7493<= not I13659;
	G7494<= not G7260;
	G7495<= not I13663;
	G7496<= not I13666;
	G7497<= not I13669;
	G7498<= not I13672;
	G7499<= not G7258;
	G7500<= not I13676;
	G7501<= not I13679;
	G7502<= not I13682;
	G7504<= not I13692;
	G7505<= not I13695;
	G7506<= not I13698;
	G7507<= not I13701;
	G7508<= not I13704;
	G7509<= not I13707;
	G7510<= not I13710;
	G7511<= not I13713;
	G7512<= not I13716;
	G7513<= not I13719;
	G7514<= not I13722;
	G7515<= not I13725;
	G7516<= not I13728;
	G7517<= not I13731;
	G7518<= not I13734;
	G7519<= not I13737;
	G7520<= not I13740;
	G7521<= not I13743;
	G7522<= not I13746;
	G7523<= not I13749;
	G7524<= not I13752;
	G7525<= not I13755;
	G7526<= not I13758;
	G7527<= not I13761;
	G7528<= not I13764;
	G7529<= not I13767;
	G7530<= not I13770;
	G7531<= not I13773;
	G7532<= not I13776;
	G7533<= not I13779;
	G7534<= not I13782;
	G7538<= not I13794;
	G7539<= not I13797;
	G7541<= not I13807;
	G7542<= not I13810;
	G7543<= not I13813;
	G7544<= not I13816;
	G7545<= not I13819;
	G7546<= not I13822;
	G7547<= not I13825;
	G7548<= not I13828;
	G7549<= not I13831;
	G7550<= not I13834;
	G7551<= not I13837;
	G7555<= not I13843;
	G7556<= not I13846;
	G7558<= not I13850;
	G7560<= not I13854;
	G7562<= not I13858;
	G7563<= not I13861;
	G7565<= not I13865;
	G7574<= not I13869;
	G7576<= not I13873;
	G7577<= not I13876;
	G7578<= not I13879;
	G7579<= not I13882;
	G7580<= not I13885;
	G7581<= not I13888;
	G7582<= not I13891;
	G7583<= not I13894;
	G7584<= not I13897;
	G7585<= not I13900;
	G7586<= not I13903;
	G7587<= not I13906;
	G7588<= not I13909;
	G7589<= not I13912;
	G7590<= not I13915;
	G7591<= not I13918;
	G7592<= not I13921;
	G7593<= not I13924;
	G7594<= not I13927;
	G7595<= not I13930;
	G7599<= not G7450;
	G7601<= not G7450;
	G7603<= not I13940;
	G7610<= not G7450;
	G7627<= not I13956;
	G7633<= not I13962;
	G7686<= not I13979;
	G7688<= not G7406;
	G7702<= not I13997;
	G7704<= not I14001;
	G7708<= not I14005;
	G7710<= not I14009;
	G7711<= not I14012;
	G7712<= not I14015;
	G7714<= not I14019;
	G7715<= not I14022;
	G7716<= not I14025;
	G7717<= not I14028;
	G7718<= not I14031;
	G7719<= not G7475;
	G7720<= not I14035;
	G7721<= not G7344;
	G7722<= not I14039;
	G7723<= not I14042;
	G7725<= not I14046;
	G7726<= not I14049;
	G7727<= not I14052;
	G7728<= not I14055;
	G7729<= not I14058;
	G7730<= not I14061;
	G7731<= not I14064;
	G7732<= not I14067;
	G7733<= not I14070;
	G7734<= not I14073;
	G7735<= not I14076;
	G7736<= not I14079;
	G7737<= not I14082;
	G7738<= not I14085;
	G7739<= not I14088;
	G7740<= not I14091;
	G7741<= not I14094;
	G7742<= not I14097;
	G7743<= not I14100;
	G7744<= not I14103;
	G7745<= not I14106;
	G7746<= not I14109;
	G7747<= not I14112;
	G7748<= not I14115;
	G7749<= not I14118;
	G7750<= not I14121;
	G7751<= not I14124;
	G7752<= not I14127;
	G7753<= not I14130;
	G7754<= not I14133;
	G7755<= not I14136;
	G7756<= not I14139;
	G7757<= not I14142;
	G7758<= not I14145;
	G7759<= not I14148;
	G7760<= not I14151;
	G7761<= not I14154;
	G7762<= not I14157;
	G7763<= not I14160;
	G7764<= not I14163;
	G7765<= not I14166;
	G7766<= not I14169;
	G7767<= not I14172;
	G7768<= not I14175;
	G7769<= not I14178;
	G7770<= not I14181;
	G7771<= not I14184;
	G7772<= not I14187;
	G7773<= not I14190;
	G7774<= not I14193;
	G7775<= not I14196;
	G7776<= not I14199;
	G7777<= not I14202;
	G7778<= not I14205;
	G7779<= not I14208;
	G7780<= not I14211;
	G7781<= not I14214;
	G7789<= not I14224;
	G7790<= not I14227;
	G7792<= not I14231;
	G7793<= not I14234;
	G7811<= not I14238;
	G7829<= not I14251;
	G7835<= not I14257;
	G7836<= not I14260;
	G7838<= not I14264;
	G7855<= not I14267;
	G7870<= not I14270;
	G7887<= not I14273;
	G7904<= not I14276;
	G7905<= not I14279;
	G7920<= not I14282;
	G7937<= not I14285;
	G7951<= not I14288;
	G7966<= not I14291;
	G7983<= not I14294;
	G7992<= not G7557;
	G7993<= not I14298;
	G8008<= not G7559;
	G8012<= not I14305;
	G8013<= not G7561;
	G8014<= not G7564;
	G8015<= not G7689;
	G8016<= not I14311;
	G8017<= not G7692;
	G8018<= not I14315;
	G8029<= not I14318;
	G8038<= not G7694;
	G8039<= not G7696;
	G8040<= not G7699;
	G8041<= not G7701;
	G8042<= not I14325;
	G8061<= not I14330;
	G8063<= not I14334;
	G8065<= not I14338;
	G8067<= not I14342;
	G8072<= not I14349;
	G8093<= not I14370;
	G8094<= not G7705;
	G8111<= not I14374;
	G8131<= not I14378;
	G8145<= not I14381;
	G8152<= not I14388;
	G8156<= not I14394;
	G8172<= not I14397;
	G8173<= not I14400;
	G8174<= not I14403;
	G8175<= not I14406;
	G8177<= not I14410;
	G8178<= not I14413;
	G8179<= not I14416;
	G8180<= not G7719;
	G8181<= not I14420;
	G8198<= not G7721;
	G8199<= not I14424;
	G8216<= not I14427;
	G8217<= not I14430;
	G8218<= not I14433;
	G8219<= not I14436;
	G8220<= not I14439;
	G8221<= not I14442;
	G8222<= not I14445;
	G8223<= not I14448;
	G8224<= not I14451;
	G8225<= not I14454;
	G8226<= not I14457;
	G8227<= not I14460;
	G8228<= not I14463;
	G8234<= not I14489;
	G8235<= not I14492;
	G8284<= not I14531;
	G8324<= not I14573;
	G8342<= not G8008;
	G8363<= not G7992;
	G8381<= not I14603;
	G8386<= not G8014;
	G8406<= not I14614;
	G8407<= not G8013;
	G8421<= not G8017;
	G8442<= not I14623;
	G8443<= not G8015;
	G8463<= not G8094;
	G8464<= not G8039;
	G8481<= not I14637;
	G8482<= not G8094;
	G8483<= not G8038;
	G8493<= not G8041;
	G8510<= not I14643;
	G8511<= not I14646;
	G8512<= not G8094;
	G8514<= not G8040;
	G8524<= not G7855;
	G8541<= not G8094;
	G8544<= not I14657;
	G8545<= not G7905;
	G8562<= not G8094;
	G8563<= not I14662;
	G8564<= not G7951;
	G8581<= not G8094;
	G8582<= not G8094;
	G8583<= not I14668;
	G8585<= not G7993;
	G8602<= not G8094;
	G8603<= not I14674;
	G8604<= not I14677;
	G8605<= not I14680;
	G8606<= not I14683;
	G8608<= not I14687;
	G8619<= not I14695;
	G8631<= not I14709;
	G8632<= not I14712;
	G8636<= not I14718;
	G8638<= not I14722;
	G8639<= not I14725;
	G8640<= not I14728;
	G8642<= not I14732;
	G8647<= not I14739;
	G8649<= not I14743;
	G8651<= not I14747;
	G8657<= not I14763;
	G8661<= not I14777;
	G8662<= not I14780;
	G8663<= not I14783;
	G8664<= not I14786;
	G8665<= not I14789;
	G8666<= not I14792;
	G8667<= not I14795;
	G8668<= not I14798;
	G8669<= not I14801;
	G8670<= not I14804;
	G8671<= not I14807;
	G8672<= not I14810;
	G8673<= not I14813;
	G8674<= not I14816;
	G8675<= not I14819;
	G8676<= not I14822;
	G8677<= not I14825;
	G8678<= not I14828;
	G8682<= not I14844;
	G8683<= not G8235;
	G8684<= not I14848;
	G8685<= not I14851;
	G8689<= not I14857;
	G8734<= not I14904;
	G8743<= not G8524;
	G8746<= not G8524;
	G8747<= not G8545;
	G8750<= not G8524;
	G8751<= not G8545;
	G8752<= not G8564;
	G8753<= not I14925;
	G8754<= not G8524;
	G8755<= not G8545;
	G8756<= not G8564;
	G8757<= not G8585;
	G8759<= not G8524;
	G8760<= not G8545;
	G8761<= not G8564;
	G8762<= not G8585;
	G8765<= not G8524;
	G8766<= not G8545;
	G8767<= not G8564;
	G8768<= not G8585;
	G8770<= not G8545;
	G8771<= not G8564;
	G8772<= not G8585;
	G8774<= not I14964;
	G8775<= not G8564;
	G8776<= not G8585;
	G8778<= not I14974;
	G8780<= not G8524;
	G8781<= not G8585;
	G8783<= not G8524;
	G8784<= not G8545;
	G8786<= not G8545;
	G8787<= not G8564;
	G8789<= not G8564;
	G8790<= not G8585;
	G8791<= not G8585;
	G8792<= not I14996;
	G8797<= not I15003;
	G8799<= not I15007;
	G8800<= not I15010;
	G8802<= not I15014;
	G8808<= not I15062;
	G8809<= not I15065;
	G8810<= not I15068;
	G8856<= not I15160;
	G8864<= not I15178;
	G8865<= not I15181;
	G8866<= not I15184;
	G8867<= not I15187;
	G8868<= not I15190;
	G8869<= not I15193;
	G8870<= not I15196;
	G8871<= not I15199;
	G8872<= not I15202;
	G8873<= not I15205;
	G8874<= not I15208;
	G8875<= not I15211;
	G8880<= not I15218;
	G8881<= not G8683;
	G8882<= not I15222;
	G8883<= not I15225;
	G8898<= not I15308;
	G8903<= not I15315;
	G8910<= not I15324;
	G8913<= not I15329;
	G8916<= not I15334;
	G8917<= not I15337;
	G8918<= not I15340;
	G8955<= not I15379;
	G8956<= not I15382;
	G8957<= not I15385;
	G8958<= not I15388;
	G8959<= not I15391;
	G8960<= not I15394;
	G8967<= not I15405;
	G8968<= not I15408;
	G8969<= not I15411;
	G8970<= not I15414;
	G8971<= not I15417;
	G8972<= not I15420;
	G8973<= not I15423;
	G8974<= not I15426;
	G8975<= not I15429;
	G8977<= not I15433;
	G9017<= not I15475;
	G9018<= not I15478;
	G9019<= not I15481;
	G9020<= not I15484;
	G9026<= not I15492;
	G9027<= not I15495;
	G9028<= not I15498;
	G9029<= not I15501;
	G9030<= not I15504;
	G9031<= not I15507;
	G9032<= not I15510;
	G9033<= not I15513;
	G9034<= not I15516;
	G9035<= not I15519;
	G9036<= not I15522;
	G9039<= not I15527;
	G9042<= not I15530;
	G9043<= not I15533;
	G9044<= not I15536;
	G9045<= not I15539;
	G9047<= not I15543;
	G9048<= not I15546;
	G9050<= not I15550;
	G9051<= not I15553;
	G9053<= not I15557;
	G9056<= not I15562;
	G9057<= not I15565;
	G9058<= not I15568;
	G9059<= not I15571;
	G9060<= not I15574;
	G9061<= not I15577;
	G9062<= not I15580;
	G9063<= not I15583;
	G9064<= not I15586;
	G9065<= not I15589;
	G9066<= not I15592;
	G9067<= not I15595;
	G9068<= not I15598;
	G9069<= not I15601;
	G9070<= not I15604;
	G9071<= not I15607;
	G9072<= not I15610;
	G9073<= not I15613;
	G9074<= not I15616;
	G9075<= not I15619;
	G9076<= not I15622;
	G9077<= not I15625;
	G9078<= not I15628;
	G9079<= not I15631;
	G9081<= not I15635;
	G9082<= not I15638;
	G9083<= not I15641;
	G9085<= not I15645;
	G9086<= not I15648;
	G9087<= not I15651;
	G9088<= not I15654;
	G9089<= not I15657;
	G9090<= not I15660;
	G9091<= not I15663;
	G9092<= not I15666;
	G9093<= not I15669;
	G9094<= not I15672;
	G9095<= not I15675;
	G9096<= not I15678;
	G9097<= not I15681;
	G9098<= not I15684;
	G9099<= not I15687;
	G9100<= not I15690;
	G9101<= not I15693;
	G9102<= not I15696;
	G9103<= not I15699;
	G9104<= not I15702;
	G9105<= not I15705;
	G9106<= not I15708;
	G9107<= not I15711;
	G9108<= not I15714;
	G9109<= not I15717;
	G9110<= not I15720;
	G9111<= not I15723;
	G9112<= not I15726;
	G9113<= not I15729;
	G9114<= not I15732;
	G9115<= not I15735;
	G9116<= not I15738;
	G9117<= not I15741;
	G9121<= not I15747;
	G9125<= not I15753;
	G9126<= not I15756;
	G9127<= not I15759;
	G9128<= not I15762;
	G9129<= not I15765;
	G9132<= not I15770;
	G9133<= not I15773;
	G9134<= not I15776;
	G9140<= not I15784;
	G9141<= not G9129;
	G9145<= not I15791;
	G9157<= not G9141;
	G9161<= not I15803;
	G9177<= not I15811;
	G9178<= not I15814;
	G9180<= not I15824;
	G9181<= not G9177;
	G9182<= not G9178;
	G9183<= not G9161;
	G9184<= not I15830;
	G9185<= not I15833;
	G9186<= not I15836;
	G9187<= not I15839;
	G9188<= not I15842;
	G9189<= not I15845;
	G9193<= not G9181;
	G9194<= not G9182;
	G9195<= not I15871;
	G9196<= not G9185;
	G9197<= not G9186;
	G9198<= not G9187;
	G9199<= not G9188;
	G9200<= not G9189;
	G9201<= not G9183;
	G9204<= not I15894;
	G9206<= not G9196;
	G9207<= not G9197;
	G9208<= not G9198;
	G9209<= not G9199;
	G9210<= not G9200;
	G9211<= not I15909;
	G9212<= not I15912;
	G9213<= not I15915;
	G9214<= not I15918;
	G9215<= not I15921;
	G9216<= not I15924;
	G9217<= not I15927;
	G9218<= not I15930;
	G9219<= not I15933;
	G9220<= not G9205;
	G9221<= not I15937;
	G9222<= not I15940;
	G9223<= not I15943;
	G9227<= not I15947;
	G9230<= not I15950;
	G9233<= not I15953;
	G9234<= not I15956;
	G9235<= not I15959;
	G9236<= not I15962;
	G9237<= not I15965;
	G9241<= not I15971;
	G9244<= not I15974;
	G9248<= not I15978;
	G9252<= not I15982;
	G9255<= not I15985;
	G9260<= not I15990;
	G9280<= not I16006;
	G9281<= not I16009;
	G9297<= not I16017;
	G9298<= not I16020;
	G9299<= not I16023;
	G9300<= not I16026;
	G9301<= not G9260;
	G9302<= not G9281;
	G9303<= not G9301;
	G9304<= not G9298;
	G9305<= not I16033;
	G9306<= not I16036;
	G9307<= not G9300;
	G9308<= not I16040;
	G9309<= not I16043;
	G9310<= not I16046;
	G9311<= not I16049;
	G9312<= not I16052;
	G9313<= not I16055;
	G9314<= not I16058;
	G9315<= not I16061;
	G9316<= not G9302;
	G9317<= not G9306;
	G9318<= not G9304;
	G9319<= not G9309;
	G9320<= not G9307;
	G9321<= not G9311;
	G9322<= not G9313;
	G9323<= not G9315;
	G9324<= not I16072;
	G9329<= not G9317;
	G9330<= not G9319;
	G9331<= not G9321;
	G9332<= not G9322;
	G9333<= not G9323;
	G9336<= not I16084;
	G9340<= not I16090;
	G9350<= not I16100;
	G9351<= not I16103;
	G9353<= not I16107;
	G9360<= not I16116;
	G9361<= not I16119;
	G9362<= not I16122;
	G9366<= not I16126;
	G9367<= not I16129;
	G9368<= not I16132;
	G9369<= not I16135;
	G9370<= not I16138;
	G9372<= not I16142;
	G9373<= not I16145;
	G9374<= not I16148;
	G9375<= not I16151;
	G9376<= not I16154;
	G9378<= not I16158;
	G9379<= not I16161;
	G9380<= not G9379;
	G9381<= not I16165;
	G9382<= not I16168;
	G9383<= not G9380;
	G9385<= not I16173;
	G9386<= not I16176;
	G9388<= not I16180;
	G9389<= not I16183;
	I5353<= not G3833;
	I5356<= not G3837;
	I5359<= not G3839;
	I5362<= not G3841;
	I5365<= not G3843;
	I5368<= not G3853;
	I5371<= not G633;
	I5374<= not G634;
	I5377<= not G635;
	I5380<= not G645;
	I5383<= not G647;
	I5386<= not G648;
	I5389<= not G690;
	I5392<= not G694;
	I5395<= not G698;
	I5398<= not G702;
	I5401<= not G723;
	I5404<= not G722;
	I5407<= not G4653;
	I5410<= not G8866;
	I5413<= not G1016;
	I5416<= not G8868;
	I5419<= not G1603;
	I5422<= not G1234;
	I5425<= not G1245;
	I5428<= not G49;
	I5432<= not G1176;
	I5435<= not G1461;
	I5466<= not G926;
	I5471<= not G1029;
	I5475<= not G1084;
	I5478<= not G1148;
	I5512<= not G557;
	I5515<= not G567;
	I5528<= not G43;
	I5531<= not G866;
	I5535<= not G48;
	I5542<= not G1272;
	I5545<= not G1276;
	I5548<= not G1280;
	I5552<= not G1284;
	I5555<= not G1288;
	I5559<= not G1292;
	I5562<= not G1300;
	I5565<= not G1296;
	I5568<= not G1409;
	I5577<= not G172;
	I5605<= not G58;
	I5609<= not G16;
	I5616<= not G979;
	I5633<= not G891;
	I5636<= not G891;
	I5646<= not G883;
	I5649<= not G1389;
	I5654<= not G921;
	I5657<= not G921;
	I5664<= not G916;
	I5667<= not G916;
	I5670<= not G941;
	I5676<= not G911;
	I5679<= not G911;
	I5682<= not G168;
	I5689<= not G906;
	I5692<= not G906;
	I5706<= not G901;
	I5709<= not G901;
	I5715<= not G896;
	I5718<= not G896;
	I5732<= not G859;
	I5747<= not G1260;
	I5751<= not G963;
	I5754<= not G966;
	I5763<= not G1207;
	I5766<= not G1254;
	I5772<= not G1240;
	I5775<= not G1240;
	I5781<= not G979;
	I5789<= not G1524;
	I5795<= not G1236;
	I5801<= not G1424;
	I5812<= not G1243;
	I5817<= not G1081;
	I5831<= not G1194;
	I5839<= not G1198;
	I5842<= not G68;
	I5847<= not G1360;
	I5852<= not G1202;
	I5855<= not G71;
	I5861<= not G1313;
	I5865<= not G1206;
	I5868<= not G74;
	I5872<= not G77;
	I5879<= not G1267;
	I5883<= not G80;
	I5889<= not G83;
	I5894<= not G86;
	I5897<= not G173;
	I5901<= not G52;
	I5908<= not G196;
	I5911<= not G216;
	I5914<= not G1097;
	I5920<= not G219;
	I5923<= not G252;
	I5926<= not G297;
	I5933<= not G1158;
	I5936<= not G222;
	I5939<= not G275;
	I5942<= not G300;
	I5945<= not G333;
	I5948<= not G378;
	I5954<= not G89;
	I5957<= not G110;
	I5960<= not G187;
	I5963<= not G225;
	I5966<= not G278;
	I5969<= not G303;
	I5972<= not G356;
	I5975<= not G381;
	I5978<= not G414;
	I5981<= not G459;
	I5984<= not G540;
	I5989<= not G1460;
	I5997<= not G114;
	I6000<= not G202;
	I6003<= not G228;
	I6006<= not G306;
	I6009<= not G359;
	I6012<= not G384;
	I6015<= not G437;
	I6018<= not G462;
	I6021<= not G495;
	I6024<= not G544;
	I6029<= not G1207;
	I6033<= not G3;
	I6036<= not G130;
	I6039<= not G207;
	I6042<= not G237;
	I6045<= not G309;
	I6048<= not G387;
	I6051<= not G440;
	I6054<= not G465;
	I6057<= not G518;
	I6060<= not G580;
	I6072<= not G1211;
	I6075<= not G2;
	I6078<= not G95;
	I6081<= not G118;
	I6084<= not G240;
	I6087<= not G318;
	I6090<= not G390;
	I6093<= not G468;
	I6096<= not G521;
	I6099<= not G584;
	I6109<= not G1214;
	I6112<= not G4;
	I6115<= not G134;
	I6118<= not G243;
	I6121<= not G321;
	I6124<= not G399;
	I6127<= not G471;
	I6130<= not G560;
	I6143<= not G1217;
	I6148<= not G5;
	I6151<= not G12;
	I6154<= not G122;
	I6157<= not G246;
	I6160<= not G324;
	I6163<= not G402;
	I6166<= not G480;
	I6178<= not G1220;
	I6183<= not G6;
	I6186<= not G138;
	I6189<= not G249;
	I6192<= not G327;
	I6195<= not G405;
	I6198<= not G483;
	I6214<= not G7;
	I6217<= not G105;
	I6220<= not G126;
	I6223<= not G330;
	I6226<= not G408;
	I6229<= not G486;
	I6239<= not G8;
	I6242<= not G1554;
	I6245<= not G142;
	I6248<= not G411;
	I6251<= not G489;
	I6254<= not G536;
	I6267<= not G100;
	I6270<= not G492;
	I6286<= not G1307;
	I6291<= not G46;
	I6294<= not G1330;
	I6299<= not G47;
	I6302<= not G1313;
	I6305<= not G1333;
	I6309<= not G1336;
	I6317<= not G1339;
	I6323<= not G1342;
	I6326<= not G1443;
	I6333<= not G1345;
	I6337<= not G1348;
	I6341<= not G1351;
	I6348<= not G1354;
	I6354<= not G1357;
	I6358<= not G13;
	I6363<= not G16;
	I6368<= not G20;
	I6371<= not G33;
	I6376<= not G38;
	I6416<= not G1794;
	I6419<= not G1799;
	I6422<= not G1805;
	I6425<= not G1811;
	I6428<= not G1818;
	I6431<= not G1825;
	I6434<= not G1830;
	I6437<= not G1784;
	I6440<= not G1806;
	I6443<= not G1774;
	I6446<= not G1812;
	I6451<= not G1895;
	I6454<= not G1868;
	I6457<= not G1886;
	I6460<= not G2104;
	I6463<= not G1769;
	I6468<= not G1917;
	I6471<= not G1923;
	I6474<= not G1941;
	I6509<= not G1684;
	I6517<= not G1687;
	I6532<= not G1694;
	I6553<= not G2246;
	I6561<= not G1715;
	I6564<= not G2073;
	I6571<= not G1711;
	I6574<= not G576;
	I6578<= not G1603;
	I6587<= not G1708;
	I6590<= not G2467;
	I6597<= not G1970;
	I6608<= not G1612;
	I6615<= not G1983;
	I6629<= not G2052;
	I6636<= not G1704;
	I6643<= not G1970;
	I6646<= not G2246;
	I6652<= not G2016;
	I6657<= not G1701;
	I6663<= not G2246;
	I6669<= not G1698;
	I6673<= not G2246;
	I6676<= not G1603;
	I6680<= not G1558;
	I6686<= not G2246;
	I6695<= not G2246;
	I6703<= not G1983;
	I6711<= not G1726;
	I6716<= not G1721;
	I6723<= not G2052;
	I6728<= not G1959;
	I6733<= not G1718;
	I6764<= not G1955;
	I6767<= not G1933;
	I6770<= not G1590;
	I6784<= not G2052;
	I6788<= not G1681;
	I6791<= not G1967;
	I6795<= not G1683;
	I6800<= not G2016;
	I6805<= not G1603;
	I6820<= not G1707;
	I6826<= not G2185;
	I6831<= not G2185;
	I6834<= not G287;
	I6839<= not G2185;
	I6849<= not G368;
	I6853<= not G2185;
	I6856<= not G449;
	I6860<= not G2185;
	I6864<= not G2528;
	I6868<= not G530;
	I6872<= not G2185;
	I6887<= not G2528;
	I6894<= not G1863;
	I6900<= not G1866;
	I6911<= not G1869;
	I6930<= not G1876;
	I6936<= not G1878;
	I6946<= not G1887;
	I6949<= not G2148;
	I6952<= not G1896;
	I6956<= not G1907;
	I6959<= not G1558;
	I6963<= not G1558;
	I6970<= not G1872;
	I6974<= not G2528;
	I7029<= not G2392;
	I7036<= not G2454;
	I7041<= not G2401;
	I7044<= not G2402;
	I7053<= not G2452;
	I7061<= not G2457;
	I7064<= not G2458;
	I7079<= not G2532;
	I7082<= not G2470;
	I7095<= not G2539;
	I7098<= not G2477;
	I7101<= not G2478;
	I7104<= not G2479;
	I7107<= not G2480;
	I7112<= not G2546;
	I7115<= not G2547;
	I7118<= not G2484;
	I7126<= not G2494;
	I7129<= not G2495;
	I7132<= not G2554;
	I7145<= not G2501;
	I7164<= not G2157;
	I7167<= not G2505;
	I7195<= not G1795;
	I7198<= not G2509;
	I7204<= not G2520;
	I7211<= not G1742;
	I7255<= not G1955;
	I7262<= not G2514;
	I7287<= not G2561;
	I7290<= not G2936;
	I7293<= not G2955;
	I7296<= not G2915;
	I7299<= not G2961;
	I7302<= not G2825;
	I7305<= not G3048;
	I7308<= not G3074;
	I7311<= not G2879;
	I7314<= not G2916;
	I7317<= not G2893;
	I7320<= not G2927;
	I7323<= not G2905;
	I7326<= not G2940;
	I7329<= not G2920;
	I7332<= not G2947;
	I7335<= not G2910;
	I7338<= not G2923;
	I7341<= not G2931;
	I7344<= not G2964;
	I7347<= not G2985;
	I7350<= not G2971;
	I7353<= not G2833;
	I7356<= not G2843;
	I7359<= not G2871;
	I7362<= not G2933;
	I7365<= not G3061;
	I7368<= not G3018;
	I7371<= not G3050;
	I7374<= not G3084;
	I7377<= not G3189;
	I7380<= not G3461;
	I7383<= not G3465;
	I7386<= not G3013;
	I7389<= not G3496;
	I7392<= not G3230;
	I7400<= not G3075;
	I7417<= not G3659;
	I7473<= not G3546;
	I7492<= not G3561;
	I7495<= not G3562;
	I7498<= not G2752;
	I7517<= not G3578;
	I7520<= not G2734;
	I7523<= not G2562;
	I7526<= not G2752;
	I7545<= not G3589;
	I7548<= not G3590;
	I7551<= not G2712;
	I7554<= not G2573;
	I7558<= not G2734;
	I7561<= not G2562;
	I7564<= not G2752;
	I7581<= not G3612;
	I7584<= not G3062;
	I7588<= not G2584;
	I7592<= not G2712;
	I7595<= not G2573;
	I7599<= not G2734;
	I7602<= not G2562;
	I7605<= not G2752;
	I7623<= not G3631;
	I7626<= not G3632;
	I7629<= not G3633;
	I7632<= not G3634;
	I7635<= not G3052;
	I7640<= not G3062;
	I7644<= not G2584;
	I7648<= not G2712;
	I7651<= not G2573;
	I7655<= not G2734;
	I7658<= not G2562;
	I7662<= not G3642;
	I7667<= not G3052;
	I7672<= not G3062;
	I7676<= not G2584;
	I7680<= not G2712;
	I7683<= not G2573;
	I7688<= not G3650;
	I7691<= not G3651;
	I7697<= not G3052;
	I7702<= not G3062;
	I7706<= not G2584;
	I7712<= not G3657;
	I7716<= not G3038;
	I7723<= not G3052;
	I7728<= not G3675;
	I7731<= not G3029;
	I7734<= not G2595;
	I7738<= not G3038;
	I7746<= not G3591;
	I7749<= not G3692;
	I7752<= not G3591;
	I7755<= not G3019;
	I7758<= not G2605;
	I7762<= not G3029;
	I7765<= not G2595;
	I7769<= not G3038;
	I7775<= not G3705;
	I7778<= not G3019;
	I7781<= not G2605;
	I7785<= not G3029;
	I7788<= not G2595;
	I7792<= not G3038;
	I7797<= not G3019;
	I7800<= not G2605;
	I7804<= not G3029;
	I7807<= not G2595;
	I7811<= not G3019;
	I7814<= not G2605;
	I7832<= not G2768;
	I7838<= not G2781;
	I7844<= not G3784;
	I7847<= not G3798;
	I7850<= not G2795;
	I7856<= not G3805;
	I7859<= not G2804;
	I7864<= not G3812;
	I7867<= not G2818;
	I7870<= not G2827;
	I7875<= not G3819;
	I7878<= not G2829;
	I7882<= not G2700;
	I7885<= not G2837;
	I7888<= not G3505;
	I7899<= not G3743;
	I7902<= not G2709;
	I7905<= not G2863;
	I7908<= not G3516;
	I7911<= not G2767;
	I7919<= not G3761;
	I7922<= not G3462;
	I7925<= not G2761;
	I7928<= not G2873;
	I7931<= not G2780;
	I7944<= not G3774;
	I7947<= not G3485;
	I7950<= not G2774;
	I7953<= not G3542;
	I7956<= not G2810;
	I7959<= not G2793;
	I7964<= not G3488;
	I7967<= not G2787;
	I7970<= not G3557;
	I7973<= not G3071;
	I7978<= not G3574;
	I7981<= not G3555;
	I7987<= not G3528;
	I8011<= not G3225;
	I8024<= not G3076;
	I8084<= not G3706;
	I8094<= not G2976;
	I8097<= not G3237;
	I8101<= not G3259;
	I8105<= not G3339;
	I8140<= not G3429;
	I8161<= not G3517;
	I8172<= not G3524;
	I8177<= not G2810;
	I8180<= not G3529;
	I8190<= not G3545;
	I8193<= not G3547;
	I8196<= not G3654;
	I8202<= not G3560;
	I8205<= not G2655;
	I8215<= not G3577;
	I8218<= not G3002;
	I8233<= not G3588;
	I8261<= not G3643;
	I8264<= not G3653;
	I8268<= not G2801;
	I8273<= not G2976;
	I8277<= not G3504;
	I8282<= not G3515;
	I8291<= not G878;
	I8308<= not G3674;
	I8315<= not G3691;
	I8333<= not G3721;
	I8351<= not G1160;
	I8354<= not G1163;
	I8357<= not G1182;
	I8360<= not G1186;
	I8373<= not G3783;
	I8428<= not G3611;
	I8446<= not G3014;
	I8449<= not G3630;
	I8452<= not G2816;
	I8477<= not G3014;
	I8480<= not G3640;
	I8483<= not G3641;
	I8486<= not G2824;
	I8517<= not G3014;
	I8520<= not G3652;
	I8543<= not G2810;
	I8565<= not G3071;
	I8665<= not G3051;
	I8706<= not G3828;
	I8709<= not G4191;
	I8712<= not G4007;
	I8715<= not G3903;
	I8718<= not G3909;
	I8721<= not G3918;
	I8724<= not G3927;
	I8727<= not G3944;
	I8730<= not G3987;
	I8733<= not G3996;
	I8736<= not G4008;
	I8739<= not G3910;
	I8742<= not G3919;
	I8745<= not G3929;
	I8748<= not G3997;
	I8751<= not G4009;
	I8754<= not G3911;
	I8757<= not G3921;
	I8760<= not G3931;
	I8763<= not G3947;
	I8766<= not G3960;
	I8769<= not G3999;
	I8772<= not G4011;
	I8775<= not G4019;
	I8778<= not G3922;
	I8781<= not G3932;
	I8784<= not G3949;
	I8787<= not G4012;
	I8790<= not G4020;
	I8793<= not G3923;
	I8796<= not G3934;
	I8799<= not G3951;
	I8802<= not G3963;
	I8805<= not G3976;
	I8808<= not G4014;
	I8811<= not G4022;
	I8814<= not G4028;
	I8817<= not G3935;
	I8820<= not G3952;
	I8823<= not G3965;
	I8826<= not G4023;
	I8829<= not G4029;
	I8832<= not G3936;
	I8835<= not G3954;
	I8838<= not G3967;
	I8841<= not G3979;
	I8844<= not G3992;
	I8847<= not G4025;
	I8850<= not G4031;
	I8853<= not G4034;
	I8856<= not G3955;
	I8859<= not G3968;
	I8862<= not G3981;
	I8865<= not G4032;
	I8868<= not G4035;
	I8871<= not G3869;
	I8874<= not G3884;
	I8877<= not G4274;
	I8880<= not G4303;
	I8883<= not G4198;
	I8886<= not G4308;
	I8889<= not G4311;
	I8892<= not G4115;
	I8895<= not G4130;
	I8898<= not G4089;
	I8901<= not G4122;
	I8904<= not G4126;
	I8907<= not G4095;
	I8910<= not G4200;
	I8913<= not G4306;
	I8916<= not G4195;
	I8919<= not G4196;
	I8922<= not G4229;
	I8925<= not G4482;
	I8928<= not G4153;
	I8932<= not G4096;
	I8935<= not G4005;
	I8945<= not G4106;
	I8949<= not G4116;
	I8952<= not G4197;
	I8962<= not G4553;
	I8966<= not G4444;
	I8971<= not G4464;
	I8974<= not G3871;
	I8977<= not G3877;
	I8980<= not G4535;
	I8983<= not G4536;
	I8986<= not G4552;
	I8989<= not G4537;
	I8994<= not G4565;
	I8998<= not G4576;
	I9001<= not G4577;
	I9005<= not G4585;
	I9009<= not G4591;
	I9014<= not G3864;
	I9018<= not G3872;
	I9021<= not G4489;
	I9025<= not G4462;
	I9034<= not G4317;
	I9050<= not G3881;
	I9053<= not G4327;
	I9064<= not G4302;
	I9076<= not G4353;
	I9081<= not G4357;
	I9084<= not G4358;
	I9089<= not G4566;
	I9095<= not G4283;
	I9103<= not G4374;
	I9111<= not G4232;
	I9116<= not G4297;
	I9123<= not G4455;
	I9126<= not G3870;
	I9129<= not G4475;
	I9132<= not G4284;
	I9136<= not G4280;
	I9139<= not G4364;
	I9142<= not G4236;
	I9145<= not G4264;
	I9148<= not G4354;
	I9158<= not G4256;
	I9162<= not G4272;
	I9177<= not G4299;
	I9209<= not G4349;
	I9217<= not G4443;
	I9250<= not G4134;
	I9258<= not G4249;
	I9271<= not G4263;
	I9301<= not G4295;
	I9310<= not G4268;
	I9325<= not G4242;
	I9333<= not G4245;
	I9336<= not G4493;
	I9341<= not G4251;
	I9344<= not G4341;
	I9347<= not G3896;
	I9350<= not G4503;
	I9360<= not G4257;
	I9363<= not G4258;
	I9366<= not G4350;
	I9369<= not G3901;
	I9372<= not G3902;
	I9393<= not G4266;
	I9396<= not G3908;
	I9407<= not G4232;
	I9416<= not G4273;
	I9419<= not G3916;
	I9422<= not G4360;
	I9425<= not G3917;
	I9440<= not G4285;
	I9443<= not G4564;
	I9446<= not G3926;
	I9457<= not G3940;
	I9460<= not G3941;
	I9463<= not G3942;
	I9466<= not G3943;
	I9484<= not G3957;
	I9493<= not G4426;
	I9496<= not G3971;
	I9499<= not G4382;
	I9502<= not G3972;
	I9505<= not G4300;
	I9512<= not G3985;
	I9515<= not G4301;
	I9520<= not G3995;
	I9525<= not G4413;
	I9528<= not G4006;
	I9531<= not G4463;
	I9539<= not G4018;
	I9543<= not G4279;
	I9555<= not G4892;
	I9558<= not G4597;
	I9561<= not G4695;
	I9564<= not G4703;
	I9567<= not G4693;
	I9570<= not G4696;
	I9573<= not G4701;
	I9576<= not G4706;
	I9579<= not G4713;
	I9582<= not G4694;
	I9585<= not G4697;
	I9588<= not G4704;
	I9591<= not G4710;
	I9594<= not G4718;
	I9597<= not G4738;
	I9600<= not G4698;
	I9603<= not G4719;
	I9606<= not G4687;
	I9609<= not G4780;
	I9612<= not G4776;
	I9615<= not G4739;
	I9618<= not G4742;
	I9621<= not G4732;
	I9624<= not G4746;
	I9627<= not G4777;
	I9630<= not G4867;
	I9633<= not G4800;
	I9636<= not G4802;
	I9639<= not G4685;
	I9642<= not G4788;
	I9645<= not G4900;
	I9648<= not G4795;
	I9651<= not G4805;
	I9654<= not G4792;
	I9657<= not G4784;
	I9660<= not G4806;
	I9663<= not G4809;
	I9666<= not G4931;
	I9669<= not G4909;
	I9672<= not G4803;
	I9675<= not G4807;
	I9678<= not G4808;
	I9681<= not G4811;
	I9684<= not G4813;
	I9687<= not G4822;
	I9752<= not G4705;
	I9760<= not G4838;
	I9774<= not G4678;
	I9782<= not G4720;
	I9785<= not G4747;
	I9788<= not G4711;
	I9791<= not G4779;
	I9794<= not G4778;
	I9804<= not G5113;
	I9819<= not G4691;
	I9823<= not G5138;
	I9834<= not G4782;
	I9837<= not G4781;
	I9840<= not G4702;
	I9845<= not G4728;
	I9850<= not G4798;
	I9884<= not G4868;
	I9889<= not G4819;
	I9892<= not G4879;
	I9907<= not G4837;
	I9910<= not G4681;
	I9918<= not G4968;
	I9929<= not G5052;
	I9935<= not G4812;
	I9938<= not G4878;
	I9974<= not G4676;
	I10028<= not G4825;
	I10032<= not G1236;
	I10046<= not G4840;
	I10125<= not G5127;
	I10128<= not G4688;
	I10135<= not G4960;
	I10151<= not G5007;
	I10154<= not G5109;
	I10157<= not G5109;
	I10160<= not G5139;
	I10166<= not G5016;
	I10169<= not G4873;
	I10172<= not G4873;
	I10177<= not G4721;
	I10180<= not G4721;
	I10183<= not G5129;
	I10186<= not G5129;
	I10190<= not G4670;
	I10193<= not G4670;
	I10204<= not G5060;
	I10207<= not G5075;
	I10236<= not G5014;
	I10243<= not G5026;
	I10247<= not G5266;
	I10250<= not G5268;
	I10253<= not G5240;
	I10256<= not G5401;
	I10259<= not G5362;
	I10262<= not G5551;
	I10265<= not G5468;
	I10268<= not G5471;
	I10271<= not G5487;
	I10274<= not G5524;
	I10277<= not G5472;
	I10280<= not G5488;
	I10283<= not G5643;
	I10286<= not G5519;
	I10289<= not G5569;
	I10292<= not G5577;
	I10295<= not G5523;
	I10343<= not G5704;
	I10347<= not G5706;
	I10350<= not G5707;
	I10353<= not G5710;
	I10356<= not G5711;
	I10366<= not G5715;
	I10369<= not G5716;
	I10373<= not G5722;
	I10377<= not G5188;
	I10380<= not G5448;
	I10384<= not G5193;
	I10387<= not G5194;
	I10390<= not G5195;
	I10393<= not G5196;
	I10397<= not G5200;
	I10400<= not G5201;
	I10403<= not G5202;
	I10406<= not G5203;
	I10409<= not G5204;
	I10412<= not G5205;
	I10415<= not G5397;
	I10418<= not G5453;
	I10421<= not G5208;
	I10424<= not G5209;
	I10427<= not G5210;
	I10430<= not G5211;
	I10433<= not G5212;
	I10436<= not G5213;
	I10439<= not G5214;
	I10442<= not G5215;
	I10445<= not G5418;
	I10448<= not G5335;
	I10451<= not G5216;
	I10454<= not G5217;
	I10457<= not G5218;
	I10460<= not G5219;
	I10463<= not G5220;
	I10466<= not G5221;
	I10469<= not G5222;
	I10472<= not G5223;
	I10475<= not G5529;
	I10479<= not G5227;
	I10482<= not G5228;
	I10485<= not G5229;
	I10488<= not G5230;
	I10491<= not G5231;
	I10494<= not G5232;
	I10497<= not G5233;
	I10500<= not G5234;
	I10503<= not G5235;
	I10506<= not G5236;
	I10509<= not G5237;
	I10512<= not G5238;
	I10516<= not G5241;
	I10519<= not G5242;
	I10522<= not G5243;
	I10525<= not G5244;
	I10528<= not G5245;
	I10532<= not G5253;
	I10535<= not G5254;
	I10538<= not G5255;
	I10541<= not G5256;
	I10545<= not G5259;
	I10548<= not G5260;
	I10552<= not G5396;
	I10555<= not G5529;
	I10558<= not G5264;
	I10561<= not G5265;
	I10565<= not G5402;
	I10569<= not G5417;
	I10574<= not G5426;
	I10579<= not G5433;
	I10582<= not G5437;
	I10587<= not G5439;
	I10592<= not G5444;
	I10605<= not G5440;
	I10608<= not G5701;
	I10614<= not G5302;
	I10617<= not G5677;
	I10639<= not G5224;
	I10643<= not G5267;
	I10646<= not G5364;
	I10649<= not G5657;
	I10675<= not G5662;
	I10678<= not G5566;
	I10681<= not G5686;
	I10684<= not G5258;
	I10687<= not G5674;
	I10690<= not G5538;
	I10694<= not G5445;
	I10702<= not G5529;
	I10705<= not G5463;
	I10708<= not G5545;
	I10716<= not G5537;
	I10719<= not G5559;
	I10739<= not G5572;
	I10752<= not G5618;
	I10758<= not G5662;
	I10761<= not G5302;
	I10766<= not G5674;
	I10770<= not G5441;
	I10773<= not G5708;
	I10776<= not G5576;
	I10780<= not G5445;
	I10783<= not G5542;
	I10786<= not G5452;
	I10796<= not G5397;
	I10801<= not G5463;
	I10804<= not G5526;
	I10807<= not G5294;
	I10810<= not G5403;
	I10815<= not G5418;
	I10826<= not G5434;
	I10829<= not G5224;
	I10842<= not G5701;
	I10862<= not G5364;
	I10882<= not G5600;
	I10896<= not G5475;
	I10914<= not G5448;
	I10919<= not G5479;
	I10930<= not G5600;
	I10933<= not G5668;
	I10937<= not G5560;
	I10940<= not G5489;
	I10946<= not G5563;
	I10949<= not G5513;
	I10962<= not G5719;
	I10965<= not G5719;
	I10969<= not G5606;
	I10973<= not G5726;
	I10976<= not G5726;
	I10987<= not G5609;
	I10998<= not G5672;
	I11001<= not G5698;
	I11004<= not G5613;
	I11008<= not G5693;
	I11011<= not G5693;
	I11014<= not G5621;
	I11018<= not G5626;
	I11021<= not G5627;
	I11025<= not G5638;
	I11028<= not G5642;
	I11031<= not G5335;
	I11034<= not G5644;
	I11037<= not G5299;
	I11040<= not G5299;
	I11043<= not G5648;
	I11047<= not G5653;
	I11050<= not G5335;
	I11055<= not G5696;
	I11060<= not G5453;
	I11066<= not G5460;
	I11069<= not G5671;
	I11086<= not G5397;
	I11090<= not G1000;
	I11129<= not G5418;
	I11132<= not G5624;
	I11191<= not G6155;
	I11194<= not G6243;
	I11197<= not G6122;
	I11200<= not G6251;
	I11203<= not G6129;
	I11206<= not G6133;
	I11209<= not G6139;
	I11212<= not G6146;
	I11215<= not G6156;
	I11218<= not G6161;
	I11221<= not G6167;
	I11224<= not G6255;
	I11227<= not G6130;
	I11230<= not G6140;
	I11233<= not G6147;
	I11236<= not G6148;
	I11239<= not G6173;
	I11242<= not G6183;
	I11245<= not G6143;
	I11248<= not G6149;
	I11251<= not G6152;
	I11254<= not G5793;
	I11257<= not G5805;
	I11260<= not G5779;
	I11263<= not G5784;
	I11266<= not G5794;
	I11269<= not G5756;
	I11272<= not G5758;
	I11275<= not G5768;
	I11278<= not G5780;
	I11281<= not G5785;
	I11284<= not G5795;
	I11287<= not G5806;
	I11290<= not G5818;
	I11293<= not G5824;
	I11296<= not G5831;
	I11299<= not G5786;
	I11302<= not G5796;
	I11305<= not G5807;
	I11308<= not G5759;
	I11311<= not G5760;
	I11314<= not G5781;
	I11317<= not G5787;
	I11320<= not G5797;
	I11323<= not G5808;
	I11326<= not G5819;
	I11329<= not G5825;
	I11332<= not G5832;
	I11335<= not G5839;
	I11338<= not G5798;
	I11341<= not G5809;
	I11344<= not G5820;
	I11347<= not G5761;
	I11350<= not G5763;
	I11353<= not G5788;
	I11356<= not G5799;
	I11359<= not G5810;
	I11362<= not G5821;
	I11365<= not G5826;
	I11368<= not G5833;
	I11371<= not G5840;
	I11374<= not G5844;
	I11377<= not G5811;
	I11380<= not G5822;
	I11383<= not G5827;
	I11386<= not G5764;
	I11389<= not G5766;
	I11392<= not G5800;
	I11395<= not G5812;
	I11398<= not G5823;
	I11401<= not G5828;
	I11404<= not G5834;
	I11407<= not G5841;
	I11410<= not G5845;
	I11413<= not G5871;
	I11416<= not G5829;
	I11419<= not G5835;
	I11422<= not G5842;
	I11425<= not G5872;
	I11428<= not G5813;
	I11431<= not G5782;
	I11434<= not G5789;
	I11437<= not G5801;
	I11440<= not G6009;
	I11443<= not G6038;
	I11446<= not G6062;
	I11449<= not G6068;
	I11452<= not G6071;
	I11455<= not G6087;
	I11458<= not G6063;
	I11461<= not G6094;
	I11464<= not G6088;
	I11467<= not G6064;
	I11470<= not G6095;
	I11473<= not G6069;
	I11476<= not G6194;
	I11479<= not G6201;
	I11482<= not G6117;
	I11485<= not G6137;
	I11488<= not G6034;
	I11491<= not G6010;
	I11494<= not G6037;
	I11497<= not G6014;
	I11500<= not G6219;
	I11503<= not G6220;
	I11506<= not G6189;
	I11512<= not G5874;
	I11515<= not G5897;
	I11522<= not G5847;
	I11525<= not G5874;
	I11533<= not G5847;
	I11556<= not G6065;
	I11559<= not G6065;
	I11562<= not G5939;
	I11569<= not G6279;
	I11586<= not G6256;
	I11591<= not G5814;
	I11596<= not G6228;
	I11607<= not G5767;
	I11622<= not G5847;
	I11627<= not G5874;
	I11633<= not G5897;
	I11638<= not G5847;
	I11641<= not G5918;
	I11645<= not G5874;
	I11648<= not G6028;
	I11652<= not G5939;
	I11656<= not G5772;
	I11659<= not G5897;
	I11662<= not G5956;
	I11666<= not G5772;
	I11669<= not G5918;
	I11672<= not G5971;
	I11677<= not G6076;
	I11680<= not G5939;
	I11683<= not G5988;
	I11686<= not G6076;
	I11689<= not G5956;
	I11693<= not G6076;
	I11696<= not G5971;
	I11701<= not G5772;
	I11704<= not G6076;
	I11707<= not G5988;
	I11710<= not G6098;
	I11714<= not G5772;
	I11718<= not G6115;
	I11722<= not G5772;
	I11725<= not G6036;
	I11729<= not G5772;
	I11732<= not G6076;
	I11736<= not G6076;
	I11740<= not G6136;
	I11744<= not G6120;
	I11747<= not G6123;
	I11764<= not G6056;
	I11773<= not G6262;
	I11778<= not G6180;
	I11781<= not G6284;
	I11787<= not G6273;
	I11790<= not G6282;
	I11793<= not G6188;
	I11796<= not G6287;
	I11800<= not G6164;
	I11803<= not G6280;
	I11806<= not G6275;
	I11809<= not G6285;
	I11815<= not G6169;
	I11818<= not G6276;
	I11821<= not G6170;
	I11824<= not G6283;
	I11827<= not G6231;
	I11832<= not G6274;
	I11835<= not G6181;
	I11838<= not G6281;
	I11848<= not G6159;
	I11851<= not G6277;
	I11855<= not G5751;
	I11858<= not G6165;
	I11861<= not G5747;
	I11864<= not G5753;
	I11867<= not G6286;
	I11870<= not G5752;
	I11880<= not G5748;
	I11884<= not G6091;
	I11887<= not G5918;
	I11890<= not G6135;
	I11894<= not G5956;
	I11897<= not G6141;
	I11900<= not G5847;
	I11903<= not G5939;
	I11908<= not G5918;
	I11912<= not G5897;
	I11917<= not G5897;
	I11920<= not G5874;
	I11923<= not G5939;
	I11926<= not G6190;
	I11929<= not G6190;
	I11933<= not G5847;
	I11936<= not G5918;
	I11939<= not G6015;
	I11942<= not G6015;
	I11945<= not G5874;
	I11948<= not G5897;
	I11951<= not G5847;
	I11955<= not G5988;
	I11958<= not G5874;
	I11961<= not G5988;
	I11964<= not G5971;
	I11967<= not G5971;
	I11971<= not G6179;
	I11974<= not G5956;
	I11978<= not G6186;
	I11981<= not G6246;
	I11984<= not G6246;
	I11987<= not G6278;
	I11991<= not G5939;
	I11994<= not G6195;
	I11998<= not G5918;
	I12003<= not G6202;
	I12008<= not G5897;
	I12011<= not G5939;
	I12022<= not G5874;
	I12025<= not G5918;
	I12038<= not G5847;
	I12041<= not G5897;
	I12044<= not G5847;
	I12059<= not G5874;
	I12062<= not G5988;
	I12065<= not G5897;
	I12068<= not G5847;
	I12085<= not G5971;
	I12088<= not G5874;
	I12091<= not G5988;
	I12098<= not G5956;
	I12101<= not G5971;
	I12108<= not G5939;
	I12111<= not G5956;
	I12117<= not G5918;
	I12120<= not G5939;
	I12124<= not G5847;
	I12128<= not G5897;
	I12131<= not G5918;
	I12135<= not G5988;
	I12138<= not G5874;
	I12141<= not G5897;
	I12145<= not G5971;
	I12148<= not G5988;
	I12151<= not G5847;
	I12154<= not G5874;
	I12158<= not G5956;
	I12161<= not G5971;
	I12164<= not G5847;
	I12167<= not G5939;
	I12170<= not G5956;
	I12173<= not G5918;
	I12176<= not G5939;
	I12187<= not G5897;
	I12190<= not G5918;
	I12193<= not G6468;
	I12196<= not G6471;
	I12199<= not G6475;
	I12202<= not G6481;
	I12205<= not G6488;
	I12208<= not G6496;
	I12211<= not G6502;
	I12214<= not G6507;
	I12217<= not G6631;
	I12220<= not G6645;
	I12223<= not G6655;
	I12226<= not G6636;
	I12229<= not G6659;
	I12232<= not G6662;
	I12235<= not G6634;
	I12238<= not G6637;
	I12241<= not G6640;
	I12244<= not G6642;
	I12247<= not G6646;
	I12250<= not G6651;
	I12253<= not G6427;
	I12256<= not G6647;
	I12259<= not G6652;
	I12262<= not G6656;
	I12265<= not G6660;
	I12268<= not G6661;
	I12271<= not G6663;
	I12274<= not G6672;
	I12277<= not G6681;
	I12280<= not G6684;
	I12283<= not G6692;
	I12286<= not G6696;
	I12289<= not G6702;
	I12292<= not G6657;
	I12295<= not G6693;
	I12298<= not G6697;
	I12301<= not G6703;
	I12304<= not G6711;
	I12307<= not G6712;
	I12310<= not G6723;
	I12313<= not G6730;
	I12316<= not G6736;
	I12319<= not G6741;
	I12322<= not G6751;
	I12325<= not G6755;
	I12328<= not G6760;
	I12331<= not G6704;
	I12334<= not G6713;
	I12337<= not G6724;
	I12340<= not G6725;
	I12343<= not G6731;
	I12346<= not G6737;
	I12349<= not G6742;
	I12352<= not G6752;
	I12355<= not G6756;
	I12358<= not G6761;
	I12361<= not G6765;
	I12364<= not G6714;
	I12367<= not G6754;
	I12370<= not G6758;
	I12373<= not G6763;
	I12376<= not G6766;
	I12379<= not G6768;
	I12382<= not G6772;
	I12385<= not G6397;
	I12388<= not G6403;
	I12391<= not G6744;
	I12394<= not G6759;
	I12397<= not G6764;
	I12400<= not G6767;
	I12403<= not G6769;
	I12406<= not G6773;
	I12409<= not G6398;
	I12412<= not G6404;
	I12415<= not G6410;
	I12418<= not G6572;
	I12421<= not G6486;
	I12424<= not G6446;
	I12427<= not G6553;
	I12430<= not G6432;
	I12433<= not G6632;
	I12436<= not G6635;
	I12439<= not G6566;
	I12442<= not G6542;
	I12445<= not G6568;
	I12448<= not G6569;
	I12451<= not G6524;
	I12454<= not G6581;
	I12457<= not G6671;
	I12460<= not G6674;
	I12463<= not G6682;
	I12466<= not G6687;
	I12469<= not G6586;
	I12472<= not G6591;
	I12475<= not G6596;
	I12478<= not G6603;
	I12481<= not G6616;
	I12484<= not G6621;
	I12487<= not G6623;
	I12490<= not G6625;
	I12493<= not G6587;
	I12496<= not G6592;
	I12499<= not G6597;
	I12502<= not G6604;
	I12505<= not G6612;
	I12508<= not G6593;
	I12511<= not G6598;
	I12514<= not G6605;
	I12517<= not G6613;
	I12520<= not G6622;
	I12523<= not G6624;
	I12526<= not G6626;
	I12529<= not G6628;
	I12532<= not G6594;
	I12535<= not G6599;
	I12538<= not G6606;
	I12541<= not G6614;
	I12544<= not G6617;
	I12547<= not G6708;
	I12558<= not G6449;
	I12561<= not G6449;
	I12564<= not G6720;
	I12567<= not G6721;
	I12571<= not G6729;
	I12582<= not G6745;
	I12586<= not G6643;
	I12592<= not G1008;
	I12609<= not G6571;
	I12629<= not G6523;
	I12632<= not G6514;
	I12635<= not G6509;
	I12639<= not G6506;
	I12643<= not G6501;
	I12646<= not G6493;
	I12649<= not G6457;
	I12652<= not G6664;
	I12655<= not G6458;
	I12659<= not G6459;
	I12666<= not G6476;
	I12669<= not G6477;
	I12672<= not G6473;
	I12675<= not G6510;
	I12678<= not G6516;
	I12681<= not G6469;
	I12684<= not G6472;
	I12687<= not G6745;
	I12690<= not G6467;
	I12696<= not G6503;
	I12699<= not G6504;
	I12702<= not G6497;
	I12708<= not G6482;
	I12712<= not G6543;
	I12717<= not G6543;
	I12722<= not G6611;
	I12725<= not G6565;
	I12731<= not G6579;
	I12737<= not G6460;
	I12742<= not G6590;
	I12748<= not G6585;
	I12753<= not G6445;
	I12757<= not G6577;
	I12760<= not G6685;
	I12763<= not G6686;
	I12768<= not G6718;
	I12771<= not G6735;
	I12776<= not G6739;
	I12779<= not G6740;
	I12782<= not G6463;
	I12806<= not G6602;
	I12810<= not G6607;
	I12813<= not G6607;
	I12826<= not G6441;
	I12829<= not G6441;
	I12839<= not G6630;
	I12866<= not G6483;
	I12877<= not G6700;
	I12881<= not G6478;
	I12885<= not G6946;
	I12888<= not G6948;
	I12891<= not G6950;
	I12894<= not G7009;
	I12897<= not G6962;
	I12900<= not G6947;
	I12903<= not G6905;
	I12906<= not G6918;
	I12909<= not G7046;
	I12912<= not G7006;
	I12915<= not G7000;
	I12918<= not G7013;
	I12921<= not G6993;
	I12924<= not G6983;
	I12927<= not G7014;
	I12930<= not G7019;
	I12933<= not G7018;
	I12936<= not G7015;
	I12939<= not G7022;
	I12942<= not G7023;
	I12945<= not G7066;
	I12948<= not G6919;
	I12958<= not G6920;
	I12961<= not G6921;
	I12965<= not G6924;
	I12968<= not G6925;
	I12973<= not G6927;
	I12976<= not G6928;
	I12980<= not G6929;
	I12983<= not G6930;
	I12986<= not G6931;
	I12989<= not G6932;
	I12993<= not G6933;
	I12996<= not G6934;
	I12999<= not G7029;
	I13009<= not G6935;
	I13012<= not G7071;
	I13023<= not G7040;
	I13028<= not G7087;
	I13031<= not G6984;
	I13035<= not G6964;
	I13039<= not G6961;
	I13042<= not G6963;
	I13045<= not G6955;
	I13048<= not G6956;
	I13051<= not G6967;
	I13054<= not G6960;
	I13057<= not G6968;
	I13060<= not G6959;
	I13063<= not G6973;
	I13066<= not G6957;
	I13072<= not G6969;
	I13075<= not G6958;
	I13084<= not G7071;
	I13088<= not G7045;
	I13092<= not G7047;
	I13099<= not G7054;
	I13103<= not G7055;
	I13106<= not G7056;
	I13109<= not G7059;
	I13112<= not G7021;
	I13118<= not G7068;
	I13122<= not G7070;
	I13126<= not G6949;
	I13131<= not G6951;
	I13134<= not G7017;
	I13137<= not G7027;
	I13140<= not G6954;
	I13144<= not G7031;
	I13147<= not G7024;
	I13152<= not G6966;
	I13157<= not G6997;
	I13161<= not G7080;
	I13164<= not G7086;
	I13173<= not G7089;
	I13185<= not G7020;
	I13189<= not G7002;
	I13193<= not G7007;
	I13196<= not G7008;
	I13199<= not G7025;
	I13203<= not G7088;
	I13209<= not G6912;
	I13225<= not G7095;
	I13228<= not G6892;
	I13231<= not G6897;
	I13234<= not G6898;
	I13238<= not G6900;
	I13241<= not G7030;
	I13244<= not G7033;
	I13247<= not G6906;
	I13250<= not G7036;
	I13255<= not G7057;
	I13258<= not G6907;
	I13261<= not G7041;
	I13264<= not G7061;
	I13267<= not G6913;
	I13271<= not G7067;
	I13274<= not G6917;
	I13277<= not G7078;
	I13281<= not G7155;
	I13284<= not G7156;
	I13287<= not G7157;
	I13290<= not G7158;
	I13293<= not G7159;
	I13296<= not G7161;
	I13299<= not G7163;
	I13302<= not G7164;
	I13305<= not G7168;
	I13308<= not G7169;
	I13311<= not G7162;
	I13314<= not G7160;
	I13317<= not G7211;
	I13320<= not G7139;
	I13323<= not G7145;
	I13326<= not G7176;
	I13329<= not G7247;
	I13332<= not G7241;
	I13335<= not G7206;
	I13338<= not G7190;
	I13341<= not G7207;
	I13344<= not G7210;
	I13347<= not G7224;
	I13350<= not G7223;
	I13353<= not G7231;
	I13356<= not G7221;
	I13359<= not G7255;
	I13362<= not G7265;
	I13365<= not G7267;
	I13369<= not G7268;
	I13373<= not G7270;
	I13383<= not G7275;
	I13388<= not G7149;
	I13403<= not G7269;
	I13407<= not G7271;
	I13410<= not G7274;
	I13413<= not G7127;
	I13416<= not G7165;
	I13419<= not G7277;
	I13422<= not G7131;
	I13425<= not G7166;
	I13428<= not G7167;
	I13432<= not G7280;
	I13435<= not G7170;
	I13438<= not G7143;
	I13441<= not G7146;
	I13444<= not G7282;
	I13447<= not G7261;
	I13451<= not G7262;
	I13454<= not G7147;
	I13457<= not G7120;
	I13460<= not G7263;
	I13463<= not G7264;
	I13466<= not G7122;
	I13469<= not G7123;
	I13472<= not G7266;
	I13475<= not G7125;
	I13478<= not G7126;
	I13481<= not G7254;
	I13484<= not G7128;
	I13487<= not G7129;
	I13490<= not G7130;
	I13493<= not G7132;
	I13496<= not G7133;
	I13499<= not G7134;
	I13502<= not G7135;
	I13506<= not G7148;
	I13509<= not G7137;
	I13512<= not G7138;
	I13515<= not G7152;
	I13518<= not G7141;
	I13524<= not G7151;
	I13527<= not G7217;
	I13533<= not G7220;
	I13537<= not G7152;
	I13541<= not G7209;
	I13544<= not G1167;
	I13547<= not G1170;
	I13550<= not G1173;
	I13559<= not G7177;
	I13562<= not G7179;
	I13565<= not G7181;
	I13570<= not G7198;
	I13574<= not G7205;
	I13577<= not G7186;
	I13580<= not G7208;
	I13583<= not G7252;
	I13595<= not G7216;
	I13605<= not G7197;
	I13610<= not G7227;
	I13613<= not G7273;
	I13617<= not G7276;
	I13622<= not G7279;
	I13628<= not G7248;
	I13631<= not G7248;
	I13635<= not G7243;
	I13646<= not G7245;
	I13649<= not G7281;
	I13653<= not G7246;
	I13656<= not G7228;
	I13659<= not G7232;
	I13663<= not G7235;
	I13666<= not G7238;
	I13669<= not G7240;
	I13672<= not G7242;
	I13676<= not G7256;
	I13679<= not G7259;
	I13682<= not G7251;
	I13692<= not G7343;
	I13695<= not G7345;
	I13698<= not G7348;
	I13701<= not G7349;
	I13704<= not G7352;
	I13707<= not G7420;
	I13710<= not G7340;
	I13713<= not G7341;
	I13716<= not G7331;
	I13719<= not G7334;
	I13722<= not G7442;
	I13725<= not G7437;
	I13728<= not G7439;
	I13731<= not G7441;
	I13734<= not G7422;
	I13737<= not G7446;
	I13740<= not G7364;
	I13743<= not G7454;
	I13746<= not G7311;
	I13749<= not G7313;
	I13752<= not G7315;
	I13755<= not G7317;
	I13758<= not G7414;
	I13761<= not G7418;
	I13764<= not G7479;
	I13767<= not G7486;
	I13770<= not G7491;
	I13773<= not G7496;
	I13776<= not G7497;
	I13779<= not G7406;
	I13782<= not G7498;
	I13794<= not G7346;
	I13797<= not G7502;
	I13807<= not G7320;
	I13810<= not G7312;
	I13813<= not G7314;
	I13816<= not G7455;
	I13819<= not G7426;
	I13822<= not G7459;
	I13825<= not G7318;
	I13828<= not G7321;
	I13831<= not G7322;
	I13834<= not G7466;
	I13837<= not G7324;
	I13843<= not G7326;
	I13846<= not G7487;
	I13850<= not G7328;
	I13854<= not G7327;
	I13858<= not G7329;
	I13861<= not G7330;
	I13865<= not G7333;
	I13869<= not G7338;
	I13873<= not G7342;
	I13876<= not G7347;
	I13879<= not G7332;
	I13882<= not G7350;
	I13885<= not G7351;
	I13888<= not G7335;
	I13891<= not G7336;
	I13894<= not G7353;
	I13897<= not G7354;
	I13900<= not G7356;
	I13903<= not G7357;
	I13906<= not G7358;
	I13909<= not G7339;
	I13912<= not G7359;
	I13915<= not G7360;
	I13918<= not G7361;
	I13921<= not G7362;
	I13924<= not G7365;
	I13927<= not G7366;
	I13930<= not G7405;
	I13940<= not G7355;
	I13956<= not G7499;
	I13962<= not G7413;
	I13979<= not G7415;
	I13997<= not G7432;
	I14001<= not G7433;
	I14005<= not G7434;
	I14009<= not G7436;
	I14012<= not G7438;
	I14015<= not G7440;
	I14019<= not G7480;
	I14022<= not G7443;
	I14025<= not G7500;
	I14028<= not G7501;
	I14031<= not G7448;
	I14035<= not G7310;
	I14039<= not G7449;
	I14042<= not G7470;
	I14046<= not G7492;
	I14049<= not G7493;
	I14052<= not G7494;
	I14055<= not G7495;
	I14058<= not G7544;
	I14061<= not G7546;
	I14064<= not G7556;
	I14067<= not G7550;
	I14070<= not G7714;
	I14073<= not G7627;
	I14076<= not G7577;
	I14079<= not G7579;
	I14082<= not G7539;
	I14085<= not G7583;
	I14088<= not G7585;
	I14091<= not G7589;
	I14094<= not G7593;
	I14097<= not G7595;
	I14100<= not G7580;
	I14103<= not G7584;
	I14106<= not G7586;
	I14109<= not G7590;
	I14112<= not G7560;
	I14115<= not G7563;
	I14118<= not G7565;
	I14121<= not G7587;
	I14124<= not G7591;
	I14127<= not G7594;
	I14130<= not G7592;
	I14133<= not G7574;
	I14136<= not G7633;
	I14139<= not G7548;
	I14142<= not G7551;
	I14145<= not G7542;
	I14148<= not G7543;
	I14151<= not G7555;
	I14154<= not G7558;
	I14157<= not G7547;
	I14160<= not G7549;
	I14163<= not G7533;
	I14166<= not G7702;
	I14169<= not G7715;
	I14172<= not G7545;
	I14175<= not G7718;
	I14178<= not G7562;
	I14181<= not G7725;
	I14184<= not G7726;
	I14187<= not G7728;
	I14190<= not G7531;
	I14193<= not G7532;
	I14196<= not G7534;
	I14199<= not G7704;
	I14202<= not G7708;
	I14205<= not G7710;
	I14208<= not G7711;
	I14211<= not G7712;
	I14214<= not G7576;
	I14224<= not G7722;
	I14227<= not G7552;
	I14231<= not G7566;
	I14234<= not G7614;
	I14238<= not G7608;
	I14251<= not G7541;
	I14257<= not G7716;
	I14260<= not G7717;
	I14264<= not G7698;
	I14267<= not G7695;
	I14270<= not G7703;
	I14273<= not G7631;
	I14276<= not G7720;
	I14279<= not G7700;
	I14282<= not G7709;
	I14285<= not G7625;
	I14288<= not G7705;
	I14291<= not G7680;
	I14294<= not G7553;
	I14298<= not G7678;
	I14305<= not G7537;
	I14311<= not G7566;
	I14315<= not G7676;
	I14318<= not G7657;
	I14325<= not G7713;
	I14330<= not G7538;
	I14334<= not G7578;
	I14338<= not G7581;
	I14342<= not G7582;
	I14349<= not G7588;
	I14370<= not G7603;
	I14374<= not G7693;
	I14378<= not G7691;
	I14381<= not G7596;
	I14388<= not G7605;
	I14394<= not G7536;
	I14397<= not G7686;
	I14400<= not G7677;
	I14403<= not G7679;
	I14406<= not G7681;
	I14410<= not G7697;
	I14413<= not G7723;
	I14416<= not G7727;
	I14420<= not G7554;
	I14424<= not G7652;
	I14427<= not G7835;
	I14430<= not G7836;
	I14433<= not G8061;
	I14436<= not G7904;
	I14439<= not G8063;
	I14442<= not G8065;
	I14445<= not G8067;
	I14448<= not G7792;
	I14451<= not G8172;
	I14454<= not G8177;
	I14457<= not G8093;
	I14460<= not G7789;
	I14463<= not G8072;
	I14489<= not G7829;
	I14492<= not G7829;
	I14531<= not G8178;
	I14573<= not G8179;
	I14603<= not G7827;
	I14614<= not G7832;
	I14623<= not G7833;
	I14637<= not G8012;
	I14643<= not G7837;
	I14646<= not G7790;
	I14657<= not G7782;
	I14662<= not G7783;
	I14668<= not G7787;
	I14674<= not G7788;
	I14677<= not G7791;
	I14680<= not G7810;
	I14683<= not G7825;
	I14687<= not G7826;
	I14695<= not G8016;
	I14709<= not G8198;
	I14712<= not G8059;
	I14718<= not G8068;
	I14722<= not G8076;
	I14725<= not G8145;
	I14728<= not G8152;
	I14732<= not G8155;
	I14739<= not G8173;
	I14743<= not G8174;
	I14747<= not G8175;
	I14763<= not G7834;
	I14777<= not G8511;
	I14780<= not G8284;
	I14783<= not G8324;
	I14786<= not G8606;
	I14789<= not G8544;
	I14792<= not G8583;
	I14795<= not G8604;
	I14798<= not G8605;
	I14801<= not G8608;
	I14804<= not G8563;
	I14807<= not G8603;
	I14810<= not G8481;
	I14813<= not G8640;
	I14816<= not G8642;
	I14819<= not G8647;
	I14822<= not G8649;
	I14825<= not G8651;
	I14828<= not G8639;
	I14844<= not G8641;
	I14848<= not G8625;
	I14851<= not G8630;
	I14857<= not G8657;
	I14904<= not G8629;
	I14925<= not G8381;
	I14964<= not G8406;
	I14974<= not G8442;
	I14996<= not G8510;
	I15003<= not G8633;
	I15007<= not G8627;
	I15010<= not G8584;
	I15014<= not G8607;
	I15062<= not G8632;
	I15065<= not G8636;
	I15068<= not G8638;
	I15160<= not G8631;
	I15178<= not G8753;
	I15181<= not G8734;
	I15184<= not G8684;
	I15187<= not G8682;
	I15190<= not G8685;
	I15193<= not G8774;
	I15196<= not G8778;
	I15199<= not G8792;
	I15202<= not G8797;
	I15205<= not G8809;
	I15208<= not G8810;
	I15211<= not G8808;
	I15218<= not G8801;
	I15222<= not G8834;
	I15225<= not G8689;
	I15308<= not G8799;
	I15315<= not G8738;
	I15324<= not G8779;
	I15329<= not G8793;
	I15334<= not G8800;
	I15337<= not G8802;
	I15340<= not G8856;
	I15379<= not G8882;
	I15382<= not G8883;
	I15385<= not G8880;
	I15388<= not G8898;
	I15391<= not G8917;
	I15394<= not G8916;
	I15405<= not G8902;
	I15408<= not G8896;
	I15411<= not G8897;
	I15414<= not G8900;
	I15417<= not G8893;
	I15420<= not G8881;
	I15423<= not G8894;
	I15426<= not G8895;
	I15429<= not G8899;
	I15433<= not G8911;
	I15475<= not G8901;
	I15478<= not G8910;
	I15481<= not G8913;
	I15484<= not G8918;
	I15492<= not G8971;
	I15495<= not G8973;
	I15498<= not G8974;
	I15501<= not G8975;
	I15504<= not G8967;
	I15507<= not G8968;
	I15510<= not G8969;
	I15513<= not G8970;
	I15516<= not G8977;
	I15519<= not G9019;
	I15522<= not G9018;
	I15527<= not G9020;
	I15530<= not G8972;
	I15533<= not G9002;
	I15536<= not G9004;
	I15539<= not G9005;
	I15543<= not G9006;
	I15546<= not G9007;
	I15550<= not G9008;
	I15553<= not G9009;
	I15557<= not G9010;
	I15562<= not G8979;
	I15565<= not G8980;
	I15568<= not G8981;
	I15571<= not G8982;
	I15574<= not G8983;
	I15577<= not G8984;
	I15580<= not G8985;
	I15583<= not G8986;
	I15586<= not G8987;
	I15589<= not G8988;
	I15592<= not G8989;
	I15595<= not G8990;
	I15598<= not G8991;
	I15601<= not G8992;
	I15604<= not G8993;
	I15607<= not G8994;
	I15610<= not G8995;
	I15613<= not G8996;
	I15616<= not G8997;
	I15619<= not G8998;
	I15622<= not G8999;
	I15625<= not G9000;
	I15628<= not G9001;
	I15631<= not G9003;
	I15635<= not G8976;
	I15638<= not G8978;
	I15641<= not G9017;
	I15645<= not G9043;
	I15648<= not G9044;
	I15651<= not G9056;
	I15654<= not G9057;
	I15657<= not G9059;
	I15660<= not G9062;
	I15663<= not G9066;
	I15666<= not G9070;
	I15669<= not G9045;
	I15672<= not G9047;
	I15675<= not G9058;
	I15678<= not G9060;
	I15681<= not G9063;
	I15684<= not G9067;
	I15687<= not G9071;
	I15690<= not G9074;
	I15693<= not G9048;
	I15696<= not G9050;
	I15699<= not G9061;
	I15702<= not G9064;
	I15705<= not G9068;
	I15708<= not G9072;
	I15711<= not G9075;
	I15714<= not G9077;
	I15717<= not G9051;
	I15720<= not G9053;
	I15723<= not G9065;
	I15726<= not G9069;
	I15729<= not G9073;
	I15732<= not G9076;
	I15735<= not G9078;
	I15738<= not G9079;
	I15741<= not G9083;
	I15747<= not G9042;
	I15753<= not G9080;
	I15756<= not G9081;
	I15759<= not G9082;
	I15762<= not G9039;
	I15765<= not G9039;
	I15770<= not G9121;
	I15773<= not G9126;
	I15776<= not G9127;
	I15784<= not G9125;
	I15791<= not G9140;
	I15803<= not G9148;
	I15811<= not G9151;
	I15814<= not G9154;
	I15824<= not G9157;
	I15830<= not G9180;
	I15833<= not G9162;
	I15836<= not G9165;
	I15839<= not G9168;
	I15842<= not G9171;
	I15845<= not G9174;
	I15871<= not G9184;
	I15894<= not G9195;
	I15909<= not G9201;
	I15912<= not G9193;
	I15915<= not G9194;
	I15918<= not G9211;
	I15921<= not G9206;
	I15924<= not G9207;
	I15927<= not G9208;
	I15930<= not G9209;
	I15933<= not G9210;
	I15937<= not G9212;
	I15940<= not G9213;
	I15943<= not G9214;
	I15947<= not G9221;
	I15950<= not G9222;
	I15953<= not G9215;
	I15956<= not G9216;
	I15959<= not G9217;
	I15962<= not G9218;
	I15965<= not G9219;
	I15971<= not G9233;
	I15974<= not G9234;
	I15978<= not G9235;
	I15982<= not G9236;
	I15985<= not G9237;
	I15990<= not G9239;
	I16006<= not G9261;
	I16009<= not G9261;
	I16017<= not G9264;
	I16020<= not G9264;
	I16023<= not G9267;
	I16026<= not G9267;
	I16033<= not G9282;
	I16036<= not G9282;
	I16040<= not G9285;
	I16043<= not G9285;
	I16046<= not G9288;
	I16049<= not G9288;
	I16052<= not G9291;
	I16055<= not G9291;
	I16058<= not G9294;
	I16061<= not G9294;
	I16072<= not G9303;
	I16084<= not G9324;
	I16090<= not G9336;
	I16100<= not G9338;
	I16103<= not G9339;
	I16107<= not G9337;
	I16116<= not G9350;
	I16119<= not G9351;
	I16122<= not G9353;
	I16126<= not G9354;
	I16129<= not G9355;
	I16132<= not G9356;
	I16135<= not G9357;
	I16138<= not G9358;
	I16142<= not G9366;
	I16145<= not G9367;
	I16148<= not G9368;
	I16151<= not G9369;
	I16154<= not G9370;
	I16158<= not G9363;
	I16161<= not G9363;
	I16165<= not G9377;
	I16168<= not G9381;
	I16173<= not G9382;
	I16176<= not G9385;
	I16180<= not G9387;
	I16183<= not G9388;
	G1714<=G1454 and G1450;
	G1725<=G1409 and G1416;
	G1728<=G1432 and G1439;
	G1733<=G1489 and G1481;
	G1739<=G803 and G799;
	G1753<=G819 and G815;
	G1834<=G933 and G929;
	G1844<=G792 and G795;
	G1898<=G959 and G955;
	G1913<=G1528 and G1532;
	G1919<=G1098 and G1087;
	G2386<=G1130 and G1092;
	G2768<=G1597 and G973;
	G2781<=G1600 and G976;
	G2827<=G1889 and G1690;
	G2889<=G1612 and G1077;
	G2912<=G1080 and G1945;
	G2935<=G1612 and G1077;
	G2949<=G822 and G1753;
	G2952<=G2474 and G2215;
	G2972<=G2397 and G2407;
	G2979<=G1494 and G1733;
	G2986<=G806 and G1739;
	G3002<=G871 and G1834;
	G3049<=G2274 and G1844;
	G3081<=G1682 and G1616;
	G3094<=G945 and G1898;
	G3188<=G2298 and G2316;
	G3190<=G1658 and G2424;
	G3222<=G1537 and G1913;
	G3226<=G1102 and G1919;
	G3229<=G1728 and G2015;
	G3258<=G2298 and G2316 and G2334 and G2354;
	G3259<=G1976 and G1960;
	G3313<=G2334 and G2316 and G2298;
	G3429<=G1454 and G1838 and G1444;
	G3466<=G936 and G2557;
	G3509<=G1637 and G1616;
	G3614<=G1134 and G2386;
	G3984<=G2403 and G3085;
	G4038<=G825 and G2949;
	G4047<=G1272 and G3503;
	G4048<=G1288 and G3513;
	G4049<=G141 and G3514;
	G4052<=G1276 and G3522;
	G4053<=G1292 and G3523;
	G4054<=G3767 and G2424;
	G4058<=G3656 and G2407;
	G4059<=G1499 and G2979;
	G4062<=G809 and G2986;
	G4066<=G1280 and G3532;
	G4067<=G133 and G3539;
	G4068<=G121 and G3540;
	G4073<=G1300 and G3567;
	G4074<=G137 and G3573;
	G4077<=G1284 and G3582;
	G4078<=G3753 and G3732 and G3712 and G3700;
	G4082<=G1296 and G3604;
	G4083<=G125 and G3610;
	G4086<=G103 and G3629;
	G4091<=G129 and G3639;
	G4097<=G2624 and G2614;
	G4098<=G985 and G3790;
	G4099<=G117 and G3647;
	G4100<=G113 and G3648;
	G4101<=G108 and G3649;
	G4107<=G2625 and G2615;
	G4108<=G782 and G3655;
	G4109<=G990 and G3790;
	G4117<=G2626 and G2616;
	G4118<=G995 and G3790;
	G4123<=G2627 and G2617;
	G4124<=G2641 and G2640;
	G4127<=G2628 and G2618;
	G4128<=G98 and G3693;
	G4129<=G2629 and G2621;
	G4131<=G2630 and G2622;
	G4132<=G2637 and G2633;
	G4133<=G2631 and G2623;
	G4135<=I7994 and I7995;
	G4138<=G2638 and G2634;
	G4139<=I8000 and I8001;
	G4142<=I8005 and I8006;
	G4145<=G2639 and G2635;
	G4147<=I8014 and I8015;
	G4150<=I8019 and I8020;
	G4154<=G1098 and G3495;
	G4155<=I8028 and I8029;
	G4158<=I8033 and I8034;
	G4159<=G1102 and G3498;
	G4163<=I8040 and I8041;
	G4166<=I8045 and I8046;
	G4167<=G2783 and G1616;
	G4168<=G1106 and G3500;
	G4169<=I8052 and I8053;
	G4172<=I8057 and I8058;
	G4175<=G1110 and G3502;
	G4176<=I8063 and I8064;
	G4180<=G1114 and G3511;
	G4181<=G1142 and G3512;
	G4182<=I8071 and I8072;
	G4185<=G2636 and G2632;
	G4186<=G1118 and G3520;
	G4187<=I8078 and I8079;
	G4190<=G1122 and G3527;
	G4192<=G1126 and G3531;
	G4193<=G145 and G2727;
	G4194<=I8089 and I8090;
	G4199<=G93 and G2769;
	G4201<=I8108 and I8109;
	G4216<=I8114 and I8115;
	G4220<=G3533 and G3549 and G3568 and G3583;
	G4224<=G2680 and G2683 and I8127;
	G4225<=G2686 and G2689 and G2692 and G2695;
	G4230<=G2683 and G3491 and I8143;
	G4236<=G3260 and G3221;
	G4238<=G2695 and G2698 and I8157;
	G4239<=G1541 and G3222;
	G4246<=G1106 and G3226;
	G4254<=G3583 and G3568 and G3549;
	G4255<=G3605 and G3644 and G3635 and I8186;
	G4268<=G2216 and G2655;
	G4269<=G2354 and G3563 and I8209;
	G4271<=G3666 and G3684;
	G4272<=G3233 and G3286;
	G4276<=G2216 and G2618;
	G4282<=G3549 and G3568;
	G4284<=G3260 and G3314;
	G4287<=G3563 and G2334 and G3579 and I8237;
	G4288<=G3563 and G3579 and G3603 and I8240;
	G4299<=G3233 and G3358;
	G4302<=G3086 and G3659 and G3124;
	G4304<=G2784 and G3779;
	G4312<=G3666 and G3684 and G3694 and G3707;
	G4314<=G3694 and G3684 and G3666;
	G4315<=G3707 and G3728 and I8288;
	G4317<=G878 and G3086 and G1857 and G3659;
	G4319<=G3728 and G3694 and G3750 and I8296;
	G4320<=G3728 and G3750 and G3768 and I8299;
	G4327<=G2959 and G1867;
	G4333<=G1087 and G2782;
	G4334<=G225 and G3097;
	G4342<=G228 and G3097;
	G4343<=G306 and G3131;
	G4351<=G309 and G3131;
	G4352<=G387 and G3160;
	G4355<=G390 and G3160;
	G4356<=G468 and G3192;
	G4361<=G471 and G3192;
	G4365<=G237 and G3097;
	G4366<=G216 and G3097;
	G4367<=G240 and G3097;
	G4368<=G318 and G3131;
	G4369<=G580 and G2845;
	G4375<=G219 and G3097;
	G4376<=G243 and G3097;
	G4377<=G297 and G3131;
	G4378<=G321 and G3131;
	G4379<=G399 and G3160;
	G4380<=G584 and G2845;
	G4383<=G222 and G3097;
	G4384<=G246 and G3097;
	G4385<=G300 and G3131;
	G4386<=G324 and G3131;
	G4387<=G378 and G3160;
	G4388<=G402 and G3160;
	G4389<=G480 and G3192;
	G4390<=G560 and G2845;
	G4391<=G249 and G3097;
	G4392<=G303 and G3131;
	G4393<=G327 and G3131;
	G4394<=G381 and G3160;
	G4395<=G405 and G3160;
	G4396<=G459 and G3192;
	G4397<=G483 and G3192;
	G4398<=G567 and G2845;
	G4400<=G1138 and G3614;
	G4403<=I8400 and I8401;
	G4407<=G252 and G3097;
	G4408<=G330 and G3131;
	G4409<=G384 and G3160;
	G4410<=G408 and G3160;
	G4411<=G462 and G3192;
	G4412<=G486 and G3192;
	G4414<=I8412 and I8413;
	G4417<=I8417 and I8418;
	G4420<=G275 and G3097;
	G4421<=G333 and G3131;
	G4422<=G411 and G3160;
	G4423<=G465 and G3192;
	G4424<=G489 and G3192;
	G4425<=G536 and G2845;
	G4427<=I8431 and I8432;
	G4430<=I8436 and I8437;
	G4433<=G278 and G3097;
	G4434<=G356 and G3131;
	G4435<=G414 and G3160;
	G4436<=G492 and G3192;
	G4437<=G540 and G2845;
	G4445<=I8455 and I8456;
	G4448<=I8460 and I8461;
	G4451<=G359 and G3131;
	G4452<=G437 and G3160;
	G4453<=G495 and G3192;
	G4454<=G544 and G2845;
	G4466<=I8490 and I8491;
	G4469<=I8495 and I8496;
	G4472<=G440 and G3160;
	G4473<=G518 and G3192;
	G4483<=I8523 and I8524;
	G4486<=I8528 and I8529;
	G4490<=G521 and G3192;
	G4491<=G557 and G2845;
	G4494<=I8546 and I8547;
	G4497<=I8551 and I8552;
	G4504<=I8568 and I8569;
	G4507<=I8573 and I8574;
	G4514<=I8588 and I8589;
	G4517<=I8593 and I8594;
	G4526<=G2642 and G741;
	G4529<=I8612 and I8613;
	G4532<=I8617 and I8618;
	G4546<=G2643 and G746;
	G4549<=I8642 and I8643;
	G4681<=G4255 and G3533;
	G4690<=G4081 and G3078;
	G4691<=G4219 and G1690;
	G4699<=G1557 and G4276;
	G4702<=G4243 and G1690;
	G4705<=G190 and G3986;
	G4707<=G812 and G4062;
	G4711<=G190 and G4072;
	G4712<=G1179 and G4276;
	G4720<=G190 and G4055;
	G4724<=G828 and G4038;
	G4728<=G190 and G4179;
	G4729<=G1504 and G4059;
	G4740<=G2242 and G4275;
	G4743<=G3518 and G4286;
	G4744<=G3525 and G4296;
	G4778<=G4169 and G1760;
	G4779<=G4176 and G1760;
	G4781<=G4182 and G1760;
	G4782<=G4187 and G1760;
	G4783<=G948 and G4527;
	G4785<=G1678 and G4202;
	G4787<=G953 and G4547;
	G4789<=G2751 and G4202;
	G4791<=G949 and G4562;
	G4793<=G3887 and G4202;
	G4794<=G954 and G4574;
	G4796<=G950 and G4584;
	G4797<=G3893 and G1616;
	G4798<=G4216 and G1760;
	G4799<=G951 and G4596;
	G4804<=G952 and G3876;
	G4814<=G150 and G4265;
	G4819<=G2573 and G2562 and I9166;
	G4823<=G4238 and G4230 and G174;
	G4825<=G4228 and G1964;
	G4826<=G1545 and G4239;
	G4830<=G4288 and G3723;
	G4832<=G1110 and G4246;
	G4837<=G2573 and G2562 and I9202;
	G4838<=G4517 and G1760;
	G4840<=G4235 and G1980;
	G4868<=G4227 and G4160;
	G4872<=G1924 and G4225 and G4224;
	G4877<=G3746 and G3723 and G4288 and G3764;
	G4878<=G2573 and G2562 and I9222;
	G4883<=G3746 and G3723 and G4288;
	G4901<=G3723 and G4288 and I9261;
	G4902<=G4304 and G2770 and G2746 and G2728;
	G4906<=G4320 and G2728;
	G4933<=G2746 and G2728 and G4320 and G2770;
	G4936<=G214 and G3888;
	G4937<=G3086 and G4309;
	G4955<=G215 and G3891;
	G4956<=G295 and G3892;
	G4957<=G2746 and G2728 and G4320;
	G4958<=G296 and G3897;
	G4959<=G376 and G3898;
	G4961<=G377 and G3904;
	G4962<=G457 and G3905;
	G4968<=G4403 and G1760;
	G4969<=G4362 and G2216;
	G5001<=G458 and G3912;
	G5005<=G2728 and G4320 and I9330;
	G5008<=G231 and G3920;
	G5017<=G211 and G3928;
	G5018<=G232 and G3930;
	G5019<=G312 and G3933;
	G5020<=G579 and G3937;
	G5029<=G212 and G3945;
	G5030<=G233 and G3946;
	G5031<=G292 and G3948;
	G5032<=G313 and G3950;
	G5033<=G393 and G3953;
	G5034<=G583 and G3956;
	G5043<=G213 and G3958;
	G5044<=G234 and G3959;
	G5045<=G293 and G3961;
	G5046<=G314 and G3962;
	G5047<=G373 and G3964;
	G5048<=G394 and G3966;
	G5049<=G474 and G3969;
	G5050<=G587 and G3970;
	G5062<=G235 and G3973;
	G5063<=G294 and G3974;
	G5064<=G315 and G3975;
	G5065<=G374 and G3977;
	G5066<=G395 and G3978;
	G5067<=G454 and G3980;
	G5068<=G475 and G3982;
	G5069<=G566 and G3983;
	G5077<=G236 and G3988;
	G5078<=G316 and G3989;
	G5079<=G375 and G3990;
	G5080<=G396 and G3991;
	G5081<=G455 and G3993;
	G5082<=G476 and G3994;
	G5089<=G273 and G3998;
	G5090<=G317 and G4000;
	G5091<=G397 and G4001;
	G5092<=G456 and G4002;
	G5093<=G477 and G4003;
	G5094<=G535 and G4004;
	G5096<=G1149 and G4400;
	G5104<=G274 and G4010;
	G5105<=G354 and G4013;
	G5106<=G398 and G4015;
	G5107<=G478 and G4016;
	G5108<=G539 and G4017;
	G5116<=G355 and G4021;
	G5117<=G435 and G4024;
	G5118<=G479 and G4026;
	G5119<=G543 and G4027;
	G5122<=G436 and G4030;
	G5123<=G516 and G4033;
	G5125<=G517 and G4036;
	G5126<=G556 and G4037;
	G5132<=I9534 and I9535;
	G5142<=G1677 and G4202;
	G5287<=G786 and G4724;
	G5298<=G1912 and G4814;
	G5313<=G4820 and G2407;
	G5314<=G1509 and G4729;
	G5334<=G4887 and G2424;
	G5425<=G1528 and G4916;
	G5428<=G775 and G4707;
	G5432<=G1537 and G4921;
	G5436<=G1541 and G4926;
	G5438<=G1545 and G4932;
	G5441<=G4870 and G3497;
	G5442<=G4679 and G4202;
	G5443<=G1549 and G4935;
	G5452<=G4876 and G3499;
	G5458<=G4686 and G1616;
	G5475<=G3801 and G5022;
	G5479<=G5141 and G5037;
	G5484<=G1037 and G5096;
	G5489<=G4912 and G5053;
	G5513<=G4889 and G5071;
	G5547<=G4814 and G1819;
	G5548<=G1549 and G4826;
	G5552<=G1114 and G4832;
	G5560<=G3390 and G5036;
	G5563<=G3390 and G5070;
	G5570<=G1759 and G4841;
	G5573<=G3011 and G4841;
	G5579<=G4090 and G4841;
	G5583<=G1775 and G4969;
	G5585<=G4741 and G4841;
	G5588<=G3028 and G4969;
	G5593<=G4110 and G4969;
	G5599<=G4745 and G4969;
	G5624<=G5140 and G2794;
	G5699<=G1667 and G4841;
	G5700<=G1638 and G4969;
	G5714<=G1532 and G4733;
	G5765<=G1695 and G5428;
	G5767<=G5344 and G3079;
	G5783<=G1897 and G5287;
	G5817<=G5395 and G3091;
	G5894<=G1118 and G5552;
	G5937<=G5562 and G2407;
	G5969<=G5564 and G2424;
	G5970<=G5605 and G2424;
	G5984<=G1041 and G5484;
	G6001<=G5540 and G2407;
	G6002<=G5539 and G2407;
	G6003<=G3716 and G5633 and I10597;
	G6005<=G5557 and G2407;
	G6006<=G5575 and G2424;
	G6013<=G5589 and G2424;
	G6021<=G5594 and G2424;
	G6022<=G5595 and G2424;
	G6039<=G1037 and G5574;
	G6040<=G1462 and G5578;
	G6041<=G5189 and G4969;
	G6042<=G1041 and G5581;
	G6043<=G1069 and G5582;
	G6044<=G1467 and G5584;
	G6045<=G1472 and G5591;
	G6046<=G1073 and G5592;
	G6047<=G1477 and G5596;
	G6049<=G1045 and G5597;
	G6052<=G1049 and G5604;
	G6053<=G1053 and G5608;
	G6054<=G1057 and G5611;
	G6055<=G5239 and G4202;
	G6056<=G3760 and G5286 and G1695;
	G6057<=G1061 and G5617;
	G6058<=G5561 and G3501;
	G6060<=G1065 and G5623;
	G6061<=G5257 and G1616;
	G6091<=G5712 and G5038;
	G6098<=G5681 and G1247;
	G6105<=G5618 and G2817;
	G6107<=G5478 and G1849;
	G6109<=G5453 and G5335;
	G6112<=G5673 and G4841 and G5541;
	G6125<=G5548 and G4202;
	G6145<=G1489 and G5705;
	G6151<=G1494 and G5709;
	G6154<=G1499 and G5713;
	G6157<=G1130 and G5717;
	G6160<=G1504 and G5718;
	G6162<=G1134 and G5724;
	G6166<=G1509 and G5725;
	G6168<=G1138 and G5191;
	G6171<=G5363 and G4841;
	G6172<=G1514 and G5192;
	G6175<=G4332 and G5614;
	G6176<=G1149 and G5198;
	G6182<=G1519 and G5199;
	G6196<=G4927 and G5615;
	G6204<=G5542 and G5294;
	G6239<=G1514 and G5314;
	G6266<=G1481 and G5285;
	G6268<=G1092 and G5309;
	G6394<=G5988 and G5494;
	G6395<=G2157 and G6007;
	G6396<=G661 and G6008;
	G6399<=G5971 and G5494;
	G6400<=G150 and G6011;
	G6401<=G5971 and G5367;
	G6402<=G665 and G6012;
	G6405<=G5956 and G5494;
	G6406<=G154 and G6018;
	G6407<=G5956 and G5367;
	G6408<=G669 and G6019;
	G6409<=G706 and G6020;
	G6411<=G5918 and G5494;
	G6412<=G158 and G6024;
	G6413<=G5939 and G5367;
	G6414<=G673 and G6025;
	G6415<=G5988 and G5367;
	G6416<=G710 and G6026;
	G6417<=G718 and G6027;
	G6418<=G5897 and G5494;
	G6419<=G162 and G6032;
	G6420<=G5918 and G5367;
	G6421<=G5847 and G5384;
	G6422<=G714 and G6033;
	G6423<=G5897 and G5384;
	G6428<=G5874 and G5494;
	G6429<=G168 and G6035;
	G6430<=G5874 and G5384;
	G6431<=G5847 and G5494;
	G6433<=G778 and G6134;
	G6434<=G855 and G6048;
	G6437<=G859 and G6050;
	G6438<=G4829 and G6051;
	G6439<=G789 and G6150;
	G6444<=G1676 and G6125;
	G6447<=G734 and G6073;
	G6448<=G5918 and G5384;
	G6456<=G6116 and G2407;
	G6460<=G6178 and G2424;
	G6462<=G6215 and G2424;
	G6464<=G6177 and G2424;
	G6474<=G6203 and G2424;
	G6487<=G5750 and G4969;
	G6541<=G6144 and G3510;
	G6554<=G5762 and G1616;
	G6567<=G6265 and G2424;
	G6574<=G1045 and G5984;
	G6577<=G6142 and G4160;
	G6578<=G6218 and G3913;
	G6582<=G1122 and G5894;
	G6611<=G3390 and G6249;
	G6629<=G6023 and G4841;
	G6633<=G5526 and G5987;
	G6638<=G174 and G5755;
	G6641<=G5939 and G5494;
	G6643<=G1860 and G5868;
	G6689<=G1519 and G6239;
	G6715<=G677 and G5843;
	G6726<=G5897 and G5367;
	G6727<=G681 and G5846;
	G6732<=G5874 and G5367;
	G6733<=G685 and G5873;
	G6738<=G5847 and G5367;
	G6743<=G730 and G5916;
	G6745<=G1872 and G6198;
	G6753<=G5939 and G5384;
	G6757<=G5874 and G5412;
	G6762<=G5847 and G5412;
	G6771<=G146 and G6004;
	G6908<=G6478 and G5246;
	G6914<=G6483 and G5246;
	G6915<=G6493 and G5246;
	G6916<=G727 and G6515;
	G6923<=G6570 and G5612;
	G6941<=G1126 and G6582;
	G6949<=G5483 and G6589;
	G6951<=G5511 and G6595;
	G6954<=G5518 and G6601;
	G6965<=G55 and G6489;
	G6966<=G6580 and G5580;
	G6970<=G5035 and G6490;
	G6971<=G6424 and G4969;
	G6972<=G5661 and G6498;
	G6974<=G3613 and G6505;
	G6976<=G4399 and G6508;
	G6979<=G5095 and G6511;
	G6990<=G799 and G6517;
	G6991<=G5689 and G6520;
	G6992<=G6610 and G3519;
	G6994<=G3658 and G6538;
	G6995<=G6435 and G1616;
	G6996<=G3678 and G6552;
	G6998<=G4474 and G6555;
	G6999<=G815 and G6556;
	G7001<=G3722 and G6562;
	G7002<=G6770 and G5054;
	G7003<=G1462 and G6689;
	G7007<=G6627 and G5072;
	G7008<=G6615 and G5083;
	G7010<=G1049 and G6574;
	G7017<=G3390 and G6706;
	G7021<=G3390 and G6673;
	G7027<=G3390 and G6698;
	G7030<=G6705 and G5723;
	G7031<=G3390 and G6717;
	G7033<=G6716 and G5190;
	G7036<=G6728 and G5197;
	G7038<=G6466 and G4841;
	G7041<=G6734 and G5206;
	G7071<=G6639 and G1872;
	G7079<=G4259 and G6677;
	G7087<=G6440 and G5311;
	G7096<=G6677 and G5101;
	G7128<=G6926 and G3047;
	G7136<=G4057 and G6953;
	G7175<=G6893 and G4841;
	G7177<=G7016 and G5586;
	G7179<=G6121 and G7035;
	G7181<=G6124 and G7039;
	G7182<=G6902 and G4969;
	G7183<=G6132 and G7042;
	G7184<=G6138 and G7043;
	G7186<=G6600 and G7044;
	G7192<=G7026 and G3526;
	G7193<=G6911 and G1616;
	G7195<=G6984 and G4226;
	G7197<=G7093 and G5055;
	G7199<=G1467 and G7003;
	G7212<=G1053 and G7010;
	G7215<=G6111 and G6984;
	G7217<=G1142 and G6941;
	G7228<=G6688 and G7090;
	G7232<=G6694 and G7091;
	G7235<=G6699 and G7094;
	G7238<=G6707 and G7098;
	G7240<=G6719 and G6894;
	G7242<=G7081 and G6899;
	G7252<=G3591 and G6977;
	G7271<=G6436 and G6922;
	G7278<=G6965 and G1745;
	G7282<=G5830 and G6939;
	G7323<=G4065 and G7171;
	G7412<=G7121 and G4841;
	G7415<=G7222 and G5603;
	G7416<=G7140 and G4969;
	G7417<=G7144 and G1616;
	G7419<=G7230 and G3530;
	G7427<=G1472 and G7199;
	G7429<=G1057 and G7212;
	G7449<=G7272 and G6901;
	G7536<=G4414 and G7367;
	G7537<=G7363 and G7411;
	G7552<=G7319 and G5749;
	G7553<=G7367 and G4135;
	G7554<=G7367 and G4139;
	G7557<=G7367 and G4147;
	G7559<=G7367 and G4155;
	G7561<=G7367 and G4163;
	G7564<=G7367 and G4172;
	G7596<=G7428 and G7028;
	G7597<=G7316 and G4841;
	G7598<=G7483 and G3466;
	G7600<=G7460 and G3466;
	G7602<=G7476 and G3466;
	G7604<=G7456 and G3466;
	G7605<=G7435 and G5607;
	G7606<=G7471 and G3466;
	G7607<=G7325 and G4969;
	G7608<=G7367 and G4169;
	G7609<=G7467 and G3466;
	G7611<=G7367 and G4507;
	G7614<=G7367 and G4176;
	G7615<=G7488 and G3466;
	G7616<=G7367 and G4517;
	G7625<=G7367 and G4182;
	G7626<=G7463 and G3466;
	G7628<=G7367 and G4532;
	G7631<=G7367 and G4187;
	G7632<=G7445 and G3548;
	G7634<=G7367 and G4549;
	G7652<=G7367 and G4194;
	G7653<=G7480 and G5754;
	G7654<=G7367 and G4142;
	G7657<=G7367 and G4201;
	G7658<=G7367 and G4150;
	G7676<=G7367 and G4216;
	G7677<=G7503 and G5073;
	G7678<=G7367 and G4158;
	G7679<=G7447 and G5084;
	G7680<=G7367 and G4166;
	G7681<=G7444 and G5099;
	G7683<=G1061 and G7429;
	G7689<=G7367 and G4417;
	G7691<=G7367 and G4427;
	G7692<=G7367 and G4430;
	G7693<=G7367 and G4445;
	G7694<=G7367 and G4448;
	G7695<=G7367 and G4466;
	G7696<=G7367 and G4469;
	G7698<=G7367 and G4483;
	G7699<=G7367 and G4486;
	G7700<=G7367 and G4494;
	G7701<=G7367 and G4497;
	G7703<=G7367 and G4504;
	G7705<=G7367 and G4514;
	G7709<=G7367 and G4529;
	G7713<=G4403 and G7367;
	G7724<=G7337 and G5938;
	G7827<=G7575 and G7173;
	G7832<=G5343 and G7599;
	G7833<=G6461 and G7601;
	G7837<=G6470 and G7610;
	G8059<=G7682 and G7032;
	G8060<=G7535 and G4841;
	G8062<=G7476 and G7634;
	G8064<=G7483 and G7634;
	G8066<=G7488 and G7634;
	G8068<=G7687 and G5610;
	G8069<=G7456 and G7634;
	G8070<=G863 and G7616;
	G8071<=G7540 and G4969;
	G8074<=G855 and G7616;
	G8075<=G7460 and G7634;
	G8076<=G7690 and G3521;
	G8077<=G859 and G7616;
	G8078<=G7463 and G7634;
	G8079<=G831 and G7658;
	G8080<=G7467 and G7634;
	G8081<=G834 and G7658;
	G8087<=G7471 and G7634;
	G8088<=G837 and G7658;
	G8089<=G840 and G7658;
	G8090<=G843 and G7658;
	G8147<=G1065 and G7683;
	G8150<=G846 and G7658;
	G8151<=G849 and G7658;
	G8153<=G852 and G7658;
	G8229<=G8180 and G5680;
	G8237<=G89 and G8131;
	G8238<=G100 and G8131;
	G8256<=G95 and G8131;
	G8257<=G146 and G8042;
	G8258<=G142 and G8111;
	G8259<=G4538 and G7855;
	G8260<=G138 and G8111;
	G8261<=G174 and G8042;
	G8262<=G4554 and G7855;
	G8263<=G4555 and G7905;
	G8264<=G105 and G8131;
	G8265<=G134 and G8111;
	G8266<=G2157 and G8042;
	G8267<=G154 and G8042;
	G8268<=G4568 and G7905;
	G8269<=G4569 and G7951;
	G8270<=G110 and G8131;
	G8271<=G130 and G8111;
	G8272<=G158 and G8042;
	G8273<=G185 and G8156;
	G8274<=G4580 and G7951;
	G8275<=G4581 and G7993;
	G8276<=G150 and G8042;
	G8277<=G162 and G8042;
	G8278<=G4589 and G7993;
	G8280<=G114 and G8111;
	G8281<=G168 and G8042;
	G8282<=G179 and G8156;
	G8283<=G267 and G7838;
	G8285<=G118 and G8111;
	G8286<=G180 and G8156;
	G8287<=G4500 and G7855;
	G8288<=G270 and G7838;
	G8289<=G348 and G7870;
	G8290<=G588 and G8181;
	G8291<=G122 and G8111;
	G8292<=G181 and G8156;
	G8293<=G4510 and G7855;
	G8294<=G281 and G7838;
	G8295<=G4512 and G7905;
	G8296<=G351 and G7870;
	G8297<=G429 and G7920;
	G8298<=G553 and G8181;
	G8299<=G591 and G8181;
	G8300<=G126 and G8111;
	G8301<=G182 and G8156;
	G8302<=G4521 and G7855;
	G8303<=G284 and G7838;
	G8304<=G4523 and G7905;
	G8305<=G362 and G7870;
	G8306<=G4525 and G7951;
	G8307<=G432 and G7920;
	G8308<=G510 and G7966;
	G8309<=G550 and G8181;
	G8310<=G573 and G8181;
	G8311<=G4540 and G7905;
	G8312<=G365 and G7870;
	G8313<=G4542 and G7951;
	G8314<=G443 and G7920;
	G8315<=G4544 and G7993;
	G8316<=G513 and G7966;
	G8317<=G547 and G8181;
	G8318<=G183 and G8156;
	G8319<=G255 and G7838;
	G8320<=G4557 and G7951;
	G8321<=G446 and G7920;
	G8322<=G4559 and G7993;
	G8323<=G524 and G7966;
	G8325<=G184 and G8156;
	G8326<=G258 and G7838;
	G8327<=G336 and G7870;
	G8328<=G4571 and G7993;
	G8329<=G527 and G7966;
	G8330<=G261 and G7838;
	G8331<=G339 and G7870;
	G8332<=G417 and G7920;
	G8333<=G563 and G8181;
	G8334<=G264 and G7838;
	G8335<=G342 and G7870;
	G8336<=G420 and G7920;
	G8337<=G498 and G7966;
	G8338<=G570 and G8181;
	G8339<=G345 and G7870;
	G8340<=G423 and G7920;
	G8341<=G501 and G7966;
	G8359<=G642 and G7793;
	G8361<=G426 and G7920;
	G8362<=G504 and G7966;
	G8377<=G507 and G7966;
	G8378<=G677 and G7887;
	G8379<=G691 and G7793;
	G8380<=G681 and G7887;
	G8382<=G685 and G7887;
	G8383<=G730 and G7937;
	G8384<=G636 and G7793;
	G8385<=G695 and G7811;
	G8403<=G639 and G7793;
	G8404<=G710 and G7937;
	G8405<=G741 and G8018;
	G8438<=G649 and G7793;
	G8439<=G699 and G7811;
	G8440<=G714 and G7937;
	G8441<=G746 and G8018;
	G8455<=G652 and G7793;
	G8456<=G703 and G7811;
	G8457<=G724 and G7811;
	G8458<=G756 and G8199;
	G8459<=G655 and G7793;
	G8460<=G757 and G8199;
	G8461<=G658 and G7793;
	G8462<=G49 and G8199;
	G8513<=G718 and G7937;
	G8542<=G661 and G7887;
	G8543<=G706 and G7887;
	G8584<=G8146 and G7034;
	G8607<=G8154 and G5616;
	G8609<=G7828 and G4969;
	G8610<=G665 and G7887;
	G8611<=G669 and G7887;
	G8612<=G673 and G7887;
	G8620<=G751 and G8199;
	G8621<=G734 and G7937;
	G8622<=G738 and G7811;
	G8623<=G755 and G8199;
	G8624<=G754 and G8199;
	G8626<=G752 and G8199;
	G8628<=G753 and G8199;
	G8643<=G547 and G8094;
	G8645<=G550 and G8094;
	G8646<=G553 and G8094;
	G8648<=G588 and G8094;
	G8650<=G591 and G8094;
	G8652<=G563 and G8094;
	G8653<=G573 and G8094;
	G8654<=G570 and G8094;
	G8660<=G1069 and G8147;
	G8686<=G3819 and G8342;
	G8687<=G3488 and G8363;
	G8688<=G3812 and G8342;
	G8690<=G3485 and G8363;
	G8691<=G3805 and G8342;
	G8692<=G3462 and G8363;
	G8693<=G3798 and G8342;
	G8695<=G2709 and G8363;
	G8696<=G3743 and G8342;
	G8697<=G3761 and G8342;
	G8698<=G3774 and G8342;
	G8700<=G3784 and G8342;
	G8701<=G2700 and G8363;
	G8702<=G2837 and G8386;
	G8703<=G3574 and G8407;
	G8704<=G2829 and G8386;
	G8705<=G2798 and G8421;
	G8708<=G3557 and G8407;
	G8709<=G2818 and G8386;
	G8710<=G2790 and G8421;
	G8711<=G3542 and G8407;
	G8712<=G2804 and G8386;
	G8713<=G2777 and G8421;
	G8714<=G2873 and G8407;
	G8715<=G2761 and G8386;
	G8716<=G3506 and G8443;
	G8717<=G2764 and G8421;
	G8718<=G2774 and G8386;
	G8719<=G2821 and G8443;
	G8720<=G3825 and G8421;
	G8721<=G2703 and G8464;
	G8722<=G2787 and G8386;
	G8723<=G2706 and G8421;
	G8724<=G3822 and G8464;
	G8725<=G3008 and G8493;
	G8726<=G2795 and G8386;
	G8727<=G2724 and G8421;
	G8728<=G3815 and G8464;
	G8729<=G2999 and G8493;
	G8730<=G2863 and G8407;
	G8731<=G2743 and G8421;
	G8732<=G3808 and G8464;
	G8733<=G2996 and G8493;
	G8735<=G2807 and G8443;
	G8736<=G3771 and G8464;
	G8737<=G2992 and G8493;
	G8738<=G8619 and G3338;
	G8739<=G3780 and G8464;
	G8740<=G2966 and G8493;
	G8741<=G3787 and G8464;
	G8742<=G2973 and G8493;
	G8744<=G3802 and G8464;
	G8745<=G2982 and G8493;
	G8748<=G2721 and G8483;
	G8749<=G2989 and G8493;
	G8764<=G8231 and G4969;
	G8779<=G8634 and G7037;
	G8793<=G8637 and G5622;
	G8813<=G255 and G8524;
	G8814<=G3880 and G8463;
	G8815<=G258 and G8524;
	G8816<=G336 and G8545;
	G8817<=G4545 and G8482;
	G8820<=G261 and G8524;
	G8821<=G339 and G8545;
	G8822<=G417 and G8564;
	G8823<=G4561 and G8512;
	G8824<=G264 and G8524;
	G8825<=G342 and G8545;
	G8826<=G420 and G8564;
	G8827<=G498 and G8585;
	G8828<=G4573 and G8541;
	G8829<=G267 and G8524;
	G8830<=G345 and G8545;
	G8831<=G423 and G8564;
	G8832<=G501 and G8585;
	G8833<=G4583 and G8562;
	G8835<=G270 and G8524;
	G8836<=G348 and G8545;
	G8837<=G426 and G8564;
	G8838<=G504 and G8585;
	G8839<=G4050 and G8581;
	G8840<=G4590 and G8582;
	G8841<=G351 and G8545;
	G8842<=G429 and G8564;
	G8843<=G507 and G8585;
	G8844<=G4056 and G8602;
	G8845<=G432 and G8564;
	G8846<=G510 and G8585;
	G8848<=G281 and G8524;
	G8849<=G513 and G8585;
	G8851<=G284 and G8524;
	G8852<=G362 and G8545;
	G8853<=G365 and G8545;
	G8854<=G443 and G8564;
	G8857<=G446 and G8564;
	G8858<=G524 and G8585;
	G8860<=G527 and G8585;
	G8876<=G8769 and G6102;
	G8877<=G8773 and G6104;
	G8878<=G8777 and G6106;
	G8879<=G8782 and G6108;
	G8892<=G8681 and G4969;
	G8901<=G8804 and G5631;
	G8911<=G8798 and G7688;
	G8912<=G8796 and G8239;
	G8914<=G8795 and G8239;
	G8915<=G8794 and G8239;
	G8919<=G4567 and G8743;
	G8920<=G4578 and G8746;
	G8921<=G4579 and G8747;
	G8922<=G4586 and G8750;
	G8923<=G4587 and G8751;
	G8924<=G4588 and G8752;
	G8925<=G4592 and G8754;
	G8926<=G4593 and G8755;
	G8927<=G4594 and G8756;
	G8928<=G4595 and G8757;
	G8929<=G3865 and G8759;
	G8930<=G3866 and G8760;
	G8931<=G3867 and G8761;
	G8932<=G3868 and G8762;
	G8933<=G4511 and G8765;
	G8934<=G3873 and G8766;
	G8935<=G3874 and G8767;
	G8936<=G3875 and G8768;
	G8937<=G4524 and G8770;
	G8938<=G3878 and G8771;
	G8939<=G3879 and G8772;
	G8940<=G4543 and G8775;
	G8941<=G3882 and G8776;
	G8942<=G4522 and G8780;
	G8943<=G4560 and G8781;
	G8944<=G4539 and G8783;
	G8945<=G4541 and G8784;
	G8946<=G4556 and G8786;
	G8947<=G4558 and G8787;
	G8948<=G4570 and G8789;
	G8949<=G4572 and G8790;
	G8950<=G4582 and G8791;
	G8951<=G8785 and G6072;
	G8952<=G8788 and G6075;
	G8953<=G8758 and G6093;
	G8954<=G8763 and G6097;
	G8961<=G8885 and G5317;
	G8962<=G8890 and G5317;
	G8963<=G8891 and G5317;
	G8976<=G8903 and G6588;
	G8978<=G8909 and G5587;
	G9012<=G8908 and G8239;
	G9013<=G8907 and G8239;
	G9014<=G8906 and G8239;
	G9015<=G8905 and G8239;
	G9016<=G8904 and G8239;
	G9021<=G8886 and G5317;
	G9022<=G8887 and G5317;
	G9023<=G8888 and G5317;
	G9024<=G8884 and G5317;
	G9025<=G8889 and G5317;
	G9037<=G8965 and G5345;
	G9038<=G8966 and G5345;
	G9080<=G9011 and G5598;
	G9084<=G8964 and G5345;
	G9118<=G9046 and G5345;
	G9119<=G9049 and G5345;
	G9120<=G9052 and G5345;
	G9130<=G9054 and G5345;
	G9131<=G9055 and G5345;
	G9142<=G9124 and G6059;
	G9143<=G9122 and G6089;
	G9144<=G9123 and G6096;
	G9146<=G9135 and G6101;
	G9147<=G9136 and G6103;
	G9158<=G9137 and G6070;
	G9159<=G9138 and G6074;
	G9160<=G9139 and G6092;
	G9226<=G9220 and G5403;
	G9238<=G4748 and G9223;
	G9240<=G9223 and G5261;
	G9247<=G4748 and G9227;
	G9251<=G4748 and G9230;
	G9258<=G9227 and G5628;
	G9259<=G9230 and G5639;
	G9270<=G4748 and G9241;
	G9271<=G4748 and G9244;
	G9272<=G4748 and G9248;
	G9273<=G4748 and G9252;
	G9274<=G4748 and G9255;
	G9275<=G9241 and G5645;
	G9276<=G9244 and G5649;
	G9277<=G9248 and G5654;
	G9278<=G9252 and G5658;
	G9279<=G9255 and G5665;
	G9327<=G9316 and G5757;
	G9328<=G9324 and G6465;
	G9334<=G9318 and G6205;
	G9335<=G9320 and G6206;
	G9343<=G9328 and G1738;
	G9344<=G9329 and G6211;
	G9345<=G9330 and G6217;
	G9346<=G9331 and G6222;
	G9347<=G9332 and G6226;
	G9348<=G9333 and G6229;
	G9349<=G9340 and G5690;
	G9359<=G4748 and G9340;
	G9371<=G9352 and G5917;
	G9384<=G9383 and G6245;
	I7994<=G3430 and G3398 and G3359 and G3341;
	I7995<=G2074 and G3287 and G2020 and G3238;
	I8000<=G3430 and G3398 and G3359 and G3341;
	I8001<=G2074 and G3287 and G2020 and G1987;
	I8005<=G3430 and G3398 and G3359 and G2106;
	I8006<=G2074 and G3287 and G2020 and G3238;
	I8014<=G3430 and G3398 and G3359 and G3341;
	I8015<=G2074 and G2057 and G3264 and G3238;
	I8019<=G3430 and G3398 and G3359 and G2106;
	I8020<=G2074 and G3287 and G2020 and G1987;
	I8028<=G3430 and G3398 and G3359 and G3341;
	I8029<=G2074 and G2057 and G3264 and G1987;
	I8033<=G3430 and G3398 and G3359 and G2106;
	I8034<=G2074 and G2057 and G3264 and G3238;
	I8040<=G3430 and G3398 and G3359 and G3341;
	I8041<=G2074 and G2057 and G2020 and G3238;
	I8045<=G3430 and G3398 and G3359 and G2106;
	I8046<=G2074 and G2057 and G3264 and G1987;
	I8052<=G2162 and G2149 and G2137 and G2106;
	I8053<=G3316 and G3287 and G3264 and G3238;
	I8057<=G3430 and G3398 and G3359 and G3341;
	I8058<=G2074 and G2057 and G2020 and G1987;
	I8063<=G2162 and G2149 and G2137 and G2106;
	I8064<=G3316 and G3287 and G3264 and G1987;
	I8071<=G2162 and G2149 and G2137 and G2106;
	I8072<=G3316 and G3287 and G2020 and G3238;
	I8078<=G2162 and G2149 and G2137 and G2106;
	I8079<=G3316 and G3287 and G2020 and G1987;
	I8089<=G2162 and G2149 and G2137 and G2106;
	I8090<=G3316 and G2057 and G2020 and G3238;
	I8108<=G2162 and G2149 and G2137 and G2106;
	I8109<=G2074 and G3287 and G3264 and G3238;
	I8114<=G2162 and G2149 and G2137 and G2106;
	I8115<=G2074 and G3287 and G3264 and G1987;
	I8127<=G2699 and G2674 and G2677;
	I8143<=G2674 and G2677 and G2680;
	I8157<=G2686 and G2689 and G2692;
	I8186<=G3778 and G3549 and G3568 and G3583;
	I8209<=G2298 and G2316 and G2334;
	I8237<=G2298 and G2316 and G2354;
	I8240<=G2298 and G2316 and G2334 and G2354;
	I8288<=G3666 and G3684 and G3694;
	I8296<=G3666 and G3684 and G3707;
	I8299<=G3666 and G3684 and G3694 and G3707;
	I8400<=G3430 and G3398 and G3359 and G3341;
	I8401<=G3316 and G3287 and G3264 and G3238;
	I8412<=G3430 and G3398 and G3359 and G3341;
	I8413<=G3316 and G3287 and G3264 and G1987;
	I8417<=G3430 and G3398 and G3359 and G2106;
	I8418<=G3316 and G3287 and G3264 and G3238;
	I8431<=G3430 and G3398 and G3359 and G3341;
	I8432<=G3316 and G3287 and G2020 and G3238;
	I8436<=G3430 and G3398 and G3359 and G2106;
	I8437<=G3316 and G3287 and G3264 and G1987;
	I8455<=G3430 and G3398 and G3359 and G3341;
	I8456<=G3316 and G3287 and G2020 and G1987;
	I8460<=G3430 and G3398 and G3359 and G2106;
	I8461<=G3316 and G3287 and G2020 and G3238;
	I8490<=G3430 and G3398 and G3359 and G3341;
	I8491<=G3316 and G2057 and G3264 and G3238;
	I8495<=G3430 and G3398 and G3359 and G2106;
	I8496<=G3316 and G3287 and G2020 and G1987;
	I8523<=G3430 and G3398 and G3359 and G3341;
	I8524<=G3316 and G2057 and G3264 and G1987;
	I8528<=G3430 and G3398 and G3359 and G2106;
	I8529<=G3316 and G2057 and G3264 and G3238;
	I8546<=G3430 and G3398 and G3359 and G3341;
	I8547<=G3316 and G2057 and G2020 and G3238;
	I8551<=G3430 and G3398 and G3359 and G2106;
	I8552<=G3316 and G2057 and G3264 and G1987;
	I8568<=G3430 and G3398 and G3359 and G3341;
	I8569<=G3316 and G2057 and G2020 and G1987;
	I8573<=G3430 and G3398 and G3359 and G2106;
	I8574<=G3316 and G2057 and G2020 and G3238;
	I8588<=G3430 and G3398 and G3359 and G3341;
	I8589<=G2074 and G3287 and G3264 and G3238;
	I8593<=G3430 and G3398 and G3359 and G2106;
	I8594<=G3316 and G2057 and G2020 and G1987;
	I8612<=G3430 and G3398 and G3359 and G3341;
	I8613<=G2074 and G3287 and G3264 and G1987;
	I8617<=G3430 and G3398 and G3359 and G2106;
	I8618<=G2074 and G3287 and G3264 and G3238;
	I8642<=G3430 and G3398 and G3359 and G2106;
	I8643<=G2074 and G3287 and G3264 and G1987;
	I9166<=G4041 and G2595 and G2584;
	I9202<=G2605 and G4044 and G2584;
	I9222<=G4041 and G4044 and G2584;
	I9261<=G3777 and G3764 and G3746;
	I9330<=G2784 and G2770 and G2746;
	I9534<=G3019 and G3029 and G3038 and G3052;
	I9535<=G3062 and G2712 and G4253 and G2752;
	I10597<=G3769 and G3754 and G3735;
	G1678<= not (I5506 and I5507);
	G1682<= not (I5520 and I5521);
	G1759<= not (I5599 and I5600);
	G1775<= not (I5620 and I5621);
	G1819<= not (I5696 and I5697);
	G1910<= not (G1435 and G1439);
	G2051<= not (G1444 and G1450);
	G2294<= not (I6065 and I6066);
	G2315<= not (I6103 and I6104);
	G2330<= not (I6134 and I6135);
	G2333<= not (G985 and G990);
	G2352<= not (I6171 and I6172);
	G2367<= not (I6202 and I6203);
	G2378<= not (I6233 and I6234);
	G2385<= not (I6258 and I6259);
	G2395<= not (I6274 and I6275);
	G2474<= not (G1405 and G1412);
	G2751<= not (I6500 and I6501);
	G2783<= not (I6523 and I6524);
	G2801<= not (I6539 and I6540);
	G2995<= not (I6740 and I6741);
	G3011<= not (I6751 and I6752);
	G3012<= not (I6758 and I6759);
	G3028<= not (I6775 and I6776);
	G3083<= not (I6814 and I6815);
	G3129<= not (I6843 and I6844);
	G3221<= not (I6877 and I6878);
	G3231<= not (G1889 and G1904);
	G3232<= not (G2298 and G2276);
	G3286<= not (I6905 and I6906);
	G3314<= not (I6917 and I6918);
	G3315<= not (I6924 and I6925);
	G3358<= not (I6940 and I6941);
	G3518<= not (I6997 and I6998);
	G3525<= not (I7010 and I7011);
	G3602<= not (I7069 and I7070);
	G3613<= not (I7086 and I7087);
	G3656<= not (I7139 and I7140);
	G3658<= not (I7149 and I7150);
	G3665<= not (I7157 and I7158);
	G3678<= not (I7173 and I7174);
	G3679<= not (I7180 and I7181);
	G3680<= not (I7187 and I7188);
	G3681<= not (G866 and G2368);
	G3706<= not (G1556 and G2510);
	G3722<= not (I7215 and I7216);
	G3767<= not (I7240 and I7241);
	G3811<= not (I7269 and I7270);
	G3818<= not (I7278 and I7279);
	G3883<= not (G2276 and G3188);
	G3886<= not (I7422 and I7423);
	G3887<= not (I7429 and I7430);
	G3889<= not (I7437 and I7438);
	G3890<= not (I7444 and I7445);
	G3893<= not (I7453 and I7454);
	G3894<= not (I7460 and I7461);
	G3895<= not (I7467 and I7468);
	G3899<= not (I7479 and I7480);
	G3900<= not (I7486 and I7487);
	G3906<= not (I7504 and I7505);
	G3907<= not (I7511 and I7512);
	G3914<= not (I7532 and I7533);
	G3915<= not (I7539 and I7540);
	G3924<= not (I7568 and I7569);
	G3925<= not (I7575 and I7576);
	G3938<= not (I7610 and I7611);
	G3939<= not (I7617 and I7618);
	G4090<= not (I7892 and I7893);
	G4110<= not (I7938 and I7939);
	G4219<= not (I8120 and I8121);
	G4227<= not (I8133 and I8134);
	G4228<= not (G1408 and G2665);
	G4231<= not (G2276 and G3258);
	G4235<= not (G1415 and G2668);
	G4237<= not (I8151 and I8152);
	G4243<= not (I8165 and I8166);
	G4244<= not (G3549 and G3533);
	G4252<= not (G2276 and G3313);
	G4256<= not (G3233 and G1444);
	G4263<= not (G3260 and G1435);
	G4294<= not (I8244 and I8245);
	G4298<= not (I8254 and I8255);
	G4305<= not (G3712 and G3700 and G3732);
	G4309<= not (G3002 and G3124 and G3659);
	G4310<= not (G3666 and G2460);
	G4313<= not (G3712 and G3700);
	G4332<= not (G3681 and G2368);
	G4359<= not (I8327 and I8328);
	G4363<= not (I8339 and I8340);
	G4399<= not (I8393 and I8394);
	G4456<= not (I8471 and I8472);
	G4474<= not (I8503 and I8504);
	G4476<= not (I8511 and I8512);
	G4492<= not (I8537 and I8538);
	G4502<= not (I8559 and I8560);
	G4513<= not (I8582 and I8583);
	G4528<= not (I8606 and I8607);
	G4548<= not (I8636 and I8637);
	G4563<= not (I8659 and I8660);
	G4575<= not (I8679 and I8680);
	G4679<= not (I8939 and I8940);
	G4686<= not (I8956 and I8957);
	G4700<= not (G2460 and G4271);
	G4714<= not (G4344 and G4335 and G4328);
	G4741<= not (I9058 and I9059);
	G4745<= not (I9070 and I9071);
	G4810<= not (I9152 and I9153);
	G4820<= not (I9170 and I9171);
	G4821<= not (G4220 and G3605);
	G4824<= not (I9182 and I9183);
	G4831<= not (G3635 and G3605 and G4220);
	G4835<= not (I9195 and I9196);
	G4836<= not (G4288 and G1879);
	G4839<= not (G1879 and G4269);
	G4869<= not (G4254 and G3533);
	G4871<= not (G3635 and G3605 and G4220 and G3644);
	G4879<= not (G2595 and G2584 and G4270 and G4281);
	G4880<= not (G4287 and G1879);
	G4881<= not (G2460 and G4315);
	G4887<= not (I9234 and I9235);
	G4889<= not (I9242 and I9243);
	G4893<= not (G2460 and G4312);
	G4905<= not (G4282 and G3533);
	G4910<= not (G2460 and G4314);
	G4911<= not (G4320 and G2044);
	G4912<= not (I9277 and I9278);
	G4954<= not (G4319 and G2460);
	G5035<= not (I9382 and I9383);
	G5095<= not (I9476 and I9477);
	G5141<= not (I9548 and I9549);
	G5189<= not (I9692 and I9693);
	G5239<= not (I9746 and I9747);
	G5257<= not (I9768 and I9769);
	G5284<= not (G4344 and G4335 and G4963);
	G5291<= not (G4344 and G5002 and G4963);
	G5305<= not (G5009 and G4335 and G4328);
	G5310<= not (G5009 and G4335 and G4963);
	G5312<= not (G5009 and G5002 and G4963);
	G5363<= not (I9827 and I9828);
	G5512<= not (G1879 and G4877);
	G5538<= not (G5132 and G1266);
	G5539<= not (I9947 and I9948);
	G5540<= not (I9954 and I9955);
	G5546<= not (I9964 and I9965);
	G5550<= not (G1879 and G4830);
	G5555<= not (I9979 and I9980);
	G5556<= not (I9986 and I9987);
	G5557<= not (I9993 and I9994);
	G5558<= not (I10000 and I10001);
	G5559<= not (G5132 and G1257);
	G5562<= not (I10010 and I10011);
	G5564<= not (I10018 and I10019);
	G5565<= not (G2044 and G4933);
	G5567<= not (G1879 and G4883);
	G5568<= not (G2044 and G4902 and G4320);
	G5575<= not (I10039 and I10040);
	G5576<= not (G4894 and G4888 and G4884);
	G5589<= not (I10061 and I10062);
	G5590<= not (G2044 and G4906);
	G5594<= not (I10072 and I10073);
	G5595<= not (I10079 and I10080);
	G5605<= not (I10093 and I10094);
	G5625<= not (G2044 and G4957);
	G5632<= not (G2276 and G4901);
	G5657<= not (G5021 and G4381);
	G5661<= not (I10143 and I10144);
	G5672<= not (G5056 and G5039 and G5023);
	G5681<= not (G5132 and G2043);
	G5686<= not (G5132 and G1263);
	G5689<= not (I10197 and I10198);
	G5697<= not (G2044 and G5005);
	G5712<= not (I10224 and I10225);
	G5747<= not (I10299 and I10300);
	G5748<= not (I10306 and I10307);
	G5750<= not (I10314 and I10315);
	G5751<= not (I10321 and I10322);
	G5752<= not (I10328 and I10329);
	G5753<= not (I10335 and I10336);
	G5762<= not (I10360 and I10361);
	G6023<= not (I10626 and I10627);
	G6119<= not (I10744 and I10745);
	G6142<= not (I10790 and I10791);
	G6153<= not (I10819 and I10820);
	G6158<= not (G3735 and G3716 and G5633 and G3754);
	G6159<= not (I10835 and I10836);
	G6163<= not (G5633 and G3716);
	G6164<= not (I10848 and I10849);
	G6165<= not (I10855 and I10856);
	G6169<= not (I10867 and I10868);
	G6170<= not (I10874 and I10875);
	G6177<= not (I10889 and I10890);
	G6178<= not (G2205 and G5568);
	G6180<= not (I10900 and I10901);
	G6181<= not (I10907 and I10908);
	G6187<= not (G5633 and G3735 and G3716);
	G6188<= not (I10924 and I10925);
	G6203<= not (I10953 and I10954);
	G6215<= not (I10981 and I10982);
	G6218<= not (I10992 and I10993);
	G6265<= not (I11079 and I11080);
	G6273<= not (I11095 and I11096);
	G6274<= not (I11102 and I11103);
	G6275<= not (I11109 and I11110);
	G6276<= not (I11116 and I11117);
	G6277<= not (I11123 and I11124);
	G6280<= not (I11136 and I11137);
	G6281<= not (I11143 and I11144);
	G6282<= not (I11150 and I11151);
	G6283<= not (I11157 and I11158);
	G6284<= not (I11164 and I11165);
	G6285<= not (I11171 and I11172);
	G6286<= not (I11178 and I11179);
	G6287<= not (I11185 and I11186);
	G6424<= not (I11550 and I11551);
	G6435<= not (I11575 and I11576);
	G6463<= not (G5918 and G5278);
	G6466<= not (I11615 and I11616);
	G6467<= not (G5956 and G5269);
	G6469<= not (G5918 and G5278);
	G6472<= not (G5971 and G5269);
	G6473<= not (G5269 and G5988);
	G6476<= not (G5939 and G5269);
	G6477<= not (G5269 and G5918);
	G6482<= not (G5269 and G5847);
	G6497<= not (G5278 and G5847);
	G6503<= not (G5269 and G5897);
	G6504<= not (G5269 and G5874);
	G6510<= not (G5278 and G5874);
	G6516<= not (G5897 and G5278);
	G6559<= not (G5814 and G6109);
	G6570<= not (I11751 and I11752);
	G6571<= not (I11758 and I11759);
	G6615<= not (I11842 and I11843);
	G6627<= not (I11874 and I11875);
	G6680<= not (G5403 and G6252);
	G6695<= not (I12016 and I12017);
	G6701<= not (I12032 and I12033);
	G6709<= not (I12052 and I12053);
	G6722<= not (I12079 and I12080);
	G6770<= not (I12180 and I12181);
	G6893<= not (I12551 and I12552);
	G6902<= not (I12576 and I12577);
	G6911<= not (I12597 and I12598);
	G7065<= not (I12833 and I12834);
	G7069<= not (G5435 and G6680);
	G7082<= not (I12853 and I12854);
	G7093<= not (I12870 and I12871);
	G7121<= not (I12952 and I12953);
	G7140<= not (I13003 and I13004);
	G7144<= not (I13017 and I13018);
	G7234<= not (G3757 and G3739 and G7050 and G3770);
	G7237<= not (G7050 and G3739);
	G7244<= not (G7050 and G3757 and G3739);
	G7257<= not (I13214 and I13215);
	G7316<= not (I13377 and I13378);
	G7325<= not (I13396 and I13397);
	G7444<= not (I13588 and I13589);
	G7447<= not (I13599 and I13600);
	G7480<= not (I13639 and I13640);
	G7503<= not (I13686 and I13687);
	G7535<= not (I13786 and I13787);
	G7540<= not (I13801 and I13802);
	G7828<= not (I14245 and I14246);
	G8231<= not (I14473 and I14474);
	G8239<= not (G8073 and G8092);
	G8627<= not (G6232 and G8091);
	G8633<= not (G8176 and G6232);
	G8681<= not (I14838 and I14839);
	G8798<= not (G6984 and G8644);
	G9179<= not (I15818 and I15819);
	G9190<= not (I15849 and I15850);
	G9191<= not (I15856 and I15857);
	G9192<= not (I15863 and I15864);
	G9202<= not (I15881 and I15882);
	G9203<= not (I15888 and I15889);
	G9205<= not (I15898 and I15899);
	I5505<= not (G1532 and G1528);
	I5506<= not (G1532 and I5505);
	I5507<= not (G1528 and I5505);
	I5519<= not (G1087 and G1098);
	I5520<= not (G1087 and I5519);
	I5521<= not (G1098 and I5519);
	I5598<= not (G1481 and G1489);
	I5599<= not (G1481 and I5598);
	I5600<= not (G1489 and I5598);
	I5619<= not (G1092 and G1130);
	I5620<= not (G1092 and I5619);
	I5621<= not (G1130 and I5619);
	I5695<= not (G1513 and G1524);
	I5696<= not (G1513 and I5695);
	I5697<= not (G1524 and I5695);
	I6064<= not (G852 and G883);
	I6065<= not (G852 and I6064);
	I6066<= not (G883 and I6064);
	I6102<= not (G849 and G921);
	I6103<= not (G849 and I6102);
	I6104<= not (G921 and I6102);
	I6133<= not (G846 and G916);
	I6134<= not (G846 and I6133);
	I6135<= not (G916 and I6133);
	I6170<= not (G843 and G911);
	I6171<= not (G843 and I6170);
	I6172<= not (G911 and I6170);
	I6201<= not (G831 and G891);
	I6202<= not (G831 and I6201);
	I6203<= not (G891 and I6201);
	I6232<= not (G834 and G896);
	I6233<= not (G834 and I6232);
	I6234<= not (G896 and I6232);
	I6257<= not (G837 and G901);
	I6258<= not (G837 and I6257);
	I6259<= not (G901 and I6257);
	I6273<= not (G840 and G906);
	I6274<= not (G840 and I6273);
	I6275<= not (G906 and I6273);
	I6499<= not (G1913 and G1537);
	I6500<= not (G1913 and I6499);
	I6501<= not (G1537 and I6499);
	I6522<= not (G1919 and G1102);
	I6523<= not (G1919 and I6522);
	I6524<= not (G1102 and I6522);
	I6538<= not (G2555 and G2557);
	I6539<= not (G2555 and I6538);
	I6540<= not (G2557 and I6538);
	I6739<= not (G195 and G1970);
	I6740<= not (G195 and I6739);
	I6741<= not (G1970 and I6739);
	I6750<= not (G1733 and G1494);
	I6751<= not (G1733 and I6750);
	I6752<= not (G1494 and I6750);
	I6757<= not (G186 and G1983);
	I6758<= not (G186 and I6757);
	I6759<= not (G1983 and I6757);
	I6774<= not (G2386 and G1134);
	I6775<= not (G2386 and I6774);
	I6776<= not (G1134 and I6774);
	I6813<= not (G210 and G2052);
	I6814<= not (G210 and I6813);
	I6815<= not (G2052 and I6813);
	I6842<= not (G205 and G2016);
	I6843<= not (G205 and I6842);
	I6844<= not (G2016 and I6842);
	I6876<= not (G1967 and G1910);
	I6877<= not (G1967 and I6876);
	I6878<= not (G1910 and I6876);
	I6904<= not (G2105 and G1838);
	I6905<= not (G2105 and I6904);
	I6906<= not (G1838 and I6904);
	I6916<= not (G2360 and G1732);
	I6917<= not (G2360 and I6916);
	I6918<= not (G1732 and I6916);
	I6923<= not (G1728 and G33);
	I6924<= not (G1728 and I6923);
	I6925<= not (G33 and I6923);
	I6939<= not (G2161 and G2051);
	I6940<= not (G2161 and I6939);
	I6941<= not (G2051 and I6939);
	I6996<= not (G2275 and G2242);
	I6997<= not (G2275 and I6996);
	I6998<= not (G2242 and I6996);
	I7009<= not (G2295 and G2333);
	I7010<= not (G2295 and I7009);
	I7011<= not (G2333 and I7009);
	I7068<= not (G1639 and G1643);
	I7069<= not (G1639 and I7068);
	I7070<= not (G1643 and I7068);
	I7085<= not (G1753 and G1918);
	I7086<= not (G1753 and I7085);
	I7087<= not (G1918 and I7085);
	I7138<= not (G2404 and G2397);
	I7139<= not (G2404 and I7138);
	I7140<= not (G2397 and I7138);
	I7148<= not (G799 and G1974);
	I7149<= not (G799 and I7148);
	I7150<= not (G1974 and I7148);
	I7156<= not (G2331 and G929);
	I7157<= not (G2331 and I7156);
	I7158<= not (G929 and I7156);
	I7172<= not (G1739 and G2006);
	I7173<= not (G1739 and I7172);
	I7174<= not (G2006 and I7172);
	I7179<= not (G2351 and G795);
	I7180<= not (G2351 and I7179);
	I7181<= not (G795 and I7179);
	I7186<= not (G2353 and G1834);
	I7187<= not (G2353 and I7186);
	I7188<= not (G1834 and I7186);
	I7214<= not (G815 and G2091);
	I7215<= not (G815 and I7214);
	I7216<= not (G2091 and I7214);
	I7239<= not (G1658 and G2134);
	I7240<= not (G1658 and I7239);
	I7241<= not (G2134 and I7239);
	I7268<= not (G2486 and G955);
	I7269<= not (G2486 and I7268);
	I7270<= not (G955 and I7268);
	I7277<= not (G2497 and G1898);
	I7278<= not (G2497 and I7277);
	I7279<= not (G1898 and I7277);
	I7421<= not (G2525 and G2703);
	I7422<= not (G2525 and I7421);
	I7423<= not (G2703 and I7421);
	I7428<= not (G3222 and G1541);
	I7429<= not (G3222 and I7428);
	I7430<= not (G1541 and I7428);
	I7436<= not (G2517 and G3822);
	I7437<= not (G2517 and I7436);
	I7438<= not (G3822 and I7436);
	I7443<= not (G2973 and G1701);
	I7444<= not (G2973 and I7443);
	I7445<= not (G1701 and I7443);
	I7452<= not (G3226 and G1106);
	I7453<= not (G3226 and I7452);
	I7454<= not (G1106 and I7452);
	I7459<= not (G2506 and G3815);
	I7460<= not (G2506 and I7459);
	I7461<= not (G3815 and I7459);
	I7466<= not (G2982 and G1704);
	I7467<= not (G2982 and I7466);
	I7468<= not (G1704 and I7466);
	I7478<= not (G2502 and G3808);
	I7479<= not (G2502 and I7478);
	I7480<= not (G3808 and I7478);
	I7485<= not (G2989 and G1708);
	I7486<= not (G2989 and I7485);
	I7487<= not (G1708 and I7485);
	I7503<= not (G2498 and G3802);
	I7504<= not (G2498 and I7503);
	I7505<= not (G3802 and I7503);
	I7510<= not (G2992 and G1711);
	I7511<= not (G2992 and I7510);
	I7512<= not (G1711 and I7510);
	I7531<= not (G2487 and G3787);
	I7532<= not (G2487 and I7531);
	I7533<= not (G3787 and I7531);
	I7538<= not (G2996 and G1715);
	I7539<= not (G2996 and I7538);
	I7540<= not (G1715 and I7538);
	I7567<= not (G2481 and G3780);
	I7568<= not (G2481 and I7567);
	I7569<= not (G3780 and I7567);
	I7574<= not (G2999 and G1718);
	I7575<= not (G2999 and I7574);
	I7576<= not (G1718 and I7574);
	I7609<= not (G2471 and G3771);
	I7610<= not (G2471 and I7609);
	I7611<= not (G3771 and I7609);
	I7616<= not (G3008 and G1721);
	I7617<= not (G3008 and I7616);
	I7618<= not (G1721 and I7616);
	I7891<= not (G2979 and G1499);
	I7892<= not (G2979 and I7891);
	I7893<= not (G1499 and I7891);
	I7937<= not (G3614 and G1138);
	I7938<= not (G3614 and I7937);
	I7939<= not (G1138 and I7937);
	I8119<= not (G1904 and G3220);
	I8120<= not (G1904 and I8119);
	I8121<= not (G3220 and I8119);
	I8132<= not (G3232 and G1646);
	I8133<= not (G3232 and I8132);
	I8134<= not (G1646 and I8132);
	I8150<= not (G3229 and G38);
	I8151<= not (G3229 and I8150);
	I8152<= not (G38 and I8150);
	I8164<= not (G1943 and G3231);
	I8165<= not (G1943 and I8164);
	I8166<= not (G3231 and I8164);
	I8243<= not (G2011 and G3506);
	I8244<= not (G2011 and I8243);
	I8245<= not (G3506 and I8243);
	I8253<= not (G2454 and G3825);
	I8254<= not (G2454 and I8253);
	I8255<= not (G3825 and I8253);
	I8326<= not (G2011 and G2721);
	I8327<= not (G2011 and I8326);
	I8328<= not (G2721 and I8326);
	I8338<= not (G2966 and G1698);
	I8339<= not (G2966 and I8338);
	I8340<= not (G1698 and I8338);
	I8392<= not (G2949 and G1925);
	I8393<= not (G2949 and I8392);
	I8394<= not (G1925 and I8392);
	I8470<= not (G2525 and G2821);
	I8471<= not (G2525 and I8470);
	I8472<= not (G2821 and I8470);
	I8502<= not (G2986 and G2038);
	I8503<= not (G2986 and I8502);
	I8504<= not (G2038 and I8502);
	I8510<= not (G2517 and G2807);
	I8511<= not (G2517 and I8510);
	I8512<= not (G2807 and I8510);
	I8536<= not (G2506 and G2798);
	I8537<= not (G2506 and I8536);
	I8538<= not (G2798 and I8536);
	I8558<= not (G2502 and G2790);
	I8559<= not (G2502 and I8558);
	I8560<= not (G2790 and I8558);
	I8581<= not (G2498 and G2777);
	I8582<= not (G2498 and I8581);
	I8583<= not (G2777 and I8581);
	I8605<= not (G2487 and G2764);
	I8606<= not (G2487 and I8605);
	I8607<= not (G2764 and I8605);
	I8635<= not (G2481 and G2743);
	I8636<= not (G2481 and I8635);
	I8637<= not (G2743 and I8635);
	I8658<= not (G2471 and G2724);
	I8659<= not (G2471 and I8658);
	I8660<= not (G2724 and I8658);
	I8678<= not (G2467 and G2706);
	I8679<= not (G2467 and I8678);
	I8680<= not (G2706 and I8678);
	I8938<= not (G4239 and G1545);
	I8939<= not (G4239 and I8938);
	I8940<= not (G1545 and I8938);
	I8955<= not (G4246 and G1110);
	I8956<= not (G4246 and I8955);
	I8957<= not (G1110 and I8955);
	I9057<= not (G4059 and G1504);
	I9058<= not (G4059 and I9057);
	I9059<= not (G1504 and I9057);
	I9069<= not (G4400 and G1149);
	I9070<= not (G4400 and I9069);
	I9071<= not (G1149 and I9069);
	I9151<= not (G3883 and G1649);
	I9152<= not (G3883 and I9151);
	I9153<= not (G1649 and I9151);
	I9169<= not (G1935 and G4244);
	I9170<= not (G1935 and I9169);
	I9171<= not (G4244 and I9169);
	I9181<= not (G4231 and G2007);
	I9182<= not (G4231 and I9181);
	I9183<= not (G2007 and I9181);
	I9194<= not (G4252 and G1652);
	I9195<= not (G4252 and I9194);
	I9196<= not (G1652 and I9194);
	I9233<= not (G4310 and G2180);
	I9234<= not (G4310 and I9233);
	I9235<= not (G2180 and I9233);
	I9241<= not (G2540 and G4305);
	I9242<= not (G2540 and I9241);
	I9243<= not (G4305 and I9241);
	I9276<= not (G2533 and G4313);
	I9277<= not (G2533 and I9276);
	I9278<= not (G4313 and I9276);
	I9381<= not (G4062 and G1908);
	I9382<= not (G4062 and I9381);
	I9383<= not (G1908 and I9381);
	I9475<= not (G4038 and G1942);
	I9476<= not (G4038 and I9475);
	I9477<= not (G1942 and I9475);
	I9547<= not (G1952 and G4307);
	I9548<= not (G1952 and I9547);
	I9549<= not (G4307 and I9547);
	I9691<= not (G5096 and G1037);
	I9692<= not (G5096 and I9691);
	I9693<= not (G1037 and I9691);
	I9745<= not (G4826 and G1549);
	I9746<= not (G4826 and I9745);
	I9747<= not (G1549 and I9745);
	I9767<= not (G4832 and G1114);
	I9768<= not (G4832 and I9767);
	I9769<= not (G1114 and I9767);
	I9826<= not (G4729 and G1509);
	I9827<= not (G4729 and I9826);
	I9828<= not (G1509 and I9826);
	I9946<= not (G2128 and G4905);
	I9947<= not (G2128 and I9946);
	I9948<= not (G4905 and I9946);
	I9953<= not (G2131 and G4831);
	I9954<= not (G2131 and I9953);
	I9955<= not (G4831 and I9953);
	I9963<= not (G1938 and G4869);
	I9964<= not (G1938 and I9963);
	I9965<= not (G4869 and I9963);
	I9978<= not (G4880 and G2092);
	I9979<= not (G4880 and I9978);
	I9980<= not (G2092 and I9978);
	I9985<= not (G4836 and G2096);
	I9986<= not (G4836 and I9985);
	I9987<= not (G2096 and I9985);
	I9992<= not (G2145 and G4871);
	I9993<= not (G2145 and I9992);
	I9994<= not (G4871 and I9992);
	I9999<= not (G4839 and G1929);
	I10000<= not (G4839 and I9999);
	I10001<= not (G1929 and I9999);
	I10009<= not (G1949 and G4821);
	I10010<= not (G1949 and I10009);
	I10011<= not (G4821 and I10009);
	I10017<= not (G4700 and G2174);
	I10018<= not (G4700 and I10017);
	I10019<= not (G2174 and I10017);
	I10038<= not (G4893 and G2202);
	I10039<= not (G4893 and I10038);
	I10040<= not (G2202 and I10038);
	I10060<= not (G4910 and G2226);
	I10061<= not (G4910 and I10060);
	I10062<= not (G2226 and I10060);
	I10071<= not (G4954 and G2253);
	I10072<= not (G4954 and I10071);
	I10073<= not (G2253 and I10071);
	I10078<= not (G4911 and G2256);
	I10079<= not (G4911 and I10078);
	I10080<= not (G2256 and I10078);
	I10092<= not (G4881 and G2177);
	I10093<= not (G4881 and I10092);
	I10094<= not (G2177 and I10092);
	I10142<= not (G4707 and G1916);
	I10143<= not (G4707 and I10142);
	I10144<= not (G1916 and I10142);
	I10196<= not (G4724 and G1958);
	I10197<= not (G4724 and I10196);
	I10198<= not (G1958 and I10196);
	I10223<= not (G2522 and G4895);
	I10224<= not (G2522 and I10223);
	I10225<= not (G4895 and I10223);
	I10298<= not (G5461 and G2562);
	I10299<= not (G5461 and I10298);
	I10300<= not (G2562 and I10298);
	I10305<= not (G5470 and G3019);
	I10306<= not (G5470 and I10305);
	I10307<= not (G3019 and I10305);
	I10313<= not (G5484 and G1041);
	I10314<= not (G5484 and I10313);
	I10315<= not (G1041 and I10313);
	I10320<= not (G5459 and G2573);
	I10321<= not (G5459 and I10320);
	I10322<= not (G2573 and I10320);
	I10327<= not (G5467 and G2562);
	I10328<= not (G5467 and I10327);
	I10329<= not (G2562 and I10327);
	I10334<= not (G5462 and G2573);
	I10335<= not (G5462 and I10334);
	I10336<= not (G2573 and I10334);
	I10359<= not (G5552 and G1118);
	I10360<= not (G5552 and I10359);
	I10361<= not (G1118 and I10359);
	I10625<= not (G5314 and G1514);
	I10626<= not (G5314 and I10625);
	I10627<= not (G1514 and I10625);
	I10743<= not (G5550 and G2100);
	I10744<= not (G5550 and I10743);
	I10745<= not (G2100 and I10743);
	I10789<= not (G5512 and G2170);
	I10790<= not (G5512 and I10789);
	I10791<= not (G2170 and I10789);
	I10818<= not (G5567 and G2039);
	I10819<= not (G5567 and I10818);
	I10820<= not (G2039 and I10818);
	I10834<= not (G5514 and G2584);
	I10835<= not (G5514 and I10834);
	I10836<= not (G2584 and I10834);
	I10847<= not (G5490 and G2595);
	I10848<= not (G5490 and I10847);
	I10849<= not (G2595 and I10847);
	I10854<= not (G5521 and G2584);
	I10855<= not (G5521 and I10854);
	I10856<= not (G2584 and I10854);
	I10866<= not (G5480 and G2605);
	I10867<= not (G5480 and I10866);
	I10868<= not (G2605 and I10866);
	I10873<= not (G5516 and G2595);
	I10874<= not (G5516 and I10873);
	I10875<= not (G2595 and I10873);
	I10888<= not (G5590 and G2259);
	I10889<= not (G5590 and I10888);
	I10890<= not (G2259 and I10888);
	I10899<= not (G5520 and G2752);
	I10900<= not (G5520 and I10899);
	I10901<= not (G2752 and I10899);
	I10906<= not (G5492 and G2605);
	I10907<= not (G5492 and I10906);
	I10908<= not (G2605 and I10906);
	I10923<= not (G5525 and G2752);
	I10924<= not (G5525 and I10923);
	I10925<= not (G2752 and I10923);
	I10952<= not (G5565 and G2340);
	I10953<= not (G5565 and I10952);
	I10954<= not (G2340 and I10952);
	I10980<= not (G5625 and G2210);
	I10981<= not (G5625 and I10980);
	I10982<= not (G2210 and I10980);
	I10991<= not (G5632 and G2389);
	I10992<= not (G5632 and I10991);
	I10993<= not (G2389 and I10991);
	I11078<= not (G5697 and G2511);
	I11079<= not (G5697 and I11078);
	I11080<= not (G2511 and I11078);
	I11094<= not (G5515 and G2734);
	I11095<= not (G5515 and I11094);
	I11096<= not (G2734 and I11094);
	I11101<= not (G5491 and G2712);
	I11102<= not (G5491 and I11101);
	I11103<= not (G2712 and I11101);
	I11108<= not (G5522 and G2734);
	I11109<= not (G5522 and I11108);
	I11110<= not (G2734 and I11108);
	I11115<= not (G5481 and G3062);
	I11116<= not (G5481 and I11115);
	I11117<= not (G3062 and I11115);
	I11122<= not (G5517 and G2712);
	I11123<= not (G5517 and I11122);
	I11124<= not (G2712 and I11122);
	I11135<= not (G5476 and G3052);
	I11136<= not (G5476 and I11135);
	I11137<= not (G3052 and I11135);
	I11142<= not (G5493 and G3062);
	I11143<= not (G5493 and I11142);
	I11144<= not (G3062 and I11142);
	I11149<= not (G5473 and G3038);
	I11150<= not (G5473 and I11149);
	I11151<= not (G3038 and I11149);
	I11156<= not (G5482 and G3052);
	I11157<= not (G5482 and I11156);
	I11158<= not (G3052 and I11156);
	I11163<= not (G5469 and G3029);
	I11164<= not (G5469 and I11163);
	I11165<= not (G3029 and I11163);
	I11170<= not (G5477 and G3038);
	I11171<= not (G5477 and I11170);
	I11172<= not (G3038 and I11170);
	I11177<= not (G5466 and G3019);
	I11178<= not (G5466 and I11177);
	I11179<= not (G3019 and I11177);
	I11184<= not (G5474 and G3029);
	I11185<= not (G5474 and I11184);
	I11186<= not (G3029 and I11184);
	I11549<= not (G5984 and G1045);
	I11550<= not (G5984 and I11549);
	I11551<= not (G1045 and I11549);
	I11574<= not (G5894 and G1122);
	I11575<= not (G5894 and I11574);
	I11576<= not (G1122 and I11574);
	I11614<= not (G6239 and G1519);
	I11615<= not (G6239 and I11614);
	I11616<= not (G1519 and I11614);
	I11750<= not (G6112 and G1486);
	I11751<= not (G6112 and I11750);
	I11752<= not (G1486 and I11750);
	I11757<= not (G1758 and G6118);
	I11758<= not (G1758 and I11757);
	I11759<= not (G6118 and I11757);
	I11841<= not (G2548 and G6158);
	I11842<= not (G2548 and I11841);
	I11843<= not (G6158 and I11841);
	I11873<= not (G2543 and G6187);
	I11874<= not (G2543 and I11873);
	I11875<= not (G6187 and I11873);
	I12015<= not (G5874 and G5847);
	I12016<= not (G5874 and I12015);
	I12017<= not (G5847 and I12015);
	I12031<= not (G5918 and G5897);
	I12032<= not (G5918 and I12031);
	I12033<= not (G5897 and I12031);
	I12051<= not (G5956 and G5939);
	I12052<= not (G5956 and I12051);
	I12053<= not (G5939 and I12051);
	I12078<= not (G5988 and G5971);
	I12079<= not (G5988 and I12078);
	I12080<= not (G5971 and I12078);
	I12179<= not (G1961 and G6163);
	I12180<= not (G1961 and I12179);
	I12181<= not (G6163 and I12179);
	I12550<= not (G6689 and G1462);
	I12551<= not (G6689 and I12550);
	I12552<= not (G1462 and I12550);
	I12575<= not (G6574 and G1049);
	I12576<= not (G6574 and I12575);
	I12577<= not (G1049 and I12575);
	I12596<= not (G6582 and G1126);
	I12597<= not (G6582 and I12596);
	I12598<= not (G1126 and I12596);
	I12832<= not (G6722 and G6709);
	I12833<= not (G6722 and I12832);
	I12834<= not (G6709 and I12832);
	I12852<= not (G6701 and G6695);
	I12853<= not (G6701 and I12852);
	I12854<= not (G6695 and I12852);
	I12869<= not (G2536 and G6618);
	I12870<= not (G2536 and I12869);
	I12871<= not (G6618 and I12869);
	I12951<= not (G7003 and G1467);
	I12952<= not (G7003 and I12951);
	I12953<= not (G1467 and I12951);
	I13002<= not (G7010 and G1053);
	I13003<= not (G7010 and I13002);
	I13004<= not (G1053 and I13002);
	I13016<= not (G6941 and G1142);
	I13017<= not (G6941 and I13016);
	I13018<= not (G1142 and I13016);
	I13213<= not (G7065 and G7082);
	I13214<= not (G7065 and I13213);
	I13215<= not (G7082 and I13213);
	I13376<= not (G7199 and G1472);
	I13377<= not (G7199 and I13376);
	I13378<= not (G1472 and I13376);
	I13395<= not (G7212 and G1057);
	I13396<= not (G7212 and I13395);
	I13397<= not (G1057 and I13395);
	I13587<= not (G2556 and G7234);
	I13588<= not (G2556 and I13587);
	I13589<= not (G7234 and I13587);
	I13598<= not (G2551 and G7244);
	I13599<= not (G2551 and I13598);
	I13600<= not (G7244 and I13598);
	I13638<= not (G7257 and G7069);
	I13639<= not (G7257 and I13638);
	I13640<= not (G7069 and I13638);
	I13685<= not (G1977 and G7237);
	I13686<= not (G1977 and I13685);
	I13687<= not (G7237 and I13685);
	I13785<= not (G7427 and G1477);
	I13786<= not (G7427 and I13785);
	I13787<= not (G1477 and I13785);
	I13800<= not (G7429 and G1061);
	I13801<= not (G7429 and I13800);
	I13802<= not (G1061 and I13800);
	I14244<= not (G7683 and G1065);
	I14245<= not (G7683 and I14244);
	I14246<= not (G1065 and I14244);
	I14472<= not (G8147 and G1069);
	I14473<= not (G8147 and I14472);
	I14474<= not (G1069 and I14472);
	I14837<= not (G8660 and G1073);
	I14838<= not (G8660 and I14837);
	I14839<= not (G1073 and I14837);
	I15817<= not (G9151 and G9148);
	I15818<= not (G9151 and I15817);
	I15819<= not (G9148 and I15817);
	I15848<= not (G9162 and G9154);
	I15849<= not (G9162 and I15848);
	I15850<= not (G9154 and I15848);
	I15855<= not (G9168 and G9165);
	I15856<= not (G9168 and I15855);
	I15857<= not (G9165 and I15855);
	I15862<= not (G9174 and G9171);
	I15863<= not (G9174 and I15862);
	I15864<= not (G9171 and I15862);
	I15880<= not (G9190 and G9179);
	I15881<= not (G9190 and I15880);
	I15882<= not (G9179 and I15880);
	I15887<= not (G9192 and G9191);
	I15888<= not (G9192 and I15887);
	I15889<= not (G9191 and I15887);
	I15897<= not (G9202 and G9203);
	I15898<= not (G9202 and I15897);
	I15899<= not (G9203 and I15897);
	G1690<=G1021 or G1025 or G1018;
	G1872<=G971 or G962 or G972 or I5757;
	G1955<=G1189 or G16;
	G2043<=G1263 or G1257;
	G2206<=G1363 or G1364 or G1365 or G1366;
	G2213<=G1367 or G1368 or G1369 or G1370;
	G2214<=G1376 or G1377 or G1378 or G1379;
	G2229<=G1371 or G1372 or G1373 or G1374;
	G2230<=G1380 or G1381 or G1382 or G1383;
	G2262<=G1384 or G1385 or G1386 or G1387;
	G2368<=I6208 or I6209;
	G2845<=G1877 or G576;
	G3097<=G1746 or G287;
	G3131<=G1749 or G368;
	G3160<=G1751 or G449;
	G3192<=G1756 or G530;
	G3339<=G1424 or G2014;
	G3541<=G1663 or G1421;
	G3760<=I7232 or I7233;
	G3986<=G202 or G3129;
	G4055<=G187 or G3012;
	G4072<=G196 or G2995;
	G4179<=G207 or G3083;
	G4249<=G3617 or G1639;
	G4264<=G2490 or G3315;
	G4280<=I8224 or I8225;
	G4283<=G3587 or G2665;
	G4295<=G2828 or G2668;
	G4297<=G3617 or G3602;
	G4364<=G2952 or G1725;
	G4374<=G1182 or G1186 or G1179 or I8363;
	G4413<=G2371 or G3285;
	G4688<=G4193 or G3190;
	G4727<=G4417 or G4172 or G4163 or I9029;
	G4734<=G4469 or G4448 or I9038;
	G4735<=G4427 or G4414 or G4403 or I9041;
	G4736<=G4532 or G4517 or I9044;
	G4737<=G4135 or G4529 or G4514 or I9047;
	G4747<=G3984 or G2912;
	G4786<=G4107 or G4097 or G4124 or I9099;
	G4790<=G4185 or G4131 or G4129 or I9107;
	G4812<=G2490 or G4237;
	G4829<=G863 or G4051;
	G4870<=G4154 or G3081;
	G4876<=G4159 or G4167;
	G4927<=G4318 or G1590;
	G5021<=G943 or G4501;
	G5036<=G4047 or G2972;
	G5040<=G3900 or G3895 or G3890 or G4363;
	G5052<=G4049 or G4054;
	G5057<=G3939 or G3925 or G3915 or G3907;
	G5070<=G4052 or G4058;
	G5138<=G4108 or G3049;
	G5140<=G4333 or G3509;
	G5188<=G5008 or G4365;
	G5193<=G5017 or G4366;
	G5194<=G5018 or G4367;
	G5195<=G5019 or G4368;
	G5196<=G5020 or G4369;
	G5200<=G5029 or G4375;
	G5201<=G5030 or G4376;
	G5202<=G5031 or G4377;
	G5203<=G5032 or G4378;
	G5204<=G5033 or G4379;
	G5205<=G5034 or G4380;
	G5208<=G5043 or G4383;
	G5209<=G5044 or G4384;
	G5210<=G5045 or G4385;
	G5211<=G5046 or G4386;
	G5212<=G5047 or G4387;
	G5213<=G5048 or G4388;
	G5214<=G5049 or G4389;
	G5215<=G5050 or G4390;
	G5216<=G5062 or G4391;
	G5217<=G5063 or G4392;
	G5218<=G5064 or G4393;
	G5219<=G5065 or G4394;
	G5220<=G5066 or G4395;
	G5221<=G5067 or G4396;
	G5222<=G5068 or G4397;
	G5223<=G5069 or G4398;
	G5227<=G5077 or G4407;
	G5228<=G5078 or G4408;
	G5229<=G5079 or G4409;
	G5230<=G5080 or G4410;
	G5231<=G5081 or G4411;
	G5232<=G5082 or G4412;
	G5233<=G5089 or G4420;
	G5234<=G5090 or G4421;
	G5235<=G5091 or G4422;
	G5236<=G5092 or G4423;
	G5237<=G5093 or G4424;
	G5238<=G5094 or G4425;
	G5241<=G5104 or G4433;
	G5242<=G5105 or G4434;
	G5243<=G5106 or G4435;
	G5244<=G5107 or G4436;
	G5245<=G5108 or G4437;
	G5253<=G5116 or G4451;
	G5254<=G5117 or G4452;
	G5255<=G5118 or G4453;
	G5256<=G5119 or G4454;
	G5259<=G5122 or G4472;
	G5260<=G5123 or G4473;
	G5264<=G5125 or G4490;
	G5265<=G5126 or G4491;
	G5317<=G4727 or G4737 or G4735;
	G5343<=G4690 or G2862;
	G5345<=G4736 or G4734;
	G5440<=G4790 or G4786;
	G5483<=G4740 or G4098;
	G5511<=G4743 or G4109;
	G5518<=G4744 or G4118;
	G5537<=G3617 or G4835;
	G5545<=G3617 or G4824;
	G5549<=G2935 or G4712;
	G5561<=G4168 or G4797;
	G5566<=G3617 or G4810;
	G5572<=G5051 or G1236;
	G5673<=G4823 or G4872;
	G5698<=G5057 or G5040;
	G5704<=G4936 or G4334;
	G5706<=G4955 or G4342;
	G5707<=G4956 or G4343;
	G5708<=G2889 or G4699;
	G5710<=G4958 or G4351;
	G5711<=G4959 or G4352;
	G5715<=G4961 or G4355;
	G5716<=G4962 or G4356;
	G5722<=G5001 or G4361;
	G5830<=G5714 or G5142;
	G6115<=G3617 or G5558;
	G6116<=G5546 or G4681;
	G6120<=G3617 or G5555;
	G6121<=G5425 or G4785;
	G6123<=G3617 or G5556;
	G6124<=G5432 or G4789;
	G6132<=G5436 or G4793;
	G6138<=G5438 or G5442;
	G6144<=G4175 or G5458;
	G6249<=G4066 or G5313;
	G6262<=G4074 or G5334;
	G6270<=G1000 or G5335 or G1909;
	G6436<=G6266 or G5699;
	G6440<=G6268 or G5700;
	G6445<=G6105 or G6107;
	G6457<=G6196 or G6209 or G4937;
	G6458<=G6184 or G6259 or G6174 or G6214;
	G6459<=G6259 or G6185 or I11603;
	G6470<=G5817 or G2934;
	G6525<=G6112 or G5547;
	G6543<=G6125 or G1553;
	G6565<=G2396 or G6131 or G1603;
	G6579<=G6098 or G1975;
	G6580<=G6039 or G6041;
	G6585<=G3617 or G6119;
	G6590<=G3617 or G6153;
	G6600<=G5443 or G6055;
	G6602<=G6058 or G3092;
	G6610<=G4180 or G6061;
	G6673<=G4053 or G5937;
	G6685<=G4067 or G5969;
	G6686<=G4068 or G5970;
	G6688<=G6145 or G5570;
	G6694<=G6151 or G5573;
	G6698<=G4073 or G6001;
	G6699<=G6154 or G5579;
	G6705<=G6157 or G5583;
	G6706<=G4077 or G6002;
	G6707<=G6160 or G5585;
	G6710<=G55 or G6264;
	G6716<=G6162 or G5588;
	G6717<=G4082 or G6005;
	G6718<=G4083 or G6006;
	G6719<=G6166 or G6171;
	G6728<=G6168 or G5593;
	G6734<=G6176 or G5599;
	G6735<=G4091 or G6013;
	G6739<=G4099 or G6021;
	G6740<=G4100 or G6022;
	G6906<=G6715 or G6726;
	G6907<=G6727 or G6732;
	G6912<=G4199 or G6567;
	G6913<=G6733 or G6738;
	G6917<=G6743 or G6753;
	G6919<=G6771 or G6394;
	G6920<=G6395 or G6399;
	G6921<=G6396 or G6401;
	G6924<=G6400 or G6405;
	G6925<=G6402 or G6407;
	G6926<=G6406 or G6411;
	G6927<=G6408 or G6413;
	G6928<=G6409 or G6415;
	G6929<=G6412 or G6418;
	G6930<=G6414 or G6420;
	G6931<=G6416 or G6421;
	G6932<=G6417 or G6423;
	G6933<=G6419 or G6428;
	G6934<=G6422 or G6430;
	G6935<=G6429 or G6431;
	G6952<=G6633 or G6204;
	G6964<=G6447 or G6448;
	G6980<=G6745 or G6028;
	G7016<=G6042 or G6487;
	G7020<=G3617 or G6578;
	G7025<=G6541 or G3095;
	G7026<=G4186 or G6554;
	G7029<=G6433 or G5765;
	G7040<=G6439 or G5783;
	G7062<=G4048 or G6456;
	G7080<=G4086 or G6462;
	G7081<=G6172 or G6629;
	G7083<=G5448 or G6267 or G6710;
	G7086<=G4101 or G6464;
	G7088<=G6638 or G6641;
	G7089<=G4128 or G6474;
	G7165<=G6434 or G6908;
	G7166<=G6437 or G6914;
	G7167<=G6438 or G6915;
	G7170<=G6916 or G6444;
	G7191<=G7071 or G6980;
	G7202<=G6028 or G7071;
	G7220<=G1304 or G7062;
	G7222<=G6049 or G6971;
	G7227<=G6992 or G3128;
	G7230<=G4190 or G6995;
	G7248<=G7079 or G5652;
	G7254<=G6923 or G5298;
	G7258<=G7083 or G5403 or I13220;
	G7272<=G6182 or G7038;
	G7337<=G7278 or G4546;
	G7363<=G7136 or G6903;
	G7421<=G6745 or G7202;
	G7426<=G1173 or G7217 or I13553;
	G7428<=G6040 or G7175;
	G7435<=G6052 or G7182;
	G7436<=G7183 or G6975;
	G7438<=G7184 or G6978;
	G7443<=G7192 or G3158;
	G7445<=G4192 or G7193;
	G7450<=G6090 or G7195;
	G7575<=G7323 or G7142;
	G7682<=G6044 or G7412;
	G7687<=G6053 or G7416;
	G7690<=G4181 or G7417;
	G7697<=G7419 or G3187;
	G7782<=G4783 or G7598;
	G7783<=G4787 or G7600;
	G7784<=G7406 or G6664 or G3492 or I14219;
	G7787<=G4791 or G7602;
	G7788<=G4794 or G7604;
	G7791<=G4796 or G7606;
	G7810<=G4799 or G7609;
	G7825<=G4801 or G7615;
	G7826<=G4804 or G7626;
	G7834<=G7724 or G6762;
	G8009<=G3591 or G7406 or G7566 or I14302;
	G8082<=G7654 or G7628 or G7611;
	G8091<=G7215 or G6452 or I14366;
	G8128<=G7566 or G6910 or G6452;
	G8146<=G6045 or G7597;
	G8154<=G6054 or G7607;
	G8155<=G7632 or G3219;
	G8176<=G7566 or G1030 or G6664 or G6452;
	G8613<=G8082 or G7616;
	G8634<=G6047 or G8060;
	G8637<=G6057 or G8071;
	G8758<=G8655 or I14932 or I14933;
	G8763<=G8232 or I14941 or I14942;
	G8769<=I14951 or I14952;
	G8773<=I14959 or I14960;
	G8777<=I14969 or I14970;
	G8782<=G8624 or G8659 or I14980;
	G8785<=G8623 or G8656 or I14985;
	G8788<=G8620 or G8658 or I14990;
	G8794<=G8153 or G8074 or G8069 or G8523;
	G8795<=G8151 or G8077 or G8075 or G8279;
	G8796<=G8150 or G8078 or G8070 or G8360;
	G8804<=G6060 or G8609;
	G8834<=G7096 or G8229;
	G8884<=G8735 or G8818 or I15232;
	G8885<=G8723 or G8806 or I15243;
	G8886<=G8727 or G8812 or I15254;
	G8887<=I15265 or G8819;
	G8888<=I15276 or G8807;
	G8889<=I15283 or I15284 or I15285;
	G8890<=I15290 or I15291 or I15292;
	G8891<=G8705 or G8811 or I15297 or I15298;
	G8893<=G8814 or G8643;
	G8894<=G8817 or G8645;
	G8895<=G8823 or G8646;
	G8896<=G8828 or G8648;
	G8897<=G8833 or G8650;
	G8899<=G8839 or G8652;
	G8900<=G8840 or G8653;
	G8902<=G8844 or G8654;
	G8904<=G8090 or G8080 or G8706;
	G8905<=G8089 or G8087 or G8694;
	G8906<=G8088 or G8062 or G8699;
	G8907<=G8081 or G8064 or G8707;
	G8908<=G8079 or G8066 or G8855;
	G8909<=G6043 or G8764;
	G8964<=G8915 or G8863 or I15400;
	G8965<=G8739 or G8742 or G8914 or G8847;
	G8966<=G8741 or G8745 or G8912 or G8850;
	G8979<=G8919 or G8813;
	G8980<=G8920 or G8815;
	G8981<=G8921 or G8816;
	G8982<=G8922 or G8820;
	G8983<=G8923 or G8821;
	G8984<=G8924 or G8822;
	G8985<=G8925 or G8824;
	G8986<=G8926 or G8825;
	G8987<=G8927 or G8826;
	G8988<=G8928 or G8827;
	G8989<=G8929 or G8829;
	G8990<=G8930 or G8830;
	G8991<=G8931 or G8831;
	G8992<=G8932 or G8832;
	G8993<=G8933 or G8835;
	G8994<=G8934 or G8836;
	G8995<=G8935 or G8837;
	G8996<=G8936 or G8838;
	G8997<=G8937 or G8841;
	G8998<=G8938 or G8842;
	G8999<=G8939 or G8843;
	G9000<=G8940 or G8845;
	G9001<=G8941 or G8846;
	G9002<=G8942 or G8848;
	G9003<=G8943 or G8849;
	G9004<=G8944 or G8851;
	G9005<=G8945 or G8852;
	G9006<=G8946 or G8853;
	G9007<=G8947 or G8854;
	G9008<=G8948 or G8857;
	G9009<=G8949 or G8858;
	G9010<=G8950 or G8860;
	G9011<=G6046 or G8892;
	G9046<=G8744 or G8749 or G9016 or G8862;
	G9049<=G8732 or G8737 or G9015 or G8861;
	G9052<=G8728 or G8733 or G9014 or G8679;
	G9054<=G8724 or G8729 or G9013 or G8680;
	G9055<=G8721 or G8725 or G9012 or G8859;
	G9122<=G8953 or G9084;
	G9123<=G8954 or G9037;
	G9124<=G8876 or G9038;
	G9135<=G8951 or G9130;
	G9136<=G8952 or G9131;
	G9137<=G8877 or G9118;
	G9138<=G8878 or G9119;
	G9139<=G8879 or G9120;
	G9148<=G9143 or G9024;
	G9151<=G9144 or G8961;
	G9154<=G9142 or G9021;
	G9162<=G9158 or G9022;
	G9165<=G9159 or G9023;
	G9168<=G9160 or G9025;
	G9171<=G9146 or G8962;
	G9174<=G9147 or G8963;
	G9239<=G7653 or G9226;
	G9261<=G9238 or G6227;
	G9264<=G9247 or G6242;
	G9267<=G9251 or G6225;
	G9282<=G9270 or G6238;
	G9285<=G9271 or G6221;
	G9288<=G9272 or G6235;
	G9291<=G9273 or G6216;
	G9294<=G9274 or G6230;
	G9337<=G9240 or G9327;
	G9338<=G9258 or G9334;
	G9339<=G9259 or G9335;
	G9352<=G9343 or G4526;
	G9354<=G9275 or G9344;
	G9355<=G9276 or G9345;
	G9356<=G9277 or G9346;
	G9357<=G9278 or G9347;
	G9358<=G9279 or G9348;
	G9363<=G9359 or G6210;
	G9377<=G9371 or G6757;
	G9387<=G9349 or G9384;
	I5757<=G969 or G970 or G966 or G963;
	I6208<=G891 or G896 or G901 or G906;
	I6209<=G911 or G916 or G921 or G883;
	I7232<=G2367 or G2352 or G2378 or G2330;
	I7233<=G2315 or G2385 or G2294 or G2395;
	I8224<=G3019 or G3029 or G3038 or G3052;
	I8225<=G3062 or G2712 or G2734 or G2752;
	I8363<=G2655 or G1163 or G1160;
	I9029<=G4504 or G4494 or G4430;
	I9038<=G4507 or G4497 or G4486;
	I9041<=G4483 or G4466 or G4445;
	I9044<=G4150 or G4142 or G4549;
	I9047<=G4155 or G4147 or G4139;
	I9099<=G4127 or G4123 or G4117;
	I9107<=G4133 or G4145 or G4138 or G4132;
	I11603<=G6193 or G6197 or G6175;
	I13220<=G58 or G6258 or G5418;
	I13553<=G1166 or G1167 or G1170;
	I14219<=G979 or G7566 or G1865;
	I14302<=G6664 or G3492 or G979;
	I14366<=G7566 or G1030 or G6664;
	I14467<=G7993 or G7966 or G7793 or G7811;
	I14468<=G7937 or G7887 or G8029 or G8018;
	I14479<=G7993 or G7966 or G7793 or G7811;
	I14480<=G7937 or G7887 or G8029 or G8018;
	I14484<=G7993 or G7966 or G7793 or G7811;
	I14485<=G7937 or G7887 or G8029 or G8018;
	I14495<=G7993 or G7966 or G7793 or G7811;
	I14496<=G7937 or G7887 or G8029 or G8018;
	I14753<=G7993 or G7966 or G7793 or G7811;
	I14754<=G7937 or G7887 or G8029 or G8018;
	I14758<=G7993 or G7966 or G7793 or G7811;
	I14759<=G7937 or G7887 or G8029 or G8018;
	I14766<=G7993 or G7966 or G7793 or G7811;
	I14767<=G7937 or G7887 or G8029 or G8018;
	I14771<=G7993 or G7966 or G7793 or G7811;
	I14772<=G7937 or G7887 or G8029 or G8018;
	I14831<=G8483 or G8464 or G8514;
	I14834<=G8483 or G8464 or G8514;
	I14932<=G8278 or G8329 or G8461 or G8382;
	I14933<=G8385 or G8404 or G8441 or G8462;
	I14941<=G8275 or G8323 or G8459 or G8380;
	I14942<=G8439 or G8440 or G8405 or G8460;
	I14951<=G8328 or G8316 or G8455 or G8378;
	I14952<=G8456 or G8513 or G8458 or G8236;
	I14959<=G8322 or G8308 or G8438 or G8612;
	I14960<=G8621 or G8622 or G8628 or G8230;
	I14969<=G8315 or G8377 or G8359 or G8611;
	I14970<=G8457 or G8383 or G8626 or G8233;
	I14980<=G8362 or G8403 or G8610;
	I14985<=G8341 or G8384 or G8542;
	I14990<=G8337 or G8379 or G8543;
	I15017<=G8131 or G8111 or G8042 or G8156;
	I15018<=G7855 or G7838 or G7905 or G7870;
	I15019<=G7951 or G7920 or G7983 or G8181;
	I15020<=G8363 or G8342 or G8407 or G8386;
	I15021<=I15017 or I15018 or I15019 or I15020;
	I15029<=G8131 or G8111 or G8042 or G8156;
	I15030<=G7855 or G7838 or G7905 or G7870;
	I15031<=G7951 or G7920 or G7983 or G8181;
	I15032<=G8363 or G8342 or G8407 or G8386;
	I15033<=I15029 or I15030 or I15031 or I15032;
	I15040<=G8131 or G8111 or G8042 or G8156;
	I15041<=G7855 or G7838 or G7905 or G7870;
	I15042<=G7951 or G7920 or G7983 or G8181;
	I15043<=G8363 or G8342 or G8407 or G8386;
	I15044<=I15040 or I15041 or I15042 or I15043;
	I15051<=G8131 or G8111 or G8042 or G8156;
	I15052<=G7855 or G7838 or G7905 or G7870;
	I15053<=G7951 or G7920 or G7983 or G8181;
	I15054<=G8363 or G8342 or G8407 or G8386;
	I15055<=I15051 or I15052 or I15053 or I15054;
	I15071<=G8131 or G8111 or G8042 or G8156;
	I15072<=G7855 or G7838 or G7905 or G7870;
	I15073<=G7951 or G7920 or G7983 or G8181;
	I15074<=G8363 or G8342 or G8407 or G8386;
	I15075<=I15071 or I15072 or I15073 or I15074;
	I15082<=G8131 or G8111 or G8042 or G8156;
	I15083<=G7855 or G7838 or G7905 or G7870;
	I15084<=G7951 or G7920 or G7983 or G8181;
	I15085<=G8363 or G8342 or G8407 or G8386;
	I15086<=I15082 or I15083 or I15084 or I15085;
	I15098<=G8131 or G8111 or G8042 or G8156;
	I15099<=G7855 or G7838 or G7905 or G7870;
	I15100<=G7951 or G7920 or G7983 or G8181;
	I15101<=G8363 or G8342 or G8407 or G8386;
	I15102<=I15098 or I15099 or I15100 or I15101;
	I15109<=G8131 or G8111 or G8042 or G8156;
	I15110<=G7855 or G7838 or G7905 or G7870;
	I15111<=G7951 or G7920 or G7983 or G8181;
	I15112<=G8363 or G8342 or G8407 or G8386;
	I15113<=I15109 or I15110 or I15111 or I15112;
	I15147<=G8483 or G8464 or G8514;
	I15152<=G8483 or G8464 or G8514;
	I15165<=G8483 or G8464 or G8514;
	I15169<=G8483 or G8464 or G8514;
	I15172<=G8483 or G8464 or G8514;
	I15175<=G8483 or G8464 or G8514;
	I15228<=G8270 or G8258 or G8281 or G8273;
	I15229<=G8262 or G8303 or G8268 or G8312;
	I15230<=G8274 or G8321 or G8298 or G8696;
	I15231<=G8701 or G8715 or G8730 or G8720;
	I15232<=I15228 or I15229 or I15230 or I15231;
	I15239<=G8264 or G8260 or G8277 or G8301;
	I15240<=G8259 or G8294 or G8263 or G8305;
	I15241<=G8269 or G8314 or G8309 or G8695;
	I15242<=G8697 or G8714 or G8718 or G8719;
	I15243<=I15239 or I15240 or I15241 or I15242;
	I15250<=G8238 or G8265 or G8272 or G8292;
	I15251<=G8302 or G8288 or G8311 or G8296;
	I15252<=G8320 or G8307 or G8317 or G8692;
	I15253<=G8698 or G8711 or G8722 or G8716;
	I15254<=I15250 or I15251 or I15252 or I15253;
	I15261<=G8256 or G8271 or G8267 or G8286;
	I15262<=G8293 or G8283 or G8304 or G8289;
	I15263<=G8313 or G8297 or G8310 or G8690;
	I15264<=G8700 or G8708 or G8726 or G8731;
	I15265<=I15261 or I15262 or I15263 or I15264;
	I15272<=G8237 or G8300 or G8261 or G8282;
	I15273<=G8287 or G8334 or G8295 or G8339;
	I15274<=G8306 or G8361 or G8299 or G8687;
	I15275<=G8693 or G8703 or G8712 or G8717;
	I15276<=I15272 or I15273 or I15274 or I15275;
	I15283<=G8291 or G8276 or G8325 or G8330;
	I15284<=G8335 or G8340 or G8290 or G8691;
	I15285<=G8709 or G8713 or G8803;
	I15290<=G8285 or G8266 or G8318 or G8326;
	I15291<=G8331 or G8336 or G8338 or G8688;
	I15292<=G8704 or G8710 or G8805;
	I15297<=G8280 or G8257 or G8319 or G8327;
	I15298<=G8332 or G8333 or G8686 or G8702;
	I15400<=G8736 or G8748 or G8740;
	G1964<= not (G1428 or G1429);
	G1980<= not (G1430 or G1431);
	G2014<= not (G1421 or G1416);
	G2521<= not (G65 or G62);
	G3225<= not (G1021 or G1025 or G1889);
	G3233<= not (G1714 or G1459);
	G3237<= not (G1444 or G1838 or G1454);
	G3260<= not (G1728 or G2490);
	G3310<= not (G936 or G2557);
	G3504<= not (G1375 or G2229 or G2213 or G2206);
	G3505<= not (G2263 or G1395);
	G3515<= not (G1388 or G2262 or G2230 or G2214);
	G3516<= not (G2282 or G1401);
	G3528<= not (G2343 or G1391);
	G3555<= not (G2359 or G1398);
	G3790<= not (G985 or G990 or G2295);
	G3885<= not (G3310 or G3466);
	G4160<= not (G1231 or G2834);
	G4232<= not (G1934 or G3591);
	G4318<= not (G3681 or G1590);
	G4349<= not (G2496 or G3310);
	G4354<= not (G1424 or G3541);
	G4676<= not (G3885 or G3094);
	G4884<= not (G4492 or G4476 or G4456 or G4294);
	G4888<= not (G4548 or G4528 or G4513 or G4502);
	G4894<= not (G4298 or G4575 or G4563);
	G5023<= not (G3894 or G3889 or G3886 or G4359);
	G5039<= not (G3924 or G3914 or G3906 or G3899);
	G5056<= not (G3556 or G2872 or G3938);
	G5614<= not (G3002 or G1590 or G4714);
	G5615<= not (G4714 or G3002);
	G5772<= not (G5428 or G1888);
	G6174<= not (G1855 or G5305);
	G6184<= not (G875 or G5291);
	G6185<= not (G5305 or G1590);
	G6193<= not (G1926 or G5310);
	G6197<= not (G875 or G866 or G1590 or G5291);
	G6209<= not (G2332 or G5305);
	G6214<= not (G878 or G5284);
	G6259<= not (G3002 or G5312);
	G6452<= not (G6270 or G2245);
	G6465<= not (G5403 or G5802 or G5769 or G5790);
	G6489<= not (G5802 or G5769 or G5790);
	G6664<= not (G5836 or G1901 or G1788);
	G6910<= not (G1011 or G1837 or G6559 or G1008);
	G7152<= not (G6253 or G7083 or G5418);
	G7209<= not (G1789 or G146 or G6984);
	G7312<= not (G7178 or G6970);
	G7314<= not (G7180 or G6972);
	G7318<= not (G7185 or G6979);
	G7321<= not (G7187 or G6990);
	G7322<= not (G7188 or G6991);
	G7324<= not (G7189 or G6994);
	G7326<= not (G7194 or G6999);
	G7328<= not (G7196 or G7001);
	G7406<= not (G7191 or G1600);
	G7566<= not (G7421 or G1597);
	G8073<= not (G7658 or G7654);
	G8092<= not (G7634 or G7628 or G7616 or G7611);
	G8230<= not (G8199 or I14467 or I14468);
	G8232<= not (G8199 or I14479 or I14480);
	G8233<= not (G8199 or I14484 or I14485);
	G8236<= not (G8199 or I14495 or I14496);
	G8279<= not (G7658 or G7616 or G8082 or G7634);
	G8360<= not (G7658 or G7616 or G8082 or G7634);
	G8523<= not (G7658 or G7616 or G8082 or G7634);
	G8625<= not (G1000 or G6573 or G1860 or G8009);
	G8629<= not (G6270 or G8009);
	G8630<= not (G6110 or G7784 or G3591 or G1864);
	G8635<= not (G1034 or G8128);
	G8641<= not (G6559 or G162 or G7784 or G3591);
	G8644<= not (G4146 or G8128);
	G8655<= not (G8199 or I14753 or I14754);
	G8656<= not (G8199 or I14758 or I14759);
	G8658<= not (G8199 or I14766 or I14767);
	G8659<= not (G8199 or I14771 or I14772);
	G8679<= not (G8493 or G8239 or I14831);
	G8680<= not (G8493 or G8239 or I14834);
	G8694<= not (G7658 or G8613 or G7634);
	G8699<= not (G7658 or G8613 or G7634);
	G8706<= not (G7658 or G8613 or G7634);
	G8707<= not (G7658 or G8613 or G7634);
	G8801<= not (G8635 or G3790);
	G8803<= not (G8443 or G8421 or I15021);
	G8805<= not (G8443 or G8421 or I15033);
	G8806<= not (G8443 or G8421 or I15044);
	G8807<= not (G8443 or G8421 or I15055);
	G8811<= not (G8443 or G8421 or I15075);
	G8812<= not (G8443 or G8421 or I15086);
	G8818<= not (G8443 or G8421 or I15102);
	G8819<= not (G8443 or G8421 or I15113);
	G8847<= not (G8493 or G8239 or I15147);
	G8850<= not (G8493 or G8239 or I15152);
	G8855<= not (G7658 or G8613 or G7634);
	G8859<= not (G8493 or G8239 or I15165);
	G8861<= not (G8493 or G8239 or I15169);
	G8862<= not (G8493 or G8239 or I15172);
	G8863<= not (G8493 or G8239 or I15175);
end RTL;
