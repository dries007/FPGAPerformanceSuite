-- File created by Bench2VHDL
-- Name: s9234
-- File: bench/s9234.bench
-- Timestamp: 2019-05-21T22:08:28.992865
--
-- Original File
-- =============
--	# s9234.1
--	# 36 inputs
--	# 39 outputs
--	# 211 D-type flipflops
--	# 3570 inverters
--	# 2027 gates (955 ANDs + 528 NANDs + 431 ORs + 113 NORs)
--	
--	INPUT(g89)
--	INPUT(g94)
--	INPUT(g98)
--	INPUT(g102)
--	INPUT(g107)
--	INPUT(g301)
--	INPUT(g306)
--	INPUT(g310)
--	INPUT(g314)
--	INPUT(g319)
--	INPUT(g557)
--	INPUT(g558)
--	INPUT(g559)
--	INPUT(g560)
--	INPUT(g561)
--	INPUT(g562)
--	INPUT(g563)
--	INPUT(g564)
--	INPUT(g705)
--	INPUT(g639)
--	INPUT(g567)
--	INPUT(g45)
--	INPUT(g42)
--	INPUT(g39)
--	INPUT(g702)
--	INPUT(g32)
--	INPUT(g38)
--	INPUT(g46)
--	INPUT(g36)
--	INPUT(g47)
--	INPUT(g40)
--	INPUT(g37)
--	INPUT(g41)
--	INPUT(g22)
--	INPUT(g44)
--	INPUT(g23)
--	
--	OUTPUT(g2584)
--	OUTPUT(g3222)
--	OUTPUT(g3600)
--	OUTPUT(g4307)
--	OUTPUT(g4321)
--	OUTPUT(g4422)
--	OUTPUT(g4809)
--	OUTPUT(g5137)
--	OUTPUT(g5468)
--	OUTPUT(g5469)
--	OUTPUT(g5692)
--	OUTPUT(g6282)
--	OUTPUT(g6284)
--	OUTPUT(g6360)
--	OUTPUT(g6362)
--	OUTPUT(g6364)
--	OUTPUT(g6366)
--	OUTPUT(g6368)
--	OUTPUT(g6370)
--	OUTPUT(g6372)
--	OUTPUT(g6374)
--	OUTPUT(g6728)
--	OUTPUT(g1290)
--	OUTPUT(g4121)
--	OUTPUT(g4108)
--	OUTPUT(g4106)
--	OUTPUT(g4103)
--	OUTPUT(g1293)
--	OUTPUT(g4099)
--	OUTPUT(g4102)
--	OUTPUT(g4109)
--	OUTPUT(g4100)
--	OUTPUT(g4112)
--	OUTPUT(g4105)
--	OUTPUT(g4101)
--	OUTPUT(g4110)
--	OUTPUT(g4104)
--	OUTPUT(g4107)
--	OUTPUT(g4098)
--	
--	g678 = DFF(g4130)
--	g332 = DFF(g6823)
--	g123 = DFF(g6940)
--	g207 = DFF(g6102)
--	g695 = DFF(g4147)
--	g461 = DFF(g4841)
--	g18 = DFF(g6725)
--	g292 = DFF(g3232)
--	g331 = DFF(g4119)
--	g689 = DFF(g4141)
--	g24 = DFF(g6726)
--	g465 = DFF(g6507)
--	g84 = DFF(g6590)
--	g291 = DFF(g3231)
--	g676 = DFF(g5330)
--	g622 = DFF(g5147)
--	g117 = DFF(g4839)
--	g278 = DFF(g6105)
--	g128 = DFF(g5138)
--	g598 = DFF(g4122)
--	g554 = DFF(g6827)
--	g496 = DFF(g6745)
--	g179 = DFF(g6405)
--	g48 = DFF(g6729)
--	g590 = DFF(g6595)
--	g551 = DFF(g6826)
--	g682 = DFF(g4134)
--	g11 = DFF(g6599)
--	g606 = DFF(g4857)
--	g188 = DFF(g6406)
--	g646 = DFF(g5148)
--	g327 = DFF(g4117)
--	g361 = DFF(g6582)
--	g289 = DFF(g3229)
--	g398 = DFF(g5700)
--	g684 = DFF(g4136)
--	g619 = DFF(g4858)
--	g208 = DFF(g5876)
--	g248 = DFF(g3239)
--	g390 = DFF(g5698)
--	g625 = DFF(g5328)
--	g681 = DFF(g4133)
--	g437 = DFF(g4847)
--	g276 = DFF(g5877)
--	g3 = DFF(g6597)
--	g323 = DFF(g4120)
--	g224 = DFF(g3235)
--	g685 = DFF(g4137)
--	g43 = DFF(g6407)
--	g157 = DFF(g5470)
--	g282 = DFF(g6841)
--	g697 = DFF(g4149)
--	g206 = DFF(g6101)
--	g449 = DFF(g4844)
--	g118 = DFF(g4113)
--	g528 = DFF(g6504)
--	g284 = DFF(g3224)
--	g426 = DFF(g4855)
--	g634 = DFF(g4424)
--	g669 = DFF(g5582)
--	g520 = DFF(g6502)
--	g281 = DFF(g6107)
--	g175 = DFF(g5472)
--	g15 = DFF(g6602)
--	g631 = DFF(g5581)
--	g69 = DFF(g6587)
--	g693 = DFF(g4145)
--	g337 = DFF(g2585)
--	g457 = DFF(g4842)
--	g486 = DFF(g2586)
--	g471 = DFF(g1291)
--	g328 = DFF(g4118)
--	g285 = DFF(g3225)
--	g418 = DFF(g4853)
--	g402 = DFF(g4849)
--	g297 = DFF(g6512)
--	g212 = DFF(g3233)
--	g410 = DFF(g4851)
--	g430 = DFF(g4856)
--	g33 = DFF(g6854)
--	g662 = DFF(g1831)
--	g453 = DFF(g4843)
--	g269 = DFF(g6510)
--	g574 = DFF(g6591)
--	g441 = DFF(g4846)
--	g664 = DFF(g1288)
--	g349 = DFF(g5478)
--	g211 = DFF(g6840)
--	g586 = DFF(g6594)
--	g571 = DFF(g5580)
--	g29 = DFF(g6853)
--	g326 = DFF(g4840)
--	g698 = DFF(g4150)
--	g654 = DFF(g5490)
--	g293 = DFF(g6511)
--	g690 = DFF(g4142)
--	g445 = DFF(g4845)
--	g374 = DFF(g5694)
--	g6 = DFF(g6722)
--	g687 = DFF(g4139)
--	g357 = DFF(g5480)
--	g386 = DFF(g5697)
--	g504 = DFF(g6498)
--	g665 = DFF(g4126)
--	g166 = DFF(g5471)
--	g541 = DFF(g6505)
--	g74 = DFF(g6588)
--	g338 = DFF(g5475)
--	g696 = DFF(g4148)
--	g516 = DFF(g6501)
--	g536 = DFF(g6506)
--	g683 = DFF(g4135)
--	g353 = DFF(g5479)
--	g545 = DFF(g6824)
--	g254 = DFF(g3240)
--	g341 = DFF(g5476)
--	g290 = DFF(g3230)
--	g2 = DFF(g6721)
--	g287 = DFF(g3227)
--	g336 = DFF(g6925)
--	g345 = DFF(g5477)
--	g628 = DFF(g5489)
--	g679 = DFF(g4131)
--	g28 = DFF(g6727)
--	g688 = DFF(g4140)
--	g283 = DFF(g6842)
--	g613 = DFF(g4423)
--	g10 = DFF(g6723)
--	g14 = DFF(g6724)
--	g680 = DFF(g4132)
--	g143 = DFF(g6401)
--	g672 = DFF(g5491)
--	g667 = DFF(g4127)
--	g366 = DFF(g6278)
--	g279 = DFF(g6106)
--	g492 = DFF(g6744)
--	g170 = DFF(g6404)
--	g686 = DFF(g4138)
--	g288 = DFF(g3228)
--	g638 = DFF(g1289)
--	g602 = DFF(g4123)
--	g642 = DFF(g4658)
--	g280 = DFF(g5878)
--	g663 = DFF(g4125)
--	g610 = DFF(g4124)
--	g148 = DFF(g5874)
--	g209 = DFF(g6103)
--	g675 = DFF(g1294)
--	g478 = DFF(g1292)
--	g122 = DFF(g4115)
--	g54 = DFF(g6584)
--	g594 = DFF(g6596)
--	g286 = DFF(g3226)
--	g489 = DFF(g2587)
--	g616 = DFF(g4657)
--	g79 = DFF(g6589)
--	g218 = DFF(g3234)
--	g242 = DFF(g3238)
--	g578 = DFF(g6592)
--	g184 = DFF(g5473)
--	g119 = DFF(g4114)
--	g668 = DFF(g6800)
--	g139 = DFF(g5141)
--	g422 = DFF(g4854)
--	g210 = DFF(g6839)
--	g394 = DFF(g5699)
--	g230 = DFF(g3236)
--	g25 = DFF(g6601)
--	g204 = DFF(g5875)
--	g658 = DFF(g4425)
--	g650 = DFF(g5329)
--	g378 = DFF(g5695)
--	g508 = DFF(g6499)
--	g548 = DFF(g6825)
--	g370 = DFF(g5693)
--	g406 = DFF(g4850)
--	g236 = DFF(g3237)
--	g500 = DFF(g6497)
--	g205 = DFF(g6100)
--	g197 = DFF(g6509)
--	g666 = DFF(g4128)
--	g114 = DFF(g4116)
--	g524 = DFF(g6503)
--	g260 = DFF(g3241)
--	g111 = DFF(g6277)
--	g131 = DFF(g5139)
--	g7 = DFF(g6598)
--	g19 = DFF(g6600)
--	g677 = DFF(g4129)
--	g582 = DFF(g6593)
--	g485 = DFF(g6801)
--	g699 = DFF(g4426)
--	g193 = DFF(g5474)
--	g135 = DFF(g5140)
--	g382 = DFF(g5696)
--	g414 = DFF(g4852)
--	g434 = DFF(g4848)
--	g266 = DFF(g4659)
--	g49 = DFF(g6583)
--	g152 = DFF(g6402)
--	g692 = DFF(g4144)
--	g277 = DFF(g6104)
--	g127 = DFF(g6941)
--	g161 = DFF(g6403)
--	g512 = DFF(g6500)
--	g532 = DFF(g6508)
--	g64 = DFF(g6586)
--	g694 = DFF(g4146)
--	g691 = DFF(g4143)
--	g1 = DFF(g6720)
--	g59 = DFF(g6585)
--	
--	I8854 = NOT(g6696)
--	g1289 = NOT(I2272)
--	I9125 = NOT(g6855)
--	I6783 = NOT(g4822)
--	I4424 = NOT(g2097)
--	g6895 = NOT(I9152)
--	g1835 = NOT(I2919)
--	I3040 = NOT(g1770)
--	g6837 = NOT(g6822)
--	I7466 = NOT(g5624)
--	I4809 = NOT(g2974)
--	g3537 = NOT(I4757)
--	g5457 = NOT(g5304)
--	g6062 = NOT(g5824)
--	g4040 = NOT(I5343)
--	I6001 = NOT(g4162)
--	g5549 = NOT(g5331)
--	I4477 = NOT(g3063)
--	g3612 = NOT(I4809)
--	I7055 = NOT(g5318)
--	g2892 = NOT(g1982)
--	I5264 = NOT(g3638)
--	I2225 = NOT(g696)
--	g4123 = NOT(I5451)
--	g4323 = NOT(g4086)
--	g908 = NOT(I1932)
--	I5933 = NOT(g4346)
--	I8252 = NOT(g6294)
--	I2473 = NOT(g971)
--	I7333 = NOT(g5386)
--	I8812 = NOT(g6688)
--	g1674 = NOT(g985)
--	I3528 = NOT(g1422)
--	I8958 = NOT(g6774)
--	I5050 = NOT(g3246)
--	g3234 = NOT(I4501)
--	I2324 = NOT(g1209)
--	g2945 = NOT(I4133)
--	g5121 = NOT(I6775)
--	g1997 = NOT(g1398)
--	g3128 = NOT(I4375)
--	I8005 = NOT(g6110)
--	g1541 = NOT(g1094)
--	g5670 = NOT(g5527)
--	g2738 = NOT(g2327)
--	g6842 = NOT(I9047)
--	g4528 = NOT(I6096)
--	g2244 = NOT(I3379)
--	g6192 = NOT(g5946)
--	g2709 = NOT(I3864)
--	g1332 = NOT(I2349)
--	g4530 = NOT(I6102)
--	g1680 = NOT(g1011)
--	g2078 = NOT(g1345)
--	g1209 = NOT(I2215)
--	I3010 = NOT(g1504)
--	g5813 = NOT(I7612)
--	I7509 = NOT(g5587)
--	I5379 = NOT(g3940)
--	g3800 = NOT(g3388)
--	g2907 = NOT(g1914)
--	g6854 = NOT(I9085)
--	g2035 = NOT(I3144)
--	g2959 = NOT(g1861)
--	g6941 = NOT(I9236)
--	g4010 = NOT(g3601)
--	I2287 = NOT(g927)
--	I4273 = NOT(g2197)
--	I8270 = NOT(g6300)
--	g5740 = NOT(I7501)
--	I5777 = NOT(g3807)
--	g2876 = NOT(g1943)
--	g873 = NOT(g306)
--	g4839 = NOT(I6525)
--	I5882 = NOT(g3871)
--	g2656 = NOT(I3800)
--	I8473 = NOT(g6485)
--	I2199 = NOT(g33)
--	g900 = NOT(I1927)
--	g6708 = NOT(I8834)
--	I2399 = NOT(g729)
--	I3278 = NOT(g1695)
--	g6520 = NOT(I8476)
--	g940 = NOT(g64)
--	I6677 = NOT(g4757)
--	g3902 = NOT(g3575)
--	g5687 = NOT(g5567)
--	g2915 = NOT(g1931)
--	g847 = NOT(g590)
--	I3235 = NOT(g1807)
--	I3343 = NOT(g1623)
--	g6431 = NOT(I8295)
--	g709 = NOT(g114)
--	g6812 = NOT(I8984)
--	I6576 = NOT(g4700)
--	g749 = NOT(I1847)
--	g3090 = NOT(I4331)
--	I9107 = NOT(g6855)
--	g2214 = NOT(I3349)
--	g4618 = NOT(g4246)
--	g6376 = NOT(g6267)
--	g4143 = NOT(I5511)
--	I6349 = NOT(g4569)
--	g4343 = NOT(g4011)
--	I5674 = NOT(g4003)
--	I8177 = NOT(g6173)
--	g2110 = NOT(g1381)
--	I3134 = NOT(g1336)
--	g6405 = NOT(I8229)
--	I3334 = NOT(g1330)
--	I7197 = NOT(g5431)
--	g4566 = NOT(g4198)
--	I7397 = NOT(g5561)
--	I4534 = NOT(g2858)
--	g1714 = NOT(g1110)
--	I4961 = NOT(g3597)
--	g2663 = NOT(g2308)
--	g3456 = NOT(g2640)
--	g5141 = NOT(I6801)
--	g922 = NOT(I1947)
--	g4693 = NOT(I6283)
--	g4134 = NOT(I5484)
--	g5570 = NOT(g5392)
--	g5860 = NOT(g5634)
--	g4334 = NOT(g3733)
--	I3804 = NOT(g2575)
--	I2207 = NOT(g7)
--	I5153 = NOT(g3330)
--	g3355 = NOT(g3100)
--	g5645 = NOT(g5537)
--	g6733 = NOT(I8891)
--	g5691 = NOT(g5568)
--	g4804 = NOT(g4473)
--	I9047 = NOT(g6838)
--	I4414 = NOT(g2090)
--	g6610 = NOT(I8696)
--	g2877 = NOT(g2434)
--	I4903 = NOT(g3223)
--	g6796 = NOT(I8958)
--	g3063 = NOT(I4288)
--	I3313 = NOT(g1337)
--	g5879 = NOT(g5770)
--	g3463 = NOT(g2682)
--	I4513 = NOT(g2765)
--	g1623 = NOT(I2578)
--	g5358 = NOT(I7012)
--	I3202 = NOT(g1812)
--	I2215 = NOT(g695)
--	g4113 = NOT(I5421)
--	g1076 = NOT(I2115)
--	g6069 = NOT(g5791)
--	I7817 = NOT(g5924)
--	g6540 = NOT(g6474)
--	I6352 = NOT(g4564)
--	I1865 = NOT(g279)
--	g4202 = NOT(I5622)
--	I6867 = NOT(g5082)
--	I5511 = NOT(g3876)
--	g5587 = NOT(I7349)
--	I8144 = NOT(g6182)
--	g1175 = NOT(g42)
--	g1375 = NOT(I2411)
--	g3118 = NOT(I4366)
--	g3318 = NOT(I4593)
--	g2464 = NOT(I3596)
--	g3872 = NOT(g3312)
--	g4494 = NOT(I6004)
--	I2870 = NOT(g1161)
--	g4518 = NOT(I6066)
--	I4288 = NOT(g2215)
--	g5615 = NOT(I7372)
--	g4567 = NOT(I6139)
--	I4382 = NOT(g2265)
--	I3776 = NOT(g2044)
--	g3057 = NOT(I4282)
--	I5600 = NOT(g3821)
--	I3593 = NOT(g1295)
--	I2825 = NOT(g1143)
--	g1285 = NOT(g852)
--	g3457 = NOT(g2653)
--	g5174 = NOT(g5099)
--	I6386 = NOT(g4462)
--	I3965 = NOT(g2268)
--	I8488 = NOT(g6426)
--	g6849 = NOT(I9074)
--	I6599 = NOT(g4823)
--	I2408 = NOT(g719)
--	g3834 = NOT(I5027)
--	g2295 = NOT(g1578)
--	g1384 = NOT(I2420)
--	g1339 = NOT(I2370)
--	g5545 = NOT(g5331)
--	I6170 = NOT(g4343)
--	I9128 = NOT(g6864)
--	g6898 = NOT(I9161)
--	g1838 = NOT(g1595)
--	g6900 = NOT(I9167)
--	g2194 = NOT(I3331)
--	g6797 = NOT(I8961)
--	g2394 = NOT(I3537)
--	I3050 = NOT(g1439)
--	I3641 = NOT(g1491)
--	I2943 = NOT(g1715)
--	I5736 = NOT(g4022)
--	g6510 = NOT(I8450)
--	I6280 = NOT(g4430)
--	g4933 = NOT(I6625)
--	g5420 = NOT(I7086)
--	g4521 = NOT(I6075)
--	g1672 = NOT(g1094)
--	I7058 = NOT(g5281)
--	I2887 = NOT(g1123)
--	I2122 = NOT(g689)
--	g1477 = NOT(g952)
--	g3232 = NOT(I4495)
--	I2228 = NOT(g15)
--	g5794 = NOT(I7593)
--	g1643 = NOT(I2608)
--	I4495 = NOT(g3022)
--	I4437 = NOT(g2108)
--	g2705 = NOT(I3858)
--	g3813 = NOT(g3258)
--	I8650 = NOT(g6529)
--	I3379 = NOT(g1647)
--	g2242 = NOT(I3373)
--	g1205 = NOT(g45)
--	I2033 = NOT(g678)
--	I5871 = NOT(g3744)
--	g774 = NOT(I1859)
--	g6819 = NOT(I8994)
--	g6694 = NOT(I8800)
--	g4379 = NOT(I5848)
--	g5905 = NOT(g5852)
--	g3519 = NOT(g2740)
--	I7856 = NOT(g5994)
--	g921 = NOT(g111)
--	g1551 = NOT(g1011)
--	g1742 = NOT(I2756)
--	I4752 = NOT(g2859)
--	g6488 = NOT(g6367)
--	g2254 = NOT(I3391)
--	I8594 = NOT(g6446)
--	g2814 = NOT(I4023)
--	g4289 = NOT(I5746)
--	g4658 = NOT(I6247)
--	I6756 = NOT(g4775)
--	g6701 = NOT(I8821)
--	I8972 = NOT(g6795)
--	I3271 = NOT(g1748)
--	I2845 = NOT(g1193)
--	g5300 = NOT(I6952)
--	g2350 = NOT(I3502)
--	I8806 = NOT(g6686)
--	I3611 = NOT(g1771)
--	I2137 = NOT(g1)
--	I8943 = NOT(g6774)
--	I2337 = NOT(g1209)
--	I2913 = NOT(g1792)
--	g1754 = NOT(I2773)
--	g6886 = NOT(I9125)
--	g2409 = NOT(g1815)
--	g894 = NOT(I1917)
--	g1273 = NOT(g839)
--	I5424 = NOT(g3725)
--	I6403 = NOT(g4492)
--	g6314 = NOT(I8044)
--	g4799 = NOT(g4485)
--	I9155 = NOT(g6882)
--	g2836 = NOT(g2509)
--	g2212 = NOT(I3343)
--	I6763 = NOT(g4780)
--	g3860 = NOT(I5081)
--	g2967 = NOT(I4166)
--	g6825 = NOT(I9008)
--	g5440 = NOT(g5266)
--	g3710 = NOT(g3029)
--	I5523 = NOT(g3840)
--	g843 = NOT(g574)
--	g1543 = NOT(g1006)
--	g4132 = NOT(I5478)
--	g6408 = NOT(g6283)
--	g4153 = NOT(I5545)
--	I6359 = NOT(g4566)
--	g6136 = NOT(I7856)
--	g2822 = NOT(I4031)
--	I8891 = NOT(g6706)
--	I8913 = NOT(g6743)
--	I2692 = NOT(g1037)
--	g6594 = NOT(I8650)
--	g946 = NOT(g361)
--	g1729 = NOT(I2731)
--	I5551 = NOT(g4059)
--	g4802 = NOT(I6470)
--	g3962 = NOT(I5214)
--	I2154 = NOT(g14)
--	I4189 = NOT(g2159)
--	I5499 = NOT(g3847)
--	g5151 = NOT(I6819)
--	g3158 = NOT(I4398)
--	g6806 = NOT(I8978)
--	I4706 = NOT(g2877)
--	g5875 = NOT(I7637)
--	g5530 = NOT(I7270)
--	I9167 = NOT(g6878)
--	I5926 = NOT(g4153)
--	g2921 = NOT(g1950)
--	g6065 = NOT(g5784)
--	I6315 = NOT(g4446)
--	I4371 = NOT(g2555)
--	g6887 = NOT(I9128)
--	I4429 = NOT(g2102)
--	g6122 = NOT(I7838)
--	g6465 = NOT(I8329)
--	g6322 = NOT(I8056)
--	g1660 = NOT(g985)
--	g1946 = NOT(I3053)
--	g6230 = NOT(g6040)
--	g5010 = NOT(I6646)
--	g4511 = NOT(I6045)
--	I6874 = NOT(g4861)
--	g2895 = NOT(g1894)
--	g6033 = NOT(g5824)
--	g2837 = NOT(g2512)
--	I2979 = NOT(g1263)
--	I3864 = NOT(g2044)
--	g5884 = NOT(g5864)
--	I8342 = NOT(g6314)
--	I2218 = NOT(g11)
--	g1513 = NOT(g878)
--	I2312 = NOT(g897)
--	I3714 = NOT(g1852)
--	I4297 = NOT(g2555)
--	I8255 = NOT(g6292)
--	I8815 = NOT(g6689)
--	g4492 = NOT(I5998)
--	I1868 = NOT(g280)
--	I7608 = NOT(g5605)
--	I5862 = NOT(g3863)
--	g1679 = NOT(g985)
--	g1378 = NOT(I2414)
--	g4714 = NOT(I6324)
--	I2293 = NOT(g971)
--	g5278 = NOT(I6937)
--	g3284 = NOT(g3019)
--	I4684 = NOT(g2687)
--	I8497 = NOT(g6481)
--	g3239 = NOT(I4516)
--	I6537 = NOT(g4711)
--	g3545 = NOT(g3085)
--	g2788 = NOT(I3983)
--	g6137 = NOT(I7859)
--	g5667 = NOT(g5524)
--	g6891 = NOT(I9140)
--	g1831 = NOT(I2907)
--	g1335 = NOT(I2358)
--	g3380 = NOT(g2831)
--	I4791 = NOT(g2814)
--	g6337 = NOT(I8089)
--	I4309 = NOT(g2525)
--	I2828 = NOT(g1193)
--	g3832 = NOT(I5023)
--	g1288 = NOT(I2269)
--	g5566 = NOT(I7318)
--	g3853 = NOT(I5068)
--	I3736 = NOT(g2460)
--	I6612 = NOT(g4660)
--	I7161 = NOT(g5465)
--	I7361 = NOT(g5566)
--	g2842 = NOT(I4050)
--	g1805 = NOT(I2854)
--	I6417 = NOT(g4617)
--	I3623 = NOT(g1491)
--	g4262 = NOT(I5713)
--	I7051 = NOT(g5219)
--	I2221 = NOT(g43)
--	g3559 = NOT(g2603)
--	g4736 = NOT(I6366)
--	g2485 = NOT(I3614)
--	I7451 = NOT(g5597)
--	I2703 = NOT(g1189)
--	I8267 = NOT(g6297)
--	g4623 = NOT(g4262)
--	g1947 = NOT(I3056)
--	I5885 = NOT(g3746)
--	I7999 = NOT(g6137)
--	g878 = NOT(g639)
--	I7146 = NOT(g5231)
--	I6330 = NOT(g4560)
--	I7346 = NOT(g5531)
--	I3871 = NOT(g2145)
--	I8329 = NOT(g6305)
--	g4375 = NOT(I5840)
--	g4871 = NOT(I6599)
--	I8761 = NOT(g6563)
--	g3204 = NOT(I4441)
--	g4722 = NOT(I6346)
--	g710 = NOT(g128)
--	I4498 = NOT(g2686)
--	g829 = NOT(g323)
--	g5113 = NOT(I6753)
--	g1632 = NOT(g760)
--	g1037 = NOT(I2067)
--	g3100 = NOT(I4347)
--	I8828 = NOT(g6661)
--	g6726 = NOT(I8872)
--	g6497 = NOT(I8411)
--	g1653 = NOT(I2630)
--	g2640 = NOT(I3782)
--	I8727 = NOT(g6536)
--	g2031 = NOT(I3140)
--	I5436 = NOT(g3729)
--	g2252 = NOT(I3385)
--	g5908 = NOT(g5753)
--	g2958 = NOT(g1861)
--	I7472 = NOT(g5626)
--	g2176 = NOT(I3319)
--	I2716 = NOT(g1115)
--	I5831 = NOT(g3842)
--	I2349 = NOT(g1160)
--	g4139 = NOT(I5499)
--	I5182 = NOT(g3271)
--	g5518 = NOT(I7258)
--	g5567 = NOT(g5418)
--	I5382 = NOT(g3952)
--	g2405 = NOT(I3543)
--	I2848 = NOT(g1193)
--	g1917 = NOT(I3016)
--	g2829 = NOT(g2491)
--	g2765 = NOT(I3946)
--	I7116 = NOT(g5299)
--	I4019 = NOT(g1841)
--	g4424 = NOT(I5923)
--	I6090 = NOT(g4393)
--	I4362 = NOT(g2555)
--	I3672 = NOT(g1656)
--	g3040 = NOT(I4255)
--	I3077 = NOT(g1439)
--	g4809 = NOT(I6485)
--	g5593 = NOT(I7355)
--	g3440 = NOT(I4678)
--	g3969 = NOT(I5233)
--	g6312 = NOT(I8040)
--	I6366 = NOT(g4569)
--	I4452 = NOT(g2117)
--	g2974 = NOT(I4173)
--	g6401 = NOT(I8217)
--	g895 = NOT(g139)
--	I6456 = NOT(g4633)
--	g4523 = NOT(I6081)
--	g1233 = NOT(I2231)
--	I6649 = NOT(g4693)
--	g4643 = NOT(g4293)
--	g5264 = NOT(g4943)
--	I9158 = NOT(g6887)
--	g1054 = NOT(g485)
--	g5160 = NOT(g5099)
--	g2796 = NOT(I3999)
--	I6355 = NOT(g4569)
--	g2473 = NOT(I3605)
--	I3099 = NOT(g1519)
--	I8576 = NOT(g6436)
--	g1770 = NOT(I2805)
--	I8866 = NOT(g6701)
--	I3304 = NOT(g1740)
--	I4486 = NOT(g3093)
--	g5521 = NOT(I7261)
--	I3499 = NOT(g1450)
--	I8716 = NOT(g6518)
--	g1725 = NOT(g1113)
--	I7596 = NOT(g5605)
--	g6727 = NOT(I8875)
--	g3875 = NOT(I5106)
--	g2324 = NOT(I3478)
--	I4504 = NOT(g2726)
--	I2119 = NOT(g688)
--	g5450 = NOT(g5292)
--	I5037 = NOT(g3705)
--	g5996 = NOT(g5824)
--	g4104 = NOT(I5394)
--	g6592 = NOT(I8644)
--	g4099 = NOT(I5379)
--	g4499 = NOT(I6015)
--	I2352 = NOT(g1161)
--	I6063 = NOT(g4381)
--	g6746 = NOT(I8916)
--	I2867 = NOT(g1143)
--	I8699 = NOT(g6573)
--	g2177 = NOT(I3322)
--	g5179 = NOT(g5099)
--	g5379 = NOT(I7035)
--	I2893 = NOT(g1236)
--	g5878 = NOT(I7646)
--	I3044 = NOT(g1257)
--	g1189 = NOT(I2196)
--	g3839 = NOT(I5040)
--	g6932 = NOT(I9217)
--	g4273 = NOT(I5728)
--	g5658 = NOT(g5512)
--	g6624 = NOT(I8730)
--	I6118 = NOT(g4406)
--	I6318 = NOT(g4447)
--	I3983 = NOT(g2276)
--	g2849 = NOT(g2577)
--	I3572 = NOT(g1295)
--	g1787 = NOT(I2835)
--	I5442 = NOT(g3731)
--	I4678 = NOT(g2670)
--	I6057 = NOT(g4379)
--	I8524 = NOT(g6496)
--	I4331 = NOT(g2555)
--	I8644 = NOT(g6526)
--	I3543 = NOT(g1461)
--	I6989 = NOT(g5307)
--	I2614 = NOT(g1123)
--	g1675 = NOT(g1101)
--	I2370 = NOT(g1123)
--	I2125 = NOT(g698)
--	g3235 = NOT(I4504)
--	g3343 = NOT(g3090)
--	I5233 = NOT(g3571)
--	I2821 = NOT(g1221)
--	g4712 = NOT(I6318)
--	g985 = NOT(g638)
--	g6576 = NOT(g6487)
--	I6549 = NOT(g4699)
--	I8258 = NOT(g6293)
--	I8818 = NOT(g6690)
--	I3534 = NOT(g1295)
--	g2245 = NOT(I3382)
--	I3729 = NOT(g2436)
--	I3961 = NOT(g1835)
--	I5454 = NOT(g3874)
--	g2291 = NOT(I3434)
--	g5997 = NOT(g5854)
--	g4534 = NOT(I6114)
--	I3927 = NOT(g2245)
--	I5532 = NOT(g3861)
--	g1684 = NOT(I2668)
--	g6699 = NOT(I8815)
--	g1639 = NOT(g815)
--	g1338 = NOT(I2367)
--	g1963 = NOT(I3074)
--	I8186 = NOT(g6179)
--	I6321 = NOT(g4559)
--	I4226 = NOT(g2525)
--	g1109 = NOT(I2137)
--	g1791 = NOT(I2845)
--	I8975 = NOT(g6791)
--	I3946 = NOT(g2256)
--	g889 = NOT(g310)
--	I2306 = NOT(g896)
--	g3792 = NOT(g3388)
--	I6625 = NOT(g4745)
--	g2819 = NOT(g2467)
--	g4014 = NOT(I5316)
--	I8426 = NOT(g6424)
--	I5412 = NOT(g4034)
--	g4660 = NOT(I6253)
--	I6253 = NOT(g4608)
--	g2088 = NOT(I3202)
--	g2923 = NOT(g1969)
--	I4173 = NOT(g2408)
--	I8614 = NOT(g6537)
--	I3513 = NOT(g1450)
--	g2488 = NOT(I3617)
--	g1759 = NOT(I2782)
--	I2756 = NOT(g1175)
--	g2701 = NOT(I3855)
--	I7190 = NOT(g5432)
--	I8821 = NOT(g6691)
--	g6524 = NOT(I8488)
--	I6740 = NOT(g4781)
--	g4513 = NOT(I6051)
--	I8984 = NOT(g6794)
--	I7501 = NOT(g5596)
--	g1957 = NOT(I3068)
--	g2215 = NOT(I3352)
--	g6119 = NOT(I7829)
--	I2904 = NOT(g1256)
--	g6319 = NOT(I8051)
--	g1049 = NOT(g266)
--	g5901 = NOT(g5753)
--	g2886 = NOT(g1966)
--	I6552 = NOT(g4702)
--	I4059 = NOT(g1878)
--	g4036 = NOT(I5337)
--	g3094 = NOT(I4337)
--	I4459 = NOT(g2134)
--	I8544 = NOT(g6453)
--	g4679 = NOT(I6269)
--	g6352 = NOT(I8110)
--	g6818 = NOT(I8991)
--	g6577 = NOT(g6488)
--	I1847 = NOT(g209)
--	I3288 = NOT(g1710)
--	g3567 = NOT(g3074)
--	I3382 = NOT(g1284)
--	g1715 = NOT(I2716)
--	g4135 = NOT(I5487)
--	I7704 = NOT(g5723)
--	g848 = NOT(g594)
--	g5092 = NOT(g4753)
--	g1498 = NOT(I2479)
--	I2763 = NOT(g1236)
--	g2870 = NOT(g2296)
--	I3022 = NOT(g1426)
--	I4261 = NOT(g1857)
--	I2391 = NOT(g774)
--	g4382 = NOT(I5857)
--	g3776 = NOT(g3466)
--	g6893 = NOT(I9146)
--	g1833 = NOT(I2913)
--	I3422 = NOT(g1641)
--	g5574 = NOT(g5407)
--	I3749 = NOT(g2484)
--	g3593 = NOT(g2997)
--	g6211 = NOT(g5992)
--	g2650 = NOT(I3794)
--	g5714 = NOT(I7475)
--	g932 = NOT(g337)
--	I8061 = NOT(g6113)
--	g4805 = NOT(g4473)
--	g4022 = NOT(I5328)
--	g1584 = NOT(g743)
--	g4422 = NOT(g4111)
--	g6599 = NOT(I8665)
--	g1539 = NOT(g878)
--	I5109 = NOT(g3710)
--	g2408 = NOT(I3546)
--	I2159 = NOT(g465)
--	I6570 = NOT(g4719)
--	g2136 = NOT(g1395)
--	I4664 = NOT(g2924)
--	I8027 = NOT(g6237)
--	I4246 = NOT(g2194)
--	g2336 = NOT(I3488)
--	g5580 = NOT(I7336)
--	g716 = NOT(I1832)
--	I3560 = NOT(g1673)
--	g736 = NOT(I1841)
--	I6525 = NOT(g4770)
--	g2768 = NOT(g2367)
--	g6370 = NOT(I8174)
--	g2594 = NOT(I3723)
--	g4798 = NOT(I6464)
--	g6325 = NOT(I8061)
--	g6821 = NOT(g6785)
--	g4560 = NOT(g4188)
--	g2806 = NOT(g2446)
--	I3632 = NOT(g1295)
--	g3450 = NOT(I4688)
--	I3037 = NOT(g1769)
--	g6939 = NOT(I9230)
--	g1052 = NOT(g668)
--	I3653 = NOT(g1305)
--	I3102 = NOT(g1426)
--	I2115 = NOT(g687)
--	I2315 = NOT(g1222)
--	I2811 = NOT(g1209)
--	g6083 = NOT(g5809)
--	g2887 = NOT(g1858)
--	I2047 = NOT(g682)
--	g6544 = NOT(I8544)
--	I6607 = NOT(g4745)
--	g4632 = NOT(g4281)
--	g5889 = NOT(g5742)
--	g5476 = NOT(I7164)
--	g2934 = NOT(g2004)
--	g2230 = NOT(I3355)
--	g4437 = NOT(I5948)
--	g4102 = NOT(I5388)
--	g4302 = NOT(g4068)
--	I5865 = NOT(g3743)
--	g6106 = NOT(I7814)
--	g4579 = NOT(g4206)
--	g4869 = NOT(g4662)
--	g6306 = NOT(I8030)
--	I3752 = NOT(g2044)
--	g5375 = NOT(I7029)
--	I8107 = NOT(g6136)
--	g4719 = NOT(I6337)
--	g1730 = NOT(g1114)
--	g3289 = NOT(g3034)
--	g1504 = NOT(I2485)
--	g3777 = NOT(g3388)
--	I6587 = NOT(g4803)
--	I8159 = NOT(g6167)
--	I6111 = NOT(g4404)
--	g3835 = NOT(I5030)
--	I6311 = NOT(g4444)
--	I8223 = NOT(g6325)
--	g2096 = NOT(I3212)
--	I9143 = NOT(g6886)
--	g3882 = NOT(I5119)
--	g1070 = NOT(g94)
--	g2550 = NOT(I3665)
--	I6615 = NOT(g4745)
--	g3271 = NOT(g3042)
--	I4671 = NOT(g2928)
--	I2880 = NOT(g1143)
--	g2845 = NOT(g2565)
--	g1897 = NOT(I2992)
--	g6622 = NOT(I8724)
--	I2537 = NOT(g971)
--	I5896 = NOT(g3879)
--	g2195 = NOT(I3334)
--	g4265 = NOT(I5716)
--	g2891 = NOT(g1884)
--	g2913 = NOT(g1925)
--	g5139 = NOT(I6795)
--	I3364 = NOT(g1648)
--	g5384 = NOT(g5220)
--	I9134 = NOT(g6864)
--	I2272 = NOT(g908)
--	g6904 = NOT(I9179)
--	g4786 = NOT(I6448)
--	g3799 = NOT(g3388)
--	g6514 = NOT(I8462)
--	g4364 = NOT(I5825)
--	I8447 = NOT(g6410)
--	I3770 = NOT(g2145)
--	I5019 = NOT(g3318)
--	I2417 = NOT(g774)
--	g6403 = NOT(I8223)
--	g5809 = NOT(I7608)
--	I7683 = NOT(g5702)
--	g6841 = NOT(I9044)
--	g3541 = NOT(g2643)
--	I2982 = NOT(g1426)
--	g1678 = NOT(I2658)
--	g4770 = NOT(I6414)
--	g1006 = NOT(I2047)
--	I2234 = NOT(g697)
--	g1331 = NOT(I2346)
--	g4296 = NOT(I5753)
--	I2128 = NOT(g18)
--	g3238 = NOT(I4513)
--	I3553 = NOT(g1305)
--	I6020 = NOT(g4176)
--	g3332 = NOT(g3079)
--	g5477 = NOT(I7167)
--	I6420 = NOT(g4618)
--	g6695 = NOT(I8803)
--	I2330 = NOT(g1122)
--	g3209 = NOT(I4452)
--	I6507 = NOT(g4644)
--	g4532 = NOT(I6108)
--	g1682 = NOT(g829)
--	g6107 = NOT(I7817)
--	I9113 = NOT(g6855)
--	I1856 = NOT(g204)
--	g1305 = NOT(I2293)
--	g6536 = NOT(I8524)
--	g3802 = NOT(g3388)
--	I5728 = NOT(g4022)
--	g2481 = NOT(I3608)
--	I7475 = NOT(g5627)
--	g931 = NOT(g54)
--	g1748 = NOT(I2763)
--	g2692 = NOT(I3840)
--	I4217 = NOT(g2163)
--	g2097 = NOT(I3215)
--	I4066 = NOT(g2582)
--	g5551 = NOT(I7295)
--	g5742 = NOT(g5686)
--	g2726 = NOT(I3886)
--	g5099 = NOT(I6737)
--	g2497 = NOT(I3626)
--	I5385 = NOT(g3962)
--	g5304 = NOT(I6956)
--	g2154 = NOT(I3271)
--	g1755 = NOT(I2776)
--	g4189 = NOT(I5597)
--	I8978 = NOT(g6792)
--	g4706 = NOT(I6308)
--	g6416 = NOT(I8258)
--	I8243 = NOT(g6286)
--	I8417 = NOT(g6420)
--	g3901 = NOT(g3575)
--	I6630 = NOT(g4745)
--	I7646 = NOT(g5774)
--	I3675 = NOT(g1491)
--	g6522 = NOT(I8482)
--	g6115 = NOT(g5879)
--	g1045 = NOT(g699)
--	I3281 = NOT(g1761)
--	I7039 = NOT(g5309)
--	I7484 = NOT(g5630)
--	g1173 = NOT(I2185)
--	I4455 = NOT(g2118)
--	I8629 = NOT(g6544)
--	g5273 = NOT(I6930)
--	I4133 = NOT(g2040)
--	g1491 = NOT(I2476)
--	g760 = NOT(I1853)
--	g2783 = NOT(I3979)
--	g4281 = NOT(I5736)
--	g3600 = NOT(I4791)
--	g2112 = NOT(I3240)
--	g1283 = NOT(g853)
--	g2312 = NOT(I3462)
--	g1369 = NOT(I2405)
--	I6750 = NOT(g4771)
--	g6654 = NOT(I8758)
--	g3714 = NOT(g3041)
--	I7583 = NOT(g5605)
--	I3684 = NOT(g1733)
--	I5006 = NOT(g3604)
--	I8800 = NOT(g6684)
--	g1059 = NOT(g702)
--	g1578 = NOT(I2552)
--	g2001 = NOT(I3112)
--	I5406 = NOT(g3976)
--	g5572 = NOT(g5399)
--	I3109 = NOT(g1504)
--	I3791 = NOT(g2044)
--	g2293 = NOT(g1567)
--	g6880 = NOT(I9107)
--	g6595 = NOT(I8653)
--	g4138 = NOT(I5496)
--	g1535 = NOT(g1088)
--	g4639 = NOT(g4289)
--	g6537 = NOT(I8527)
--	g5543 = NOT(g5331)
--	I3808 = NOT(g2125)
--	I7276 = NOT(g5375)
--	I5487 = NOT(g3881)
--	I2355 = NOT(g1177)
--	g4109 = NOT(I5409)
--	g4309 = NOT(g4074)
--	g2828 = NOT(g2488)
--	g2830 = NOT(g2494)
--	g2727 = NOT(g2324)
--	g4808 = NOT(g4473)
--	I2964 = NOT(g1257)
--	g821 = NOT(I1880)
--	g6612 = NOT(I8702)
--	g5534 = NOT(I7276)
--	g5729 = NOT(I7494)
--	I6666 = NOT(g4740)
--	I9179 = NOT(g6875)
--	g1415 = NOT(g1246)
--	g4707 = NOT(I6311)
--	g6417 = NOT(I8261)
--	I7404 = NOT(g5541)
--	g3076 = NOT(I4309)
--	I8512 = NOT(g6441)
--	g3889 = NOT(g3575)
--	I6528 = NOT(g4815)
--	g1664 = NOT(I2643)
--	g1246 = NOT(I2237)
--	g6234 = NOT(g6057)
--	I3575 = NOT(g1305)
--	g5885 = NOT(g5865)
--	g6328 = NOT(I8066)
--	g1203 = NOT(I2207)
--	I5445 = NOT(g4040)
--	g5946 = NOT(g5729)
--	g6542 = NOT(I8538)
--	g6330 = NOT(I8070)
--	g1721 = NOT(I2721)
--	I5091 = NOT(g3242)
--	I8056 = NOT(g6109)
--	g2932 = NOT(g1998)
--	I8456 = NOT(g6417)
--	g5903 = NOT(g5753)
--	I3833 = NOT(g2266)
--	I2318 = NOT(g1236)
--	g4715 = NOT(I6327)
--	I2367 = NOT(g1161)
--	I1924 = NOT(g663)
--	g6800 = NOT(I8966)
--	I5169 = NOT(g3593)
--	I6410 = NOT(g4473)
--	g4098 = NOT(I5376)
--	g3500 = NOT(g2647)
--	g4498 = NOT(I6012)
--	I2057 = NOT(g685)
--	g1502 = NOT(g709)
--	I5059 = NOT(g3259)
--	I5920 = NOT(g4228)
--	I2457 = NOT(g1253)
--	I3584 = NOT(g1678)
--	I5868 = NOT(g3864)
--	I2989 = NOT(g1519)
--	I2193 = NOT(g693)
--	g5436 = NOT(I7116)
--	g3384 = NOT(g2834)
--	g1940 = NOT(I3047)
--	g2576 = NOT(I3687)
--	g2866 = NOT(g1905)
--	g5135 = NOT(I6783)
--	g2716 = NOT(I3871)
--	g3838 = NOT(I5037)
--	I7906 = NOT(g5912)
--	I3268 = NOT(g1656)
--	I3019 = NOT(g1755)
--	g3424 = NOT(I4671)
--	g5382 = NOT(I7042)
--	I5793 = NOT(g3803)
--	I3419 = NOT(g1287)
--	g6902 = NOT(I9173)
--	I6143 = NOT(g4237)
--	I6343 = NOT(g4458)
--	g846 = NOT(g586)
--	g1671 = NOT(g985)
--	g5805 = NOT(I7604)
--	I5415 = NOT(g3723)
--	g6512 = NOT(I8456)
--	I3452 = NOT(g1450)
--	g4162 = NOT(I5562)
--	g5022 = NOT(I6666)
--	g1030 = NOT(I2057)
--	I8279 = NOT(g6307)
--	g3231 = NOT(I4492)
--	g6490 = NOT(g6371)
--	I2321 = NOT(g898)
--	g6823 = NOT(I9002)
--	g3477 = NOT(g2692)
--	g6166 = NOT(I7892)
--	g6366 = NOT(I8162)
--	I6334 = NOT(g4454)
--	I8872 = NOT(g6695)
--	g2241 = NOT(I3370)
--	g1564 = NOT(g1030)
--	I7892 = NOT(g5916)
--	I3086 = NOT(g1439)
--	g6529 = NOT(I8503)
--	I8843 = NOT(g6658)
--	g6649 = NOT(I8745)
--	I6555 = NOT(g4703)
--	g1741 = NOT(I2753)
--	I6792 = NOT(g5097)
--	g3104 = NOT(I4351)
--	I3385 = NOT(g1318)
--	g2524 = NOT(I3647)
--	g2644 = NOT(I3788)
--	I8834 = NOT(g6661)
--	g6698 = NOT(I8812)
--	g1638 = NOT(g754)
--	g839 = NOT(g567)
--	I6621 = NOT(g4745)
--	g2119 = NOT(g1391)
--	I5502 = NOT(g3853)
--	g1108 = NOT(I2134)
--	I3025 = NOT(g1439)
--	I2552 = NOT(g971)
--	g5437 = NOT(I7119)
--	g4385 = NOT(I5862)
--	I3425 = NOT(g1274)
--	I9092 = NOT(g6855)
--	I4441 = NOT(g2109)
--	g2818 = NOT(g2464)
--	g2867 = NOT(g1908)
--	g1883 = NOT(g1797)
--	g5579 = NOT(I7333)
--	I7478 = NOT(g5628)
--	g4425 = NOT(I5926)
--	I7035 = NOT(g5150)
--	I5388 = NOT(g3969)
--	I7517 = NOT(g5593)
--	g2893 = NOT(g1985)
--	g5752 = NOT(I7509)
--	I8232 = NOT(g6332)
--	g5917 = NOT(I7683)
--	I6567 = NOT(g4715)
--	g6720 = NOT(I8854)
--	I3678 = NOT(g1690)
--	g2975 = NOT(I4176)
--	I5030 = NOT(g3242)
--	I3331 = NOT(g1631)
--	g1861 = NOT(I2967)
--	g6367 = NOT(I8165)
--	g1048 = NOT(g492)
--	I5430 = NOT(g3727)
--	g2599 = NOT(I3729)
--	g5042 = NOT(I6672)
--	g1711 = NOT(I2712)
--	I3635 = NOT(g1305)
--	g6652 = NOT(I8752)
--	g5442 = NOT(g5270)
--	g1055 = NOT(g269)
--	I2570 = NOT(g1222)
--	I2860 = NOT(g1177)
--	g6057 = NOT(g5824)
--	g4131 = NOT(I5475)
--	I4743 = NOT(g2594)
--	I3105 = NOT(g1439)
--	g2170 = NOT(I3301)
--	g2370 = NOT(I3522)
--	g4406 = NOT(I5913)
--	g6193 = NOT(g5957)
--	g1333 = NOT(I2352)
--	g2125 = NOT(I3255)
--	I8552 = NOT(g6455)
--	g1774 = NOT(I2817)
--	g4766 = NOT(I6406)
--	g4105 = NOT(I5397)
--	g1846 = NOT(I2940)
--	g5054 = NOT(g4816)
--	g4801 = NOT(g4487)
--	g6834 = NOT(g6821)
--	g4487 = NOT(I5991)
--	I7110 = NOT(g5291)
--	g3534 = NOT(I4752)
--	I5910 = NOT(g3750)
--	g5770 = NOT(g5645)
--	I3755 = NOT(g2125)
--	g5296 = NOT(I6946)
--	I8687 = NOT(g6568)
--	I6933 = NOT(g5124)
--	g2544 = NOT(I3662)
--	g6598 = NOT(I8662)
--	I5609 = NOT(g3893)
--	I4474 = NOT(g3052)
--	I2358 = NOT(g1176)
--	g3014 = NOT(I4217)
--	g6121 = NOT(I7835)
--	I7002 = NOT(g5308)
--	g766 = NOT(I1856)
--	g3885 = NOT(I5124)
--	g4226 = NOT(g4050)
--	g2106 = NOT(g1378)
--	g2306 = NOT(g1743)
--	I3373 = NOT(g1320)
--	g2790 = NOT(g2413)
--	g6232 = NOT(g6048)
--	I5217 = NOT(g3673)
--	I8570 = NOT(g6433)
--	I8860 = NOT(g6699)
--	I4480 = NOT(g3073)
--	g1994 = NOT(I3105)
--	g1290 = NOT(I2275)
--	I2275 = NOT(g909)
--	g6938 = NOT(I9227)
--	I5466 = NOT(g3787)
--	g4173 = NOT(I5577)
--	I8710 = NOT(g6517)
--	g2461 = NOT(I3593)
--	I7590 = NOT(g5605)
--	I3602 = NOT(g1491)
--	I3007 = NOT(g1439)
--	g2756 = NOT(g2353)
--	g2622 = NOT(I3764)
--	I3059 = NOT(g1519)
--	I3578 = NOT(g1484)
--	I3868 = NOT(g2125)
--	g5888 = NOT(g5731)
--	g1256 = NOT(g838)
--	g6519 = NOT(I8473)
--	I6289 = NOT(g4433)
--	I9024 = NOT(g6803)
--	I5448 = NOT(g3960)
--	I3767 = NOT(g2125)
--	g5787 = NOT(g5685)
--	g2904 = NOT(g1991)
--	g6552 = NOT(I8552)
--	g6606 = NOT(I8684)
--	g2446 = NOT(I3581)
--	I5333 = NOT(g3491)
--	I2284 = NOT(g922)
--	g1381 = NOT(I2417)
--	g4718 = NOT(I6334)
--	g4767 = NOT(g4601)
--	I3261 = NOT(g1783)
--	g1847 = NOT(I2943)
--	I4688 = NOT(g3207)
--	I5774 = NOT(g3807)
--	I9077 = NOT(g6845)
--	I8659 = NOT(g6523)
--	g4535 = NOT(g4173)
--	I4976 = NOT(g3575)
--	g1685 = NOT(I2671)
--	g2145 = NOT(I3268)
--	I8506 = NOT(g6483)
--	g2841 = NOT(g2541)
--	g4582 = NOT(g4210)
--	g3022 = NOT(I4229)
--	g2391 = NOT(I3534)
--	g6586 = NOT(I8626)
--	g952 = NOT(I2029)
--	g1263 = NOT(g846)
--	g964 = NOT(g357)
--	I2420 = NOT(g791)
--	g2695 = NOT(I3843)
--	g2637 = NOT(I3779)
--	g1950 = NOT(I3059)
--	g5138 = NOT(I6792)
--	g4227 = NOT(g4059)
--	I7295 = NOT(g5439)
--	g5791 = NOT(I7590)
--	g3798 = NOT(g3388)
--	I9104 = NOT(g6864)
--	g5309 = NOT(g5063)
--	g2159 = NOT(I3284)
--	g6570 = NOT(I8594)
--	g4246 = NOT(I5692)
--	I6132 = NOT(g4219)
--	I8174 = NOT(g6173)
--	g6525 = NOT(I8491)
--	g6710 = NOT(I8840)
--	I5418 = NOT(g4036)
--	I6680 = NOT(g4713)
--	g4721 = NOT(I6343)
--	g1631 = NOT(I2588)
--	g2416 = NOT(I3556)
--	g3095 = NOT(I4340)
--	g3037 = NOT(I4252)
--	I3502 = NOT(g1295)
--	g1257 = NOT(g845)
--	g1101 = NOT(I2125)
--	I2204 = NOT(g694)
--	I2630 = NOT(g1143)
--	I5493 = NOT(g3834)
--	I8180 = NOT(g6176)
--	I4220 = NOT(g2164)
--	I7966 = NOT(g6166)
--	I8591 = NOT(g6448)
--	g2315 = NOT(I3465)
--	g5957 = NOT(g5866)
--	g6879 = NOT(I9104)
--	g6607 = NOT(I8687)
--	I6558 = NOT(g4705)
--	g4502 = NOT(I6020)
--	g5049 = NOT(I6685)
--	I9044 = NOT(g6836)
--	g927 = NOT(I1958)
--	I1942 = NOT(g664)
--	I4023 = NOT(g2315)
--	g3719 = NOT(g3053)
--	g6506 = NOT(I8438)
--	g5575 = NOT(g5411)
--	I8420 = NOT(g6422)
--	I3388 = NOT(g1324)
--	g2874 = NOT(g1849)
--	g3752 = NOT(I4935)
--	I5397 = NOT(g3932)
--	I3028 = NOT(g1504)
--	g4188 = NOT(I5594)
--	g6587 = NOT(I8629)
--	g4388 = NOT(I5871)
--	I5421 = NOT(g3724)
--	I3428 = NOT(g1825)
--	I2973 = NOT(g1687)
--	I7254 = NOT(g5458)
--	I7814 = NOT(g5922)
--	I3247 = NOT(g1791)
--	g3042 = NOT(I4261)
--	g6615 = NOT(I8707)
--	I7150 = NOT(g5355)
--	I4327 = NOT(g2525)
--	g4428 = NOT(I5933)
--	g3786 = NOT(g3388)
--	g5584 = NOT(I7346)
--	g5539 = NOT(g5331)
--	g5896 = NOT(g5753)
--	g1673 = NOT(I2653)
--	g6374 = NOT(I8186)
--	I3826 = NOT(g2145)
--	g3364 = NOT(g3114)
--	g3233 = NOT(I4498)
--	I8515 = NOT(g6492)
--	g4564 = NOT(g4192)
--	g3054 = NOT(I4279)
--	I5562 = NOT(g4002)
--	I4303 = NOT(g1897)
--	g2612 = NOT(I3752)
--	I8300 = NOT(g6299)
--	g6284 = NOT(I8002)
--	g2243 = NOT(I3376)
--	g3770 = NOT(I4961)
--	I9014 = NOT(g6820)
--	I3638 = NOT(g1484)
--	g1772 = NOT(I2811)
--	I5723 = NOT(g3942)
--	g4741 = NOT(I6371)
--	g6591 = NOT(I8641)
--	g5052 = NOT(I6692)
--	g6832 = NOT(I9021)
--	g4910 = NOT(I6612)
--	I2648 = NOT(g980)
--	g2234 = NOT(I3367)
--	g6853 = NOT(I9082)
--	g1890 = NOT(g1359)
--	I3883 = NOT(g2574)
--	g6420 = NOT(I8270)
--	I4240 = NOT(g2165)
--	g2330 = NOT(g1777)
--	g4108 = NOT(I5406)
--	g4609 = NOT(I6182)
--	g6507 = NOT(I8441)
--	g4308 = NOT(I5777)
--	g1011 = NOT(I2050)
--	g1734 = NOT(g952)
--	I3758 = NOT(g2041)
--	g5086 = NOT(g4732)
--	g897 = NOT(g41)
--	I8040 = NOT(g6142)
--	g951 = NOT(g84)
--	I8969 = NOT(g6797)
--	g2800 = NOT(g2430)
--	g5730 = NOT(I7497)
--	g2554 = NOT(I3669)
--	g4758 = NOT(I6382)
--	I2839 = NOT(g1123)
--	I3861 = NOT(g1834)
--	g6905 = NOT(I9182)
--	g3029 = NOT(I4240)
--	I3711 = NOT(g1848)
--	I9182 = NOT(g6879)
--	g3787 = NOT(I4986)
--	g2213 = NOT(I3346)
--	g5897 = NOT(g5731)
--	g5025 = NOT(g4814)
--	g6515 = NOT(g6408)
--	g4861 = NOT(I6587)
--	g5425 = NOT(I7091)
--	I4347 = NOT(g2555)
--	I2172 = NOT(g691)
--	I2278 = NOT(g917)
--	g4711 = NOT(I6315)
--	g6100 = NOT(I7796)
--	I4681 = NOT(g2947)
--	g1480 = NOT(g985)
--	g2902 = NOT(g1899)
--	I8875 = NOT(g6697)
--	I2143 = NOT(g2)
--	I2343 = NOT(g1177)
--	I6139 = NOT(g4222)
--	g4133 = NOT(I5481)
--	g3297 = NOT(g3046)
--	g2512 = NOT(I3638)
--	g2090 = NOT(I3206)
--	g4846 = NOT(I6546)
--	I2134 = NOT(g705)
--	I6795 = NOT(g5022)
--	I6737 = NOT(g4662)
--	I2334 = NOT(g1193)
--	I6809 = NOT(g5051)
--	I5743 = NOT(g4022)
--	g5331 = NOT(I6995)
--	I5890 = NOT(g3878)
--	I3509 = NOT(g1461)
--	g3963 = NOT(I5217)
--	g3791 = NOT(g3388)
--	I8884 = NOT(g6704)
--	I5505 = NOT(g3860)
--	g1688 = NOT(I2688)
--	I6672 = NOT(g4752)
--	g4780 = NOT(I6434)
--	g6040 = NOT(g5824)
--	g1857 = NOT(I2961)
--	I6231 = NOT(g4350)
--	I3662 = NOT(g1688)
--	g4509 = NOT(I6039)
--	g5087 = NOT(g4736)
--	I9095 = NOT(g6855)
--	g5801 = NOT(I7600)
--	g2155 = NOT(I3274)
--	I9208 = NOT(g6922)
--	g4662 = NOT(g4640)
--	I3093 = NOT(g1426)
--	g965 = NOT(I2033)
--	I3493 = NOT(g1461)
--	I3816 = NOT(g2580)
--	g1326 = NOT(g894)
--	I8235 = NOT(g6312)
--	I6099 = NOT(g4398)
--	I8282 = NOT(g6309)
--	g3049 = NOT(I4270)
--	g6528 = NOT(I8500)
--	g1760 = NOT(I2785)
--	g4493 = NOT(I6001)
--	g6351 = NOT(I8107)
--	I1850 = NOT(g210)
--	g6875 = NOT(I9092)
--	g834 = NOT(g341)
--	I8988 = NOT(g6787)
--	g6530 = NOT(I8506)
--	g3575 = NOT(I4777)
--	g5045 = NOT(I6677)
--	I8693 = NOT(g6570)
--	g6655 = NOT(I8761)
--	g5445 = NOT(g5274)
--	I5713 = NOT(g4022)
--	g3604 = NOT(I4799)
--	I8548 = NOT(g6454)
--	g5491 = NOT(I7193)
--	g3498 = NOT(g2634)
--	g4381 = NOT(I5854)
--	g4847 = NOT(I6549)
--	g2118 = NOT(I3247)
--	g2619 = NOT(I3761)
--	I8555 = NOT(g6456)
--	g2367 = NOT(I3519)
--	g2872 = NOT(g1922)
--	g1608 = NOT(I2570)
--	g1220 = NOT(I2221)
--	g4700 = NOT(I6292)
--	g6410 = NOT(I8240)
--	I9164 = NOT(g6885)
--	g4397 = NOT(I5890)
--	I9233 = NOT(g6938)
--	I2776 = NOT(g1192)
--	I7640 = NOT(g5773)
--	g5407 = NOT(I7073)
--	g6884 = NOT(I9119)
--	I2593 = NOT(g1177)
--	g5059 = NOT(I6697)
--	g5920 = NOT(I7692)
--	g6839 = NOT(I9038)
--	g2457 = NOT(I3587)
--	g5578 = NOT(g5425)
--	I6444 = NOT(g4503)
--	I6269 = NOT(g4655)
--	g1423 = NOT(I2442)
--	g923 = NOT(g332)
--	I5857 = NOT(g3740)
--	I7176 = NOT(g5437)
--	g1588 = NOT(g798)
--	I8113 = NOT(g6147)
--	g5582 = NOT(I7342)
--	g1161 = NOT(I2182)
--	g6278 = NOT(I7966)
--	g2686 = NOT(I3830)
--	g6372 = NOT(I8180)
--	g3162 = NOT(I4402)
--	g5261 = NOT(I6918)
--	g3019 = NOT(I4226)
--	I4294 = NOT(g2525)
--	I6543 = NOT(g4718)
--	g6618 = NOT(I8716)
--	g1665 = NOT(g985)
--	I7829 = NOT(g5926)
--	I3723 = NOT(g2158)
--	g6143 = NOT(I7865)
--	g4562 = NOT(I6132)
--	g6235 = NOT(g6062)
--	g2598 = NOT(I3726)
--	g3052 = NOT(I4273)
--	g1327 = NOT(I2334)
--	I2521 = NOT(g1063)
--	I3301 = NOT(g1730)
--	g5415 = NOT(I7081)
--	g3452 = NOT(g2625)
--	g6282 = NOT(I7996)
--	I2050 = NOT(g683)
--	I5400 = NOT(g3963)
--	g6566 = NOT(I8582)
--	I8494 = NOT(g6428)
--	I4501 = NOT(g2705)
--	I6534 = NOT(g4706)
--	I8518 = NOT(g6494)
--	I3605 = NOT(g1681)
--	g4723 = NOT(I6349)
--	I8567 = NOT(g6432)
--	g4101 = NOT(I5385)
--	g6134 = NOT(I7852)
--	g5664 = NOT(g5521)
--	g2625 = NOT(I3767)
--	I7270 = NOT(g5352)
--	g2232 = NOT(I3361)
--	g6548 = NOT(I8548)
--	I6927 = NOT(g5124)
--	g3086 = NOT(I4327)
--	I2724 = NOT(g1220)
--	g2253 = NOT(I3388)
--	I2179 = NOT(g293)
--	g3486 = NOT(g2869)
--	g2813 = NOT(g2457)
--	I2379 = NOT(g1123)
--	g1696 = NOT(I2700)
--	I7073 = NOT(g5281)
--	I7796 = NOT(g5917)
--	I6885 = NOT(g4872)
--	I6414 = NOT(g4497)
--	g3504 = NOT(g2675)
--	I6946 = NOT(g5124)
--	g1732 = NOT(I2738)
--	g3881 = NOT(I5116)
--	g2740 = NOT(I3909)
--	I2658 = NOT(g1001)
--	I3441 = NOT(g1502)
--	I7069 = NOT(g5281)
--	g3070 = NOT(I4297)
--	I8264 = NOT(g6296)
--	g6621 = NOT(I8721)
--	I2835 = NOT(g1209)
--	I7469 = NOT(g5625)
--	g3897 = NOT(g3251)
--	I5023 = NOT(g3263)
--	g1472 = NOT(g952)
--	g1043 = NOT(g486)
--	I5977 = NOT(g4319)
--	I8521 = NOT(g6495)
--	I6036 = NOT(g4370)
--	I8641 = NOT(g6524)
--	I2611 = NOT(g1209)
--	g893 = NOT(g23)
--	g2687 = NOT(I3833)
--	I8450 = NOT(g6412)
--	I3669 = NOT(g1739)
--	g1116 = NOT(I2154)
--	g2586 = NOT(I3711)
--	I3531 = NOT(g1593)
--	I5451 = NOT(g3967)
--	I6182 = NOT(g4249)
--	g6518 = NOT(I8470)
--	g6567 = NOT(I8585)
--	I8724 = NOT(g6533)
--	I6382 = NOT(g4460)
--	g996 = NOT(I2041)
--	g3331 = NOT(g3076)
--	I3890 = NOT(g2145)
--	g4772 = NOT(I6420)
--	g5247 = NOT(g4900)
--	g4531 = NOT(I6105)
--	I5633 = NOT(g3768)
--	I8878 = NOT(g6710)
--	g1681 = NOT(I2663)
--	I3505 = NOT(g1305)
--	g6593 = NOT(I8647)
--	g3766 = NOT(I4955)
--	g1533 = NOT(g878)
--	g5564 = NOT(g5382)
--	I5103 = NOT(g3440)
--	g2525 = NOT(I3650)
--	g3801 = NOT(g3388)
--	g3487 = NOT(g2622)
--	g1914 = NOT(I3013)
--	I5696 = NOT(g3942)
--	g2691 = NOT(g2317)
--	g4011 = NOT(g3486)
--	I6798 = NOT(g5042)
--	g4856 = NOT(I6576)
--	g5741 = NOT(g5602)
--	I2802 = NOT(g1204)
--	I3074 = NOT(g1426)
--	I3474 = NOT(g1450)
--	I5753 = NOT(g4022)
--	g5638 = NOT(I7397)
--	g6160 = NOT(g5926)
--	g3226 = NOT(I4477)
--	I5508 = NOT(g3867)
--	g6360 = NOT(I8144)
--	g6933 = NOT(I9220)
--	I5944 = NOT(g4356)
--	g2962 = NOT(g2008)
--	g6521 = NOT(I8479)
--	I9098 = NOT(g6864)
--	g2158 = NOT(I3281)
--	I5472 = NOT(g3846)
--	I8981 = NOT(g6793)
--	g2506 = NOT(I3632)
--	I3080 = NOT(g1519)
--	I8674 = NOT(g6521)
--	g1820 = NOT(I2880)
--	I5043 = NOT(g3247)
--	I6495 = NOT(g4607)
--	g1936 = NOT(g1756)
--	I6437 = NOT(g4501)
--	g3173 = NOT(I4410)
--	I6102 = NOT(g4399)
--	I6302 = NOT(g4440)
--	I8997 = NOT(g6790)
--	g1117 = NOT(g32)
--	I8541 = NOT(g6452)
--	g1317 = NOT(I2306)
--	g3491 = NOT(g2608)
--	g2587 = NOT(I3714)
--	I6579 = NOT(g4798)
--	I5116 = NOT(g3259)
--	I7852 = NOT(g5993)
--	I5316 = NOT(g3557)
--	g6724 = NOT(I8866)
--	I3569 = NOT(g1789)
--	g2111 = NOT(g1384)
--	g2275 = NOT(I3422)
--	g5466 = NOT(I7146)
--	I8332 = NOT(g6306)
--	g4713 = NOT(I6321)
--	I7701 = NOT(g5720)
--	g3369 = NOT(I4646)
--	I8153 = NOT(g6185)
--	g3007 = NOT(g2197)
--	g2615 = NOT(I3755)
--	g6878 = NOT(I9101)
--	I2864 = NOT(g1177)
--	g4569 = NOT(I6143)
--	g5571 = NOT(g5395)
--	g5861 = NOT(g5636)
--	g3868 = NOT(g3491)
--	g2174 = NOT(I3313)
--	g3459 = NOT(g2664)
--	g815 = NOT(I1877)
--	g1775 = NOT(g952)
--	g5448 = NOT(g5278)
--	g1922 = NOT(I3025)
--	g835 = NOT(g345)
--	g5711 = NOT(I7472)
--	g6835 = NOT(I9028)
--	g1581 = NOT(g910)
--	g6882 = NOT(I9113)
--	I6042 = NOT(g4374)
--	g1060 = NOT(g107)
--	g2284 = NOT(I3431)
--	I6786 = NOT(g4824)
--	g1460 = NOT(I2457)
--	g5774 = NOT(I7517)
--	g4857 = NOT(I6579)
--	g3793 = NOT(g3491)
--	g6611 = NOT(I8699)
--	g2591 = NOT(I3720)
--	g3015 = NOT(I4220)
--	g3227 = NOT(I4480)
--	g1739 = NOT(I2749)
--	I6054 = NOT(g4194)
--	g5538 = NOT(g5331)
--	I6296 = NOT(g4436)
--	I4646 = NOT(g2602)
--	I2623 = NOT(g1161)
--	g4126 = NOT(I5460)
--	g5509 = NOT(I7251)
--	g4400 = NOT(I5899)
--	g1937 = NOT(I3044)
--	g6541 = NOT(I8535)
--	I9185 = NOT(g6877)
--	I2476 = NOT(g971)
--	I7336 = NOT(g5534)
--	I8600 = NOT(g6451)
--	g2931 = NOT(g1988)
--	g4760 = NOT(I6386)
--	g1294 = NOT(I2287)
--	I1877 = NOT(g283)
--	g6332 = NOT(I8074)
--	g5067 = NOT(g4801)
--	g1190 = NOT(I2199)
--	I2175 = NOT(g25)
--	g6353 = NOT(I8113)
--	g5994 = NOT(g5873)
--	I3608 = NOT(g1461)
--	g2905 = NOT(g1994)
--	I6012 = NOT(g4167)
--	g6744 = NOT(I8910)
--	I3779 = NOT(g2125)
--	g6802 = NOT(I8972)
--	g2628 = NOT(I3770)
--	g1156 = NOT(I2175)
--	g2515 = NOT(I3641)
--	g5493 = NOT(I7197)
--	I7065 = NOT(g5281)
--	g5256 = NOT(g5077)
--	I6706 = NOT(g4731)
--	g4220 = NOT(I5644)
--	g3940 = NOT(I5177)
--	I6371 = NOT(g4569)
--	I4276 = NOT(g2170)
--	g4423 = NOT(I5920)
--	I3161 = NOT(g1270)
--	I3361 = NOT(g1331)
--	g5381 = NOT(I7039)
--	g3388 = NOT(I4667)
--	I9131 = NOT(g6855)
--	I6956 = NOT(g5124)
--	g6901 = NOT(I9170)
--	I5460 = NOT(g3771)
--	I5597 = NOT(g3821)
--	I8623 = NOT(g6542)
--	g3216 = NOT(I4459)
--	I3665 = NOT(g1824)
--	g5685 = NOT(g5552)
--	g6511 = NOT(I8453)
--	I8476 = NOT(g6457)
--	I2424 = NOT(g719)
--	g743 = NOT(I1844)
--	g862 = NOT(g319)
--	g2973 = NOT(I4170)
--	g1954 = NOT(I3065)
--	g3030 = NOT(I4243)
--	g1250 = NOT(g123)
--	I5739 = NOT(g3942)
--	g1363 = NOT(I2399)
--	I4986 = NOT(g3638)
--	I3999 = NOT(g1837)
--	g3247 = NOT(g2973)
--	g4127 = NOT(I5463)
--	I3346 = NOT(g1327)
--	g5950 = NOT(g5730)
--	g1053 = NOT(g197)
--	g2040 = NOT(g1738)
--	g6600 = NOT(I8668)
--	g6574 = NOT(g6484)
--	I2231 = NOT(g465)
--	I1844 = NOT(g208)
--	g2440 = NOT(I3575)
--	g3564 = NOT(g2618)
--	g6714 = NOT(g6670)
--	I2643 = NOT(g965)
--	g4146 = NOT(I5520)
--	I5668 = NOT(g3828)
--	g4633 = NOT(g4284)
--	I8285 = NOT(g6310)
--	I5840 = NOT(g3732)
--	I8500 = NOT(g6431)
--	g791 = NOT(I1865)
--	g4103 = NOT(I5391)
--	g6580 = NOT(g6491)
--	I7859 = NOT(g6032)
--	g5631 = NOT(g5536)
--	g3638 = NOT(g3108)
--	g5723 = NOT(I7484)
--	I9173 = NOT(g6876)
--	I3240 = NOT(g1460)
--	g4732 = NOT(I6362)
--	g3108 = NOT(I4354)
--	g3308 = NOT(g3060)
--	I6759 = NOT(g4778)
--	g2875 = NOT(g1940)
--	g4753 = NOT(I6377)
--	g4508 = NOT(I6036)
--	g917 = NOT(I1942)
--	I8809 = NOT(g6687)
--	I7342 = NOT(g5579)
--	g6623 = NOT(I8727)
--	g6076 = NOT(g5797)
--	I7081 = NOT(g5281)
--	g6889 = NOT(I9134)
--	g5751 = NOT(I7506)
--	I3316 = NOT(g1344)
--	g3589 = NOT(g3094)
--	I7481 = NOT(g5629)
--	I3034 = NOT(g1519)
--	g3466 = NOT(I4706)
--	g2410 = NOT(I3550)
--	I7692 = NOT(g5711)
--	I3434 = NOT(g1627)
--	I4516 = NOT(g2777)
--	I7497 = NOT(g5687)
--	g4116 = NOT(I5430)
--	g6375 = NOT(I8189)
--	g2884 = NOT(g1957)
--	I2044 = NOT(g681)
--	g3571 = NOT(g3084)
--	g2839 = NOT(g2535)
--	g3861 = NOT(I5084)
--	g6722 = NOT(I8860)
--	g4034 = NOT(I5333)
--	I7960 = NOT(g5925)
--	g852 = NOT(g634)
--	I2269 = NOT(g899)
--	g6651 = NOT(I8749)
--	g3448 = NOT(I4684)
--	g4565 = NOT(g4195)
--	I3681 = NOT(g1821)
--	I5053 = NOT(g3710)
--	g3455 = NOT(g2637)
--	g6285 = NOT(I8005)
--	g4147 = NOT(I5523)
--	g6500 = NOT(I8420)
--	g2172 = NOT(I3307)
--	I2712 = NOT(g1203)
--	I9227 = NOT(g6937)
--	I5568 = NOT(g3897)
--	g4533 = NOT(I6111)
--	g3846 = NOT(I5053)
--	g2618 = NOT(I3758)
--	I3596 = NOT(g1305)
--	g2667 = NOT(I3811)
--	g1683 = NOT(g1017)
--	g2343 = NOT(I3493)
--	g5168 = NOT(g5099)
--	I3013 = NOT(g1519)
--	g6339 = NOT(I8093)
--	g3196 = NOT(I4433)
--	g4914 = NOT(g4816)
--	g3803 = NOT(I5002)
--	g4210 = NOT(I5630)
--	I7267 = NOT(g5458)
--	g1894 = NOT(I2989)
--	I5157 = NOT(g3454)
--	g6838 = NOT(I9035)
--	I9203 = NOT(g6921)
--	I2961 = NOT(g1731)
--	g6424 = NOT(I8282)
--	g2134 = NOT(I3258)
--	I6362 = NOT(g4569)
--	g1735 = NOT(I2745)
--	I8273 = NOT(g6301)
--	g6809 = NOT(I8981)
--	g5890 = NOT(g5753)
--	g1782 = NOT(I2828)
--	I4340 = NOT(g1935)
--	I6452 = NOT(g4629)
--	I5929 = NOT(g4152)
--	g1661 = NOT(g1076)
--	I8044 = NOT(g6252)
--	g2555 = NOT(I3672)
--	g6231 = NOT(g6044)
--	g5011 = NOT(I6649)
--	I8444 = NOT(g6421)
--	g3067 = NOT(I4294)
--	I2414 = NOT(g784)
--	g729 = NOT(I1838)
--	g5411 = NOT(I7077)
--	g6523 = NOT(I8485)
--	g861 = NOT(g179)
--	I2946 = NOT(g1587)
--	g2792 = NOT(g2416)
--	g1627 = NOT(I2584)
--	g4117 = NOT(I5433)
--	g1292 = NOT(I2281)
--	I5626 = NOT(g3914)
--	g3093 = NOT(I4334)
--	g898 = NOT(g47)
--	g1998 = NOT(I3109)
--	g1646 = NOT(I2617)
--	g5992 = NOT(g5869)
--	g4601 = NOT(g4191)
--	g1084 = NOT(g98)
--	g6104 = NOT(I7808)
--	g854 = NOT(g646)
--	g1039 = NOT(g662)
--	g1484 = NOT(I2473)
--	I3581 = NOT(g1491)
--	g6499 = NOT(I8417)
--	g1439 = NOT(I2449)
--	I9028 = NOT(g6806)
--	I8961 = NOT(g6778)
--	g4775 = NOT(I6425)
--	I6470 = NOT(g4473)
--	g5573 = NOT(g5403)
--	g3847 = NOT(I5056)
--	g5480 = NOT(I7176)
--	I6425 = NOT(g4619)
--	I2831 = NOT(g1209)
--	g2494 = NOT(I3623)
--	I2182 = NOT(g692)
--	g2518 = NOT(I3644)
--	g1583 = NOT(g1001)
--	g1702 = NOT(g1107)
--	I2382 = NOT(g719)
--	I8414 = NOT(g6418)
--	g3263 = NOT(g3015)
--	I8946 = NOT(g6778)
--	g1919 = NOT(I3022)
--	I2805 = NOT(g1205)
--	I2916 = NOT(g1643)
--	g2776 = NOT(g2378)
--	I2749 = NOT(g1209)
--	g4784 = NOT(I6444)
--	g6044 = NOT(g5824)
--	g1276 = NOT(g847)
--	I4402 = NOT(g2283)
--	I3294 = NOT(g1720)
--	I3840 = NOT(g2125)
--	I6406 = NOT(g4473)
--	I5475 = NOT(g3852)
--	g6572 = NOT(I8600)
--	I4762 = NOT(g2862)
--	I7349 = NOT(g5532)
--	I6635 = NOT(g4745)
--	g2264 = NOT(I3405)
--	g6712 = NOT(g6676)
--	g851 = NOT(g606)
--	I6766 = NOT(g4783)
--	I6087 = NOT(g4392)
--	I6105 = NOT(g4400)
--	g6543 = NOT(I8541)
--	g4840 = NOT(I6528)
--	I6305 = NOT(g4441)
--	I6801 = NOT(g5045)
--	g2360 = NOT(g1793)
--	g2933 = NOT(I4123)
--	g3723 = NOT(I4903)
--	g1647 = NOT(I2620)
--	g4190 = NOT(I5600)
--	I5526 = NOT(g3848)
--	I5998 = NOT(g4157)
--	I8335 = NOT(g6308)
--	I8831 = NOT(g6665)
--	I9217 = NOT(g6931)
--	g1546 = NOT(g1101)
--	I2873 = NOT(g1161)
--	I2037 = NOT(g679)
--	g6534 = NOT(I8518)
--	g6729 = NOT(I8881)
--	g3605 = NOT(I4802)
--	I5084 = NOT(g3593)
--	I5603 = NOT(g3893)
--	g2996 = NOT(I4189)
--	I2653 = NOT(g996)
--	I5484 = NOT(g3875)
--	I3942 = NOT(g1833)
--	g1503 = NOT(g878)
--	I5439 = NOT(g3730)
--	I8916 = NOT(g6742)
--	g1925 = NOT(I3028)
--	I8749 = NOT(g6560)
--	g2179 = NOT(I3328)
--	g6014 = NOT(g5824)
--	g6885 = NOT(I9122)
--	I6045 = NOT(g4375)
--	g4704 = NOT(I6302)
--	g6414 = NOT(I8252)
--	I5702 = NOT(g3845)
--	g1320 = NOT(I2315)
--	g3041 = NOT(I4258)
--	g5383 = NOT(I7045)
--	g5924 = NOT(I7704)
--	g5220 = NOT(g4903)
--	I7119 = NOT(g5303)
--	g6903 = NOT(I9176)
--	g2777 = NOT(I3965)
--	g3441 = NOT(I4681)
--	g2835 = NOT(g2506)
--	I3053 = NOT(g1407)
--	I1958 = NOT(g702)
--	g4250 = NOT(I5702)
--	g6513 = NOT(I8459)
--	g913 = NOT(g658)
--	I6283 = NOT(g4613)
--	I7258 = NOT(g5458)
--	I5952 = NOT(g4367)
--	g4810 = NOT(I6488)
--	g2882 = NOT(g1854)
--	I7352 = NOT(g5533)
--	g3673 = NOT(g3075)
--	I2442 = NOT(g872)
--	g1789 = NOT(I2839)
--	g6036 = NOT(g5824)
--	I8632 = NOT(g6548)
--	I2364 = NOT(g1143)
--	g980 = NOT(I2037)
--	I8653 = NOT(g6531)
--	g1771 = NOT(I2808)
--	g3772 = NOT(g3466)
--	I6582 = NOT(g4765)
--	g5051 = NOT(I6689)
--	g2981 = NOT(g2179)
--	I8579 = NOT(g6438)
--	I8869 = NOT(g6694)
--	I4489 = NOT(g2975)
--	g3458 = NOT(g2656)
--	g865 = NOT(g188)
--	I2296 = NOT(g893)
--	g3890 = NOT(g3575)
--	g2997 = NOT(I4192)
--	I6015 = NOT(g4170)
--	g2541 = NOT(I3659)
--	I8752 = NOT(g6514)
--	I4471 = NOT(g3040)
--	I7170 = NOT(g5435)
--	g6422 = NOT(I8276)
--	g2353 = NOT(I3505)
--	g4929 = NOT(I6621)
--	I4955 = NOT(g3673)
--	I3626 = NOT(g1684)
--	g2744 = NOT(g2336)
--	g909 = NOT(I1935)
--	g1738 = NOT(g1108)
--	g2802 = NOT(g2437)
--	g3074 = NOT(I4303)
--	g949 = NOT(g79)
--	g1991 = NOT(I3102)
--	g6560 = NOT(I8564)
--	I5320 = NOT(g3559)
--	g4626 = NOT(g4270)
--	g1340 = NOT(I2373)
--	I2029 = NOT(g677)
--	I9021 = NOT(g6812)
--	g3480 = NOT(g2986)
--	g1690 = NOT(I2692)
--	g6653 = NOT(I8755)
--	g6102 = NOT(I7802)
--	I2281 = NOT(g900)
--	I7061 = NOT(g5281)
--	I7187 = NOT(g5387)
--	g6579 = NOT(g6490)
--	g5116 = NOT(g4810)
--	I5987 = NOT(g4224)
--	g5316 = NOT(I6976)
--	g1656 = NOT(I2635)
--	I6689 = NOT(g4758)
--	g5434 = NOT(I7110)
--	g2574 = NOT(I3681)
--	g2864 = NOT(g1887)
--	g4778 = NOT(I6430)
--	g855 = NOT(g650)
--	g5147 = NOT(I6809)
--	I3782 = NOT(g2145)
--	g4894 = NOT(g4813)
--	I2745 = NOT(g1249)
--	I8189 = NOT(g6179)
--	I4229 = NOT(g2284)
--	I6430 = NOT(g4620)
--	g3976 = NOT(I5252)
--	I2791 = NOT(g1236)
--	I6247 = NOT(g4609)
--	I7514 = NOT(g5590)
--	I2309 = NOT(g1236)
--	I9101 = NOT(g6855)
--	g1110 = NOT(I2140)
--	I8888 = NOT(g6708)
--	g2580 = NOT(I3691)
--	g5210 = NOT(I6874)
--	g6786 = NOT(I8946)
--	I6564 = NOT(g4712)
--	I8171 = NOT(g6170)
--	I2808 = NOT(g1161)
--	I8429 = NOT(g6425)
--	g5596 = NOT(I7358)
--	g6164 = NOT(g5926)
--	g6364 = NOT(I8156)
--	g6233 = NOT(g6052)
--	I5991 = NOT(g4226)
--	I2707 = NOT(g1190)
--	g4292 = NOT(g4059)
--	I7695 = NOT(g5714)
--	I7637 = NOT(g5751)
--	g2968 = NOT(g2179)
--	I5078 = NOT(g3719)
--	g1824 = NOT(I2890)
--	g4526 = NOT(I6090)
--	I5478 = NOT(g3859)
--	g1236 = NOT(I2234)
--	I7107 = NOT(g5277)
--	I5907 = NOT(g3883)
--	g6725 = NOT(I8869)
--	g1762 = NOT(I2791)
--	g2889 = NOT(g1975)
--	I6108 = NOT(g4403)
--	g4603 = NOT(I6170)
--	g6532 = NOT(I8512)
--	I6308 = NOT(g4443)
--	I5517 = NOT(g3885)
--	I9041 = NOT(g6835)
--	I2449 = NOT(g971)
--	g4439 = NOT(I5952)
--	g5117 = NOT(I6763)
--	g6553 = NOT(I8555)
--	g4850 = NOT(I6558)
--	I8684 = NOT(g6567)
--	I5876 = NOT(g3870)
--	I8745 = NOT(g6513)
--	g2175 = NOT(I3316)
--	g2871 = NOT(g1919)
--	I2604 = NOT(g1222)
--	g3183 = NOT(I4420)
--	g2722 = NOT(I3883)
--	I4462 = NOT(g2135)
--	I8309 = NOT(g6304)
--	g1556 = NOT(g878)
--	I6066 = NOT(g4382)
--	g3779 = NOT(g3466)
--	g1222 = NOT(I2225)
--	g4702 = NOT(I6296)
--	g6412 = NOT(I8246)
--	g896 = NOT(g22)
--	g3023 = NOT(g2215)
--	I7251 = NOT(g5458)
--	g1928 = NOT(I3031)
--	I7811 = NOT(g5921)
--	g6706 = NOT(I8828)
--	g5922 = NOT(I7698)
--	I8707 = NOT(g6520)
--	g1064 = NOT(g102)
--	I2584 = NOT(g839)
--	I5214 = NOT(g3567)
--	g6888 = NOT(I9131)
--	g1899 = NOT(I2998)
--	I6048 = NOT(g4376)
--	g5581 = NOT(I7339)
--	I6448 = NOT(g4626)
--	g6371 = NOT(I8177)
--	g4276 = NOT(I5731)
--	I4249 = NOT(g2525)
--	g5597 = NOT(I7361)
--	I3004 = NOT(g1426)
--	I1825 = NOT(g361)
--	g4561 = NOT(g4189)
--	g2838 = NOT(g2515)
--	I3647 = NOT(g1747)
--	g3451 = NOT(g2615)
--	I2162 = NOT(g197)
--	g1563 = NOT(g1006)
--	I9011 = NOT(g6819)
--	I4192 = NOT(g1847)
--	g2809 = NOT(I4019)
--	I3764 = NOT(g2044)
--	g5784 = NOT(I7583)
--	I3546 = NOT(g1586)
--	I5002 = NOT(g3612)
--	g4527 = NOT(I6093)
--	g4404 = NOT(I5907)
--	g1295 = NOT(I2290)
--	g4647 = NOT(g4296)
--	g3346 = NOT(I4623)
--	I5236 = NOT(g3545)
--	g2672 = NOT(I3816)
--	g2231 = NOT(I3358)
--	g4764 = NOT(I6400)
--	g5995 = NOT(g5824)
--	I9074 = NOT(g6844)
--	g5479 = NOT(I7173)
--	g2643 = NOT(I3785)
--	I6780 = NOT(g4825)
--	g6745 = NOT(I8913)
--	g1394 = NOT(g1206)
--	g4503 = NOT(I6023)
--	I7612 = NOT(g5605)
--	g1731 = NOT(I2735)
--	I2728 = NOT(g1232)
--	g1557 = NOT(g1017)
--	g2634 = NOT(I3776)
--	g1966 = NOT(I3077)
--	g4224 = NOT(g4046)
--	I5556 = NOT(g4059)
--	I2185 = NOT(g29)
--	g2104 = NOT(g1372)
--	g2099 = NOT(g1366)
--	g3240 = NOT(I4519)
--	I2385 = NOT(g784)
--	g6707 = NOT(I8831)
--	g1471 = NOT(I2464)
--	g4120 = NOT(I5442)
--	I4031 = NOT(g1846)
--	g4320 = NOT(g4011)
--	I4252 = NOT(g2555)
--	I3617 = NOT(g1305)
--	I3906 = NOT(g2234)
--	I6093 = NOT(g4394)
--	I8162 = NOT(g6189)
--	g3043 = NOT(I4264)
--	g971 = NOT(g658)
--	I5899 = NOT(g3748)
--	I4176 = NOT(g2268)
--	I6816 = NOT(g5111)
--	I3516 = NOT(g1295)
--	g2754 = NOT(g2347)
--	g4617 = NOT(g4242)
--	g3034 = NOT(I4249)
--	g1254 = NOT(g152)
--	g1814 = NOT(I2873)
--	g6575 = NOT(g6486)
--	g4516 = NOT(I6060)
--	g6715 = NOT(g6673)
--	g4771 = NOT(I6417)
--	g2044 = NOT(I3161)
--	I6685 = NOT(g4716)
--	g5250 = NOT(g4929)
--	g6604 = NOT(I8678)
--	g1038 = NOT(g127)
--	I6397 = NOT(g4473)
--	g6498 = NOT(I8414)
--	g1773 = NOT(I2814)
--	I2131 = NOT(g24)
--	g5432 = NOT(I7104)
--	g4299 = NOT(I5756)
--	g6833 = NOT(I9024)
--	I8730 = NOT(g6535)
--	g5453 = NOT(g5296)
--	I4270 = NOT(g2555)
--	g2862 = NOT(I4066)
--	I2635 = NOT(g1055)
--	g2712 = NOT(g2320)
--	I8881 = NOT(g6711)
--	I5394 = NOT(g4016)
--	g1769 = NOT(I2802)
--	g3914 = NOT(I5153)
--	g6584 = NOT(I8620)
--	I1859 = NOT(g277)
--	g6539 = NOT(I8531)
--	g6896 = NOT(I9155)
--	g1836 = NOT(I2922)
--	g5568 = NOT(g5423)
--	I8070 = NOT(g6116)
--	I5731 = NOT(g3942)
--	I8470 = NOT(g6461)
--	I8897 = NOT(g6707)
--	g1918 = NOT(I3019)
--	I3244 = NOT(g1772)
--	I7490 = NOT(g5583)
--	I4980 = NOT(g3546)
--	g5912 = NOT(g5853)
--	I4324 = NOT(g1918)
--	I3140 = NOT(g1317)
--	g2961 = NOT(g1861)
--	I5071 = NOT(g3263)
--	I3340 = NOT(g1282)
--	I5705 = NOT(g3942)
--	g6162 = NOT(g5926)
--	I3478 = NOT(g1450)
--	g6362 = NOT(I8150)
--	g6419 = NOT(I8267)
--	I6723 = NOT(g4761)
--	g4140 = NOT(I5502)
--	g6052 = NOT(g5824)
--	g2927 = NOT(g1979)
--	I5948 = NOT(g4360)
--	I9220 = NOT(g6930)
--	g2885 = NOT(g1963)
--	I7355 = NOT(g5535)
--	I8678 = NOT(g6565)
--	I2445 = NOT(g971)
--	g2660 = NOT(I3804)
--	g2946 = NOT(g2296)
--	g938 = NOT(g59)
--	g4435 = NOT(I5944)
--	I2373 = NOT(g1143)
--	g4517 = NOT(I6063)
--	I7698 = NOT(g5717)
--	I3656 = NOT(g1484)
--	g3601 = NOT(I4794)
--	I2491 = NOT(g821)
--	g2903 = NOT(g1902)
--	I8635 = NOT(g6552)
--	g6728 = NOT(I8878)
--	g6486 = NOT(g6363)
--	I2169 = NOT(g269)
--	g942 = NOT(g69)
--	g6730 = NOT(I8884)
--	I9161 = NOT(g6880)
--	g3775 = NOT(g3388)
--	g6504 = NOT(I8432)
--	g3922 = NOT(I5157)
--	I7463 = NOT(g5622)
--	I2578 = NOT(g1209)
--	g6385 = NOT(g6271)
--	g6881 = NOT(I9110)
--	I5409 = NOT(g3980)
--	g2036 = NOT(g1764)
--	g706 = NOT(I1825)
--	I6441 = NOT(g4624)
--	g4915 = NOT(g4669)
--	g2178 = NOT(I3325)
--	g2436 = NOT(I3569)
--	g2679 = NOT(I3823)
--	g6070 = NOT(g5824)
--	g2378 = NOT(I3525)
--	g3060 = NOT(I4285)
--	I3310 = NOT(g1640)
--	g6897 = NOT(I9158)
--	g1837 = NOT(I2925)
--	I8755 = NOT(g6561)
--	g3460 = NOT(g2667)
--	I8226 = NOT(g6328)
--	g6425 = NOT(I8285)
--	g2135 = NOT(I3261)
--	I4510 = NOT(g2753)
--	I9146 = NOT(g6890)
--	g4110 = NOT(I5412)
--	I7167 = NOT(g5434)
--	I7318 = NOT(g5452)
--	I4291 = NOT(g2241)
--	g5894 = NOT(g5731)
--	g2805 = NOT(g2443)
--	g910 = NOT(I1938)
--	g1788 = NOT(g985)
--	g2422 = NOT(I3560)
--	I6772 = NOT(g4788)
--	I7193 = NOT(g5466)
--	I8491 = NOT(g6480)
--	g3079 = NOT(I4312)
--	I6531 = NOT(g4704)
--	g4402 = NOT(g4017)
--	g784 = NOT(I1862)
--	g1249 = NOT(I2240)
--	g4824 = NOT(g4615)
--	g837 = NOT(g353)
--	g5661 = NOT(g5518)
--	g3840 = NOT(I5043)
--	g719 = NOT(I1835)
--	I3590 = NOT(g1781)
--	g6406 = NOT(I8232)
--	g5475 = NOT(I7161)
--	I7686 = NOT(g5705)
--	g1842 = NOT(g1612)
--	I2721 = NOT(g1219)
--	g1192 = NOT(g44)
--	I8459 = NOT(g6427)
--	g6105 = NOT(I7811)
--	g6087 = NOT(g5813)
--	g6801 = NOT(I8969)
--	g6305 = NOT(I8027)
--	g5292 = NOT(I6942)
--	I8767 = NOT(g6619)
--	g6487 = NOT(g6365)
--	I3556 = NOT(g1484)
--	g3501 = NOT(g2650)
--	I3222 = NOT(g1790)
--	I8535 = NOT(g6447)
--	g4657 = NOT(I6244)
--	I8582 = NOT(g6439)
--	g1854 = NOT(I2958)
--	I9116 = NOT(g6864)
--	I8261 = NOT(g6298)
--	g5084 = NOT(g4727)
--	g4222 = NOT(I5654)
--	g2437 = NOT(I3572)
--	g2653 = NOT(I3797)
--	I6992 = NOT(g5151)
--	I1932 = NOT(g667)
--	g2102 = NOT(I3222)
--	g5439 = NOT(g5261)
--	I3785 = NOT(g2346)
--	I2940 = NOT(g1653)
--	I5837 = NOT(g3850)
--	g2869 = NOT(g2433)
--	I2388 = NOT(g878)
--	I6573 = NOT(g4721)
--	I3563 = NOT(g1461)
--	g5702 = NOT(I7463)
--	I8246 = NOT(g6290)
--	g1219 = NOT(I2218)
--	g1640 = NOT(I2601)
--	g2752 = NOT(g2343)
--	g6373 = NOT(I8183)
--	g3363 = NOT(g3110)
--	g6491 = NOT(g6373)
--	g5919 = NOT(I7689)
--	I2671 = NOT(g1017)
--	g1812 = NOT(I2867)
--	I8721 = NOT(g6534)
--	I2428 = NOT(g774)
--	g4563 = NOT(g4190)
--	g3053 = NOT(I4276)
--	g1176 = NOT(I2190)
--	g2265 = NOT(I3408)
--	g3453 = NOT(g2628)
--	g6283 = NOT(I7999)
--	g6369 = NOT(I8171)
--	g2042 = NOT(I3155)
--	g6602 = NOT(I8674)
--	I5249 = NOT(g3589)
--	g6407 = NOT(I8235)
--	g6578 = NOT(g6489)
--	g4844 = NOT(I6540)
--	g2164 = NOT(I3291)
--	g1286 = NOT(g854)
--	g2364 = NOT(I3516)
--	g2233 = NOT(I3364)
--	g4194 = NOT(I5612)
--	g1911 = NOT(I3010)
--	g4394 = NOT(I5885)
--	g6535 = NOT(I8521)
--	I6976 = NOT(g5136)
--	g3912 = NOT(g3505)
--	I2741 = NOT(g1222)
--	g5527 = NOT(I7267)
--	g6582 = NOT(I8614)
--	I8940 = NOT(g6783)
--	g4731 = NOT(I6359)
--	I2910 = NOT(g1645)
--	I3071 = NOT(g1504)
--	g5647 = NOT(g5509)
--	I3705 = NOT(g2316)
--	I3471 = NOT(g1450)
--	g2296 = NOT(I3441)
--	g1733 = NOT(I2741)
--	I2638 = NOT(g1123)
--	g1270 = NOT(g844)
--	g5546 = NOT(g5388)
--	I5854 = NOT(g3857)
--	I4465 = NOT(g2945)
--	g6015 = NOT(g5857)
--	g4705 = NOT(I6305)
--	g6415 = NOT(I8255)
--	I6126 = NOT(g4240)
--	I6400 = NOT(g4473)
--	g4242 = NOT(I5686)
--	I2883 = NOT(g1143)
--	I8671 = NOT(g6519)
--	g5925 = NOT(I7707)
--	I8030 = NOT(g6239)
--	I4433 = NOT(g2103)
--	g1324 = NOT(I2327)
--	I5708 = NOT(g3942)
--	I5520 = NOT(g3835)
--	g6721 = NOT(I8857)
--	I5640 = NOT(g3770)
--	g5120 = NOT(I6772)
--	I8564 = NOT(g6429)
--	g2706 = NOT(I3861)
--	I5252 = NOT(g3546)
--	I3773 = NOT(g2524)
--	g1177 = NOT(I2193)
--	g4150 = NOT(I5532)
--	I2165 = NOT(g690)
--	g1206 = NOT(I2212)
--	g4350 = NOT(g4010)
--	g2888 = NOT(g1972)
--	I7358 = NOT(g5565)
--	I4195 = NOT(g2173)
--	g2029 = NOT(I3134)
--	I7506 = NOT(g5584)
--	I5376 = NOT(g4014)
--	g2171 = NOT(I3304)
--	I4337 = NOT(g1934)
--	I8910 = NOT(g6730)
--	g2787 = NOT(g2405)
--	g6502 = NOT(I8426)
--	g2956 = NOT(g1861)
--	I6023 = NOT(g4151)
--	I8638 = NOT(g6553)
--	g1287 = NOT(g855)
--	g2675 = NOT(I3819)
--	I3836 = NOT(g1832)
--	I3212 = NOT(g1806)
--	I7587 = NOT(g5605)
--	g6940 = NOT(I9233)
--	g4769 = NOT(g4606)
--	g1849 = NOT(I2949)
--	g3778 = NOT(g3388)
--	g6188 = NOT(g5950)
--	I2196 = NOT(g3)
--	g5299 = NOT(I6949)
--	g1781 = NOT(I2825)
--	I6051 = NOT(g4185)
--	g1898 = NOT(I2995)
--	g3782 = NOT(g3388)
--	I8217 = NOT(g6319)
--	I8758 = NOT(g6562)
--	I8066 = NOT(g6114)
--	g5892 = NOT(g5742)
--	I6327 = NOT(g4451)
--	g6428 = NOT(I8290)
--	g3075 = NOT(I4306)
--	g4229 = NOT(g4059)
--	g2109 = NOT(I3235)
--	I7284 = NOT(g5383)
--	I4255 = NOT(g2179)
--	I6346 = NOT(g4563)
--	I8165 = NOT(g6189)
--	g4822 = NOT(g4614)
--	g1291 = NOT(I2278)
--	I5124 = NOT(g3719)
--	I2067 = NOT(g686)
--	g6564 = NOT(I8576)
--	I5324 = NOT(g3466)
--	I7832 = NOT(g5943)
--	g6826 = NOT(I9011)
--	I5469 = NOT(g3838)
--	I2290 = NOT(g971)
--	g1344 = NOT(I2379)
--	I4354 = NOT(g1953)
--	g5140 = NOT(I6798)
--	I5177 = NOT(g3267)
--	g3084 = NOT(I4321)
--	g5478 = NOT(I7170)
--	g1819 = NOT(I2877)
--	I6753 = NOT(g4772)
--	g2957 = NOT(g1861)
--	I8803 = NOT(g6685)
--	g1088 = NOT(I2119)
--	g1852 = NOT(I2952)
--	I6072 = NOT(g4385)
--	g6609 = NOT(I8693)
--	g5435 = NOT(I7113)
--	g6308 = NOT(I8034)
--	I3062 = NOT(g1776)
--	g5082 = NOT(g4723)
--	g2449 = NOT(I3584)
--	I3620 = NOT(g1484)
--	I3462 = NOT(g1450)
--	I8538 = NOT(g6450)
--	g2575 = NOT(I3684)
--	g2865 = NOT(g2296)
--	g6883 = NOT(I9116)
--	g5876 = NOT(I7640)
--	g4837 = NOT(g4473)
--	I8509 = NOT(g6437)
--	I2700 = NOT(g1173)
--	g2604 = NOT(I3736)
--	I4267 = NOT(g2525)
--	g2098 = NOT(g1363)
--	I4312 = NOT(g2555)
--	g4620 = NOT(g4251)
--	g4462 = NOT(I5977)
--	g6589 = NOT(I8635)
--	g945 = NOT(g536)
--	I8662 = NOT(g6525)
--	I3788 = NOT(g2554)
--	g6466 = NOT(I8332)
--	g5915 = NOT(I7679)
--	g3952 = NOT(I5182)
--	I6434 = NOT(g4622)
--	I8467 = NOT(g6457)
--	I8994 = NOT(g6789)
--	I8290 = NOT(g6291)
--	g1114 = NOT(I2150)
--	g6165 = NOT(g5926)
--	g6571 = NOT(I8597)
--	g6365 = NOT(I8159)
--	g2584 = NOT(I3705)
--	g4788 = NOT(I6452)
--	g6048 = NOT(g5824)
--	I1841 = NOT(g207)
--	g6711 = NOT(I8843)
--	I8093 = NOT(g6122)
--	g5110 = NOT(I6740)
--	g4249 = NOT(I5699)
--	g5310 = NOT(g5067)
--	I3298 = NOT(g1725)
--	g1825 = NOT(I2893)
--	g6827 = NOT(I9014)
--	g1650 = NOT(I2627)
--	I3485 = NOT(g1450)
--	g3527 = NOT(I4743)
--	g809 = NOT(I1874)
--	I6697 = NOT(g4722)
--	g4842 = NOT(I6534)
--	g849 = NOT(g598)
--	g2268 = NOT(I3419)
--	g4192 = NOT(I5606)
--	g4392 = NOT(I5879)
--	g3546 = NOT(g3095)
--	g4485 = NOT(I5987)
--	I2817 = NOT(g1222)
--	g5824 = NOT(g5631)
--	g1336 = NOT(I2361)
--	g6803 = NOT(I8975)
--	g3970 = NOT(I5236)
--	g1594 = NOT(g1143)
--	g4854 = NOT(I6570)
--	g6538 = NOT(g6469)
--	g1972 = NOT(I3083)
--	I5923 = NOT(g4299)
--	g6509 = NOT(I8447)
--	g1806 = NOT(I2857)
--	g5877 = NOT(I7643)
--	g5590 = NOT(I7352)
--	g1943 = NOT(I3050)
--	I3708 = NOT(g1946)
--	g3224 = NOT(I4471)
--	g2086 = NOT(I3198)
--	g2728 = NOT(I3890)
--	I3031 = NOT(g1504)
--	I4468 = NOT(g2583)
--	g3320 = NOT(g3067)
--	g6067 = NOT(g5788)
--	g1887 = NOT(I2982)
--	I3431 = NOT(g1275)
--	g1122 = NOT(I2162)
--	g6418 = NOT(I8264)
--	g6467 = NOT(I8335)
--	g1322 = NOT(I2321)
--	g4520 = NOT(I6072)
--	g1934 = NOT(I3037)
--	I2041 = NOT(g680)
--	I3376 = NOT(g1328)
--	g4431 = NOT(I5938)
--	g4252 = NOT(I5708)
--	I1874 = NOT(g282)
--	I3405 = NOT(g1321)
--	g3906 = NOT(g3575)
--	g2470 = NOT(I3602)
--	g3789 = NOT(g3388)
--	g5064 = NOT(I6706)
--	g2025 = NOT(g1276)
--	g6493 = NOT(g6375)
--	g5899 = NOT(g5753)
--	I6775 = NOT(g4790)
--	g4376 = NOT(I5843)
--	g4405 = NOT(I5910)
--	g3771 = NOT(I4964)
--	I5825 = NOT(g3914)
--	g872 = NOT(g143)
--	g1550 = NOT(g996)
--	I6060 = NOT(g4380)
--	g4286 = NOT(I5743)
--	g4765 = NOT(I6403)
--	I1880 = NOT(g276)
--	I4198 = NOT(g2276)
--	g3299 = NOT(g3049)
--	g5563 = NOT(g5381)
--	I4398 = NOT(g2086)
--	g4911 = NOT(I6615)
--	I3733 = NOT(g2031)
--	g6700 = NOT(I8818)
--	g1395 = NOT(I2428)
--	g1891 = NOT(I2986)
--	g1337 = NOT(I2364)
--	g5237 = NOT(g5083)
--	g3892 = NOT(g3575)
--	g2678 = NOT(g2312)
--	I3225 = NOT(g1813)
--	g6421 = NOT(I8273)
--	I2890 = NOT(g1123)
--	I8585 = NOT(g6442)
--	I5594 = NOT(g3821)
--	g4270 = NOT(I5723)
--	I7372 = NOT(g5493)
--	g1807 = NOT(I2860)
--	g4225 = NOT(g4059)
--	g2682 = NOT(I3826)
--	g2766 = NOT(g2361)
--	I6995 = NOT(g5220)
--	I1935 = NOT(g666)
--	g2087 = NOT(g1352)
--	g2105 = NOT(g1375)
--	I6937 = NOT(g5124)
--	I7143 = NOT(g5323)
--	I8441 = NOT(g6419)
--	g2801 = NOT(I4003)
--	I2411 = NOT(g736)
--	g5089 = NOT(I6723)
--	g5489 = NOT(I7187)
--	I5065 = NOT(g3714)
--	g4124 = NOT(I5454)
--	g714 = NOT(g131)
--	I3540 = NOT(g1670)
--	g4980 = NOT(g4678)
--	g2748 = NOT(I3923)
--	g6562 = NOT(I8570)
--	I3206 = NOT(g1823)
--	g5705 = NOT(I7466)
--	I2992 = NOT(g1741)
--	g3478 = NOT(g2695)
--	g1142 = NOT(I2169)
--	g2755 = NOT(g2350)
--	I4258 = NOT(g2169)
--	g5242 = NOT(g5085)
--	I8168 = NOT(g6170)
--	g6723 = NOT(I8863)
--	g1255 = NOT(g161)
--	I5033 = NOT(g3527)
--	g6101 = NOT(I7799)
--	g6817 = NOT(I8988)
--	I5433 = NOT(g3728)
--	g4206 = NOT(I5626)
--	g3082 = NOT(I4315)
--	g3482 = NOT(g2713)
--	I8531 = NOT(g6444)
--	g1692 = NOT(I2696)
--	g6605 = NOT(I8681)
--	g1726 = NOT(I2728)
--	g3876 = NOT(I5109)
--	g2173 = NOT(I3310)
--	I6942 = NOT(g5124)
--	g2091 = NOT(g1355)
--	I5496 = NOT(g3839)
--	g1960 = NOT(I3071)
--	g2491 = NOT(I3620)
--	g5150 = NOT(I6816)
--	g4849 = NOT(I6555)
--	g2169 = NOT(I3298)
--	g2283 = NOT(I3428)
--	I7113 = NOT(g5295)
--	I8411 = NOT(g6415)
--	I5337 = NOT(g3564)
--	I5913 = NOT(g3751)
--	g2602 = NOT(g2061)
--	g6585 = NOT(I8623)
--	g2007 = NOT(g1411)
--	g5773 = NOT(I7514)
--	g4399 = NOT(I5896)
--	I3797 = NOT(g2125)
--	I6250 = NOT(g4514)
--	g2059 = NOT(g1402)
--	g2920 = NOT(g1947)
--	I4170 = NOT(g2157)
--	g4781 = NOT(I6437)
--	g6441 = NOT(I8309)
--	I8074 = NOT(g6118)
--	g2767 = NOT(g2364)
--	g4900 = NOT(I6607)
--	g1783 = NOT(I2831)
--	g3110 = NOT(I4358)
--	I4821 = NOT(g2877)
--	I2688 = NOT(g1030)
--	I2857 = NOT(g1161)
--	g2535 = NOT(I3653)
--	I3291 = NOT(g1714)
--	g1979 = NOT(I3090)
--	g1112 = NOT(g336)
--	g1267 = NOT(g843)
--	I7494 = NOT(g5691)
--	g4510 = NOT(I6042)
--	I3144 = NOT(g1319)
--	g5918 = NOT(I7686)
--	g1001 = NOT(I2044)
--	g3002 = NOT(g2215)
--	I8573 = NOT(g6435)
--	I8863 = NOT(g6700)
--	I4483 = NOT(g3082)
--	g1293 = NOT(I2284)
--	g6368 = NOT(I8168)
--	g4144 = NOT(I5514)
--	I8713 = NOT(g6522)
--	I7593 = NOT(g5605)
--	I3819 = NOT(g2044)
--	g3236 = NOT(I4507)
--	g1329 = NOT(I2340)
--	I3694 = NOT(g1811)
--	g1761 = NOT(I2788)
--	g857 = NOT(g170)
--	g5993 = NOT(g5872)
--	g6531 = NOT(I8509)
--	I5081 = NOT(g3589)
--	I3923 = NOT(g2581)
--	I4306 = NOT(g1898)
--	I2760 = NOT(g1193)
--	g2664 = NOT(I3808)
--	I5481 = NOT(g3866)
--	I3488 = NOT(g1295)
--	g6743 = NOT(I8907)
--	g6890 = NOT(I9137)
--	g1830 = NOT(I2904)
--	I5692 = NOT(g3942)
--	I7264 = NOT(g5458)
--	g4852 = NOT(I6564)
--	g6505 = NOT(I8435)
--	I3215 = NOT(g1820)
--	g1221 = NOT(g46)
--	g6411 = NOT(I8243)
--	g6734 = NOT(I8894)
--	g3222 = NOT(I4465)
--	I3886 = NOT(g2215)
--	I8857 = NOT(g6698)
--	g1703 = NOT(I2707)
--	I2608 = NOT(g1143)
--	g5921 = NOT(I7695)
--	g4215 = NOT(I5637)
--	I2779 = NOT(g1038)
--	I7996 = NOT(g6137)
--	g6074 = NOT(g5794)
--	g3064 = NOT(I4291)
--	g3785 = NOT(g3466)
--	g1624 = NOT(I2581)
--	g1953 = NOT(I3062)
--	I4003 = NOT(g2284)
--	g5895 = NOT(g5742)
--	g4114 = NOT(I5424)
--	g4314 = NOT(g4080)
--	I2588 = NOT(g1193)
--	I3650 = NOT(g1650)
--	g6080 = NOT(g5805)
--	I2361 = NOT(g1075)
--	g6573 = NOT(I8603)
--	I4391 = NOT(g2275)
--	g6713 = NOT(g6679)
--	I3408 = NOT(g1644)
--	g3237 = NOT(I4510)
--	I7835 = NOT(g5926)
--	I2327 = NOT(g1222)
--	g6569 = NOT(I8591)
--	g2030 = NOT(I3137)
--	g5788 = NOT(I7587)
--	g2430 = NOT(I3563)
--	I2346 = NOT(g1193)
--	g4136 = NOT(I5490)
--	I8183 = NOT(g6176)
--	I4223 = NOT(g2176)
--	I8220 = NOT(g6322)
--	g4768 = NOT(I6410)
--	g1848 = NOT(I2946)
--	I9140 = NOT(g6888)
--	g2826 = NOT(g2481)
--	g1699 = NOT(I2703)
--	g1747 = NOT(I2760)
--	g838 = NOT(g564)
--	I6075 = NOT(g4386)
--	I2696 = NOT(g1156)
--	I4757 = NOT(g2861)
--	I7799 = NOT(g5918)
--	I3065 = NOT(g1426)
--	g3557 = NOT(g2598)
--	I5746 = NOT(g4022)
--	g4806 = NOT(g4473)
--	g5392 = NOT(I7058)
--	I8423 = NOT(g6423)
--	I9035 = NOT(g6812)
--	I6949 = NOT(g5050)
--	g4943 = NOT(I6635)
--	I3465 = NOT(g1724)
--	I3322 = NOT(g1333)
--	I9082 = NOT(g6849)
--	g3705 = NOT(g3014)
--	I8588 = NOT(g6443)
--	I4522 = NOT(g2801)
--	I2753 = NOT(g1174)
--	g842 = NOT(g571)
--	I6292 = NOT(g4434)
--	I4315 = NOT(g2245)
--	g3242 = NOT(g3083)
--	g4122 = NOT(I5448)
--	g4228 = NOT(I5668)
--	g4322 = NOT(I5793)
--	I2240 = NOT(g19)
--	I1938 = NOT(g332)
--	g2108 = NOT(I3232)
--	g2609 = NOT(I3749)
--	I6646 = NOT(g4687)
--	g2308 = NOT(I3452)
--	I8665 = NOT(g6527)
--	I8051 = NOT(g6108)
--	I7153 = NOT(g5358)
--	g2883 = NOT(g1954)
--	I6084 = NOT(g4391)
--	I6039 = NOT(g4182)
--	I5068 = NOT(g3571)
--	I3096 = NOT(g1439)
--	g1644 = NOT(I2611)
--	I3496 = NOT(g1326)
--	g715 = NOT(g135)
--	I3550 = NOT(g1295)
--	I7802 = NOT(g5920)
--	g5708 = NOT(I7469)
--	g1119 = NOT(I2159)
--	g1319 = NOT(I2312)
--	g2066 = NOT(g1341)
--	g3150 = NOT(I4391)
--	g5219 = NOT(I6885)
--	I3137 = NOT(g1315)
--	I8103 = NOT(g6134)
--	I3395 = NOT(g1286)
--	I3337 = NOT(g1338)
--	g4496 = NOT(I6008)
--	g1352 = NOT(I2391)
--	I9110 = NOT(g6864)
--	g1577 = NOT(g1001)
--	g4550 = NOT(I6126)
--	g3773 = NOT(g3466)
--	g4845 = NOT(I6543)
--	I4537 = NOT(g2877)
--	I8696 = NOT(g6569)
--	g2165 = NOT(I3294)
--	g5958 = NOT(g5818)
--	I2147 = NOT(g6)
--	g6608 = NOT(I8690)
--	g4195 = NOT(I5615)
--	g4137 = NOT(I5493)
--	g830 = NOT(g338)
--	I5716 = NOT(g3942)
--	g3769 = NOT(g3622)
--	I9002 = NOT(g6802)
--	g2827 = NOT(g2485)
--	I6952 = NOT(g5124)
--	I5848 = NOT(g3856)
--	g3836 = NOT(I5033)
--	g3212 = NOT(I4455)
--	g6423 = NOT(I8279)
--	I4243 = NOT(g1853)
--	g2333 = NOT(I3485)
--	I8240 = NOT(g6287)
--	g1975 = NOT(I3086)
--	I5699 = NOT(g3844)
--	g4807 = NOT(g4473)
--	I9236 = NOT(g6939)
--	g3967 = NOT(I5223)
--	I6561 = NOT(g4707)
--	g6588 = NOT(I8632)
--	I4935 = NOT(g3369)
--	I2596 = NOT(g985)
--	g6161 = NOT(g5926)
--	g1274 = NOT(g856)
--	g6361 = NOT(I8147)
--	g1426 = NOT(I2445)
--	g2196 = NOT(I3337)
--	I7600 = NOT(g5605)
--	g2803 = NOT(g2440)
--	I6004 = NOT(g4159)
--	g3229 = NOT(I4486)
--	I6986 = NOT(g5230)
--	g6051 = NOT(g5824)
--	g5270 = NOT(I6927)
--	g804 = NOT(I1871)
--	I3255 = NOT(g1650)
--	g2538 = NOT(I3656)
--	g1325 = NOT(I2330)
--	g1821 = NOT(I2883)
--	g844 = NOT(g578)
--	I3481 = NOT(g1461)
--	I8034 = NOT(g6242)
--	g4142 = NOT(I5508)
--	g4248 = NOT(I5696)
--	g2509 = NOT(I3635)
--	I6546 = NOT(g4692)
--	I3726 = NOT(g2030)
--	g4815 = NOT(I6495)
--	I5644 = NOT(g4059)
--	I8147 = NOT(g6182)
--	g5124 = NOT(I6780)
--	g6103 = NOT(I7805)
--	I5119 = NOT(g3714)
--	g4692 = NOT(I6280)
--	g2467 = NOT(I3599)
--	I8681 = NOT(g6566)
--	g4726 = NOT(I6352)
--	g5469 = NOT(I7153)
--	g4154 = NOT(I5548)
--	I2601 = NOT(g1161)
--	g6696 = NOT(I8806)
--	g1636 = NOT(I2593)
--	g3921 = NOT(g3512)
--	g5540 = NOT(I7284)
--	I5577 = NOT(g4022)
--	g1106 = NOT(I2128)
--	g6732 = NOT(I8888)
--	g853 = NOT(g642)
--	g2256 = NOT(I3395)
--	g1790 = NOT(I2842)
--	I2922 = NOT(g1774)
--	g6508 = NOT(I8444)
--	I5893 = NOT(g3747)
--	I3979 = NOT(g1836)
--	I2581 = NOT(g946)
--	I3112 = NOT(g1439)
--	g1461 = NOT(I2460)
--	g3462 = NOT(g2679)
--	g1756 = NOT(I2779)
--	g2381 = NOT(I3528)
--	I6789 = NOT(g4871)
--	g4783 = NOT(I6441)
--	g6043 = NOT(g5824)
--	I7871 = NOT(g6097)
--	I2460 = NOT(g952)
--	I3001 = NOT(g1267)
--	g4112 = NOT(I5418)
--	g4218 = NOT(I5640)
--	g2197 = NOT(I3340)
--	g4267 = NOT(I5720)
--	I4166 = NOT(g2390)
--	g2397 = NOT(I3540)
--	I4366 = NOT(g2244)
--	g5199 = NOT(I6867)
--	g5399 = NOT(I7065)
--	g1046 = NOT(g489)
--	I3761 = NOT(g2505)
--	g3788 = NOT(g3466)
--	g6034 = NOT(g5824)
--	g6434 = NOT(I8300)
--	g6565 = NOT(I8579)
--	I6299 = NOT(g4438)
--	g4293 = NOT(I5750)
--	g4129 = NOT(I5469)
--	g5797 = NOT(I7596)
--	I3830 = NOT(g2179)
--	I2995 = NOT(g1742)
--	g6147 = NOT(I7871)
--	g1345 = NOT(I2382)
--	g1841 = NOT(I2929)
--	g6347 = NOT(I8103)
--	I1832 = NOT(g143)
--	I2479 = NOT(g1049)
--	I7339 = NOT(g5540)
--	g1191 = NOT(g38)
--	I2668 = NOT(g1011)
--	g1391 = NOT(I2424)
--	I1853 = NOT(g211)
--	g3192 = NOT(I4429)
--	g6533 = NOT(I8515)
--	g3085 = NOT(I4324)
--	I3746 = NOT(g2035)
--	I7838 = NOT(g5947)
--	g4727 = NOT(I6355)
--	I4964 = NOT(g3673)
--	g3485 = NOT(g2986)
--	I2190 = NOT(g297)
--	g1695 = NOT(g1106)
--	g6697 = NOT(I8809)
--	g1637 = NOT(I2596)
--	g1107 = NOT(I2131)
--	g2631 = NOT(I3773)
--	g6596 = NOT(I8656)
--	g3854 = NOT(I5071)
--	I5106 = NOT(g3247)
--	I8597 = NOT(g6445)
--	g2817 = NOT(g2461)
--	I6244 = NOT(g4519)
--	I7077 = NOT(g5281)
--	g4703 = NOT(I6299)
--	g6413 = NOT(I8249)
--	I5790 = NOT(g3803)
--	g1858 = NOT(I2964)
--	I6078 = NOT(g4387)
--	I6340 = NOT(g4561)
--	I7643 = NOT(g5752)
--	I3068 = NOT(g1439)
--	g5923 = NOT(I7701)
--	I9038 = NOT(g6833)
--	I3468 = NOT(g1802)
--	I4279 = NOT(g2230)
--	I5756 = NOT(g3922)
--	g6820 = NOT(I8997)
--	g4624 = NOT(g4265)
--	I6959 = NOT(g5089)
--	I5622 = NOT(g3914)
--	g3219 = NOT(I4462)
--	I5027 = NOT(g3267)
--	I4318 = NOT(g2171)
--	I7634 = NOT(g5727)
--	I5427 = NOT(g3726)
--	g3031 = NOT(I4246)
--	g1115 = NOT(g40)
--	g6117 = NOT(g5880)
--	g1315 = NOT(I2296)
--	g1811 = NOT(I2864)
--	g1642 = NOT(g809)
--	I8479 = NOT(g6482)
--	g2585 = NOT(I3708)
--	I7104 = NOT(g5273)
--	I5904 = NOT(g3749)
--	I8668 = NOT(g6530)
--	g5886 = NOT(g5753)
--	I8840 = NOT(g6657)
--	g2041 = NOT(I3152)
--	g6601 = NOT(I8671)
--	I5514 = NOT(g3882)
--	I3349 = NOT(g1334)
--	I2053 = NOT(g684)
--	g5114 = NOT(I6756)
--	I5403 = NOT(g3970)
--	g5314 = NOT(I6972)
--	I2453 = NOT(g952)
--	g1654 = NOT(g878)
--	g4716 = NOT(I6330)
--	g4149 = NOT(I5529)
--	g6922 = NOT(I9203)
--	I8156 = NOT(g6167)
--	I3198 = NOT(g1819)
--	I3855 = NOT(g2550)
--	I5391 = NOT(g3975)
--	g3911 = NOT(I5148)
--	g6581 = NOT(g6493)
--	g4848 = NOT(I6552)
--	I5637 = NOT(g3914)
--	g1880 = NOT(g1603)
--	g4198 = NOT(I5618)
--	g4699 = NOT(I6289)
--	g6597 = NOT(I8659)
--	g4855 = NOT(I6573)
--	g4398 = NOT(I5893)
--	g2772 = NOT(I3961)
--	I4321 = NOT(g1917)
--	g5136 = NOT(I6786)
--	g3225 = NOT(I4474)
--	I5223 = NOT(g3537)
--	g2743 = NOT(g2333)
--	g6784 = NOT(I8940)
--	g2890 = NOT(g1875)
--	g3073 = NOT(I4300)
--	g1978 = NOT(g1387)
--	g3796 = NOT(g3388)
--	g1017 = NOT(I2053)
--	I2929 = NOT(g1659)
--	g798 = NOT(I1868)
--	g2505 = NOT(I3629)
--	I3644 = NOT(g1685)
--	g3124 = NOT(I4371)
--	g1935 = NOT(I3040)
--	g3980 = NOT(I5264)
--	g2856 = NOT(g2010)
--	g2734 = NOT(I3902)
--	I8432 = NOT(g6411)
--	I3319 = NOT(g1636)
--	g1982 = NOT(I3093)
--	g754 = NOT(I1850)
--	g4524 = NOT(I6084)
--	g836 = NOT(g349)
--	I8453 = NOT(g6414)
--	g6840 = NOT(I9041)
--	I4519 = NOT(g2788)
--	g4644 = NOT(I6231)
--	I3152 = NOT(g1322)
--	I3258 = NOT(g1760)
--	g3540 = NOT(I4762)
--	I3352 = NOT(g1285)
--	g1328 = NOT(I2337)
--	g5887 = NOT(g5742)
--	g4119 = NOT(I5439)
--	g5465 = NOT(I7143)
--	g1542 = NOT(g878)
--	g1330 = NOT(I2343)
--	g3177 = NOT(I4414)
--	I3717 = NOT(g2154)
--	g5230 = NOT(I6895)
--	g845 = NOT(g582)
--	g4152 = NOT(I5542)
--	g6501 = NOT(I8423)
--	g4577 = NOT(g4202)
--	g4717 = NOT(g4465)
--	g5433 = NOT(I7107)
--	I5654 = NOT(g3742)
--	I6930 = NOT(g5017)
--	g2863 = NOT(g2296)
--	I6464 = NOT(g4562)
--	I3599 = NOT(g1484)
--	g2713 = NOT(I3868)
--	I3274 = NOT(g1773)
--	g4386 = NOT(I5865)
--	g3199 = NOT(g1861)
--	g5550 = NOT(g5331)
--	I3614 = NOT(g1295)
--	g3781 = NOT(I4976)
--	I3370 = NOT(g1805)
--	g5137 = NOT(I6789)
--	g5395 = NOT(I7061)
--	g5891 = NOT(g5731)
--	g3898 = NOT(g3575)
--	g3900 = NOT(g3575)
--	I3325 = NOT(g1340)
--	g4426 = NOT(I5929)
--	I2735 = NOT(g1118)
--	g3797 = NOT(g3388)
--	I9085 = NOT(g6850)
--	g1902 = NOT(I3001)
--	g6163 = NOT(g5926)
--	g4614 = NOT(g4308)
--	I2782 = NOT(g1177)
--	I7679 = NOT(g5726)
--	g6363 = NOT(I8153)
--	g4370 = NOT(I5831)
--	I8626 = NOT(g6543)
--	g3510 = NOT(g2709)
--	I5612 = NOT(g3910)
--	g6032 = NOT(g5770)
--	g4125 = NOT(I5457)
--	g2688 = NOT(I3836)
--	g2857 = NOT(I4059)
--	g3291 = NOT(g3037)
--	I3083 = NOT(g1426)
--	g2976 = NOT(g2197)
--	g1823 = NOT(I2887)
--	I2949 = NOT(g1263)
--	g1366 = NOT(I2402)
--	g5266 = NOT(I6923)
--	I2627 = NOT(g1053)
--	g1056 = NOT(g89)
--	g6568 = NOT(I8588)
--	I5328 = NOT(g3502)
--	g1529 = NOT(g1076)
--	I7805 = NOT(g5923)
--	I5542 = NOT(g3984)
--	I2998 = NOT(g1257)
--	g1649 = NOT(g985)
--	g1348 = NOT(I2385)
--	g3259 = NOT(g2996)
--	I4358 = NOT(g2525)
--	g5248 = NOT(g4911)
--	g4636 = NOT(g4286)
--	g1355 = NOT(I2394)
--	g4106 = NOT(I5400)
--	g5255 = NOT(g4933)
--	g3852 = NOT(I5065)
--	I9031 = NOT(g6809)
--	g2760 = NOT(I3942)
--	g3488 = NOT(g2728)
--	I8894 = NOT(g6709)
--	g4790 = NOT(I6456)
--	g5692 = NOT(I7451)
--	I4587 = NOT(g2962)
--	g5097 = NOT(I6733)
--	g5726 = NOT(I7487)
--	g4187 = NOT(I5591)
--	I9176 = NOT(g6881)
--	g4387 = NOT(I5868)
--	I9005 = NOT(g6817)
--	g1063 = NOT(g675)
--	g3886 = NOT(g3346)
--	g4622 = NOT(g4252)
--	g2608 = NOT(I3746)
--	I2919 = NOT(g1787)
--	g2779 = NOT(g2394)
--	g4904 = NOT(g4812)
--	g3114 = NOT(I4362)
--	I2952 = NOT(g1594)
--	g1279 = NOT(g848)
--	g4514 = NOT(I6054)
--	g1720 = NOT(g1111)
--	g4003 = NOT(g3441)
--	g1118 = NOT(g36)
--	I3391 = NOT(g1646)
--	g1318 = NOT(I2309)
--	g4403 = NOT(I5904)
--	I5490 = NOT(g3832)
--	g5112 = NOT(I6750)
--	g2588 = NOT(I3717)
--	g4145 = NOT(I5517)
--	g4841 = NOT(I6531)
--	I8603 = NOT(g6449)
--	g2361 = NOT(I3513)
--	I6769 = NOT(g4786)
--	g4763 = NOT(I6397)
--	g4191 = NOT(I5603)
--	g4391 = NOT(I5876)
--	I5056 = NOT(g3567)
--	I2986 = NOT(g1504)
--	I3307 = NOT(g1339)
--	g1193 = NOT(I2204)
--	I5529 = NOT(g3854)
--	I4420 = NOT(g2096)
--	I5148 = NOT(g3450)
--	g3136 = NOT(I4382)
--	g2327 = NOT(I3481)
--	I6918 = NOT(g5124)
--	I4507 = NOT(g2739)
--	g5329 = NOT(I6989)
--	g1549 = NOT(g878)
--	g4107 = NOT(I5403)
--	I7042 = NOT(g5310)
--	g947 = NOT(g74)
--	g6894 = NOT(I9149)
--	g1834 = NOT(I2916)
--	I4794 = NOT(g2814)
--	g4307 = NOT(I5774)
--	I5851 = NOT(g3739)
--	g4536 = NOT(I6118)
--	I3858 = NOT(g2197)
--	I8702 = NOT(g6572)
--	g2346 = NOT(I3496)
--	g6735 = NOT(I8897)
--	I3016 = NOT(g1754)
--	I2970 = NOT(g1504)
--	g5727 = NOT(I7490)
--	I7164 = NOT(g5433)
--	g2103 = NOT(I3225)
--	g858 = NOT(g301)
--	I2925 = NOT(g1762)
--	g4858 = NOT(I6582)
--	I3522 = NOT(g1664)
--	g4016 = NOT(I5320)
--	I3115 = NOT(g1519)
--	I3251 = NOT(g1471)
--	I3811 = NOT(g2145)
--	I8276 = NOT(g6303)
--	g1321 = NOT(I2318)
--	I3047 = NOT(g1426)
--	g1670 = NOT(I2648)
--	g3228 = NOT(I4483)
--	g3465 = NOT(g2986)
--	g3322 = NOT(g3070)
--	I5463 = NOT(g3783)
--	g3230 = NOT(I4489)
--	g4522 = NOT(I6078)
--	g4115 = NOT(I5427)
--	g2753 = NOT(I3927)
--	g4251 = NOT(I5705)
--	g1232 = NOT(I2228)
--	I4300 = NOT(g2234)
--	g6526 = NOT(I8494)
--	g1813 = NOT(I2870)
--	I8527 = NOT(g6440)
--	I8647 = NOT(g6528)
--	I2617 = NOT(g1193)
--	I5720 = NOT(g4022)
--	g2043 = NOT(I3158)
--	g6039 = NOT(g5824)
--	I8764 = NOT(g6564)
--	g2443 = NOT(I3578)
--	g6484 = NOT(g6361)
--	g3096 = NOT(I4343)
--	g5468 = NOT(I7150)
--	g1519 = NOT(I2491)
--	g1740 = NOT(g1116)
--	I7012 = NOT(g5316)
--	g6850 = NOT(I9077)
--	I6895 = NOT(g5010)
--	I1835 = NOT(g205)
--	g3845 = NOT(I5050)
--	I5843 = NOT(g3851)
--	g2316 = NOT(I3468)
--	I3537 = NOT(g1305)
--	I8503 = NOT(g6434)
--	g1552 = NOT(g1030)
--	I5457 = NOT(g3766)
--	g2565 = NOT(I3675)
--	g6583 = NOT(I8617)
--	g850 = NOT(g602)
--	g5576 = NOT(g5415)
--	g4537 = NOT(g4410)
--	I7029 = NOT(g5149)
--	g2347 = NOT(I3499)
--	I5686 = NOT(g3942)
--	I4123 = NOT(g2043)
--	g3807 = NOT(I5006)
--	g1586 = NOT(g1052)
--	g3859 = NOT(I5078)
--	g6276 = NOT(I7960)
--	g4612 = NOT(g4320)
--	g2914 = NOT(g1928)
--	g6616 = NOT(I8710)
--	I3629 = NOT(g1759)
--	g6561 = NOT(I8567)
--	I3328 = NOT(g1273)
--	I2738 = NOT(g1236)
--	I8617 = NOT(g6539)
--	g1341 = NOT(I2376)
--	g2413 = NOT(I3553)
--	I4351 = NOT(g2233)
--	g3342 = NOT(g3086)
--	g4128 = NOT(I5466)
--	g1710 = NOT(g1109)
--	g4629 = NOT(g4276)
--	I6485 = NOT(g4603)
--	g6527 = NOT(I8497)
--	g6404 = NOT(I8226)
--	g4328 = NOT(g4092)
--	I2140 = NOT(g28)
--	g1645 = NOT(I2614)
--	I2340 = NOT(g1142)
--	g4130 = NOT(I5472)
--	I5938 = NOT(g4351)
--	I7963 = NOT(g6276)
--	I3800 = NOT(g2145)
--	g3481 = NOT(g2612)
--	I2907 = NOT(g1498)
--	g2820 = NOT(g2470)
--	g2936 = NOT(g2026)
--	g5524 = NOT(I7264)
--	g6503 = NOT(I8429)
--	g3354 = NOT(g3096)
--	I4410 = NOT(g2088)
--	I7808 = NOT(g5919)
--	g2117 = NOT(I3244)
--	g3960 = NOT(I5204)
--	g2317 = NOT(I3471)
--	g5119 = NOT(I6769)
--	g6925 = NOT(I9208)
--	I7707 = NOT(g5701)
--	I5606 = NOT(g3821)
--	g1659 = NOT(I2638)
--	g1358 = NOT(g1119)
--	g5352 = NOT(I7002)
--	g5577 = NOT(g5420)
--	g4213 = NOT(I5633)
--	g5717 = NOT(I7478)
--	I3902 = NOT(g2576)
--	g6120 = NOT(I7832)
--	g2922 = NOT(g1960)
--	g1587 = NOT(g1123)
--	I6812 = NOT(g5110)
--	I8991 = NOT(g6788)
--	g3783 = NOT(I4980)
--	g1111 = NOT(I2143)
--	I3090 = NOT(g1504)
--	I9008 = NOT(g6818)
--	g5893 = NOT(g5753)
--	g1275 = NOT(g842)
--	g6277 = NOT(I7963)
--	g2581 = NOT(I3694)
--	I3823 = NOT(g2125)
--	g3267 = NOT(g3030)
--	I4667 = NOT(g2908)
--	g3312 = NOT(I4587)
--	I7865 = NOT(g6095)
--	I4343 = NOT(g2525)
--	g2060 = NOT(g1369)
--	g6617 = NOT(I8713)
--	g6906 = NOT(I9185)
--	g5975 = NOT(g5821)
--	g4512 = NOT(I6048)
--	I4282 = NOT(g2525)
--	g2460 = NOT(I3590)
--	I7604 = NOT(g5605)
--	I8907 = NOT(g6702)
--	I3056 = NOT(g1519)
--	g3001 = NOT(I4198)
--	g1174 = NOT(g37)
--	g4823 = NOT(I6507)
--	I2663 = NOT(g1006)
--	g4166 = NOT(I5568)
--	g6516 = NOT(g6409)
--	g5274 = NOT(I6933)
--	I8435 = NOT(g6413)
--	I3148 = NOT(g1595)
--	I8690 = NOT(g6571)
--	g1985 = NOT(I3096)
--	I4334 = NOT(g2256)
--	I8482 = NOT(g6461)
--	g2739 = NOT(I3906)
--	g3761 = NOT(g3605)
--	I3155 = NOT(g1612)
--	I3355 = NOT(g1608)
--	I2402 = NOT(g774)
--	g4529 = NOT(I6099)
--	g1284 = NOT(g851)
--	g4148 = NOT(I5526)
--	I6733 = NOT(g4773)
--	I8656 = NOT(g6532)
--	g3830 = NOT(I5019)
--	I9122 = NOT(g6864)
--	g2079 = NOT(g1348)
--	g4155 = NOT(I5551)
--	g4851 = NOT(I6561)
--	g6892 = NOT(I9143)
--	g1832 = NOT(I2910)
--	I9230 = NOT(g6936)
--	g1853 = NOT(I2955)
--	g2840 = NOT(g2538)
--	I2877 = NOT(g1123)
--	I5879 = NOT(g3745)
--	g5544 = NOT(g5331)
--	g2390 = NOT(I3531)
--	I6324 = NOT(g4450)
--	g1559 = NOT(g965)
--	I6069 = NOT(g4213)
--	I8110 = NOT(g6143)
--	g4463 = NOT(g4364)
--	g943 = NOT(g496)
--	g1931 = NOT(I3034)
--	g6709 = NOT(I8837)
--	g3932 = NOT(I5169)
--	I6540 = NOT(g4714)
--	I3720 = NOT(g2155)
--	g6078 = NOT(g5801)
--	I1871 = NOT(g281)
--	I6377 = NOT(g4569)
--	g5061 = NOT(I6701)
--	g6478 = NOT(I8342)
--	I2464 = NOT(g850)
--	I3367 = NOT(g1283)
--	g5387 = NOT(I7051)
--	I9137 = NOT(g6864)
--	g1905 = NOT(I3004)
--	I8002 = NOT(g6110)
--	g866 = NOT(g314)
--	I2785 = NOT(g1222)
--	I7086 = NOT(g5281)
--	I5615 = NOT(g3914)
--	g6035 = NOT(g5824)
--	g4720 = NOT(I6340)
--	I3843 = NOT(g2145)
--	g4118 = NOT(I5436)
--	g4619 = NOT(g4248)
--	g6517 = NOT(I8467)
--	g1204 = NOT(g39)
--	g3677 = NOT(g3140)
--	g6876 = NOT(I9095)
--	g4843 = NOT(I6537)
--	g3866 = NOT(I5091)
--	g2954 = NOT(g2381)
--	I4593 = NOT(g2966)
--	g5046 = NOT(I6680)
--	g2163 = NOT(I3288)
--	g6656 = NOT(I8764)
--	g4193 = NOT(I5609)
--	I2237 = NOT(g465)
--	g2032 = NOT(g1749)
--	g4393 = NOT(I5882)
--	I5545 = NOT(g3814)
--	g5403 = NOT(I7069)
--	I1838 = NOT(g206)
--	g3848 = NOT(I5059)
--	I5591 = NOT(g3821)
--	I4264 = NOT(g2212)
--	I2394 = NOT(g719)
--	g5391 = NOT(I7055)
--	g2568 = NOT(I3678)
--	I2731 = NOT(g1117)
--	I4050 = NOT(g2059)
--	g3241 = NOT(I4522)
--	g2912 = NOT(g2001)
--	g4121 = NOT(I5445)
--	g1969 = NOT(I3080)
--	I3232 = NOT(g1782)
--	g4321 = NOT(I5790)
--	g5307 = NOT(I6959)
--	g2157 = NOT(I3278)
--	g5536 = NOT(g5467)
--	g2357 = NOT(I3509)
--	g1123 = NOT(I2165)
--	g1323 = NOT(I2324)
--	g4625 = NOT(g4267)
--	I3909 = NOT(g2044)
--	g4232 = NOT(I5674)
--	g6402 = NOT(I8220)
--	g6824 = NOT(I9005)
--	g1666 = NOT(g1088)
--	g4938 = NOT(I6630)
--	I6819 = NOT(g5019)
--	g6236 = NOT(g6070)
--	I3519 = NOT(g1305)
--	I8295 = NOT(g6295)
--	I2955 = NOT(g1729)
--	I7487 = NOT(g5684)
--	g856 = NOT(g654)
--	I6923 = NOT(g5124)
--	g1528 = NOT(g878)
--	I5204 = NOT(g3534)
--	I5630 = NOT(g3914)
--	I6488 = NOT(g4603)
--	g1351 = NOT(I2388)
--	g1648 = NOT(I2623)
--	I2814 = NOT(g1222)
--	g1875 = NOT(I2970)
--	g4519 = NOT(I6069)
--	g5115 = NOT(I6759)
--	g6590 = NOT(I8638)
--	g5251 = NOT(g5069)
--	g6877 = NOT(I9098)
--	g3258 = NOT(I4537)
--	I4777 = NOT(g2962)
--	I6701 = NOT(g4726)
--	g5315 = NOT(g5116)
--	g3867 = NOT(I5094)
--	I2150 = NOT(g10)
--	g1655 = NOT(g985)
--	g6657 = NOT(I8767)
--	g4606 = NOT(g4193)
--	I3687 = NOT(g1814)
--	I8089 = NOT(g6120)
--	I2773 = NOT(g1191)
--	g5874 = NOT(I7634)
--	g1410 = NOT(g1233)
--	I8966 = NOT(g6796)
--	I5750 = NOT(g4022)
--	I7045 = NOT(g5167)
--	I6114 = NOT(g4405)
--	g3975 = NOT(I5249)
--	I7173 = NOT(g5436)
--	g1884 = NOT(I2979)
--	I7091 = NOT(g5281)
--	g6899 = NOT(I9164)
--	I4799 = NOT(g2967)
--	I2212 = NOT(g123)
--	g929 = NOT(g49)
--	g6785 = NOT(I8943)
--	g5880 = NOT(g5824)
--	I5040 = NOT(g3271)
--	I2967 = NOT(g1682)
--	g5537 = NOT(g5385)
--	g2778 = NOT(g2391)
--	I1862 = NOT(g278)
--	I3525 = NOT(g1461)
--	g3370 = NOT(g3124)
--	g2894 = NOT(g1891)
--	I7007 = NOT(g5314)
--	g1372 = NOT(I2408)
--	g4141 = NOT(I5505)
--	g6563 = NOT(I8573)
--	I6008 = NOT(g4163)
--	I3691 = NOT(g1732)
--	g4525 = NOT(I6087)
--	g1143 = NOT(I2172)
--	g3984 = NOT(g3564)
--	I8150 = NOT(g6185)
--	g1282 = NOT(g849)
--	I8438 = NOT(g6416)
--	g3083 = NOT(I4318)
--	g1988 = NOT(I3099)
--	I4802 = NOT(g2877)
--	I6972 = NOT(g5135)
--	g3483 = NOT(g2716)
--	I7261 = NOT(g5458)
--	g6194 = NOT(I7906)
--	g1334 = NOT(I2355)
--	I3158 = NOT(g1829)
--	I3659 = NOT(g1491)
--	I3358 = NOT(g1323)
--	g5328 = NOT(I6986)
--	I1927 = NOT(g665)
--	g6489 = NOT(g6369)
--	g5542 = NOT(g5331)
--	g5330 = NOT(I6992)
--	g3306 = NOT(g3057)
--	g2998 = NOT(I4195)
--	g4158 = NOT(I5556)
--	g4659 = NOT(I6250)
--	g1555 = NOT(I2521)
--	g3790 = NOT(g3388)
--	I3587 = NOT(g1461)
--	g1792 = NOT(I2848)
--	g2603 = NOT(I3733)
--	g2039 = NOT(I3148)
--	g3187 = NOT(I4424)
--	g2484 = NOT(I3611)
--	g3387 = NOT(I4664)
--	g3461 = NOT(g2986)
--	g4587 = NOT(g4215)
--	I6033 = NOT(g4179)
--	g5554 = NOT(g5455)
--	g3622 = NOT(I4821)
--	g4111 = NOT(I5415)
--	I8229 = NOT(g6330)
--	I9149 = NOT(g6884)
--	I2620 = NOT(g1177)
--	g1113 = NOT(I2147)
--	I4492 = NOT(g3001)
--	g4615 = NOT(g4322)
--	g2583 = NOT(g1830)
--	g3904 = NOT(g3575)
--	g3200 = NOT(I4437)
--	I6096 = NOT(g4397)
--	g3046 = NOT(I4267)
--	g899 = NOT(I1924)
--	g4374 = NOT(I5837)
--	I3284 = NOT(g1702)
--	g2919 = NOT(g1937)
--	g1908 = NOT(I3007)
--	I2788 = NOT(g1236)
--	g1094 = NOT(I2122)
--	I5618 = NOT(g3821)
--	g2952 = NOT(g2381)
--	I6337 = NOT(g4455)
--	I5343 = NOT(g3599)
--	g2276 = NOT(I3425)
--	g1567 = NOT(I2537)
--	g4284 = NOT(I5739)
--	g5512 = NOT(I7254)
--	g4545 = NOT(g4416)
--	g5090 = NOT(g4741)
--	g6409 = NOT(g6285)
--	g5490 = NOT(I7190)
--	I7689 = NOT(g5708)
--	g4380 = NOT(I5851)
--	I2842 = NOT(g1177)
--	g1776 = NOT(I2821)
--	g1593 = NOT(g1054)
--	g2004 = NOT(I3115)
--	g4853 = NOT(I6567)
--	g6836 = NOT(I9031)
--	I2485 = NOT(g766)
--	I3794 = NOT(g2044)
--	g2986 = NOT(g2010)
--	g4020 = NOT(I5324)
--	g6212 = NOT(I7910)
--	I5548 = NOT(g4059)
--	g5456 = NOT(g5300)
--	g2647 = NOT(I3791)
--	I8837 = NOT(g6665)
--	g5148 = NOT(I6812)
--	g5649 = NOT(I7404)
--	g4507 = NOT(I6033)
--	g3223 = NOT(I4468)
--	I4623 = NOT(g2962)
--	I1947 = NOT(g699)
--	g2764 = NOT(g2357)
--	I8620 = NOT(g6541)
--	I8462 = NOT(g6430)
--	I9119 = NOT(g6855)
--	I2854 = NOT(g1236)
--	g4559 = NOT(g4187)
--	g5155 = NOT(g5099)
--	g5355 = NOT(I7007)
--	I9152 = NOT(g6889)
--	g3016 = NOT(I4223)
--	g6229 = NOT(g6036)
--	g1160 = NOT(I2179)
--	g5260 = NOT(g4938)
--	I6081 = NOT(g4388)
--	I4375 = NOT(g2254)
--	g6822 = NOT(g6786)
--	g1641 = NOT(I2604)
--	g3251 = NOT(I4534)
--	I6692 = NOT(g4720)
--	g1450 = NOT(I2453)
--	g5063 = NOT(g4799)
--	I7910 = NOT(g5905)
--	I8249 = NOT(g6289)
--	g4628 = NOT(g4273)
--	g4515 = NOT(I6057)
--	g2120 = NOT(I3251)
--	I4285 = NOT(g2555)
--	g2320 = NOT(I3474)
--	g4100 = NOT(I5382)
--	g1724 = NOT(I2724)
--	g3874 = NOT(I5103)
--	I2958 = NOT(g1257)
--	I5094 = NOT(g3705)
--	I2376 = NOT(g729)
--	I8485 = NOT(g6479)
--	g5720 = NOT(I7481)
--	I2405 = NOT(g1112)
--	g2906 = NOT(g1911)
--	g2789 = NOT(g2410)
--	g1878 = NOT(I2973)
--	g5118 = NOT(I6766)
--	I9170 = NOT(g6883)
--	I1917 = NOT(g48)
--	
--	g2771 = AND(g2497, g1975)
--	g6620 = AND(g6516, g6117)
--	g5193 = AND(g532, g4967)
--	I5360 = AND(g3532, g3536, g3539, g3544)
--	g5598 = AND(g5046, g5509)
--	g6249 = AND(g1332, g5892)
--	g4666 = AND(g4630, g4627)
--	g3629 = AND(g2809, g2738)
--	g3328 = AND(g2701, g1894)
--	g6085 = AND(g1161, g5731)
--	g4351 = AND(g166, g3776)
--	g4648 = AND(g4407, g79)
--	g5232 = AND(g548, g4980)
--	g2340 = AND(g1398, g1387)
--	g5938 = AND(g5114, g5791)
--	g5909 = AND(g5787, g3384)
--	g1802 = AND(g89, g1064)
--	g3554 = AND(g2941, g179)
--	g4410 = AND(g3903, g1474)
--	g6640 = AND(g1612, g6549)
--	g4172 = AND(g3930, g1366)
--	g4372 = AND(g406, g3790)
--	g3512 = AND(g2928, g1764)
--	g3490 = AND(g353, g2959)
--	g4667 = AND(g4653, g4651)
--	g3166 = AND(g2042, g1233)
--	g3366 = AND(g248, g2893)
--	g6829 = AND(g6806, g5958)
--	g3649 = AND(g3104, g2764)
--	g6911 = AND(g6904, g6902)
--	g3155 = AND(g248, g2461)
--	g3698 = AND(g2284, g2835)
--	g6270 = AND(g1726, g6062)
--	g4792 = AND(g1417, g4471)
--	g6473 = AND(g2036, g6397, g1628)
--	g4621 = AND(g3953, g4364)
--	g5158 = AND(g504, g4993)
--	g6124 = AND(g5705, g5958)
--	g6324 = AND(g3880, g6212)
--	g6469 = AND(g2121, g2032, g6394)
--	g3279 = AND(g2599, g2612)
--	g3619 = AND(g2449, g3057)
--	g3167 = AND(g1883, g921)
--	g5311 = AND(g5013, g4468)
--	g3367 = AND(g2809, g1960)
--	g3652 = AND(g2544, g3096)
--	g3843 = AND(g2856, g945, g3533)
--	g4593 = AND(g4277, g947)
--	g3686 = AND(g2256, g2819)
--	g5180 = AND(g414, g4950)
--	g5380 = AND(g188, g5264)
--	g4160 = AND(g3923, g1345)
--	g3321 = AND(g2252, g2713)
--	g2089 = AND(g1123, g1578)
--	g6245 = AND(g1329, g5889)
--	g4360 = AND(g184, g3785)
--	g3670 = AND(g2234, g2792)
--	g3625 = AND(g2619, g2320)
--	g6291 = AND(g5210, g6161)
--	g4050 = AND(I5359, I5360)
--	g5559 = AND(g5024, g5453)
--	g6144 = AND(g3183, g5997)
--	g6344 = AND(g6272, g6080)
--	g2948 = AND(g2137, g1595)
--	g6259 = AND(g1699, g6044)
--	g4179 = AND(g390, g3902)
--	g2955 = AND(g2381, g297)
--	g6088 = AND(g1143, g5753)
--	g6852 = AND(g6847, g2295)
--	g6923 = AND(g6918, g6917)
--	g5515 = AND(g590, g5364)
--	g1499 = AND(g1101, g1094)
--	g4835 = AND(g4533, g4530)
--	g3687 = AND(g2245, g2820)
--	g4271 = AND(g2121, g1749, g4004)
--	g4611 = AND(g3985, g119, g4300)
--	g3341 = AND(g2998, g2709)
--	g6650 = AND(g6580, g6235)
--	g4541 = AND(g631, g4199)
--	g3645 = AND(g2497, g3090)
--	g5123 = AND(g4670, g1936)
--	g3691 = AND(g2268, g2828)
--	g4209 = AND(g3816, g865)
--	g4353 = AND(g3989, g3332)
--	g6336 = AND(g6246, g6065)
--	g6768 = AND(g6750, g3477)
--	g4744 = AND(g3434, g4582)
--	g3659 = AND(g2672, g2361)
--	g5351 = AND(g5326, g3459)
--	g3358 = AND(g2842, g1369)
--	g5648 = AND(g4507, g5545)
--	g6934 = AND(g6932, g3605)
--	g3275 = AND(g2172, g2615)
--	g3311 = AND(g218, g2872)
--	g5410 = AND(g378, g5274)
--	g3615 = AND(g2422, g3046)
--	g2062 = AND(g1499, g1666)
--	g3374 = AND(g2809, g1969)
--	g4600 = AND(g4054, g4289)
--	g6096 = AND(g1193, g5753)
--	g1436 = AND(g834, g830)
--	g5172 = AND(g441, g4877)
--	g3180 = AND(g260, g2506)
--	g5618 = AND(g5506, g4933)
--	g5143 = AND(g157, g5099)
--	g6913 = AND(g6900, g6898)
--	g5235 = AND(g554, g4980)
--	g4580 = AND(g706, g4262)
--	g2085 = AND(g1123, g1567)
--	g6266 = AND(g1721, g6057)
--	g5555 = AND(g5014, g5442)
--	g2941 = AND(g2166, g170)
--	g6248 = AND(g465, g5894)
--	g6342 = AND(g6264, g6076)
--	g5621 = AND(g5508, g4943)
--	g3628 = AND(g2449, g3070)
--	g6255 = AND(g1335, g5895)
--	g6081 = AND(g1177, g5731)
--	g3630 = AND(g3167, g1756)
--	g6692 = AND(g6616, g6615)
--	g3300 = AND(g2232, g2682)
--	g6154 = AND(g3219, g6015)
--	g6354 = AND(g5866, g6193)
--	g4184 = AND(g3934, g2136)
--	g5494 = AND(g5443, g3455)
--	g4384 = AND(g414, g3797)
--	g4339 = AND(g3971, g3289)
--	g4838 = AND(g4648, g84)
--	g3123 = AND(g230, g2391)
--	g3323 = AND(g2253, g2716)
--	g4672 = AND(g4635, g4631)
--	g2733 = AND(g2422, g1943)
--	g3666 = AND(g3128, g2787)
--	g6129 = AND(g5717, g5975)
--	g6329 = AND(g3888, g6212)
--	g2073 = AND(g1088, g1499)
--	g5360 = AND(g4431, g5160)
--	g6828 = AND(g6803, g5958)
--	g5050 = AND(g4285, g4807)
--	g3351 = AND(g2760, g1931)
--	g6830 = AND(g6809, g5975)
--	g3648 = AND(g2722, g2343)
--	g3655 = AND(g2197, g2768)
--	g1706 = AND(g766, g719, g729)
--	g6068 = AND(g5824, g1726)
--	g4044 = AND(g410, g3388)
--	g6468 = AND(g2032, g6394, g1609)
--	g3172 = AND(g2449, g2491)
--	g3278 = AND(g2175, g2628)
--	g3372 = AND(g254, g2905)
--	g2781 = AND(g2544, g1982)
--	g3618 = AND(g3016, g2712)
--	g3667 = AND(g2245, g2789)
--	g3143 = AND(g242, g2437)
--	g3282 = AND(g131, g2863)
--	g6716 = AND(g6682, g932)
--	g6149 = AND(g3200, g5997)
--	g3693 = AND(g2256, g2830)
--	g3134 = AND(g230, g2413)
--	g3334 = AND(g236, g2883)
--	g6848 = AND(g3741, g328, g6843)
--	g5153 = AND(g492, g4904)
--	g5209 = AND(g560, g5025)
--	g5353 = AND(g5327, g3463)
--	g6241 = AND(g1325, g5887)
--	g1808 = AND(g706, g49)
--	g3113 = AND(g224, g2364)
--	g5558 = AND(g5018, g5450)
--	g6644 = AND(g6575, g6230)
--	g6152 = AND(g3212, g6015)
--	g6258 = AND(g512, g5899)
--	g4178 = AND(g3959, g2110)
--	g1575 = AND(g980, g965)
--	g4378 = AND(g410, g3792)
--	g4831 = AND(g4528, g4524)
--	g4182 = AND(g394, g3904)
--	g5492 = AND(g5441, g3452)
--	g5600 = AND(g5502, g4900)
--	g6614 = AND(g932, g6556)
--	g4947 = AND(g184, g4741)
--	g3360 = AND(g2783, g1947)
--	g6125 = AND(g5708, g5975)
--	g1419 = AND(g613, g918)
--	g3641 = AND(g2644, g2333)
--	g4873 = AND(g4838, g4173)
--	g4037 = AND(g2896, g3388)
--	g3724 = AND(g117, g3251)
--	g4495 = AND(g3913, g4292)
--	g3379 = AND(g3104, g1988)
--	g5175 = AND(g5094, g1384)
--	g3658 = AND(g3118, g2776)
--	g6061 = AND(g5824, g1711)
--	g5500 = AND(g5430, g5074)
--	g3611 = AND(g2370, g3037)
--	g2137 = AND(g760, g1638)
--	g4042 = AND(g406, g3388)
--	g5184 = AND(g453, g4877)
--	g4442 = AND(g4239, g2882)
--	g4164 = AND(g3958, g2091)
--	g2807 = AND(g2568, g2001)
--	g5424 = AND(g390, g5296)
--	g6145 = AND(g3187, g6015)
--	g2859 = AND(g2112, g1649)
--	g3997 = AND(g1250, g3425, g2849)
--	g4054 = AND(g3694, g69)
--	g6345 = AND(g6273, g6083)
--	g3132 = AND(g2306, g1206)
--	g3680 = AND(g2245, g2805)
--	g6637 = AND(g1842, g6549)
--	g3353 = AND(g3162, g2921)
--	g2142 = AND(g1793, g1777)
--	g2255 = AND(g1706, g736)
--	g6159 = AND(g3177, g6015)
--	g2081 = AND(g1094, g1546)
--	g3558 = AND(g338, g3199)
--	g5499 = AND(g5451, g3462)
--	g4389 = AND(g449, g3798)
--	g4171 = AND(g3956, g2104)
--	g6315 = AND(g3849, g6194)
--	g4371 = AND(g461, g3789)
--	g4429 = AND(g923, g4253, g2936)
--	g4787 = AND(g2937, g4628)
--	g6047 = AND(g5824, g1692)
--	g6874 = AND(g6873, g2060)
--	g2267 = AND(g1716, g791)
--	g5444 = AND(g4545, g5256, g1574)
--	g5269 = AND(g557, g5025)
--	g1407 = AND(g301, g866)
--	g4684 = AND(g4584, g1341)
--	g4791 = AND(g3936, g4636)
--	g6243 = AND(g500, g5890)
--	g6935 = AND(g6933, g3622)
--	g2746 = AND(g2473, g1954)
--	g4759 = AND(g536, g4500)
--	g6128 = AND(g5590, g5958)
--	g5414 = AND(g382, g5278)
--	g6130 = AND(g5720, g5958)
--	g5660 = AND(g4509, g5549)
--	g3375 = AND(g260, g2912)
--	g4449 = AND(g4266, g2887)
--	g3651 = AND(g3064, g2766)
--	g4865 = AND(g4776, g1849)
--	g2953 = AND(g2381, g293)
--	g2068 = AND(g1541, g1546)
--	g3285 = AND(g2195, g2653)
--	g4833 = AND(g4521, g4516)
--	g5178 = AND(g516, g4993)
--	g5679 = AND(g74, g5576)
--	g5378 = AND(g179, g5260)
--	g3339 = AND(g2734, g1914)
--	g1689 = AND(g766, g719)
--	g5182 = AND(g520, g4993)
--	g2699 = AND(g2397, g1905)
--	g2747 = AND(g2449, g1957)
--	g6090 = AND(g1161, g5742)
--	g4362 = AND(g3996, g3355)
--	g3672 = AND(g3136, g2800)
--	g4052 = AND(g418, g3388)
--	g3643 = AND(g2518, g3086)
--	g4452 = AND(g3820, g4227)
--	g6056 = AND(g5824, g1699)
--	g1826 = AND(g714, g710)
--	g6148 = AND(g3196, g6015)
--	g6348 = AND(g5869, g6211)
--	g5560 = AND(g5044, g5456)
--	g3634 = AND(g2179, g2744)
--	g6155 = AND(g2588, g5997)
--	g6851 = AND(g6846, g2293)
--	g3551 = AND(g2937, g938)
--	g3099 = AND(g218, g2350)
--	g3304 = AND(g2857, g1513)
--	g4486 = AND(g716, g4195)
--	g3499 = AND(g357, g2961)
--	g4730 = AND(g1423, g4565)
--	g5632 = AND(g4494, g5538)
--	g5095 = AND(g4794, g951)
--	g6260 = AND(g1703, g6048)
--	g4185 = AND(g398, g3906)
--	g1609 = AND(g760, g754)
--	g5495 = AND(g5444, g3456)
--	g2577 = AND(g1743, g1797, g1793, g1138)
--	g3613 = AND(g2604, g2312)
--	g6619 = AND(g6515, g6115)
--	g6318 = AND(g3865, g6212)
--	g2026 = AND(g1359, g1402, g1398, g901)
--	g5164 = AND(g437, g4877)
--	g5364 = AND(g574, g5194)
--	g5233 = AND(g551, g4980)
--	g2821 = AND(g1890, g910)
--	g3729 = AND(g327, g3441)
--	g5454 = AND(g5256, g4549)
--	g5553 = AND(g5012, g5440)
--	g6321 = AND(g3873, g6212)
--	g3660 = AND(g2568, g3110)
--	g6625 = AND(g2121, g1595, g6538)
--	g4045 = AND(g3425, g123)
--	g4445 = AND(g4235, g1854)
--	g6253 = AND(g508, g5896)
--	g4373 = AND(g4001, g3370)
--	g5189 = AND(g528, g4993)
--	g4491 = AND(g3554, g4215)
--	g6909 = AND(g6896, g6894)
--	g4169 = AND(g3966, g2099)
--	g5171 = AND(g406, g4950)
--	g4369 = AND(g3999, g3364)
--	g3679 = AND(g2245, g2803)
--	g4602 = AND(g4407, g4293)
--	g5371 = AND(g152, g5248)
--	g3378 = AND(g3136, g2932)
--	g5429 = AND(g398, g5304)
--	g4407 = AND(g4054, g74)
--	g5956 = AND(g5783, g5425)
--	g4868 = AND(g4774, g2891)
--	g5675 = AND(g64, g5574)
--	g3135 = AND(g2370, g2416)
--	g4459 = AND(g4245, g1899)
--	g3335 = AND(g230, g2884)
--	g3831 = AND(g2330, g3425)
--	g3182 = AND(g2473, g2512)
--	g3288 = AND(g2631, g2634)
--	g3382 = AND(g3136, g2934)
--	g4793 = AND(g4277, g4639)
--	g4015 = AND(g445, g3388)
--	g2107 = AND(g1583, g1543)
--	g6141 = AND(g3173, g5997)
--	g6341 = AND(g6261, g6074)
--	g6645 = AND(g6576, g6231)
--	g3632 = AND(g3043, g2743)
--	g3437 = AND(g837, g2853)
--	g3653 = AND(g2215, g2767)
--	g5201 = AND(g4859, g5084)
--	g3208 = AND(g895, g2551)
--	g3302 = AND(g212, g2867)
--	g6158 = AND(g2594, g6015)
--	g5449 = AND(g4545, g5246)
--	g5604 = AND(g5059, g5521)
--	g5098 = AND(g4021, g4837)
--	g5498 = AND(g5449, g3460)
--	g1585 = AND(g1017, g1011)
--	g6275 = AND(g1735, g6070)
--	g6311 = AND(g3837, g6194)
--	g4671 = AND(g4645, g4641)
--	g4247 = AND(g1764, g4007, g1628)
--	g3454 = AND(g2933, g1660)
--	g4826 = AND(g4209, g4463)
--	g5162 = AND(g5088, g2105)
--	g5362 = AND(g4437, g5174)
--	g3296 = AND(g3054, g2650)
--	g5419 = AND(g386, g5292)
--	g3725 = AND(g118, g3251)
--	g2935 = AND(g2291, g1788)
--	g5452 = AND(g5315, g4612)
--	g6559 = AND(g1612, g6474)
--	g5728 = AND(g5623, g3889)
--	g5486 = AND(g386, g5331)
--	g5185 = AND(g524, g4993)
--	g3171 = AND(g248, g2488)
--	g3371 = AND(g260, g2904)
--	g6628 = AND(g2138, g1612, g6540)
--	g4165 = AND(g3927, g1352)
--	g4048 = AND(g414, g3388)
--	g4448 = AND(g3815, g4225)
--	g3281 = AND(g2178, g2640)
--	g4827 = AND(g4520, g4515)
--	g4333 = AND(g3964, g3284)
--	I2566 = AND(g749, g743, g736)
--	g2166 = AND(g1633, g161)
--	g3684 = AND(g2268, g2817)
--	g4396 = AND(g422, g3801)
--	g3338 = AND(g3162, g2914)
--	g2056 = AND(g1672, g1675)
--	g5406 = AND(g374, g5270)
--	g3309 = AND(g2243, g2695)
--	g5635 = AND(g4498, g5542)
--	g5682 = AND(g84, g5578)
--	g5487 = AND(g390, g5331)
--	g6123 = AND(g5702, g5958)
--	g6323 = AND(g3877, g6194)
--	g3759 = AND(g2644, g3498)
--	g5226 = AND(g672, g5054)
--	g6151 = AND(g3209, g5997)
--	g3449 = AND(g128, g2946)
--	g6648 = AND(g6579, g6234)
--	g5173 = AND(g512, g4993)
--	g5373 = AND(g161, g5250)
--	g4181 = AND(g3939, g1381)
--	g2720 = AND(g2422, g1919)
--	g4685 = AND(g4591, g2079)
--	g5169 = AND(g5093, g1375)
--	g5369 = AND(g143, g5247)
--	g5602 = AND(g594, g5515)
--	g2834 = AND(g1263, g1257, g1270, I4040)
--	g3362 = AND(g3031, g2740)
--	g6343 = AND(g6268, g6078)
--	g2121 = AND(g1632, g754)
--	g2670 = AND(g2029, g1503)
--	g6693 = AND(g6618, g6617)
--	g1633 = AND(g716, g152)
--	g6334 = AND(g3858, g6212)
--	g3728 = AND(g326, g3441)
--	g6555 = AND(g1838, g6469)
--	g3730 = AND(g328, g3441)
--	g2909 = AND(g606, g2092)
--	g4041 = AND(g461, g3388)
--	g3425 = AND(g2296, g3208)
--	g6313 = AND(g3841, g6194)
--	g5940 = AND(g5115, g5794)
--	g4673 = AND(g4656, g4654)
--	g5188 = AND(g1043, g4894)
--	g6908 = AND(g6907, g3886)
--	g5216 = AND(g563, g5025)
--	g6094 = AND(g1177, g5753)
--	g4168 = AND(g3925, g1355)
--	g4368 = AND(g3998, g3363)
--	g5671 = AND(g54, g5572)
--	g3678 = AND(g2256, g2802)
--	g5428 = AND(g394, g5300)
--	g4058 = AND(g3424, g1246)
--	g3635 = AND(g2473, g3079)
--	g2860 = AND(g710, g2296)
--	g3682 = AND(g2772, g2430)
--	g3305 = AND(g2960, g2296)
--	g5910 = AND(g5816, g5667)
--	g3755 = AND(g2604, g3481)
--	g2659 = AND(g1686, g2296)
--	g5883 = AND(g5824, g3752)
--	g3373 = AND(g3118, g2927)
--	g5217 = AND(g4866, g5092)
--	g4863 = AND(g4777, g2874)
--	g3283 = AND(g2609, g2622)
--	g3602 = AND(g2688, g2663)
--	I2574 = AND(g804, g798, g791)
--	g5165 = AND(g508, g4993)
--	g6777 = AND(g6762, g3488)
--	g3718 = AND(g1743, g3140, g1157)
--	g3767 = AND(g2706, g3504)
--	g4688 = AND(g1474, g4568)
--	g1784 = AND(g858, g889)
--	g2853 = AND(g836, g2021)
--	g6799 = AND(g4948, g6782)
--	g2794 = AND(g2544, g1994)
--	g3203 = AND(g2497, g2565)
--	g6132 = AND(g3752, g5880)
--	g6238 = AND(g528, g5886)
--	g6153 = AND(g3216, g5997)
--	g4183 = AND(g3965, g1391)
--	g4383 = AND(g453, g3796)
--	g6558 = AND(g1842, g6474)
--	g5181 = AND(g449, g4877)
--	g3689 = AND(g3162, g2826)
--	g4588 = AND(g2419, g4273)
--	g5197 = AND(g465, g4967)
--	g4161 = AND(g3931, g2087)
--	g4361 = AND(g3995, g3354)
--	g3671 = AND(g2760, g2405)
--	g4051 = AND(g449, g3388)
--	g6092 = AND(g1123, g5731)
--	g4346 = AND(g157, g3773)
--	g2323 = AND(g471, g1358)
--	g5562 = AND(g5228, g5457)
--	g3910 = AND(g3546, g1049)
--	g3609 = AND(g2706, g2678)
--	g6262 = AND(g516, g5901)
--	g6736 = AND(g6712, g754, g5237)
--	g3758 = AND(g545, g3461)
--	g4043 = AND(g457, g3388)
--	g3365 = AND(g254, g2892)
--	g5441 = AND(g4537, g5251, g1558)
--	g5673 = AND(g59, g5573)
--	g4347 = AND(g3986, g3320)
--	g3133 = AND(g236, g2410)
--	g3333 = AND(g2264, g2728)
--	g3774 = AND(g3016, g3510)
--	g4697 = AND(g4589, g1363)
--	g3780 = AND(g3043, g3519)
--	g6737 = AND(g6714, g760, g5237)
--	g6077 = AND(g5824, g1735)
--	g3662 = AND(g2544, g3114)
--	g6643 = AND(g6574, g6229)
--	g3290 = AND(g2213, g2664)
--	g6634 = AND(g1595, g6545)
--	g3816 = AND(g3434, g861)
--	g2113 = AND(g1576, g1535)
--	g6099 = AND(g1222, g5753)
--	g6304 = AND(g5915, g6165)
--	g3181 = AND(g254, g2509)
--	g3381 = AND(g3128, g1998)
--	g3685 = AND(g2256, g2818)
--	g3700 = AND(g2276, g2837)
--	g3421 = AND(g622, g2846)
--	g5569 = AND(g5348, g3772)
--	g4460 = AND(g4218, g1539)
--	g4597 = AND(g3694, g4286)
--	g6613 = AND(g932, g6554)
--	g4739 = AND(g2850, g4579)
--	g6269 = AND(g524, g5908)
--	g4937 = AND(g166, g4732)
--	g4668 = AND(g4642, g4638)
--	g3631 = AND(g2631, g2324)
--	g2160 = AND(g1624, g929)
--	g4390 = AND(g418, g3799)
--	g3301 = AND(g218, g2866)
--	g4501 = AND(g4250, g1671)
--	g4156 = AND(g3926, g2078)
--	g4356 = AND(g175, g3779)
--	g4942 = AND(g175, g4736)
--	g5183 = AND(g418, g4950)
--	g4163 = AND(g374, g3892)
--	g5023 = AND(g3935, g4804)
--	g4363 = AND(g402, g3786)
--	g4032 = AND(g441, g3388)
--	g4053 = AND(g3387, g1415)
--	g4453 = AND(g4238, g1858)
--	g5161 = AND(g5095, g4535)
--	g3669 = AND(g2234, g2790)
--	g5361 = AND(g4435, g5168)
--	g3368 = AND(g2822, g2923)
--	g6135 = AND(g5584, g5958)
--	g5665 = AND(g361, g5570)
--	g6831 = AND(g6812, g5975)
--	g5451 = AND(g5251, g4544)
--	g6288 = AND(g5615, g6160)
--	g4157 = AND(g3830, g1533)
--	g4357 = AND(g3990, g3342)
--	g5146 = AND(g184, g5099)
--	g6916 = AND(g6903, g6901)
--	g5633 = AND(g4496, g5539)
--	g3505 = AND(g2924, g1749)
--	g6749 = AND(g6735, g6734)
--	g6798 = AND(g4946, g6781)
--	g5944 = AND(g5778, g5403)
--	g5240 = AND(g293, g4915)
--	g5043 = AND(g3941, g4805)
--	g5443 = AND(g4537, g5251, g2307)
--	g6302 = AND(g5740, g6164)
--	g6719 = AND(g4518, g6665)
--	g2092 = AND(g642, g1570)
--	g4683 = AND(g4585, g2066)
--	g5681 = AND(g79, g5577)
--	g3688 = AND(g2783, g2457)
--	g4735 = AND(g2018, g4577)
--	g6265 = AND(g520, g5903)
--	g4782 = AND(g1624, g4623)
--	g4661 = AND(g4637, g4634)
--	g4949 = AND(g193, g4753)
--	g3326 = AND(g2734, g1891)
--	g6770 = AND(g6754, g3482)
--	g3760 = AND(g548, g3465)
--	g5936 = AND(g5113, g5788)
--	g4039 = AND(g402, g3388)
--	g5317 = AND(g148, g4869)
--	g3383 = AND(g3128, g2004)
--	g5601 = AND(g5052, g5518)
--	g3608 = AND(g2599, g2308)
--	g3924 = AND(g3505, g471)
--	g4583 = AND(g1808, g4267)
--	g3161 = AND(g2397, g2470)
--	g2339 = AND(g1603, g197)
--	g3361 = AND(g3150, g1950)
--	g4616 = AND(g4231, g3761)
--	g3665 = AND(g2748, g2378)
--	g3127 = AND(g224, g2394)
--	g3327 = AND(g2772, g2906)
--	g3146 = AND(g2370, g2446)
--	g3633 = AND(g2497, g3076)
--	g5937 = AND(g5775, g5392)
--	g3103 = AND(g212, g2353)
--	g3303 = AND(g2722, g2890)
--	g5668 = AND(g49, g5571)
--	g6338 = AND(g6251, g6067)
--	g5190 = AND(g426, g4950)
--	g5501 = AND(g5454, g3478)
--	g2551 = AND(g715, g1826)
--	g5156 = AND(g434, g4877)
--	g5356 = AND(g5265, g1902)
--	g4277 = AND(g3936, g942)
--	g5942 = AND(g5117, g5797)
--	g4789 = AND(g3551, g4632)
--	g3316 = AND(g2748, g2894)
--	g3434 = AND(g2850, g857)
--	g5954 = AND(g5121, g5813)
--	g5163 = AND(g402, g4950)
--	g6098 = AND(g1209, g5753)
--	g3147 = AND(g2419, g59)
--	g5363 = AND(g4439, g5179)
--	g3681 = AND(g2234, g2806)
--	g5053 = AND(g4599, g4808)
--	g3697 = AND(g2796, g2481)
--	g5157 = AND(g496, g4904)
--	g5357 = AND(g398, g5220)
--	g4244 = AND(g1749, g4004, g1609)
--	g4340 = AND(g3972, g3291)
--	g3936 = AND(g3551, g940)
--	g3117 = AND(g218, g2367)
--	g3317 = AND(g2722, g2895)
--	g4035 = AND(g437, g3388)
--	g918 = AND(g610, g602)
--	g6086 = AND(g1143, g5742)
--	g4214 = AND(g1822, g4045)
--	g1620 = AND(g1056, g1084)
--	g3784 = AND(g114, g3251)
--	g2916 = AND(g1030, g2113)
--	g3479 = AND(g345, g2957)
--	g6131 = AND(g5593, g5975)
--	g3668 = AND(g2568, g3124)
--	g6331 = AND(g3891, g6212)
--	g4236 = AND(g654, g3907)
--	g3294 = AND(g139, g2870)
--	g5949 = AND(g5119, g5805)
--	g3190 = AND(g260, g2535)
--	g6766 = AND(g6750, g2986)
--	g3156 = AND(g242, g2464)
--	g3356 = AND(g248, g2888)
--	g5646 = AND(g4502, g5544)
--	g2873 = AND(g1845, g1861)
--	g6748 = AND(g6733, g6732)
--	g5603 = AND(g5504, g4911)
--	g5484 = AND(g378, g5331)
--	g4928 = AND(g148, g4723)
--	g3704 = AND(g2276, g2841)
--	g4464 = AND(g4272, g1937)
--	g4785 = AND(g2160, g4625)
--	g6091 = AND(g1161, g5753)
--	g3810 = AND(g625, g3421)
--	g5952 = AND(g5120, g5809)
--	g5616 = AND(g5505, g4929)
--	g6718 = AND(g4511, g6661)
--	g6767 = AND(g6754, g2986)
--	g3157 = AND(g2422, g2467)
--	g3357 = AND(g242, g2889)
--	g4489 = AND(g2166, g4206)
--	g2770 = AND(g2518, g1972)
--	g4471 = AND(g4253, g332)
--	g5503 = AND(g366, g5384)
--	g3626 = AND(g3031, g2727)
--	g4038 = AND(g430, g3388)
--	g5617 = AND(g5061, g5524)
--	g3683 = AND(g3150, g2813)
--	g4836 = AND(g4527, g4523)
--	g2138 = AND(g1639, g809)
--	g3661 = AND(g2234, g2778)
--	g6247 = AND(g504, g5893)
--	g3627 = AND(g2473, g3067)
--	g5945 = AND(g5118, g5801)
--	g2808 = AND(g2009, g1581)
--	g3292 = AND(g2214, g2667)
--	g3646 = AND(g2179, g2756)
--	g2759 = AND(g2473, g1966)
--	g6910 = AND(g6892, g6891)
--	g3603 = AND(g2370, g3019)
--	g3484 = AND(g349, g2958)
--	g5482 = AND(g370, g5331)
--	g3702 = AND(g2284, g2839)
--	g6066 = AND(g5824, g1721)
--	g5214 = AND(g562, g5025)
--	g3616 = AND(g2397, g3049)
--	g6055 = AND(g5824, g1696)
--	g6133 = AND(g5723, g5975)
--	g5663 = AND(g4513, g5550)
--	g6333 = AND(g3896, g6212)
--	g2419 = AND(g1808, g54)
--	g3764 = AND(g551, g3480)
--	g5402 = AND(g370, g5266)
--	g5236 = AND(g269, g4915)
--	g4708 = AND(g578, g4541)
--	g5556 = AND(g5015, g5445)
--	g4219 = AND(g3911, g1655)
--	g3277 = AND(g2174, g2625)
--	g3617 = AND(g2609, g2317)
--	g6093 = AND(g1177, g5742)
--	g2897 = AND(g1030, g2062)
--	g6256 = AND(g1696, g6040)
--	g4176 = AND(g386, g3901)
--	g6816 = AND(g6784, g3346)
--	g4829 = AND(g4526, g4522)
--	g6263 = AND(g1711, g6052)
--	g5194 = AND(g586, g4874)
--	g3709 = AND(g2284, g2845)
--	g5557 = AND(g5016, g5448)
--	g3340 = AND(g2772, g2915)
--	g6631 = AND(g1838, g6545)
--	g3907 = AND(g650, g3522)
--	g4177 = AND(g3933, g1372)
--	g5948 = AND(g5779, g5407)
--	g4377 = AND(g457, g3791)
--	g3690 = AND(g2276, g2827)
--	g5955 = AND(g5782, g5420)
--	g5350 = AND(g5325, g3453)
--	g4199 = AND(g628, g3810)
--	g5438 = AND(g5224, g3769)
--	g2868 = AND(g1316, g1861)
--	g3310 = AND(g224, g2871)
--	g4797 = AND(g4593, g4643)
--	g5212 = AND(g561, g5025)
--	g3663 = AND(g2215, g2779)
--	g2793 = AND(g2568, g1991)
--	g2015 = AND(g616, g1419)
--	g4344 = AND(g3981, g3306)
--	g5229 = AND(g545, g4980)
--	g6772 = AND(g6746, g3312)
--	g3762 = AND(g2672, g3500)
--	g4694 = AND(g1481, g4578)
--	g3657 = AND(g2734, g2357)
--	g2721 = AND(g2397, g1922)
--	g4488 = AND(g1633, g4202)
--	g4701 = AND(g4596, g1378)
--	g3928 = AND(g3512, g478)
--	g6474 = AND(g2138, g2036, g6397)
--	g3899 = AND(g323, g3441)
--	g3464 = AND(g341, g2956)
--	g5620 = AND(g5507, g4938)
--	g4870 = AND(g4779, g1884)
--	g3295 = AND(g2660, g2647)
--	g2671 = AND(g2263, g2296)
--	g1576 = AND(g1101, g1094)
--	g3844 = AND(g3540, g1665)
--	g1716 = AND(g821, g774, g784)
--	g3089 = AND(g212, g2336)
--	g3731 = AND(g331, g3441)
--	g3489 = AND(g2607, g1861)
--	g5192 = AND(g1046, g4894)
--	g5485 = AND(g382, g5331)
--	g5941 = AND(g5777, g5399)
--	g4230 = AND(g3756, g1861)
--	g6126 = AND(g5711, g5958)
--	g6326 = AND(g3833, g6194)
--	g4033 = AND(g426, g3388)
--	g3814 = AND(g913, g3546)
--	g2758 = AND(g2497, g1963)
--	g3350 = AND(g3150, g1928)
--	g2861 = AND(g2120, g1654)
--	g6924 = AND(g6920, g6919)
--	g5176 = AND(g410, g4950)
--	g4395 = AND(g445, g3800)
--	g5376 = AND(g170, g5255)
--	g5911 = AND(g5817, g5670)
--	g2846 = AND(g619, g2015)
--	g6127 = AND(g5714, g5975)
--	g6327 = AND(g3884, g6212)
--	g5225 = AND(g669, g5054)
--	g4342 = AND(g3978, g3299)
--	g6146 = AND(g3192, g5997)
--	g6346 = AND(g6274, g6087)
--	g2018 = AND(g1423, g1254)
--	g4354 = AND(g437, g3777)
--	I5352 = AND(g3529, g3531, g3535, g3538)
--	g5177 = AND(g445, g4877)
--	g6240 = AND(g4205, g5888)
--	g3620 = AND(g2422, g3060)
--	g1027 = AND(g598, g567)
--	g2685 = AND(g2370, g1887)
--	g2700 = AND(g2370, g1908)
--	g2021 = AND(g835, g1436)
--	g6316 = AND(g3855, g6194)
--	g5898 = AND(g5800, g5647)
--	g4401 = AND(g426, g3802)
--	g1514 = AND(g1017, g1011)
--	g5900 = AND(g5804, g5658)
--	g2950 = AND(g2156, g1612)
--	g4761 = AND(g4567, g1674)
--	g5245 = AND(g297, g4915)
--	g1763 = AND(g478, g1119)
--	g4828 = AND(g4510, g4508)
--	g3298 = AND(g2231, g2679)
--	g4830 = AND(g4529, g4525)
--	g5144 = AND(g166, g5099)
--	g4592 = AND(g3147, g4281)
--	g6914 = AND(g6895, g6893)
--	g2101 = AND(g1001, g1543)
--	g5488 = AND(g394, g5331)
--	g4932 = AND(g157, g4727)
--	g1416 = AND(g913, g266)
--	g5701 = AND(g5683, g3813)
--	g6317 = AND(g3862, g6194)
--	g5215 = AND(g4864, g5090)
--	g5951 = AND(g5780, g5411)
--	g4677 = AND(g4652, g4646)
--	g3176 = AND(g2422, g2494)
--	g3376 = AND(g3104, g1979)
--	g3286 = AND(g2196, g2656)
--	g3765 = AND(g554, g3485)
--	g4349 = AND(g441, g3775)
--	g6060 = AND(g5824, g1703)
--	g1595 = AND(g729, g719, g766, I2566)
--	I5359 = AND(g3518, g3521, g3526, g3530)
--	g3610 = AND(g2397, g3034)
--	g6739 = AND(g6715, g815, g5242)
--	g1612 = AND(g784, g774, g821, I2574)
--	g3324 = AND(g230, g2875)
--	g6079 = AND(g1236, g5753)
--	g5122 = AND(g193, g4662)
--	g3377 = AND(g3118, g2931)
--	g4352 = AND(g3988, g3331)
--	g4867 = AND(g4811, g3872)
--	g6156 = AND(g2591, g6015)
--	g3287 = AND(g135, g2865)
--	g5096 = AND(g4794, g4647)
--	g4186 = AND(g3973, g1395)
--	g5496 = AND(g5446, g3457)
--	g6250 = AND(g1692, g6036)
--	g4170 = AND(g382, g3900)
--	g4280 = AND(g2138, g1764, g4007)
--	g3144 = AND(g236, g2440)
--	g3344 = AND(g242, g2885)
--	g5142 = AND(g148, g5099)
--	g3819 = AND(g964, g3437)
--	g6912 = AND(g6899, g6897)
--	g3694 = AND(g3147, g64)
--	g6157 = AND(g3158, g5997)
--	g5481 = AND(g366, g5331)
--	g3701 = AND(g2268, g2838)
--	g5497 = AND(g5447, g3458)
--	g5154 = AND(g500, g4993)
--	g5354 = AND(g5249, g2903)
--	g4461 = AND(g4241, g2919)
--	g4756 = AND(g3816, g4587)
--	g4046 = AND(I5351, I5352)
--	g5218 = AND(g564, g5025)
--	g3650 = AND(g2660, g2347)
--	g4345 = AND(g3982, g3308)
--	g3336 = AND(g2760, g1911)
--	g3768 = AND(g3448, g1528)
--	g4159 = AND(g370, g3890)
--	g4359 = AND(g434, g3782)
--	g3806 = AND(g3384, g2024)
--	g4416 = AND(g3905, g1481)
--	g3887 = AND(g3276, g1861)
--	g3122 = AND(g2435, g1394)
--	g2732 = AND(g2449, g1940)
--	g4047 = AND(g453, g3388)
--	g6646 = AND(g6577, g6232)
--	g3433 = AND(g1359, g2831, g905)
--	g5953 = AND(g5781, g5415)
--	g6084 = AND(g1123, g5753)
--	g6603 = AND(g6581, g6236)
--	g4874 = AND(g582, g4708)
--	g5677 = AND(g69, g5575)
--	g3195 = AND(g2473, g2541)
--	g3337 = AND(g2796, g2913)
--	I4040 = AND(g1279, g2025, g1267)
--	g5149 = AND(g4910, g1480)
--	g5349 = AND(g5324, g3451)
--	g5198 = AND(g558, g5025)
--	g5398 = AND(g366, g5261)
--	g1570 = AND(g634, g1027)
--	g6647 = AND(g6578, g6233)
--	g1691 = AND(g821, g774)
--	g3692 = AND(g2268, g2829)
--	g3726 = AND(g119, g3251)
--	g3154 = AND(g2039, g1410)
--	g4800 = AND(g4648, g4296)
--	g5152 = AND(g430, g4950)
--	g6320 = AND(g3869, g6194)
--	g5211 = AND(g4860, g5086)
--	g5186 = AND(g422, g4950)
--	g5599 = AND(g5049, g5512)
--	g4490 = AND(g2941, g4210)
--	g3293 = AND(g212, g2864)
--	g6771 = AND(g6758, g3483)
--	g3329 = AND(g2748, g2907)
--	g5170 = AND(g5091, g2111)
--	g4456 = AND(g3829, g4229)
--	g6299 = AND(g5530, g6163)
--	g4348 = AND(g3987, g3322)
--	g3727 = AND(g122, g3251)
--	g2937 = AND(g2160, g931)
--	g4355 = AND(g430, g3778)
--	g5939 = AND(g5776, g5395)
--	g2294 = AND(g1716, g791, g798)
--	g4698 = AND(g4586, g2106)
--	g5483 = AND(g374, g5331)
--	g3703 = AND(g2284, g2840)
--	g6738 = AND(g6713, g809, g5242)
--	g2156 = AND(g815, g1642)
--	g6244 = AND(g4759, g5891)
--	g2356 = AND(g1603, g269)
--	g6140 = AND(g5587, g5975)
--	g3953 = AND(g3554, g188)
--	g6340 = AND(g6257, g6069)
--	g5187 = AND(g457, g4877)
--	g1628 = AND(g815, g809)
--	g4167 = AND(g378, g3898)
--	g6082 = AND(g1123, g5742)
--	g4367 = AND(g193, g3788)
--	g4872 = AND(g4760, g1549)
--	g4057 = AND(g422, g3388)
--	g5904 = AND(g5812, g5664)
--	g5200 = AND(g559, g5025)
--	g4457 = AND(g4261, g2902)
--	g5446 = AND(g4537, g5241)
--	g3349 = AND(g2783, g1925)
--	g2053 = AND(g1094, g1675)
--	g5145 = AND(g175, g5099)
--	g6915 = AND(g6906, g6905)
--	g4834 = AND(g4534, g4531)
--	g4686 = AND(g4590, g1348)
--	g5191 = AND(g461, g4877)
--	g3699 = AND(g2276, g2836)
--	g4598 = AND(g1978, g4253)
--	g5637 = AND(g4499, g5543)
--	g5159 = AND(g536, g4967)
--	g5359 = AND(g4428, g5155)
--	g4253 = AND(g1861, g3819)
--	g3644 = AND(g2197, g2755)
--	g3319 = AND(g2688, g2675)
--	g3352 = AND(g2796, g2920)
--	g5047 = AND(g3954, g4806)
--	g5447 = AND(g4545, g5256, g2311)
--	g4687 = AND(g4493, g1542)
--	g3186 = AND(g2449, g2515)
--	g3170 = AND(g254, g2485)
--	g3614 = AND(g2998, g2691)
--	g3325 = AND(g224, g2876)
--	g4341 = AND(g3977, g3297)
--	g2782 = AND(g2518, g1985)
--	g6295 = AND(g5379, g6162)
--	g3280 = AND(g2177, g2637)
--	g5017 = AND(g4784, g1679)
--	g4691 = AND(g4581, g2098)
--	g5935 = AND(g5112, g5784)
--	g2949 = AND(g830, g1861)
--	I5351 = AND(g3511, g3517, g3520, g3525)
--	g5234 = AND(g197, g4915)
--	g3636 = AND(g2701, g2327)
--	g2292 = AND(g1706, g736, g743)
--	g6089 = AND(g1143, g5731)
--	g6731 = AND(g6717, g4427)
--	g6557 = AND(g1595, g6469)
--	g4358 = AND(g3991, g3343)
--	g2084 = AND(g1577, g1563)
--	g2850 = AND(g2018, g1255)
--	g5213 = AND(g4862, g5087)
--	g6254 = AND(g532, g5897)
--	g6150 = AND(g3204, g6015)
--	g5902 = AND(g5808, g5661)
--	g3145 = AND(g2397, g2443)
--	g3345 = AND(g236, g2886)
--	g6773 = AND(g6762, g2986)
--	g3763 = AND(g3064, g3501)
--	g3191 = AND(g2497, g2538)
--	g4180 = AND(g3929, g2119)
--	g5166 = AND(g541, g4967)
--	g3637 = AND(g2822, g2752)
--	g4832 = AND(g4517, g4512)
--	g6769 = AND(g6758, g2986)
--	g3307 = AND(g2242, g2692)
--	g3359 = AND(g2822, g2922)
--	g4794 = AND(g4593, g949)
--	g3757 = AND(g2619, g3487)
--	g3522 = AND(g646, g2909)
--	g3315 = AND(g2701, g1875)
--	g3642 = AND(g3054, g2754)
--	g3654 = AND(g2518, g3100)
--	g5619 = AND(g5064, g5527)
--	g5167 = AND(g5011, g1556)
--	
--	g3880 = OR(g3658, g3665)
--	g4440 = OR(g4371, g4038)
--	g3978 = OR(g3655, g3117)
--	g6788 = OR(g3760, g6767)
--	g3935 = OR(g3464, g2868)
--	g3982 = OR(g3663, g3127)
--	I8376 = OR(g6315, g6126, g6129, g6146)
--	g5625 = OR(g5495, g3281)
--	g6298 = OR(g6255, g6093)
--	g6485 = OR(I8393, I8394, I8395)
--	g4655 = OR(g4368, g3660)
--	g6252 = OR(g5905, g2381)
--	g6176 = OR(g6068, g6033)
--	I8377 = OR(g6150, g6324, g5180, g5181)
--	g6286 = OR(g6238, g6079)
--	g3851 = OR(g3681, g3146)
--	g3964 = OR(g3634, g3089)
--	g5659 = OR(g5551, g5398)
--	g2928 = OR(g2100, g1582)
--	g6287 = OR(g6241, g6082)
--	g3989 = OR(g3679, g3144)
--	g5374 = OR(g5215, g4947)
--	g3971 = OR(g3644, g3099)
--	g6781 = OR(g6718, g6748)
--	g3598 = OR(g2808, g2821)
--	g4641 = OR(g4347, g3627)
--	g4450 = OR(g4389, g4047)
--	g3740 = OR(g3335, g2747)
--	I8136 = OR(g6015, g6212, g4950, g4877)
--	g5628 = OR(g5498, g3292)
--	g5630 = OR(g5501, g3309)
--	g6114 = OR(g5904, g5604)
--	g5323 = OR(g5098, g4802)
--	g5666 = OR(g5555, g5406)
--	I8137 = OR(g4894, g4904, g4993, g4967)
--	I8395 = OR(g5182, g5200, g6280)
--	g3879 = OR(g3704, g3195)
--	I9057 = OR(g6320, g6828, g6830, g6153)
--	g4092 = OR(g3311, g2721)
--	I8081 = OR(g4894, g4904, g4993, g4967)
--	g4864 = OR(g4744, g4490)
--	g6845 = OR(I9064, I9065, I9066)
--	g5372 = OR(g5213, g4942)
--	g5693 = OR(g5632, g5481)
--	g5804 = OR(g5371, g5603)
--	g6142 = OR(g5909, g3806)
--	I8129 = OR(g4915, g5025)
--	g6481 = OR(I8367, I8368, I8369, I8370)
--	g4651 = OR(g4357, g3643)
--	g4285 = OR(g3490, g3887)
--	g4500 = OR(g4243, g2010)
--	g5202 = OR(g4904, g4914, g4894)
--	g3750 = OR(g3372, g2794)
--	g6267 = OR(g2953, g5884)
--	g4231 = OR(g3997, g4000)
--	g6676 = OR(g6631, g6555)
--	g6293 = OR(g6244, g6085)
--	g4205 = OR(g3843, g541)
--	g4634 = OR(g4341, g3615)
--	I8349 = OR(I8345, I8346, I8347, I8348)
--	g6703 = OR(g6692, g4831)
--	g3884 = OR(g3666, g3671)
--	g4444 = OR(g4378, g4042)
--	g4862 = OR(g4739, g4489)
--	I8119 = OR(g5202, g4993, g4967, g4980)
--	g3988 = OR(g3678, g3143)
--	g5674 = OR(g5558, g5419)
--	g6747 = OR(g6614, g6731)
--	g6855 = OR(g6851, g2085)
--	I8211 = OR(g4915, g5025)
--	I8386 = OR(g6152, g6327, g5183, g5177)
--	g5680 = OR(g5562, g5429)
--	g4946 = OR(g4830, g4833)
--	I8370 = OR(g5214, g6358)
--	g4436 = OR(g4359, g4035)
--	I8387 = OR(g5178, g5209, g6281)
--	g6274 = OR(g5682, g5956)
--	g6426 = OR(g6288, g6119)
--	g6170 = OR(g6061, g6014)
--	g3996 = OR(g3691, g3171)
--	I8345 = OR(g6326, g6135, g6140, g6157)
--	g5623 = OR(g5503, g5357)
--	g6483 = OR(I8385, I8386, I8387)
--	g4653 = OR(g4361, g3652)
--	g3878 = OR(g3703, g3191)
--	g6790 = OR(g3765, g6773)
--	I8359 = OR(g5232, g5236, g5216, g5226)
--	g4752 = OR(g4452, g4155)
--	g6461 = OR(g6353, g6351)
--	g3981 = OR(g3661, g3123)
--	g5024 = OR(g4793, g4600)
--	g4233 = OR(g3912, g471)
--	g4454 = OR(g4395, g4051)
--	g5672 = OR(g5557, g5414)
--	g5077 = OR(g1612, g4694)
--	g5231 = OR(g5048, g672)
--	g6307 = OR(g6262, g6096)
--	g3744 = OR(g3345, g2759)
--	g6251 = OR(g5668, g5939)
--	g6447 = OR(g6340, g5938)
--	I8128 = OR(g5202, g4993, g4967, g4980)
--	g3864 = OR(g3693, g3176)
--	g5044 = OR(g4797, g4602)
--	g4745 = OR(g4468, g4569)
--	g6272 = OR(g5679, g5953)
--	g5014 = OR(g4785, g4583)
--	g3871 = OR(g3701, g3186)
--	I7970 = OR(g6015, g6212, g4950, g4877)
--	I8348 = OR(g5229, g5234, g5218, g5225)
--	g6554 = OR(g6337, g6466)
--	I7987 = OR(g6194, g5958, g5975, g5997)
--	g5916 = OR(g5728, g3781)
--	I8118 = OR(g6015, g6212, g4950, g4877)
--	I8367 = OR(g6313, g6124, g6127, g6144)
--	g6456 = OR(g6346, g5954)
--	I8393 = OR(g6317, g6130, g6133, g6151)
--	g4086 = OR(g3310, g2720)
--	g1589 = OR(g1059, g1045)
--	g6118 = OR(g5911, g5619)
--	g6167 = OR(g6056, g6039)
--	g3862 = OR(g3632, g3641)
--	g6457 = OR(g6352, g6347)
--	g4635 = OR(g4342, g3616)
--	g6549 = OR(g6473, g4247)
--	g6686 = OR(g6259, g6645)
--	g5532 = OR(g5350, g3278)
--	g6670 = OR(g6557, g6634, g4410, g2948)
--	g5012 = OR(g4782, g4580)
--	g4059 = OR(g3466, g3425)
--	g5281 = OR(g5074, g5124)
--	I8358 = OR(g5192, g5153, g5158, g5197)
--	g6687 = OR(g6260, g6646)
--	g3749 = OR(g3371, g2793)
--	g5808 = OR(g5373, g5616)
--	g6691 = OR(g6275, g6603)
--	g3873 = OR(g3649, g3657)
--	g3869 = OR(g3642, g3650)
--	g6659 = OR(g6634, g6631)
--	g4430 = OR(g4349, g4015)
--	g6239 = OR(g2339, g6073)
--	g6545 = OR(g6468, g4244)
--	g4638 = OR(g4345, g3620)
--	g6794 = OR(g6777, g3333)
--	g6931 = OR(g6741, g6929)
--	g3990 = OR(g3684, g3155)
--	g5385 = OR(g3992, g5318)
--	g3888 = OR(g3672, g3682)
--	g5470 = OR(g5359, g5142)
--	g6300 = OR(g6253, g6091)
--	g4455 = OR(g4396, g4052)
--	g6750 = OR(g6670, g6625, g6736)
--	g5678 = OR(g5560, g5428)
--	g3745 = OR(g3356, g2770)
--	g6440 = OR(g6336, g5935)
--	g3865 = OR(g3637, g3648)
--	g3833 = OR(g3602, g3608)
--	g4021 = OR(g3558, g2949)
--	g3896 = OR(g3689, g3697)
--	g5535 = OR(g5353, g3300)
--	g5015 = OR(g4787, g4588)
--	g4631 = OR(g4340, g3611)
--	g5246 = OR(g5077, g2080)
--	g6792 = OR(g6770, g3321)
--	I7980 = OR(g5202, g4993, g4967, g4980)
--	I8360 = OR(I8356, I8357, I8358, I8359)
--	g4441 = OR(g4372, g4039)
--	g6113 = OR(g5902, g5601)
--	g5388 = OR(g5318, g1589, g3491)
--	I8379 = OR(g5212, g6357)
--	g5430 = OR(g5161, g4873)
--	g4458 = OR(g4401, g4057)
--	g3748 = OR(g3366, g2782)
--	g6264 = OR(g5675, g5948)
--	g4074 = OR(g3301, g2699)
--	g6450 = OR(g6341, g5940)
--	g4080 = OR(g3302, g2700)
--	g5066 = OR(g4668, g4672)
--	g6179 = OR(g6077, g6051)
--	I8209 = OR(g6015, g6212, g4950, g4877)
--	g6289 = OR(g6240, g6081)
--	g6658 = OR(g6132, g6620)
--	g6271 = OR(g2955, g5885)
--	g5662 = OR(g5553, g5402)
--	g5018 = OR(g4791, g4597)
--	I7972 = OR(g4915, g5025)
--	g5467 = OR(g3868, g5318, g3992)
--	g5816 = OR(g5378, g5620)
--	g5700 = OR(g5663, g5488)
--	g4451 = OR(g4390, g4048)
--	g6864 = OR(g6852, g2089)
--	g5817 = OR(g5380, g5621)
--	g3883 = OR(g3709, g3203)
--	g5605 = OR(g3575, g5500)
--	I9059 = OR(g5185, g5198, g6279)
--	g4443 = OR(g4377, g4041)
--	g4434 = OR(g4355, g4033)
--	g5669 = OR(g5556, g5410)
--	g5368 = OR(g5201, g4932)
--	I7979 = OR(g6015, g6212, g4950, g4877)
--	g5531 = OR(g5349, g3275)
--	g5458 = OR(g3466, g5311)
--	g6795 = OR(g4867, g6772)
--	g4936 = OR(g4827, g4828)
--	g5074 = OR(g4792, g4598)
--	g5474 = OR(g5363, g5146)
--	g6926 = OR(g6798, g6923)
--	g6754 = OR(g6676, g6625, g6737)
--	g6273 = OR(g5681, g5955)
--	g6444 = OR(g6338, g5936)
--	I8378 = OR(g5173, g5166, g5235, g5245)
--	I8135 = OR(g6194, g5958, g5975, g5997)
--	g5326 = OR(g5069, g4410, g3012)
--	I9066 = OR(g5189, g5269, g6400)
--	g6927 = OR(g6799, g6924)
--	g3751 = OR(g3375, g2807)
--	g6660 = OR(g6640, g6637)
--	g6679 = OR(g6637, g6558)
--	I8208 = OR(g6194, g5958, g5975, g5997)
--	g6182 = OR(g6047, g6034)
--	g5327 = OR(g5077, g4416, g3028)
--	g3743 = OR(g3344, g2758)
--	g3856 = OR(g3686, g3157)
--	g5303 = OR(g5053, g4768)
--	g5696 = OR(g5637, g5484)
--	g3992 = OR(g1555, g3559)
--	g5472 = OR(g5361, g5144)
--	g3863 = OR(g3692, g3172)
--	g6437 = OR(g6302, g6121)
--	g6917 = OR(g6909, g6910)
--	g3857 = OR(g3687, g3161)
--	g5533 = OR(g5351, g3290)
--	g5697 = OR(g5646, g5485)
--	g5013 = OR(g4826, g4621)
--	g4627 = OR(g4333, g3603)
--	g6454 = OR(g6344, g5949)
--	g6296 = OR(g6247, g6088)
--	g4646 = OR(g4353, g3635)
--	I8138 = OR(g4980, g4915, g5025, g5054)
--	g6189 = OR(g6060, g6035)
--	g3977 = OR(g3653, g3113)
--	I9058 = OR(g6156, g6331, g5190, g5164)
--	g6787 = OR(g3758, g6766)
--	g5060 = OR(g3491, g4819)
--	g6297 = OR(g6248, g6089)
--	g3999 = OR(g3699, g3181)
--	g6684 = OR(g6250, g6643)
--	I7978 = OR(g6194, g5958, g5975, g5997)
--	g6109 = OR(g5900, g5599)
--	g6791 = OR(g6768, g3307)
--	g6309 = OR(g6265, g6098)
--	g3732 = OR(g3324, g2732)
--	g3533 = OR(g3154, g3166)
--	I8385 = OR(g6316, g6128, g6131, g6149)
--	g6268 = OR(g5677, g5951)
--	g3820 = OR(g3287, g2671)
--	g6452 = OR(g6342, g5942)
--	g5626 = OR(g5496, g3285)
--	g4656 = OR(g4369, g3662)
--	g6185 = OR(g6055, g5995)
--	g3739 = OR(g3334, g2746)
--	I7989 = OR(g5202, g4993, g4967, g4980)
--	g3995 = OR(g3690, g3170)
--	I8369 = OR(g5165, g5159, g5233, g5240)
--	I7971 = OR(g5202, g4993, g4967, g4980)
--	g5627 = OR(g5497, g3286)
--	g6682 = OR(g6478, g6624, g6623)
--	g3942 = OR(g3215, g3575)
--	g5583 = OR(g5569, g4020)
--	g6173 = OR(g6066, g6043)
--	g3954 = OR(g3484, g3489)
--	g6920 = OR(g6915, g6916)
--	g6261 = OR(g5673, g5944)
--	g6793 = OR(g6771, g3323)
--	g4948 = OR(g4834, g4836)
--	g6246 = OR(g5665, g5937)
--	g5224 = OR(g5123, g3630)
--	g5277 = OR(g5023, g4763)
--	g4438 = OR(g4363, g4037)
--	g4773 = OR(g4495, g4220)
--	g6689 = OR(g6266, g6648)
--	g3998 = OR(g3698, g3180)
--	I8774 = OR(g6655, g6653, g6651, g6649)
--	g3850 = OR(g3680, g3145)
--	g6108 = OR(g5898, g5598)
--	g6758 = OR(g6673, g6628, g6738)
--	g2896 = OR(g2323, g1763)
--	g6455 = OR(g6345, g5952)
--	g3986 = OR(g3667, g3133)
--	g6846 = OR(g5860, g6834)
--	g3503 = OR(g3122, g3132)
--	I7969 = OR(g6194, g5958, g5975, g5997)
--	g4941 = OR(g4829, g4832)
--	g6290 = OR(g6245, g6086)
--	g3987 = OR(g3669, g3134)
--	g6847 = OR(g5861, g6837)
--	g6685 = OR(g6256, g6644)
--	g5295 = OR(g5047, g4766)
--	g4473 = OR(g3575, g4253)
--	g3991 = OR(g3685, g3156)
--	I7988 = OR(g6015, g6212, g4950, g4877)
--	g5471 = OR(g5360, g5143)
--	I8368 = OR(g6148, g6321, g5176, g5184)
--	g6257 = OR(g5671, g5941)
--	g6301 = OR(g6254, g6092)
--	g6673 = OR(g6559, g6640, g4416, g2950)
--	I8080 = OR(g6015, g6212, g4950, g4877)
--	g6669 = OR(g6613, g4679)
--	g3877 = OR(g3651, g3659)
--	I8126 = OR(g6194, g5958, g5975, g5997)
--	g5062 = OR(g4661, g4666)
--	g6480 = OR(I8360, g6359)
--	I8779 = OR(g6605, g6656, g6654, g6652)
--	g6688 = OR(g6263, g6647)
--	g5085 = OR(g4694, g4280)
--	I7981 = OR(g4915, g5025)
--	I8127 = OR(g6015, g6212, g4950, g4877)
--	g4433 = OR(g4354, g4032)
--	I8346 = OR(g6159, g6334, g5163, g5191)
--	g5812 = OR(g5376, g5618)
--	g4859 = OR(g4730, g4486)
--	g6665 = OR(I8778, I8779)
--	g5473 = OR(g5362, g5145)
--	I8347 = OR(g5188, g5157, g5154, g5193)
--	g6303 = OR(g6258, g6094)
--	g5069 = OR(g1595, g4688)
--	I9064 = OR(g6323, g6829, g6831, g6155)
--	g4497 = OR(g4166, g3784)
--	I8210 = OR(g5202, g4993, g4967, g4980)
--	g5377 = OR(g5217, g4949)
--	g3837 = OR(g3609, g3613)
--	g6116 = OR(g5910, g5617)
--	I8117 = OR(g6194, g5958, g5975, g5997)
--	g4001 = OR(g3702, g3190)
--	g3842 = OR(g3670, g3135)
--	g5291 = OR(g5043, g4764)
--	g3941 = OR(g3479, g2873)
--	g5694 = OR(g5633, g5482)
--	g6936 = OR(g5438, g6935)
--	g4068 = OR(g3293, g2685)
--	I8079 = OR(g6194, g5958, g5975, g5997)
--	g4468 = OR(g4214, g3831)
--	g4866 = OR(g4756, g4491)
--	g3829 = OR(g3294, g3305)
--	I8356 = OR(g6311, g6123, g6125, g6141)
--	g3733 = OR(g3325, g2733)
--	g6937 = OR(g4616, g6934)
--	g6479 = OR(I8349, g6335)
--	g6294 = OR(g6249, g6090)
--	g5065 = OR(g4667, g4671)
--	g5228 = OR(g5096, g4800)
--	I8357 = OR(g6145, g6318, g5171, g5187)
--	g3849 = OR(g3618, g3625)
--	g6704 = OR(g6660, g492)
--	g4599 = OR(g3499, g4230)
--	g6453 = OR(g6343, g5945)
--	g4544 = OR(g4410, g2995)
--	I8778 = OR(g6612, g6611, g6609, g6607)
--	g2924 = OR(g2095, g1573)
--	g4427 = OR(g4373, g3668)
--	g4446 = OR(g4383, g4043)
--	g3870 = OR(g3700, g3182)
--	g6683 = OR(g6465, g6622, g6621)
--	g5676 = OR(g5559, g5424)
--	g4637 = OR(g4344, g3619)
--	g3972 = OR(g3646, g3103)
--	g6782 = OR(g6719, g6749)
--	g6661 = OR(I8773, I8774)
--	g4757 = OR(g4456, g4158)
--	g6292 = OR(g6243, g6084)
--	g4811 = OR(g4429, g4432)
--	g4642 = OR(g4348, g3628)
--	g4447 = OR(g4384, g4044)
--	g5624 = OR(g5494, g3280)
--	g5068 = OR(g4673, g4677)
--	g4654 = OR(g4362, g3654)
--	g3891 = OR(g3683, g3688)
--	g3913 = OR(g3449, g2860)
--	I7990 = OR(g4915, g5025)
--	g6702 = OR(g6659, g496)
--	g6919 = OR(g6912, g6914)
--	I8120 = OR(g4915, g5025)
--	g4243 = OR(g4053, g4058)
--	g5699 = OR(g5660, g5487)
--	g5241 = OR(g5069, g2067)
--	g4234 = OR(g3921, g478)
--	g3815 = OR(g3282, g2659)
--	g5386 = OR(g5227, g669)
--	g6789 = OR(g3764, g6769)
--	I8082 = OR(g4980, g4915, g5025, g5054)
--	g5370 = OR(g5211, g4937)
--	g3828 = OR(g3304, g1351)
--	I9065 = OR(g6158, g6333, g5152, g5156)
--	g3746 = OR(g3357, g2771)
--	g5083 = OR(g4688, g4271)
--	g6907 = OR(g6874, g3358)
--	g5622 = OR(g5492, g3277)
--	g6690 = OR(g6270, g6650)
--	g6482 = OR(I8376, I8377, I8378, I8379)
--	g4652 = OR(g4358, g3645)
--	g4549 = OR(g4416, g3013)
--	g3747 = OR(g3365, g2781)
--	g3855 = OR(g3626, g3631)
--	g5695 = OR(g5635, g5483)
--	g6110 = OR(g5883, g5996)
--	g6310 = OR(g6269, g6099)
--	g5016 = OR(g4789, g4592)
--	g6762 = OR(g6679, g6628, g6739)
--	g4740 = OR(g4448, g4154)
--	I8394 = OR(g6154, g6329, g5186, g5172)
--	g6556 = OR(g6339, g6467)
--	g6930 = OR(g6740, g6928)
--	g3599 = OR(g2935, g1637)
--	g3821 = OR(g2951, g3466)
--	g4860 = OR(g4735, g4488)
--	g6237 = OR(g5912, g2381)
--	g4645 = OR(g4352, g3633)
--	g6844 = OR(I9057, I9058, I9059)
--	I8773 = OR(g6610, g6608, g6606, g6604)
--	g5629 = OR(g5499, g3298)
--	g4607 = OR(g4232, g3899)
--	g6705 = OR(g6693, g4835)
--	g5800 = OR(g5369, g5600)
--	g6242 = OR(g2356, g6075)
--	g3841 = OR(g3614, g3617)
--	g6918 = OR(g6911, g6913)
--	g5348 = OR(g5317, g5122)
--	g3858 = OR(g3629, g3636)
--	g5698 = OR(g5648, g5486)
--	g4630 = OR(g4339, g3610)
--	g6921 = OR(g6908, g6816)
--	g5367 = OR(g5199, g4928)
--	
--	g1777 = NAND(g1060, g102, g89)
--	I7217 = NAND(g152, I7216)
--	I7571 = NAND(g5678, I7569)
--	g5686 = NAND(g5546, g1017, g1551, g2916)
--	I2073 = NAND(g15, I2072)
--	I2796 = NAND(g804, I2795)
--	g948 = NAND(I2014, I2015)
--	I4205 = NAND(g743, I4203)
--	I3875 = NAND(g285, I3874)
--	g3330 = NAND(g1815, g1797, g3109)
--	g4151 = NAND(I5536, I5537)
--	g2435 = NAND(g1138, g1777, g1157)
--	I5658 = NAND(g3983, I5657)
--	g1558 = NAND(I2527, I2528)
--	I4444 = NAND(g2092, g606)
--	I5271 = NAND(g3710, I5269)
--	I2898 = NAND(g1027, I2897)
--	I2797 = NAND(g798, I2795)
--	I2245 = NAND(g567, I2244)
--	I3988 = NAND(g291, g2544)
--	g1574 = NAND(I2543, I2544)
--	g3529 = NAND(g3200, g2215, g2976, g2968)
--	I1963 = NAND(g242, I1961)
--	I5209 = NAND(g3271, I5207)
--	I7562 = NAND(g74, g5676)
--	g5506 = NAND(I7231, I7232)
--	g5111 = NAND(I6744, I6745)
--	I4182 = NAND(g2292, g749)
--	I6186 = NAND(g4301, I6185)
--	I7441 = NAND(g594, I7439)
--	I6026 = NAND(g4223, g4221)
--	I2768 = NAND(g743, I2766)
--	I3933 = NAND(g288, g2473)
--	g5853 = NAND(g5638, g2053, g1076)
--	g2731 = NAND(I3894, I3895)
--	g5507 = NAND(I7238, I7239)
--	g2966 = NAND(I4160, I4161)
--	I2934 = NAND(g1436, I2933)
--	I3179 = NAND(g736, I3177)
--	I6187 = NAND(g3955, I6185)
--	I6027 = NAND(g4223, I6026)
--	g2009 = NAND(g901, g1387, g905)
--	I4233 = NAND(g2267, g798)
--	g2769 = NAND(I3953, I3954)
--	g1044 = NAND(I2081, I2082)
--	g4674 = NAND(g4550, g1514, g2107, g2897)
--	I7569 = NAND(g79, g5678)
--	I6391 = NAND(g4504, I6390)
--	g3525 = NAND(g3192, g3002, g2197, g2179)
--	g4680 = NAND(g4550, g1514, g1006, g2897)
--	I2081 = NAND(g25, I2080)
--	I8195 = NAND(g471, I8194)
--	g1534 = NAND(I2498, I2499)
--	I2497 = NAND(g1042, g1036)
--	g939 = NAND(I1987, I1988)
--	I5269 = NAND(g3705, g3710)
--	g3985 = NAND(g1138, g3718, g2142)
--	g1036 = NAND(I2061, I2062)
--	I2676 = NAND(g131, I2674)
--	g1749 = NAND(I2767, I2768)
--	g6097 = NAND(g2954, g5857)
--	g6783 = NAND(g6747, g5068, g5066)
--	g5776 = NAND(I7528, I7529)
--	I7434 = NAND(g5554, I7432)
--	g1042 = NAND(I2073, I2074)
--	I7210 = NAND(g5367, I7208)
--	g3530 = NAND(g3204, g3023, g2197, g2179)
--	I6964 = NAND(g586, I6962)
--	I5208 = NAND(g3267, I5207)
--	I5302 = NAND(g3505, I5300)
--	g5777 = NAND(I7535, I7536)
--	g4613 = NAND(I6195, I6196)
--	I2544 = NAND(g774, I2542)
--	g1138 = NAND(g102, g98)
--	I1994 = NAND(g504, g218)
--	I4445 = NAND(g2092, I4444)
--	I2061 = NAND(g7, I2060)
--	I5189 = NAND(g3593, I5187)
--	g4903 = NAND(g4717, g858)
--	I3178 = NAND(g1706, I3177)
--	I4920 = NAND(g3522, I4919)
--	g2951 = NAND(g2142, g1797)
--	g3518 = NAND(g3177, g3023, g3007, g2981)
--	I2003 = NAND(g500, g212)
--	g6717 = NAND(g6669, g5065, g5062)
--	I3916 = NAND(g2449, I3914)
--	g5864 = NAND(g5649, g1529, g1088, g2068)
--	g2008 = NAND(g866, g873, g1784)
--	I5309 = NAND(g3512, I5307)
--	I7432 = NAND(g111, g5554)
--	I4203 = NAND(g2255, g743)
--	g3521 = NAND(g3187, g3023, g3007, g2179)
--	I5759 = NAND(g3836, g3503)
--	I6962 = NAND(g4874, g586)
--	I6659 = NAND(g4762, g3541)
--	I4940 = NAND(g3437, I4939)
--	I2935 = NAND(g345, I2933)
--	g2266 = NAND(I3412, I3413)
--	I2542 = NAND(g821, g774)
--	I3412 = NAND(g1419, I3411)
--	I3189 = NAND(g1716, I3188)
--	g5634 = NAND(g5563, g4767)
--	I3990 = NAND(g2544, I3988)
--	g2960 = NAND(I4151, I4152)
--	g5926 = NAND(g5741, g639)
--	g3511 = NAND(g3158, g3002, g2976, g2968)
--	I7439 = NAND(g5515, g594)
--	I2090 = NAND(g33, I2089)
--	g5862 = NAND(g5649, g1529, g1535, g2068)
--	I9050 = NAND(g6832, g3598)
--	I5766 = NAND(g3961, g3957)
--	g1582 = NAND(g784, g774, g821)
--	g1793 = NAND(g94, g1084)
--	g3968 = NAND(I5227, I5228)
--	I7527 = NAND(g49, g5662)
--	I5226 = NAND(g3259, g3263)
--	g4049 = NAND(g3677, g3425)
--	I7224 = NAND(g161, I7223)
--	I5767 = NAND(g3961, I5766)
--	I5535 = NAND(g3907, g654)
--	I5227 = NAND(g3259, I5226)
--	g5947 = NAND(g5821, g2944)
--	g3742 = NAND(I4920, I4921)
--	g5873 = NAND(g5649, g1017, g1564, g2113)
--	g4504 = NAND(I6027, I6028)
--	I7244 = NAND(g188, g5377)
--	g5869 = NAND(g5649, g1076, g2081)
--	I5188 = NAND(g3589, I5187)
--	g3983 = NAND(I5270, I5271)
--	g4678 = NAND(g2897, g2101, g1514, g4550)
--	g6843 = NAND(I9051, I9052)
--	g3961 = NAND(I5208, I5209)
--	I5308 = NAND(g478, I5307)
--	I2506 = NAND(g1047, g1044)
--	I3445 = NAND(g1689, g729)
--	g2061 = NAND(I3169, I3170)
--	I3169 = NAND(g1540, I3168)
--	g6740 = NAND(g6703, g6457, g4936)
--	I7556 = NAND(g69, I7555)
--	g4007 = NAND(I5308, I5309)
--	I5196 = NAND(g3567, I5195)
--	I7563 = NAND(g74, I7562)
--	g5684 = NAND(I7440, I7441)
--	I2507 = NAND(g1047, I2506)
--	I1995 = NAND(g504, I1994)
--	g2307 = NAND(I3446, I3447)
--	I7237 = NAND(g179, g5374)
--	g2858 = NAND(g1815, g2577)
--	g2757 = NAND(I3934, I3935)
--	I6744 = NAND(g4708, I6743)
--	I4183 = NAND(g2292, I4182)
--	I7557 = NAND(g5674, I7555)
--	I2300 = NAND(g830, I2299)
--	I3188 = NAND(g1716, g791)
--	g5865 = NAND(g5649, g1088, g1076, g2068)
--	I5197 = NAND(g3571, I5195)
--	I4161 = NAND(g619, I4159)
--	I3741 = NAND(g349, I3739)
--	g5019 = NAND(I6660, I6661)
--	I5257 = NAND(g3714, g3719)
--	g3532 = NAND(g3212, g2215, g3007, g2981)
--	I2528 = NAND(g719, I2526)
--	I5301 = NAND(g471, I5300)
--	g1743 = NAND(g1064, g94)
--	g1411 = NAND(g314, g873)
--	g3012 = NAND(I4204, I4205)
--	g5504 = NAND(I7217, I7218)
--	I6175 = NAND(g4236, g571)
--	I3455 = NAND(g1691, g784)
--	I6500 = NAND(g4504, I6499)
--	g1573 = NAND(g729, g719, g766)
--	I3846 = NAND(g284, g2370)
--	I4210 = NAND(g2294, g804)
--	g4803 = NAND(I6474, I6475)
--	g3109 = NAND(g2360, g1064)
--	g2698 = NAND(I3847, I3848)
--	g3957 = NAND(I5196, I5197)
--	I6499 = NAND(g4504, g3541)
--	g4816 = NAND(g996, g4550, g1518, g2073)
--	I3847 = NAND(g284, I3846)
--	I7520 = NAND(g361, g5659)
--	I4784 = NAND(g622, I4782)
--	I1952 = NAND(g524, I1951)
--	g3539 = NAND(g2591, g2215, g2197, g2981)
--	I8202 = NAND(g478, I8201)
--	I1986 = NAND(g508, g224)
--	I2933 = NAND(g1436, g345)
--	I5760 = NAND(g3836, I5759)
--	g4301 = NAND(I5767, I5768)
--	I1970 = NAND(g516, I1969)
--	I7225 = NAND(g5370, I7223)
--	I6660 = NAND(g4762, I6659)
--	g5502 = NAND(I7209, I7210)
--	I3168 = NAND(g1540, g1534)
--	I1987 = NAND(g508, I1986)
--	g1316 = NAND(I2300, I2301)
--	I2674 = NAND(g710, g131)
--	g4669 = NAND(g4550, g1017, g1680, g2897)
--	I3411 = NAND(g1419, g616)
--	I7245 = NAND(g188, I7244)
--	g2607 = NAND(I3740, I3741)
--	g5308 = NAND(I6963, I6964)
--	g2311 = NAND(I3456, I3457)
--	g3535 = NAND(g3216, g2215, g2197, g2968)
--	g5455 = NAND(g2330, g5311)
--	I4782 = NAND(g2846, g622)
--	I9052 = NAND(g3598, I9050)
--	I3126 = NAND(g1279, I3125)
--	I3400 = NAND(g135, I3398)
--	I4526 = NAND(g2909, g646)
--	g5780 = NAND(I7556, I7557)
--	g3246 = NAND(I4527, I4528)
--	g3502 = NAND(g1411, g1402, g2795)
--	g4608 = NAND(I6176, I6177)
--	I4919 = NAND(g3522, g650)
--	g2100 = NAND(g1588, g804, g791)
--	I7230 = NAND(g170, g5372)
--	I7433 = NAND(g111, I7432)
--	I3127 = NAND(g1276, I3125)
--	g3028 = NAND(I4234, I4235)
--	I2795 = NAND(g804, g798)
--	I5784 = NAND(g628, I5782)
--	I4527 = NAND(g2909, I4526)
--	I7550 = NAND(g5672, I7548)
--	I4546 = NAND(g2853, I4545)
--	I6745 = NAND(g582, I6743)
--	I5294 = NAND(g625, I5292)
--	I6963 = NAND(g4874, I6962)
--	g3741 = NAND(g901, g3433, g2340)
--	g1157 = NAND(g89, g107)
--	I2499 = NAND(g1036, I2497)
--	g937 = NAND(I1979, I1980)
--	g4472 = NAND(g3380, g4253)
--	g2010 = NAND(g1473, g1470, g1459)
--	g928 = NAND(I1962, I1963)
--	I7097 = NAND(g5194, g574)
--	I4547 = NAND(g353, I4545)
--	I3697 = NAND(g1570, g642)
--	I3914 = NAND(g287, g2449)
--	I2543 = NAND(g821, I2542)
--	I3413 = NAND(g616, I3411)
--	I7218 = NAND(g5368, I7216)
--	I7312 = NAND(g5364, I7311)
--	g3538 = NAND(g2588, g2215, g2197, g2179)
--	g5505 = NAND(I7224, I7225)
--	g1075 = NAND(I2109, I2110)
--	I2014 = NAND(g532, I2013)
--	g2804 = NAND(I4009, I4010)
--	g6742 = NAND(g6683, g932, g6716)
--	I6185 = NAND(g4301, g3955)
--	g5863 = NAND(g5649, g1076, g1535, g2068)
--	I3739 = NAND(g2021, g349)
--	I2022 = NAND(g528, I2021)
--	I5782 = NAND(g3810, g628)
--	I7576 = NAND(g84, g5680)
--	g5688 = NAND(g5546, g1585, g2084, g2916)
--	g5857 = NAND(g5638, g1552, g1017, g2062)
--	I3190 = NAND(g791, I3188)
--	I5292 = NAND(g3421, g625)
--	g1764 = NAND(I2796, I2797)
--	I3954 = NAND(g2497, I3952)
--	g5779 = NAND(I7549, I7550)
--	I7577 = NAND(g84, I7576)
--	I5647 = NAND(g3974, g3968)
--	g3531 = NAND(g3209, g2215, g2976, g2179)
--	I1980 = NAND(g230, I1978)
--	g5508 = NAND(I7245, I7246)
--	I4150 = NAND(g2551, g139)
--	g6873 = NAND(g6848, g3621)
--	g6095 = NAND(g2952, g5854)
--	I4009 = NAND(g292, I4008)
--	I2675 = NAND(g710, I2674)
--	g926 = NAND(I1952, I1953)
--	I3894 = NAND(g286, I3893)
--	I4212 = NAND(g804, I4210)
--	g5565 = NAND(I7312, I7313)
--	I6028 = NAND(g4221, I6026)
--	I2109 = NAND(g602, I2108)
--	I5244 = NAND(g3247, I5242)
--	g1402 = NAND(g310, g866, g873)
--	I4921 = NAND(g650, I4919)
--	I7536 = NAND(g5666, I7534)
--	I7223 = NAND(g161, g5370)
--	I2498 = NAND(g1042, I2497)
--	I1951 = NAND(g524, g248)
--	I7522 = NAND(g5659, I7520)
--	I3952 = NAND(g289, g2497)
--	g5775 = NAND(I7521, I7522)
--	I8201 = NAND(g478, g6192)
--	g2024 = NAND(I3126, I3127)
--	g2795 = NAND(g1997, g866)
--	g4004 = NAND(I5301, I5302)
--	I6196 = NAND(g631, I6194)
--	I3970 = NAND(g290, g2518)
--	I4941 = NAND(g357, I4939)
--	I5657 = NAND(g3983, g3979)
--	I7542 = NAND(g59, I7541)
--	I2897 = NAND(g1027, g634)
--	I2682 = NAND(g918, I2681)
--	I2766 = NAND(g749, g743)
--	g3013 = NAND(I4211, I4212)
--	I5242 = NAND(g3242, g3247)
--	I7529 = NAND(g5662, I7527)
--	g1822 = NAND(g1070, g1084)
--	I3876 = NAND(g2397, I3874)
--	I2091 = NAND(g29, I2089)
--	I3915 = NAND(g287, I3914)
--	I9051 = NAND(g6832, I9050)
--	I2767 = NAND(g749, I2766)
--	I1979 = NAND(g512, I1978)
--	g3597 = NAND(I4783, I4784)
--	g2831 = NAND(g2007, g862, g1784)
--	g5683 = NAND(I7433, I7434)
--	g5778 = NAND(I7542, I7543)
--	I2015 = NAND(g260, I2013)
--	g930 = NAND(I1970, I1971)
--	g5782 = NAND(I7570, I7571)
--	g4002 = NAND(I5293, I5294)
--	I2246 = NAND(g598, I2244)
--	I6743 = NAND(g4708, g582)
--	I7549 = NAND(g64, I7548)
--	g2947 = NAND(g1411, g2026)
--	g4762 = NAND(I6391, I6392)
--	g2095 = NAND(g1584, g749, g736)
--	g944 = NAND(I2004, I2005)
--	I6474 = NAND(g4541, I6473)
--	I7232 = NAND(g5372, I7230)
--	I1953 = NAND(g248, I1951)
--	g2719 = NAND(I3875, I3876)
--	I8203 = NAND(g6192, I8201)
--	I4008 = NAND(g292, g2568)
--	g4237 = NAND(g4049, g4017)
--	g1829 = NAND(I2898, I2899)
--	g901 = NAND(g314, g310)
--	g941 = NAND(I1995, I1996)
--	I7570 = NAND(g79, I7569)
--	I2108 = NAND(g602, g610)
--	g1540 = NAND(I2507, I2508)
--	g4814 = NAND(g4550, g1575, g1550, g2073)
--	I7311 = NAND(g5364, g590)
--	I5270 = NAND(g3705, I5269)
--	g2745 = NAND(I3915, I3916)
--	g1797 = NAND(g98, g1064, g1070)
--	g2791 = NAND(I3989, I3990)
--	I7239 = NAND(g5374, I7237)
--	g3526 = NAND(g3196, g3023, g2197, g2981)
--	g6741 = NAND(g6705, g6461, g4941)
--	I8196 = NAND(g6188, I8194)
--	I3895 = NAND(g2422, I3893)
--	I4783 = NAND(g2846, I4782)
--	I2021 = NAND(g528, g254)
--	g905 = NAND(g301, g319)
--	g3276 = NAND(I4546, I4547)
--	g6774 = NAND(g6754, g6750)
--	I5207 = NAND(g3267, g3271)
--	I2301 = NAND(g341, I2299)
--	I5259 = NAND(g3719, I5257)
--	I7440 = NAND(g5515, I7439)
--	I7528 = NAND(g49, I7527)
--	g4640 = NAND(g4402, g1056)
--	g4812 = NAND(g4550, g1560, g1559, g2073)
--	g1845 = NAND(I2934, I2935)
--	g6397 = NAND(I8202, I8203)
--	I5768 = NAND(g3957, I5766)
--	I1978 = NAND(g512, g230)
--	g4610 = NAND(I6186, I6187)
--	I5228 = NAND(g3263, I5226)
--	I2074 = NAND(g11, I2072)
--	g3140 = NAND(g2409, g1060, g1620)
--	I6390 = NAND(g4504, g4610)
--	I3177 = NAND(g1706, g736)
--	I4152 = NAND(g139, I4150)
--	I6501 = NAND(g3541, I6499)
--	I7548 = NAND(g64, g5672)
--	g1815 = NAND(g102, g1070)
--	I7555 = NAND(g69, g5674)
--	g3517 = NAND(g3173, g3002, g2976, g2179)
--	I2080 = NAND(g25, g19)
--	I4211 = NAND(g2294, I4210)
--	I3399 = NAND(g1826, I3398)
--	I5195 = NAND(g3567, g3571)
--	I7313 = NAND(g590, I7311)
--	g2582 = NAND(I3698, I3699)
--	I4939 = NAND(g3437, g357)
--	g950 = NAND(I2022, I2023)
--	g4819 = NAND(I6500, I6501)
--	I7521 = NAND(g361, I7520)
--	I2023 = NAND(g254, I2021)
--	I4446 = NAND(g606, I4444)
--	I5783 = NAND(g3810, I5782)
--	g2940 = NAND(g197, g2381)
--	g4825 = NAND(g4472, g4465)
--	I5293 = NAND(g3421, I5292)
--	I5761 = NAND(g3503, I5759)
--	I1971 = NAND(g236, I1969)
--	I3972 = NAND(g2518, I3970)
--	I4159 = NAND(g2015, g619)
--	I6661 = NAND(g3541, I6659)
--	g1398 = NAND(g306, g889)
--	I6475 = NAND(g578, I6473)
--	I3934 = NAND(g288, I3933)
--	I7541 = NAND(g59, g5669)
--	I2508 = NAND(g1044, I2506)
--	g5854 = NAND(g5638, g1683, g1552, g2062)
--	g4465 = NAND(g319, g4253)
--	I2072 = NAND(g15, g11)
--	I7238 = NAND(g179, I7237)
--	g3955 = NAND(I5188, I5189)
--	I7209 = NAND(g143, I7208)
--	g5431 = NAND(I7098, I7099)
--	I2681 = NAND(g918, g613)
--	I2013 = NAND(g532, g260)
--	I4234 = NAND(g2267, I4233)
--	g2780 = NAND(I3971, I3972)
--	g2067 = NAND(I3178, I3179)
--	I1962 = NAND(g520, I1961)
--	I5258 = NAND(g3714, I5257)
--	g1387 = NAND(g862, g314, g301)
--	I2060 = NAND(g7, g3)
--	g5781 = NAND(I7563, I7564)
--	g2263 = NAND(I3399, I3400)
--	g4221 = NAND(I5648, I5649)
--	g1359 = NAND(g866, g306)
--	I7231 = NAND(g170, I7230)
--	I3953 = NAND(g289, I3952)
--	I5187 = NAND(g3589, g3593)
--	g5852 = NAND(g5638, g2053, g1661)
--	g3520 = NAND(g3183, g3002, g2197, g2968)
--	g1047 = NAND(I2090, I2091)
--	I7099 = NAND(g574, I7097)
--	I3848 = NAND(g2370, I3846)
--	I3699 = NAND(g642, I3697)
--	I3398 = NAND(g1826, g135)
--	I1969 = NAND(g516, g236)
--	I5307 = NAND(g478, g3512)
--	g3974 = NAND(I5243, I5244)
--	I5536 = NAND(g3907, I5535)
--	g1417 = NAND(g873, g889)
--	I7543 = NAND(g5669, I7541)
--	g5943 = NAND(g5818, g2940)
--	I7534 = NAND(g54, g5666)
--	g4319 = NAND(I5783, I5784)
--	I3893 = NAND(g286, g2422)
--	g2080 = NAND(I3189, I3190)
--	I2683 = NAND(g613, I2681)
--	I5537 = NAND(g654, I5535)
--	I3170 = NAND(g1534, I3168)
--	I3125 = NAND(g1279, g1276)
--	I5243 = NAND(g3242, I5242)
--	I1988 = NAND(g224, I1986)
--	I6194 = NAND(g4199, g631)
--	g3207 = NAND(I4445, I4446)
--	I2526 = NAND(g766, g719)
--	g6929 = NAND(g4536, g6927)
--	g3215 = NAND(g2340, g1402)
--	I3446 = NAND(g1689, I3445)
--	I7208 = NAND(g143, g5367)
--	g5783 = NAND(I7577, I7578)
--	I4545 = NAND(g2853, g353)
--	I2004 = NAND(g500, I2003)
--	I2527 = NAND(g766, I2526)
--	I5649 = NAND(g3968, I5647)
--	g6778 = NAND(g6762, g6758)
--	g1686 = NAND(I2675, I2676)
--	g4223 = NAND(I5658, I5659)
--	I1996 = NAND(g218, I1994)
--	I3447 = NAND(g729, I3445)
--	I4204 = NAND(g2255, I4203)
--	I3874 = NAND(g285, g2397)
--	g2944 = NAND(g269, g2381)
--	g1253 = NAND(I2245, I2246)
--	g2434 = NAND(g1064, g1070, g1620)
--	I2299 = NAND(g830, g341)
--	g5866 = NAND(g5649, g1529, g2081)
--	g1687 = NAND(I2682, I2683)
--	I3935 = NAND(g2473, I3933)
--	g4017 = NAND(g107, g3425)
--	I4528 = NAND(g646, I4526)
--	I2244 = NAND(g567, g598)
--	I4151 = NAND(g2551, I4150)
--	I6392 = NAND(g4610, I6390)
--	I4010 = NAND(g2568, I4008)
--	I2082 = NAND(g19, I2080)
--	g5818 = NAND(g5638, g2056, g1666, g1661)
--	g3979 = NAND(I5258, I5259)
--	I6176 = NAND(g4236, I6175)
--	I4235 = NAND(g798, I4233)
--	I2110 = NAND(g610, I2108)
--	I7098 = NAND(g5194, I7097)
--	I3456 = NAND(g1691, I3455)
--	g5821 = NAND(g5638, g2056, g1076, g1666)
--	I3698 = NAND(g1570, I3697)
--	g2995 = NAND(I4183, I4184)
--	I6473 = NAND(g4541, g578)
--	I5659 = NAND(g3979, I5657)
--	g5636 = NAND(g5564, g4769)
--	I6177 = NAND(g571, I6175)
--	I2899 = NAND(g634, I2897)
--	I3457 = NAND(g784, I3455)
--	I3989 = NAND(g291, I3988)
--	I3971 = NAND(g290, I3970)
--	I4160 = NAND(g2015, I4159)
--	I2089 = NAND(g33, g29)
--	g4670 = NAND(g4611, g3528)
--	g4813 = NAND(g4550, g965, g1560, g2073)
--	I3740 = NAND(g2021, I3739)
--	I8194 = NAND(g471, g6188)
--	I5300 = NAND(g471, g3505)
--	g3893 = NAND(g3664, g3656, g3647)
--	g6928 = NAND(g4532, g6926)
--	I7578 = NAND(g5680, I7576)
--	I7535 = NAND(g54, I7534)
--	I1961 = NAND(g520, g242)
--	g3544 = NAND(g2594, g2215, g2197, g2179)
--	g6394 = NAND(I8195, I8196)
--	I5648 = NAND(g3974, I5647)
--	I7246 = NAND(g5377, I7244)
--	g3756 = NAND(I4940, I4941)
--	I2062 = NAND(g3, I2060)
--	I6195 = NAND(g4199, I6194)
--	I7216 = NAND(g152, g5368)
--	g3536 = NAND(g3219, g2215, g3007, g2179)
--	I7564 = NAND(g5676, I7562)
--	g4300 = NAND(I5760, I5761)
--	I4184 = NAND(g749, I4182)
--	I2005 = NAND(g212, I2003)
--	g5318 = NAND(g676, g5060)
--	g5872 = NAND(g5649, g1557, g1564, g2113)
--	
--	g5552 = NOR(g5354, g5356)
--	g4235 = NOR(g3780, g3362)
--	g6073 = NOR(g197, g5862)
--	g4776 = NOR(g4449, g4453)
--	g4777 = NOR(g4457, g4459)
--	g4238 = NOR(g3755, g3279)
--	g6433 = NOR(g6385, g3733, g4092, g4314)
--	g6496 = NOR(g952, g6354)
--	g1422 = NOR(g1039, g913)
--	g3931 = NOR(g3353, g3361)
--	g1560 = NOR(g996, g980)
--	g3905 = NOR(g3512, g478)
--	g5094 = NOR(g4685, g4686)
--	g3973 = NOR(g3368, g3374)
--	g3528 = NOR(g1802, g3167)
--	g5541 = NOR(g5388, g1880)
--	g3621 = NOR(g1407, g2842)
--	g1449 = NOR(g489, g1048)
--	g3965 = NOR(g3359, g3367)
--	g3933 = NOR(g3327, g3336)
--	g6280 = NOR(I7978, I7979, I7980, I7981)
--	g2433 = NOR(g1418, g1449)
--	g1470 = NOR(g937, g930, g928)
--	g6427 = NOR(g6376, g4086, g4074, g4068)
--	g6446 = NOR(g6385, g4334, g4092, g4314)
--	g6359 = NOR(I8135, I8136, I8137, I8138)
--	g1459 = NOR(g926, g950, g948)
--	g4584 = NOR(g4164, g4168)
--	g3926 = NOR(g3338, g3350)
--	g6279 = NOR(I7969, I7970, I7971, I7972)
--	g5265 = NOR(g4863, g4865)
--	g3927 = NOR(g3382, g3383)
--	g3903 = NOR(g3505, g471)
--	g1418 = NOR(g486, g943)
--	g4578 = NOR(g4234, g3928)
--	g4261 = NOR(g3762, g3295)
--	g6358 = NOR(I8126, I8127, I8128, I8129)
--	g4589 = NOR(g4180, g4183)
--	g1474 = NOR(g760, g754)
--	g3956 = NOR(g3337, g3349)
--	g4774 = NOR(g4442, g4445)
--	g5091 = NOR(g4698, g4701)
--	g4950 = NOR(g1472, g4680)
--	g5227 = NOR(g5019, g3559)
--	g4585 = NOR(g4171, g4177)
--	g6494 = NOR(g952, g6348)
--	g5048 = NOR(g4819, g3491, g3559)
--	g3664 = NOR(g2804, g2791, g2780)
--	g4000 = NOR(g1250, g3425)
--	g5418 = NOR(g5162, g5169)
--	g5093 = NOR(g4683, g4684)
--	g4779 = NOR(g4461, g4464)
--	g6492 = NOR(g6348, g1734)
--	g4240 = NOR(g1589, g1879, g3793)
--	g4596 = NOR(g4184, g4186)
--	g1603 = NOR(g1039, g658)
--	g2908 = NOR(g536, g2010, g541)
--	g4581 = NOR(g4156, g4160)
--	g5423 = NOR(g5170, g5175)
--	g4432 = NOR(g923, g4253)
--	g6436 = NOR(g6385, g3733, g4328, g4080)
--	g4568 = NOR(g4233, g3924)
--	g6335 = NOR(I8079, I8080, I8081, I8082)
--	g5753 = NOR(g1477, g5688)
--	g6495 = NOR(g6354, g1775)
--	g6442 = NOR(g6376, g4323, g4074, g4302)
--	g6429 = NOR(g6376, g4086, g4074, g4302)
--	g6281 = NOR(I7987, I7988, I7989, I7990)
--	g6449 = NOR(g6385, g4334, g4328, g4080)
--	g4590 = NOR(g4169, g4172)
--	g4877 = NOR(g952, g4680)
--	g6445 = NOR(g6376, g4323, g4309, g4068)
--	g5561 = NOR(g5391, g1589, g3793, g1880)
--	g3929 = NOR(g3373, g3376)
--	g1473 = NOR(g944, g941, g939)
--	g4967 = NOR(g4674, g952)
--	g6430 = NOR(g6385, g3733, g4092, g4080)
--	g4993 = NOR(g4674, g1477)
--	g6448 = NOR(g6376, g4323, g4309, g4302)
--	g3647 = NOR(g2731, g2719, g2698)
--	g3925 = NOR(g3303, g3315)
--	g5731 = NOR(g952, g5688)
--	g3959 = NOR(g3352, g3360)
--	g1481 = NOR(g815, g809)
--	g3656 = NOR(g2769, g2757, g2745)
--	g4245 = NOR(g3759, g3288)
--	g3930 = NOR(g3317, g3328)
--	g5249 = NOR(g4868, g4870)
--	g3966 = NOR(g3329, g3339)
--	g6400 = NOR(I8208, I8209, I8210, I8211)
--	g4266 = NOR(g3757, g3283)
--	g6451 = NOR(g6385, g4334, g4328, g4314)
--	g5324 = NOR(g5069, g4410, g766)
--	g6443 = NOR(g6385, g4334, g4092, g4080)
--	g5088 = NOR(g4691, g4697)
--	g3958 = NOR(g3316, g3326)
--	g4241 = NOR(g3774, g3341)
--	g6432 = NOR(g6376, g4086, g4309, g4068)
--	g6357 = NOR(I8117, I8118, I8119, I8120)
--	g3923 = NOR(g3378, g3381)
--	g6075 = NOR(g269, g5863)
--	g3934 = NOR(g3377, g3379)
--	g6439 = NOR(g6385, g3733, g4328, g4314)
--	g4272 = NOR(g3767, g3319)
--	g1879 = NOR(g1603, g1416)
--	g5325 = NOR(g5077, g4416, g821)
--	g6435 = NOR(g6376, g4086, g4309, g4302)
--	g4586 = NOR(g4161, g4165)
--	g3939 = NOR(g3340, g3351)
--	g6438 = NOR(g6376, g4323, g4074, g4068)
--	g1518 = NOR(g980, g965)
--	g4239 = NOR(g3763, g3296)
--	g4591 = NOR(g4178, g4181)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s9234 is
	port (
		CLK: in std_logic;
		G22: in std_logic;
		G23: in std_logic;
		G32: in std_logic;
		G36: in std_logic;
		G37: in std_logic;
		G38: in std_logic;
		G39: in std_logic;
		G40: in std_logic;
		G41: in std_logic;
		G42: in std_logic;
		G44: in std_logic;
		G45: in std_logic;
		G46: in std_logic;
		G47: in std_logic;
		G89: in std_logic;
		G94: in std_logic;
		G98: in std_logic;
		G102: in std_logic;
		G107: in std_logic;
		G301: in std_logic;
		G306: in std_logic;
		G310: in std_logic;
		G314: in std_logic;
		G319: in std_logic;
		G557: in std_logic;
		G558: in std_logic;
		G559: in std_logic;
		G560: in std_logic;
		G561: in std_logic;
		G562: in std_logic;
		G563: in std_logic;
		G564: in std_logic;
		G567: in std_logic;
		G639: in std_logic;
		G702: in std_logic;
		G705: in std_logic;
		G1290: out std_logic;
		G1293: out std_logic;
		G2584: out std_logic;
		G3222: out std_logic;
		G3600: out std_logic;
		G4098: out std_logic;
		G4099: out std_logic;
		G4100: out std_logic;
		G4101: out std_logic;
		G4102: out std_logic;
		G4103: out std_logic;
		G4104: out std_logic;
		G4105: out std_logic;
		G4106: out std_logic;
		G4107: out std_logic;
		G4108: out std_logic;
		G4109: out std_logic;
		G4110: out std_logic;
		G4112: out std_logic;
		G4121: out std_logic;
		G4307: out std_logic;
		G4321: out std_logic;
		G4422: out std_logic;
		G4809: out std_logic;
		G5137: out std_logic;
		G5468: out std_logic;
		G5469: out std_logic;
		G5692: out std_logic;
		G6282: out std_logic;
		G6284: out std_logic;
		G6360: out std_logic;
		G6362: out std_logic;
		G6364: out std_logic;
		G6366: out std_logic;
		G6368: out std_logic;
		G6370: out std_logic;
		G6372: out std_logic;
		G6374: out std_logic;
		G6728: out std_logic
	);
end entity;

architecture RTL of s9234 is
	attribute dont_touch: boolean;

	signal G1: std_logic; attribute dont_touch of G1: signal is true;
	signal G2: std_logic; attribute dont_touch of G2: signal is true;
	signal G3: std_logic; attribute dont_touch of G3: signal is true;
	signal G6: std_logic; attribute dont_touch of G6: signal is true;
	signal G7: std_logic; attribute dont_touch of G7: signal is true;
	signal G10: std_logic; attribute dont_touch of G10: signal is true;
	signal G11: std_logic; attribute dont_touch of G11: signal is true;
	signal G14: std_logic; attribute dont_touch of G14: signal is true;
	signal G15: std_logic; attribute dont_touch of G15: signal is true;
	signal G18: std_logic; attribute dont_touch of G18: signal is true;
	signal G19: std_logic; attribute dont_touch of G19: signal is true;
	signal G24: std_logic; attribute dont_touch of G24: signal is true;
	signal G25: std_logic; attribute dont_touch of G25: signal is true;
	signal G28: std_logic; attribute dont_touch of G28: signal is true;
	signal G29: std_logic; attribute dont_touch of G29: signal is true;
	signal G33: std_logic; attribute dont_touch of G33: signal is true;
	signal G43: std_logic; attribute dont_touch of G43: signal is true;
	signal G48: std_logic; attribute dont_touch of G48: signal is true;
	signal G49: std_logic; attribute dont_touch of G49: signal is true;
	signal G54: std_logic; attribute dont_touch of G54: signal is true;
	signal G59: std_logic; attribute dont_touch of G59: signal is true;
	signal G64: std_logic; attribute dont_touch of G64: signal is true;
	signal G69: std_logic; attribute dont_touch of G69: signal is true;
	signal G74: std_logic; attribute dont_touch of G74: signal is true;
	signal G79: std_logic; attribute dont_touch of G79: signal is true;
	signal G84: std_logic; attribute dont_touch of G84: signal is true;
	signal G111: std_logic; attribute dont_touch of G111: signal is true;
	signal G114: std_logic; attribute dont_touch of G114: signal is true;
	signal G117: std_logic; attribute dont_touch of G117: signal is true;
	signal G118: std_logic; attribute dont_touch of G118: signal is true;
	signal G119: std_logic; attribute dont_touch of G119: signal is true;
	signal G122: std_logic; attribute dont_touch of G122: signal is true;
	signal G123: std_logic; attribute dont_touch of G123: signal is true;
	signal G127: std_logic; attribute dont_touch of G127: signal is true;
	signal G128: std_logic; attribute dont_touch of G128: signal is true;
	signal G131: std_logic; attribute dont_touch of G131: signal is true;
	signal G135: std_logic; attribute dont_touch of G135: signal is true;
	signal G139: std_logic; attribute dont_touch of G139: signal is true;
	signal G143: std_logic; attribute dont_touch of G143: signal is true;
	signal G148: std_logic; attribute dont_touch of G148: signal is true;
	signal G152: std_logic; attribute dont_touch of G152: signal is true;
	signal G157: std_logic; attribute dont_touch of G157: signal is true;
	signal G161: std_logic; attribute dont_touch of G161: signal is true;
	signal G166: std_logic; attribute dont_touch of G166: signal is true;
	signal G170: std_logic; attribute dont_touch of G170: signal is true;
	signal G175: std_logic; attribute dont_touch of G175: signal is true;
	signal G179: std_logic; attribute dont_touch of G179: signal is true;
	signal G184: std_logic; attribute dont_touch of G184: signal is true;
	signal G188: std_logic; attribute dont_touch of G188: signal is true;
	signal G193: std_logic; attribute dont_touch of G193: signal is true;
	signal G197: std_logic; attribute dont_touch of G197: signal is true;
	signal G204: std_logic; attribute dont_touch of G204: signal is true;
	signal G205: std_logic; attribute dont_touch of G205: signal is true;
	signal G206: std_logic; attribute dont_touch of G206: signal is true;
	signal G207: std_logic; attribute dont_touch of G207: signal is true;
	signal G208: std_logic; attribute dont_touch of G208: signal is true;
	signal G209: std_logic; attribute dont_touch of G209: signal is true;
	signal G210: std_logic; attribute dont_touch of G210: signal is true;
	signal G211: std_logic; attribute dont_touch of G211: signal is true;
	signal G212: std_logic; attribute dont_touch of G212: signal is true;
	signal G218: std_logic; attribute dont_touch of G218: signal is true;
	signal G224: std_logic; attribute dont_touch of G224: signal is true;
	signal G230: std_logic; attribute dont_touch of G230: signal is true;
	signal G236: std_logic; attribute dont_touch of G236: signal is true;
	signal G242: std_logic; attribute dont_touch of G242: signal is true;
	signal G248: std_logic; attribute dont_touch of G248: signal is true;
	signal G254: std_logic; attribute dont_touch of G254: signal is true;
	signal G260: std_logic; attribute dont_touch of G260: signal is true;
	signal G266: std_logic; attribute dont_touch of G266: signal is true;
	signal G269: std_logic; attribute dont_touch of G269: signal is true;
	signal G276: std_logic; attribute dont_touch of G276: signal is true;
	signal G277: std_logic; attribute dont_touch of G277: signal is true;
	signal G278: std_logic; attribute dont_touch of G278: signal is true;
	signal G279: std_logic; attribute dont_touch of G279: signal is true;
	signal G280: std_logic; attribute dont_touch of G280: signal is true;
	signal G281: std_logic; attribute dont_touch of G281: signal is true;
	signal G282: std_logic; attribute dont_touch of G282: signal is true;
	signal G283: std_logic; attribute dont_touch of G283: signal is true;
	signal G284: std_logic; attribute dont_touch of G284: signal is true;
	signal G285: std_logic; attribute dont_touch of G285: signal is true;
	signal G286: std_logic; attribute dont_touch of G286: signal is true;
	signal G287: std_logic; attribute dont_touch of G287: signal is true;
	signal G288: std_logic; attribute dont_touch of G288: signal is true;
	signal G289: std_logic; attribute dont_touch of G289: signal is true;
	signal G290: std_logic; attribute dont_touch of G290: signal is true;
	signal G291: std_logic; attribute dont_touch of G291: signal is true;
	signal G292: std_logic; attribute dont_touch of G292: signal is true;
	signal G293: std_logic; attribute dont_touch of G293: signal is true;
	signal G297: std_logic; attribute dont_touch of G297: signal is true;
	signal G323: std_logic; attribute dont_touch of G323: signal is true;
	signal G326: std_logic; attribute dont_touch of G326: signal is true;
	signal G327: std_logic; attribute dont_touch of G327: signal is true;
	signal G328: std_logic; attribute dont_touch of G328: signal is true;
	signal G331: std_logic; attribute dont_touch of G331: signal is true;
	signal G332: std_logic; attribute dont_touch of G332: signal is true;
	signal G336: std_logic; attribute dont_touch of G336: signal is true;
	signal G337: std_logic; attribute dont_touch of G337: signal is true;
	signal G338: std_logic; attribute dont_touch of G338: signal is true;
	signal G341: std_logic; attribute dont_touch of G341: signal is true;
	signal G345: std_logic; attribute dont_touch of G345: signal is true;
	signal G349: std_logic; attribute dont_touch of G349: signal is true;
	signal G353: std_logic; attribute dont_touch of G353: signal is true;
	signal G357: std_logic; attribute dont_touch of G357: signal is true;
	signal G361: std_logic; attribute dont_touch of G361: signal is true;
	signal G366: std_logic; attribute dont_touch of G366: signal is true;
	signal G370: std_logic; attribute dont_touch of G370: signal is true;
	signal G374: std_logic; attribute dont_touch of G374: signal is true;
	signal G378: std_logic; attribute dont_touch of G378: signal is true;
	signal G382: std_logic; attribute dont_touch of G382: signal is true;
	signal G386: std_logic; attribute dont_touch of G386: signal is true;
	signal G390: std_logic; attribute dont_touch of G390: signal is true;
	signal G394: std_logic; attribute dont_touch of G394: signal is true;
	signal G398: std_logic; attribute dont_touch of G398: signal is true;
	signal G402: std_logic; attribute dont_touch of G402: signal is true;
	signal G406: std_logic; attribute dont_touch of G406: signal is true;
	signal G410: std_logic; attribute dont_touch of G410: signal is true;
	signal G414: std_logic; attribute dont_touch of G414: signal is true;
	signal G418: std_logic; attribute dont_touch of G418: signal is true;
	signal G422: std_logic; attribute dont_touch of G422: signal is true;
	signal G426: std_logic; attribute dont_touch of G426: signal is true;
	signal G430: std_logic; attribute dont_touch of G430: signal is true;
	signal G434: std_logic; attribute dont_touch of G434: signal is true;
	signal G437: std_logic; attribute dont_touch of G437: signal is true;
	signal G441: std_logic; attribute dont_touch of G441: signal is true;
	signal G445: std_logic; attribute dont_touch of G445: signal is true;
	signal G449: std_logic; attribute dont_touch of G449: signal is true;
	signal G453: std_logic; attribute dont_touch of G453: signal is true;
	signal G457: std_logic; attribute dont_touch of G457: signal is true;
	signal G461: std_logic; attribute dont_touch of G461: signal is true;
	signal G465: std_logic; attribute dont_touch of G465: signal is true;
	signal G471: std_logic; attribute dont_touch of G471: signal is true;
	signal G478: std_logic; attribute dont_touch of G478: signal is true;
	signal G485: std_logic; attribute dont_touch of G485: signal is true;
	signal G486: std_logic; attribute dont_touch of G486: signal is true;
	signal G489: std_logic; attribute dont_touch of G489: signal is true;
	signal G492: std_logic; attribute dont_touch of G492: signal is true;
	signal G496: std_logic; attribute dont_touch of G496: signal is true;
	signal G500: std_logic; attribute dont_touch of G500: signal is true;
	signal G504: std_logic; attribute dont_touch of G504: signal is true;
	signal G508: std_logic; attribute dont_touch of G508: signal is true;
	signal G512: std_logic; attribute dont_touch of G512: signal is true;
	signal G516: std_logic; attribute dont_touch of G516: signal is true;
	signal G520: std_logic; attribute dont_touch of G520: signal is true;
	signal G524: std_logic; attribute dont_touch of G524: signal is true;
	signal G528: std_logic; attribute dont_touch of G528: signal is true;
	signal G532: std_logic; attribute dont_touch of G532: signal is true;
	signal G536: std_logic; attribute dont_touch of G536: signal is true;
	signal G541: std_logic; attribute dont_touch of G541: signal is true;
	signal G545: std_logic; attribute dont_touch of G545: signal is true;
	signal G548: std_logic; attribute dont_touch of G548: signal is true;
	signal G551: std_logic; attribute dont_touch of G551: signal is true;
	signal G554: std_logic; attribute dont_touch of G554: signal is true;
	signal G571: std_logic; attribute dont_touch of G571: signal is true;
	signal G574: std_logic; attribute dont_touch of G574: signal is true;
	signal G578: std_logic; attribute dont_touch of G578: signal is true;
	signal G582: std_logic; attribute dont_touch of G582: signal is true;
	signal G586: std_logic; attribute dont_touch of G586: signal is true;
	signal G590: std_logic; attribute dont_touch of G590: signal is true;
	signal G594: std_logic; attribute dont_touch of G594: signal is true;
	signal G598: std_logic; attribute dont_touch of G598: signal is true;
	signal G602: std_logic; attribute dont_touch of G602: signal is true;
	signal G606: std_logic; attribute dont_touch of G606: signal is true;
	signal G610: std_logic; attribute dont_touch of G610: signal is true;
	signal G613: std_logic; attribute dont_touch of G613: signal is true;
	signal G616: std_logic; attribute dont_touch of G616: signal is true;
	signal G619: std_logic; attribute dont_touch of G619: signal is true;
	signal G622: std_logic; attribute dont_touch of G622: signal is true;
	signal G625: std_logic; attribute dont_touch of G625: signal is true;
	signal G628: std_logic; attribute dont_touch of G628: signal is true;
	signal G631: std_logic; attribute dont_touch of G631: signal is true;
	signal G634: std_logic; attribute dont_touch of G634: signal is true;
	signal G638: std_logic; attribute dont_touch of G638: signal is true;
	signal G642: std_logic; attribute dont_touch of G642: signal is true;
	signal G646: std_logic; attribute dont_touch of G646: signal is true;
	signal G650: std_logic; attribute dont_touch of G650: signal is true;
	signal G654: std_logic; attribute dont_touch of G654: signal is true;
	signal G658: std_logic; attribute dont_touch of G658: signal is true;
	signal G662: std_logic; attribute dont_touch of G662: signal is true;
	signal G663: std_logic; attribute dont_touch of G663: signal is true;
	signal G664: std_logic; attribute dont_touch of G664: signal is true;
	signal G665: std_logic; attribute dont_touch of G665: signal is true;
	signal G666: std_logic; attribute dont_touch of G666: signal is true;
	signal G667: std_logic; attribute dont_touch of G667: signal is true;
	signal G668: std_logic; attribute dont_touch of G668: signal is true;
	signal G669: std_logic; attribute dont_touch of G669: signal is true;
	signal G672: std_logic; attribute dont_touch of G672: signal is true;
	signal G675: std_logic; attribute dont_touch of G675: signal is true;
	signal G676: std_logic; attribute dont_touch of G676: signal is true;
	signal G677: std_logic; attribute dont_touch of G677: signal is true;
	signal G678: std_logic; attribute dont_touch of G678: signal is true;
	signal G679: std_logic; attribute dont_touch of G679: signal is true;
	signal G680: std_logic; attribute dont_touch of G680: signal is true;
	signal G681: std_logic; attribute dont_touch of G681: signal is true;
	signal G682: std_logic; attribute dont_touch of G682: signal is true;
	signal G683: std_logic; attribute dont_touch of G683: signal is true;
	signal G684: std_logic; attribute dont_touch of G684: signal is true;
	signal G685: std_logic; attribute dont_touch of G685: signal is true;
	signal G686: std_logic; attribute dont_touch of G686: signal is true;
	signal G687: std_logic; attribute dont_touch of G687: signal is true;
	signal G688: std_logic; attribute dont_touch of G688: signal is true;
	signal G689: std_logic; attribute dont_touch of G689: signal is true;
	signal G690: std_logic; attribute dont_touch of G690: signal is true;
	signal G691: std_logic; attribute dont_touch of G691: signal is true;
	signal G692: std_logic; attribute dont_touch of G692: signal is true;
	signal G693: std_logic; attribute dont_touch of G693: signal is true;
	signal G694: std_logic; attribute dont_touch of G694: signal is true;
	signal G695: std_logic; attribute dont_touch of G695: signal is true;
	signal G696: std_logic; attribute dont_touch of G696: signal is true;
	signal G697: std_logic; attribute dont_touch of G697: signal is true;
	signal G698: std_logic; attribute dont_touch of G698: signal is true;
	signal G699: std_logic; attribute dont_touch of G699: signal is true;
	signal G706: std_logic; attribute dont_touch of G706: signal is true;
	signal G709: std_logic; attribute dont_touch of G709: signal is true;
	signal G710: std_logic; attribute dont_touch of G710: signal is true;
	signal G714: std_logic; attribute dont_touch of G714: signal is true;
	signal G715: std_logic; attribute dont_touch of G715: signal is true;
	signal G716: std_logic; attribute dont_touch of G716: signal is true;
	signal G719: std_logic; attribute dont_touch of G719: signal is true;
	signal G729: std_logic; attribute dont_touch of G729: signal is true;
	signal G736: std_logic; attribute dont_touch of G736: signal is true;
	signal G743: std_logic; attribute dont_touch of G743: signal is true;
	signal G749: std_logic; attribute dont_touch of G749: signal is true;
	signal G754: std_logic; attribute dont_touch of G754: signal is true;
	signal G760: std_logic; attribute dont_touch of G760: signal is true;
	signal G766: std_logic; attribute dont_touch of G766: signal is true;
	signal G774: std_logic; attribute dont_touch of G774: signal is true;
	signal G784: std_logic; attribute dont_touch of G784: signal is true;
	signal G791: std_logic; attribute dont_touch of G791: signal is true;
	signal G798: std_logic; attribute dont_touch of G798: signal is true;
	signal G804: std_logic; attribute dont_touch of G804: signal is true;
	signal G809: std_logic; attribute dont_touch of G809: signal is true;
	signal G815: std_logic; attribute dont_touch of G815: signal is true;
	signal G821: std_logic; attribute dont_touch of G821: signal is true;
	signal G829: std_logic; attribute dont_touch of G829: signal is true;
	signal G830: std_logic; attribute dont_touch of G830: signal is true;
	signal G834: std_logic; attribute dont_touch of G834: signal is true;
	signal G835: std_logic; attribute dont_touch of G835: signal is true;
	signal G836: std_logic; attribute dont_touch of G836: signal is true;
	signal G837: std_logic; attribute dont_touch of G837: signal is true;
	signal G838: std_logic; attribute dont_touch of G838: signal is true;
	signal G839: std_logic; attribute dont_touch of G839: signal is true;
	signal G842: std_logic; attribute dont_touch of G842: signal is true;
	signal G843: std_logic; attribute dont_touch of G843: signal is true;
	signal G844: std_logic; attribute dont_touch of G844: signal is true;
	signal G845: std_logic; attribute dont_touch of G845: signal is true;
	signal G846: std_logic; attribute dont_touch of G846: signal is true;
	signal G847: std_logic; attribute dont_touch of G847: signal is true;
	signal G848: std_logic; attribute dont_touch of G848: signal is true;
	signal G849: std_logic; attribute dont_touch of G849: signal is true;
	signal G850: std_logic; attribute dont_touch of G850: signal is true;
	signal G851: std_logic; attribute dont_touch of G851: signal is true;
	signal G852: std_logic; attribute dont_touch of G852: signal is true;
	signal G853: std_logic; attribute dont_touch of G853: signal is true;
	signal G854: std_logic; attribute dont_touch of G854: signal is true;
	signal G855: std_logic; attribute dont_touch of G855: signal is true;
	signal G856: std_logic; attribute dont_touch of G856: signal is true;
	signal G857: std_logic; attribute dont_touch of G857: signal is true;
	signal G858: std_logic; attribute dont_touch of G858: signal is true;
	signal G861: std_logic; attribute dont_touch of G861: signal is true;
	signal G862: std_logic; attribute dont_touch of G862: signal is true;
	signal G865: std_logic; attribute dont_touch of G865: signal is true;
	signal G866: std_logic; attribute dont_touch of G866: signal is true;
	signal G872: std_logic; attribute dont_touch of G872: signal is true;
	signal G873: std_logic; attribute dont_touch of G873: signal is true;
	signal G878: std_logic; attribute dont_touch of G878: signal is true;
	signal G889: std_logic; attribute dont_touch of G889: signal is true;
	signal G893: std_logic; attribute dont_touch of G893: signal is true;
	signal G894: std_logic; attribute dont_touch of G894: signal is true;
	signal G895: std_logic; attribute dont_touch of G895: signal is true;
	signal G896: std_logic; attribute dont_touch of G896: signal is true;
	signal G897: std_logic; attribute dont_touch of G897: signal is true;
	signal G898: std_logic; attribute dont_touch of G898: signal is true;
	signal G899: std_logic; attribute dont_touch of G899: signal is true;
	signal G900: std_logic; attribute dont_touch of G900: signal is true;
	signal G901: std_logic; attribute dont_touch of G901: signal is true;
	signal G905: std_logic; attribute dont_touch of G905: signal is true;
	signal G908: std_logic; attribute dont_touch of G908: signal is true;
	signal G909: std_logic; attribute dont_touch of G909: signal is true;
	signal G910: std_logic; attribute dont_touch of G910: signal is true;
	signal G913: std_logic; attribute dont_touch of G913: signal is true;
	signal G917: std_logic; attribute dont_touch of G917: signal is true;
	signal G918: std_logic; attribute dont_touch of G918: signal is true;
	signal G921: std_logic; attribute dont_touch of G921: signal is true;
	signal G922: std_logic; attribute dont_touch of G922: signal is true;
	signal G923: std_logic; attribute dont_touch of G923: signal is true;
	signal G926: std_logic; attribute dont_touch of G926: signal is true;
	signal G927: std_logic; attribute dont_touch of G927: signal is true;
	signal G928: std_logic; attribute dont_touch of G928: signal is true;
	signal G929: std_logic; attribute dont_touch of G929: signal is true;
	signal G930: std_logic; attribute dont_touch of G930: signal is true;
	signal G931: std_logic; attribute dont_touch of G931: signal is true;
	signal G932: std_logic; attribute dont_touch of G932: signal is true;
	signal G937: std_logic; attribute dont_touch of G937: signal is true;
	signal G938: std_logic; attribute dont_touch of G938: signal is true;
	signal G939: std_logic; attribute dont_touch of G939: signal is true;
	signal G940: std_logic; attribute dont_touch of G940: signal is true;
	signal G941: std_logic; attribute dont_touch of G941: signal is true;
	signal G942: std_logic; attribute dont_touch of G942: signal is true;
	signal G943: std_logic; attribute dont_touch of G943: signal is true;
	signal G944: std_logic; attribute dont_touch of G944: signal is true;
	signal G945: std_logic; attribute dont_touch of G945: signal is true;
	signal G946: std_logic; attribute dont_touch of G946: signal is true;
	signal G947: std_logic; attribute dont_touch of G947: signal is true;
	signal G948: std_logic; attribute dont_touch of G948: signal is true;
	signal G949: std_logic; attribute dont_touch of G949: signal is true;
	signal G950: std_logic; attribute dont_touch of G950: signal is true;
	signal G951: std_logic; attribute dont_touch of G951: signal is true;
	signal G952: std_logic; attribute dont_touch of G952: signal is true;
	signal G964: std_logic; attribute dont_touch of G964: signal is true;
	signal G965: std_logic; attribute dont_touch of G965: signal is true;
	signal G971: std_logic; attribute dont_touch of G971: signal is true;
	signal G980: std_logic; attribute dont_touch of G980: signal is true;
	signal G985: std_logic; attribute dont_touch of G985: signal is true;
	signal G996: std_logic; attribute dont_touch of G996: signal is true;
	signal G1001: std_logic; attribute dont_touch of G1001: signal is true;
	signal G1006: std_logic; attribute dont_touch of G1006: signal is true;
	signal G1011: std_logic; attribute dont_touch of G1011: signal is true;
	signal G1017: std_logic; attribute dont_touch of G1017: signal is true;
	signal G1027: std_logic; attribute dont_touch of G1027: signal is true;
	signal G1030: std_logic; attribute dont_touch of G1030: signal is true;
	signal G1036: std_logic; attribute dont_touch of G1036: signal is true;
	signal G1037: std_logic; attribute dont_touch of G1037: signal is true;
	signal G1038: std_logic; attribute dont_touch of G1038: signal is true;
	signal G1039: std_logic; attribute dont_touch of G1039: signal is true;
	signal G1042: std_logic; attribute dont_touch of G1042: signal is true;
	signal G1043: std_logic; attribute dont_touch of G1043: signal is true;
	signal G1044: std_logic; attribute dont_touch of G1044: signal is true;
	signal G1045: std_logic; attribute dont_touch of G1045: signal is true;
	signal G1046: std_logic; attribute dont_touch of G1046: signal is true;
	signal G1047: std_logic; attribute dont_touch of G1047: signal is true;
	signal G1048: std_logic; attribute dont_touch of G1048: signal is true;
	signal G1049: std_logic; attribute dont_touch of G1049: signal is true;
	signal G1052: std_logic; attribute dont_touch of G1052: signal is true;
	signal G1053: std_logic; attribute dont_touch of G1053: signal is true;
	signal G1054: std_logic; attribute dont_touch of G1054: signal is true;
	signal G1055: std_logic; attribute dont_touch of G1055: signal is true;
	signal G1056: std_logic; attribute dont_touch of G1056: signal is true;
	signal G1059: std_logic; attribute dont_touch of G1059: signal is true;
	signal G1060: std_logic; attribute dont_touch of G1060: signal is true;
	signal G1063: std_logic; attribute dont_touch of G1063: signal is true;
	signal G1064: std_logic; attribute dont_touch of G1064: signal is true;
	signal G1070: std_logic; attribute dont_touch of G1070: signal is true;
	signal G1075: std_logic; attribute dont_touch of G1075: signal is true;
	signal G1076: std_logic; attribute dont_touch of G1076: signal is true;
	signal G1084: std_logic; attribute dont_touch of G1084: signal is true;
	signal G1088: std_logic; attribute dont_touch of G1088: signal is true;
	signal G1094: std_logic; attribute dont_touch of G1094: signal is true;
	signal G1101: std_logic; attribute dont_touch of G1101: signal is true;
	signal G1106: std_logic; attribute dont_touch of G1106: signal is true;
	signal G1107: std_logic; attribute dont_touch of G1107: signal is true;
	signal G1108: std_logic; attribute dont_touch of G1108: signal is true;
	signal G1109: std_logic; attribute dont_touch of G1109: signal is true;
	signal G1110: std_logic; attribute dont_touch of G1110: signal is true;
	signal G1111: std_logic; attribute dont_touch of G1111: signal is true;
	signal G1112: std_logic; attribute dont_touch of G1112: signal is true;
	signal G1113: std_logic; attribute dont_touch of G1113: signal is true;
	signal G1114: std_logic; attribute dont_touch of G1114: signal is true;
	signal G1115: std_logic; attribute dont_touch of G1115: signal is true;
	signal G1116: std_logic; attribute dont_touch of G1116: signal is true;
	signal G1117: std_logic; attribute dont_touch of G1117: signal is true;
	signal G1118: std_logic; attribute dont_touch of G1118: signal is true;
	signal G1119: std_logic; attribute dont_touch of G1119: signal is true;
	signal G1122: std_logic; attribute dont_touch of G1122: signal is true;
	signal G1123: std_logic; attribute dont_touch of G1123: signal is true;
	signal G1138: std_logic; attribute dont_touch of G1138: signal is true;
	signal G1142: std_logic; attribute dont_touch of G1142: signal is true;
	signal G1143: std_logic; attribute dont_touch of G1143: signal is true;
	signal G1156: std_logic; attribute dont_touch of G1156: signal is true;
	signal G1157: std_logic; attribute dont_touch of G1157: signal is true;
	signal G1160: std_logic; attribute dont_touch of G1160: signal is true;
	signal G1161: std_logic; attribute dont_touch of G1161: signal is true;
	signal G1173: std_logic; attribute dont_touch of G1173: signal is true;
	signal G1174: std_logic; attribute dont_touch of G1174: signal is true;
	signal G1175: std_logic; attribute dont_touch of G1175: signal is true;
	signal G1176: std_logic; attribute dont_touch of G1176: signal is true;
	signal G1177: std_logic; attribute dont_touch of G1177: signal is true;
	signal G1189: std_logic; attribute dont_touch of G1189: signal is true;
	signal G1190: std_logic; attribute dont_touch of G1190: signal is true;
	signal G1191: std_logic; attribute dont_touch of G1191: signal is true;
	signal G1192: std_logic; attribute dont_touch of G1192: signal is true;
	signal G1193: std_logic; attribute dont_touch of G1193: signal is true;
	signal G1203: std_logic; attribute dont_touch of G1203: signal is true;
	signal G1204: std_logic; attribute dont_touch of G1204: signal is true;
	signal G1205: std_logic; attribute dont_touch of G1205: signal is true;
	signal G1206: std_logic; attribute dont_touch of G1206: signal is true;
	signal G1209: std_logic; attribute dont_touch of G1209: signal is true;
	signal G1219: std_logic; attribute dont_touch of G1219: signal is true;
	signal G1220: std_logic; attribute dont_touch of G1220: signal is true;
	signal G1221: std_logic; attribute dont_touch of G1221: signal is true;
	signal G1222: std_logic; attribute dont_touch of G1222: signal is true;
	signal G1232: std_logic; attribute dont_touch of G1232: signal is true;
	signal G1233: std_logic; attribute dont_touch of G1233: signal is true;
	signal G1236: std_logic; attribute dont_touch of G1236: signal is true;
	signal G1246: std_logic; attribute dont_touch of G1246: signal is true;
	signal G1249: std_logic; attribute dont_touch of G1249: signal is true;
	signal G1250: std_logic; attribute dont_touch of G1250: signal is true;
	signal G1253: std_logic; attribute dont_touch of G1253: signal is true;
	signal G1254: std_logic; attribute dont_touch of G1254: signal is true;
	signal G1255: std_logic; attribute dont_touch of G1255: signal is true;
	signal G1256: std_logic; attribute dont_touch of G1256: signal is true;
	signal G1257: std_logic; attribute dont_touch of G1257: signal is true;
	signal G1263: std_logic; attribute dont_touch of G1263: signal is true;
	signal G1267: std_logic; attribute dont_touch of G1267: signal is true;
	signal G1270: std_logic; attribute dont_touch of G1270: signal is true;
	signal G1273: std_logic; attribute dont_touch of G1273: signal is true;
	signal G1274: std_logic; attribute dont_touch of G1274: signal is true;
	signal G1275: std_logic; attribute dont_touch of G1275: signal is true;
	signal G1276: std_logic; attribute dont_touch of G1276: signal is true;
	signal G1279: std_logic; attribute dont_touch of G1279: signal is true;
	signal G1282: std_logic; attribute dont_touch of G1282: signal is true;
	signal G1283: std_logic; attribute dont_touch of G1283: signal is true;
	signal G1284: std_logic; attribute dont_touch of G1284: signal is true;
	signal G1285: std_logic; attribute dont_touch of G1285: signal is true;
	signal G1286: std_logic; attribute dont_touch of G1286: signal is true;
	signal G1287: std_logic; attribute dont_touch of G1287: signal is true;
	signal G1288: std_logic; attribute dont_touch of G1288: signal is true;
	signal G1289: std_logic; attribute dont_touch of G1289: signal is true;
	signal G1291: std_logic; attribute dont_touch of G1291: signal is true;
	signal G1292: std_logic; attribute dont_touch of G1292: signal is true;
	signal G1294: std_logic; attribute dont_touch of G1294: signal is true;
	signal G1295: std_logic; attribute dont_touch of G1295: signal is true;
	signal G1305: std_logic; attribute dont_touch of G1305: signal is true;
	signal G1315: std_logic; attribute dont_touch of G1315: signal is true;
	signal G1316: std_logic; attribute dont_touch of G1316: signal is true;
	signal G1317: std_logic; attribute dont_touch of G1317: signal is true;
	signal G1318: std_logic; attribute dont_touch of G1318: signal is true;
	signal G1319: std_logic; attribute dont_touch of G1319: signal is true;
	signal G1320: std_logic; attribute dont_touch of G1320: signal is true;
	signal G1321: std_logic; attribute dont_touch of G1321: signal is true;
	signal G1322: std_logic; attribute dont_touch of G1322: signal is true;
	signal G1323: std_logic; attribute dont_touch of G1323: signal is true;
	signal G1324: std_logic; attribute dont_touch of G1324: signal is true;
	signal G1325: std_logic; attribute dont_touch of G1325: signal is true;
	signal G1326: std_logic; attribute dont_touch of G1326: signal is true;
	signal G1327: std_logic; attribute dont_touch of G1327: signal is true;
	signal G1328: std_logic; attribute dont_touch of G1328: signal is true;
	signal G1329: std_logic; attribute dont_touch of G1329: signal is true;
	signal G1330: std_logic; attribute dont_touch of G1330: signal is true;
	signal G1331: std_logic; attribute dont_touch of G1331: signal is true;
	signal G1332: std_logic; attribute dont_touch of G1332: signal is true;
	signal G1333: std_logic; attribute dont_touch of G1333: signal is true;
	signal G1334: std_logic; attribute dont_touch of G1334: signal is true;
	signal G1335: std_logic; attribute dont_touch of G1335: signal is true;
	signal G1336: std_logic; attribute dont_touch of G1336: signal is true;
	signal G1337: std_logic; attribute dont_touch of G1337: signal is true;
	signal G1338: std_logic; attribute dont_touch of G1338: signal is true;
	signal G1339: std_logic; attribute dont_touch of G1339: signal is true;
	signal G1340: std_logic; attribute dont_touch of G1340: signal is true;
	signal G1341: std_logic; attribute dont_touch of G1341: signal is true;
	signal G1344: std_logic; attribute dont_touch of G1344: signal is true;
	signal G1345: std_logic; attribute dont_touch of G1345: signal is true;
	signal G1348: std_logic; attribute dont_touch of G1348: signal is true;
	signal G1351: std_logic; attribute dont_touch of G1351: signal is true;
	signal G1352: std_logic; attribute dont_touch of G1352: signal is true;
	signal G1355: std_logic; attribute dont_touch of G1355: signal is true;
	signal G1358: std_logic; attribute dont_touch of G1358: signal is true;
	signal G1359: std_logic; attribute dont_touch of G1359: signal is true;
	signal G1363: std_logic; attribute dont_touch of G1363: signal is true;
	signal G1366: std_logic; attribute dont_touch of G1366: signal is true;
	signal G1369: std_logic; attribute dont_touch of G1369: signal is true;
	signal G1372: std_logic; attribute dont_touch of G1372: signal is true;
	signal G1375: std_logic; attribute dont_touch of G1375: signal is true;
	signal G1378: std_logic; attribute dont_touch of G1378: signal is true;
	signal G1381: std_logic; attribute dont_touch of G1381: signal is true;
	signal G1384: std_logic; attribute dont_touch of G1384: signal is true;
	signal G1387: std_logic; attribute dont_touch of G1387: signal is true;
	signal G1391: std_logic; attribute dont_touch of G1391: signal is true;
	signal G1394: std_logic; attribute dont_touch of G1394: signal is true;
	signal G1395: std_logic; attribute dont_touch of G1395: signal is true;
	signal G1398: std_logic; attribute dont_touch of G1398: signal is true;
	signal G1402: std_logic; attribute dont_touch of G1402: signal is true;
	signal G1407: std_logic; attribute dont_touch of G1407: signal is true;
	signal G1410: std_logic; attribute dont_touch of G1410: signal is true;
	signal G1411: std_logic; attribute dont_touch of G1411: signal is true;
	signal G1415: std_logic; attribute dont_touch of G1415: signal is true;
	signal G1416: std_logic; attribute dont_touch of G1416: signal is true;
	signal G1417: std_logic; attribute dont_touch of G1417: signal is true;
	signal G1418: std_logic; attribute dont_touch of G1418: signal is true;
	signal G1419: std_logic; attribute dont_touch of G1419: signal is true;
	signal G1422: std_logic; attribute dont_touch of G1422: signal is true;
	signal G1423: std_logic; attribute dont_touch of G1423: signal is true;
	signal G1426: std_logic; attribute dont_touch of G1426: signal is true;
	signal G1436: std_logic; attribute dont_touch of G1436: signal is true;
	signal G1439: std_logic; attribute dont_touch of G1439: signal is true;
	signal G1449: std_logic; attribute dont_touch of G1449: signal is true;
	signal G1450: std_logic; attribute dont_touch of G1450: signal is true;
	signal G1459: std_logic; attribute dont_touch of G1459: signal is true;
	signal G1460: std_logic; attribute dont_touch of G1460: signal is true;
	signal G1461: std_logic; attribute dont_touch of G1461: signal is true;
	signal G1470: std_logic; attribute dont_touch of G1470: signal is true;
	signal G1471: std_logic; attribute dont_touch of G1471: signal is true;
	signal G1472: std_logic; attribute dont_touch of G1472: signal is true;
	signal G1473: std_logic; attribute dont_touch of G1473: signal is true;
	signal G1474: std_logic; attribute dont_touch of G1474: signal is true;
	signal G1477: std_logic; attribute dont_touch of G1477: signal is true;
	signal G1480: std_logic; attribute dont_touch of G1480: signal is true;
	signal G1481: std_logic; attribute dont_touch of G1481: signal is true;
	signal G1484: std_logic; attribute dont_touch of G1484: signal is true;
	signal G1491: std_logic; attribute dont_touch of G1491: signal is true;
	signal G1498: std_logic; attribute dont_touch of G1498: signal is true;
	signal G1499: std_logic; attribute dont_touch of G1499: signal is true;
	signal G1502: std_logic; attribute dont_touch of G1502: signal is true;
	signal G1503: std_logic; attribute dont_touch of G1503: signal is true;
	signal G1504: std_logic; attribute dont_touch of G1504: signal is true;
	signal G1513: std_logic; attribute dont_touch of G1513: signal is true;
	signal G1514: std_logic; attribute dont_touch of G1514: signal is true;
	signal G1518: std_logic; attribute dont_touch of G1518: signal is true;
	signal G1519: std_logic; attribute dont_touch of G1519: signal is true;
	signal G1528: std_logic; attribute dont_touch of G1528: signal is true;
	signal G1529: std_logic; attribute dont_touch of G1529: signal is true;
	signal G1533: std_logic; attribute dont_touch of G1533: signal is true;
	signal G1534: std_logic; attribute dont_touch of G1534: signal is true;
	signal G1535: std_logic; attribute dont_touch of G1535: signal is true;
	signal G1539: std_logic; attribute dont_touch of G1539: signal is true;
	signal G1540: std_logic; attribute dont_touch of G1540: signal is true;
	signal G1541: std_logic; attribute dont_touch of G1541: signal is true;
	signal G1542: std_logic; attribute dont_touch of G1542: signal is true;
	signal G1543: std_logic; attribute dont_touch of G1543: signal is true;
	signal G1546: std_logic; attribute dont_touch of G1546: signal is true;
	signal G1549: std_logic; attribute dont_touch of G1549: signal is true;
	signal G1550: std_logic; attribute dont_touch of G1550: signal is true;
	signal G1551: std_logic; attribute dont_touch of G1551: signal is true;
	signal G1552: std_logic; attribute dont_touch of G1552: signal is true;
	signal G1555: std_logic; attribute dont_touch of G1555: signal is true;
	signal G1556: std_logic; attribute dont_touch of G1556: signal is true;
	signal G1557: std_logic; attribute dont_touch of G1557: signal is true;
	signal G1558: std_logic; attribute dont_touch of G1558: signal is true;
	signal G1559: std_logic; attribute dont_touch of G1559: signal is true;
	signal G1560: std_logic; attribute dont_touch of G1560: signal is true;
	signal G1563: std_logic; attribute dont_touch of G1563: signal is true;
	signal G1564: std_logic; attribute dont_touch of G1564: signal is true;
	signal G1567: std_logic; attribute dont_touch of G1567: signal is true;
	signal G1570: std_logic; attribute dont_touch of G1570: signal is true;
	signal G1573: std_logic; attribute dont_touch of G1573: signal is true;
	signal G1574: std_logic; attribute dont_touch of G1574: signal is true;
	signal G1575: std_logic; attribute dont_touch of G1575: signal is true;
	signal G1576: std_logic; attribute dont_touch of G1576: signal is true;
	signal G1577: std_logic; attribute dont_touch of G1577: signal is true;
	signal G1578: std_logic; attribute dont_touch of G1578: signal is true;
	signal G1581: std_logic; attribute dont_touch of G1581: signal is true;
	signal G1582: std_logic; attribute dont_touch of G1582: signal is true;
	signal G1583: std_logic; attribute dont_touch of G1583: signal is true;
	signal G1584: std_logic; attribute dont_touch of G1584: signal is true;
	signal G1585: std_logic; attribute dont_touch of G1585: signal is true;
	signal G1586: std_logic; attribute dont_touch of G1586: signal is true;
	signal G1587: std_logic; attribute dont_touch of G1587: signal is true;
	signal G1588: std_logic; attribute dont_touch of G1588: signal is true;
	signal G1589: std_logic; attribute dont_touch of G1589: signal is true;
	signal G1593: std_logic; attribute dont_touch of G1593: signal is true;
	signal G1594: std_logic; attribute dont_touch of G1594: signal is true;
	signal G1595: std_logic; attribute dont_touch of G1595: signal is true;
	signal G1603: std_logic; attribute dont_touch of G1603: signal is true;
	signal G1608: std_logic; attribute dont_touch of G1608: signal is true;
	signal G1609: std_logic; attribute dont_touch of G1609: signal is true;
	signal G1612: std_logic; attribute dont_touch of G1612: signal is true;
	signal G1620: std_logic; attribute dont_touch of G1620: signal is true;
	signal G1623: std_logic; attribute dont_touch of G1623: signal is true;
	signal G1624: std_logic; attribute dont_touch of G1624: signal is true;
	signal G1627: std_logic; attribute dont_touch of G1627: signal is true;
	signal G1628: std_logic; attribute dont_touch of G1628: signal is true;
	signal G1631: std_logic; attribute dont_touch of G1631: signal is true;
	signal G1632: std_logic; attribute dont_touch of G1632: signal is true;
	signal G1633: std_logic; attribute dont_touch of G1633: signal is true;
	signal G1636: std_logic; attribute dont_touch of G1636: signal is true;
	signal G1637: std_logic; attribute dont_touch of G1637: signal is true;
	signal G1638: std_logic; attribute dont_touch of G1638: signal is true;
	signal G1639: std_logic; attribute dont_touch of G1639: signal is true;
	signal G1640: std_logic; attribute dont_touch of G1640: signal is true;
	signal G1641: std_logic; attribute dont_touch of G1641: signal is true;
	signal G1642: std_logic; attribute dont_touch of G1642: signal is true;
	signal G1643: std_logic; attribute dont_touch of G1643: signal is true;
	signal G1644: std_logic; attribute dont_touch of G1644: signal is true;
	signal G1645: std_logic; attribute dont_touch of G1645: signal is true;
	signal G1646: std_logic; attribute dont_touch of G1646: signal is true;
	signal G1647: std_logic; attribute dont_touch of G1647: signal is true;
	signal G1648: std_logic; attribute dont_touch of G1648: signal is true;
	signal G1649: std_logic; attribute dont_touch of G1649: signal is true;
	signal G1650: std_logic; attribute dont_touch of G1650: signal is true;
	signal G1653: std_logic; attribute dont_touch of G1653: signal is true;
	signal G1654: std_logic; attribute dont_touch of G1654: signal is true;
	signal G1655: std_logic; attribute dont_touch of G1655: signal is true;
	signal G1656: std_logic; attribute dont_touch of G1656: signal is true;
	signal G1659: std_logic; attribute dont_touch of G1659: signal is true;
	signal G1660: std_logic; attribute dont_touch of G1660: signal is true;
	signal G1661: std_logic; attribute dont_touch of G1661: signal is true;
	signal G1664: std_logic; attribute dont_touch of G1664: signal is true;
	signal G1665: std_logic; attribute dont_touch of G1665: signal is true;
	signal G1666: std_logic; attribute dont_touch of G1666: signal is true;
	signal G1670: std_logic; attribute dont_touch of G1670: signal is true;
	signal G1671: std_logic; attribute dont_touch of G1671: signal is true;
	signal G1672: std_logic; attribute dont_touch of G1672: signal is true;
	signal G1673: std_logic; attribute dont_touch of G1673: signal is true;
	signal G1674: std_logic; attribute dont_touch of G1674: signal is true;
	signal G1675: std_logic; attribute dont_touch of G1675: signal is true;
	signal G1678: std_logic; attribute dont_touch of G1678: signal is true;
	signal G1679: std_logic; attribute dont_touch of G1679: signal is true;
	signal G1680: std_logic; attribute dont_touch of G1680: signal is true;
	signal G1681: std_logic; attribute dont_touch of G1681: signal is true;
	signal G1682: std_logic; attribute dont_touch of G1682: signal is true;
	signal G1683: std_logic; attribute dont_touch of G1683: signal is true;
	signal G1684: std_logic; attribute dont_touch of G1684: signal is true;
	signal G1685: std_logic; attribute dont_touch of G1685: signal is true;
	signal G1686: std_logic; attribute dont_touch of G1686: signal is true;
	signal G1687: std_logic; attribute dont_touch of G1687: signal is true;
	signal G1688: std_logic; attribute dont_touch of G1688: signal is true;
	signal G1689: std_logic; attribute dont_touch of G1689: signal is true;
	signal G1690: std_logic; attribute dont_touch of G1690: signal is true;
	signal G1691: std_logic; attribute dont_touch of G1691: signal is true;
	signal G1692: std_logic; attribute dont_touch of G1692: signal is true;
	signal G1695: std_logic; attribute dont_touch of G1695: signal is true;
	signal G1696: std_logic; attribute dont_touch of G1696: signal is true;
	signal G1699: std_logic; attribute dont_touch of G1699: signal is true;
	signal G1702: std_logic; attribute dont_touch of G1702: signal is true;
	signal G1703: std_logic; attribute dont_touch of G1703: signal is true;
	signal G1706: std_logic; attribute dont_touch of G1706: signal is true;
	signal G1710: std_logic; attribute dont_touch of G1710: signal is true;
	signal G1711: std_logic; attribute dont_touch of G1711: signal is true;
	signal G1714: std_logic; attribute dont_touch of G1714: signal is true;
	signal G1715: std_logic; attribute dont_touch of G1715: signal is true;
	signal G1716: std_logic; attribute dont_touch of G1716: signal is true;
	signal G1720: std_logic; attribute dont_touch of G1720: signal is true;
	signal G1721: std_logic; attribute dont_touch of G1721: signal is true;
	signal G1724: std_logic; attribute dont_touch of G1724: signal is true;
	signal G1725: std_logic; attribute dont_touch of G1725: signal is true;
	signal G1726: std_logic; attribute dont_touch of G1726: signal is true;
	signal G1729: std_logic; attribute dont_touch of G1729: signal is true;
	signal G1730: std_logic; attribute dont_touch of G1730: signal is true;
	signal G1731: std_logic; attribute dont_touch of G1731: signal is true;
	signal G1732: std_logic; attribute dont_touch of G1732: signal is true;
	signal G1733: std_logic; attribute dont_touch of G1733: signal is true;
	signal G1734: std_logic; attribute dont_touch of G1734: signal is true;
	signal G1735: std_logic; attribute dont_touch of G1735: signal is true;
	signal G1738: std_logic; attribute dont_touch of G1738: signal is true;
	signal G1739: std_logic; attribute dont_touch of G1739: signal is true;
	signal G1740: std_logic; attribute dont_touch of G1740: signal is true;
	signal G1741: std_logic; attribute dont_touch of G1741: signal is true;
	signal G1742: std_logic; attribute dont_touch of G1742: signal is true;
	signal G1743: std_logic; attribute dont_touch of G1743: signal is true;
	signal G1747: std_logic; attribute dont_touch of G1747: signal is true;
	signal G1748: std_logic; attribute dont_touch of G1748: signal is true;
	signal G1749: std_logic; attribute dont_touch of G1749: signal is true;
	signal G1754: std_logic; attribute dont_touch of G1754: signal is true;
	signal G1755: std_logic; attribute dont_touch of G1755: signal is true;
	signal G1756: std_logic; attribute dont_touch of G1756: signal is true;
	signal G1759: std_logic; attribute dont_touch of G1759: signal is true;
	signal G1760: std_logic; attribute dont_touch of G1760: signal is true;
	signal G1761: std_logic; attribute dont_touch of G1761: signal is true;
	signal G1762: std_logic; attribute dont_touch of G1762: signal is true;
	signal G1763: std_logic; attribute dont_touch of G1763: signal is true;
	signal G1764: std_logic; attribute dont_touch of G1764: signal is true;
	signal G1769: std_logic; attribute dont_touch of G1769: signal is true;
	signal G1770: std_logic; attribute dont_touch of G1770: signal is true;
	signal G1771: std_logic; attribute dont_touch of G1771: signal is true;
	signal G1772: std_logic; attribute dont_touch of G1772: signal is true;
	signal G1773: std_logic; attribute dont_touch of G1773: signal is true;
	signal G1774: std_logic; attribute dont_touch of G1774: signal is true;
	signal G1775: std_logic; attribute dont_touch of G1775: signal is true;
	signal G1776: std_logic; attribute dont_touch of G1776: signal is true;
	signal G1777: std_logic; attribute dont_touch of G1777: signal is true;
	signal G1781: std_logic; attribute dont_touch of G1781: signal is true;
	signal G1782: std_logic; attribute dont_touch of G1782: signal is true;
	signal G1783: std_logic; attribute dont_touch of G1783: signal is true;
	signal G1784: std_logic; attribute dont_touch of G1784: signal is true;
	signal G1787: std_logic; attribute dont_touch of G1787: signal is true;
	signal G1788: std_logic; attribute dont_touch of G1788: signal is true;
	signal G1789: std_logic; attribute dont_touch of G1789: signal is true;
	signal G1790: std_logic; attribute dont_touch of G1790: signal is true;
	signal G1791: std_logic; attribute dont_touch of G1791: signal is true;
	signal G1792: std_logic; attribute dont_touch of G1792: signal is true;
	signal G1793: std_logic; attribute dont_touch of G1793: signal is true;
	signal G1797: std_logic; attribute dont_touch of G1797: signal is true;
	signal G1802: std_logic; attribute dont_touch of G1802: signal is true;
	signal G1805: std_logic; attribute dont_touch of G1805: signal is true;
	signal G1806: std_logic; attribute dont_touch of G1806: signal is true;
	signal G1807: std_logic; attribute dont_touch of G1807: signal is true;
	signal G1808: std_logic; attribute dont_touch of G1808: signal is true;
	signal G1811: std_logic; attribute dont_touch of G1811: signal is true;
	signal G1812: std_logic; attribute dont_touch of G1812: signal is true;
	signal G1813: std_logic; attribute dont_touch of G1813: signal is true;
	signal G1814: std_logic; attribute dont_touch of G1814: signal is true;
	signal G1815: std_logic; attribute dont_touch of G1815: signal is true;
	signal G1819: std_logic; attribute dont_touch of G1819: signal is true;
	signal G1820: std_logic; attribute dont_touch of G1820: signal is true;
	signal G1821: std_logic; attribute dont_touch of G1821: signal is true;
	signal G1822: std_logic; attribute dont_touch of G1822: signal is true;
	signal G1823: std_logic; attribute dont_touch of G1823: signal is true;
	signal G1824: std_logic; attribute dont_touch of G1824: signal is true;
	signal G1825: std_logic; attribute dont_touch of G1825: signal is true;
	signal G1826: std_logic; attribute dont_touch of G1826: signal is true;
	signal G1829: std_logic; attribute dont_touch of G1829: signal is true;
	signal G1830: std_logic; attribute dont_touch of G1830: signal is true;
	signal G1831: std_logic; attribute dont_touch of G1831: signal is true;
	signal G1832: std_logic; attribute dont_touch of G1832: signal is true;
	signal G1833: std_logic; attribute dont_touch of G1833: signal is true;
	signal G1834: std_logic; attribute dont_touch of G1834: signal is true;
	signal G1835: std_logic; attribute dont_touch of G1835: signal is true;
	signal G1836: std_logic; attribute dont_touch of G1836: signal is true;
	signal G1837: std_logic; attribute dont_touch of G1837: signal is true;
	signal G1838: std_logic; attribute dont_touch of G1838: signal is true;
	signal G1841: std_logic; attribute dont_touch of G1841: signal is true;
	signal G1842: std_logic; attribute dont_touch of G1842: signal is true;
	signal G1845: std_logic; attribute dont_touch of G1845: signal is true;
	signal G1846: std_logic; attribute dont_touch of G1846: signal is true;
	signal G1847: std_logic; attribute dont_touch of G1847: signal is true;
	signal G1848: std_logic; attribute dont_touch of G1848: signal is true;
	signal G1849: std_logic; attribute dont_touch of G1849: signal is true;
	signal G1852: std_logic; attribute dont_touch of G1852: signal is true;
	signal G1853: std_logic; attribute dont_touch of G1853: signal is true;
	signal G1854: std_logic; attribute dont_touch of G1854: signal is true;
	signal G1857: std_logic; attribute dont_touch of G1857: signal is true;
	signal G1858: std_logic; attribute dont_touch of G1858: signal is true;
	signal G1861: std_logic; attribute dont_touch of G1861: signal is true;
	signal G1875: std_logic; attribute dont_touch of G1875: signal is true;
	signal G1878: std_logic; attribute dont_touch of G1878: signal is true;
	signal G1879: std_logic; attribute dont_touch of G1879: signal is true;
	signal G1880: std_logic; attribute dont_touch of G1880: signal is true;
	signal G1883: std_logic; attribute dont_touch of G1883: signal is true;
	signal G1884: std_logic; attribute dont_touch of G1884: signal is true;
	signal G1887: std_logic; attribute dont_touch of G1887: signal is true;
	signal G1890: std_logic; attribute dont_touch of G1890: signal is true;
	signal G1891: std_logic; attribute dont_touch of G1891: signal is true;
	signal G1894: std_logic; attribute dont_touch of G1894: signal is true;
	signal G1897: std_logic; attribute dont_touch of G1897: signal is true;
	signal G1898: std_logic; attribute dont_touch of G1898: signal is true;
	signal G1899: std_logic; attribute dont_touch of G1899: signal is true;
	signal G1902: std_logic; attribute dont_touch of G1902: signal is true;
	signal G1905: std_logic; attribute dont_touch of G1905: signal is true;
	signal G1908: std_logic; attribute dont_touch of G1908: signal is true;
	signal G1911: std_logic; attribute dont_touch of G1911: signal is true;
	signal G1914: std_logic; attribute dont_touch of G1914: signal is true;
	signal G1917: std_logic; attribute dont_touch of G1917: signal is true;
	signal G1918: std_logic; attribute dont_touch of G1918: signal is true;
	signal G1919: std_logic; attribute dont_touch of G1919: signal is true;
	signal G1922: std_logic; attribute dont_touch of G1922: signal is true;
	signal G1925: std_logic; attribute dont_touch of G1925: signal is true;
	signal G1928: std_logic; attribute dont_touch of G1928: signal is true;
	signal G1931: std_logic; attribute dont_touch of G1931: signal is true;
	signal G1934: std_logic; attribute dont_touch of G1934: signal is true;
	signal G1935: std_logic; attribute dont_touch of G1935: signal is true;
	signal G1936: std_logic; attribute dont_touch of G1936: signal is true;
	signal G1937: std_logic; attribute dont_touch of G1937: signal is true;
	signal G1940: std_logic; attribute dont_touch of G1940: signal is true;
	signal G1943: std_logic; attribute dont_touch of G1943: signal is true;
	signal G1946: std_logic; attribute dont_touch of G1946: signal is true;
	signal G1947: std_logic; attribute dont_touch of G1947: signal is true;
	signal G1950: std_logic; attribute dont_touch of G1950: signal is true;
	signal G1953: std_logic; attribute dont_touch of G1953: signal is true;
	signal G1954: std_logic; attribute dont_touch of G1954: signal is true;
	signal G1957: std_logic; attribute dont_touch of G1957: signal is true;
	signal G1960: std_logic; attribute dont_touch of G1960: signal is true;
	signal G1963: std_logic; attribute dont_touch of G1963: signal is true;
	signal G1966: std_logic; attribute dont_touch of G1966: signal is true;
	signal G1969: std_logic; attribute dont_touch of G1969: signal is true;
	signal G1972: std_logic; attribute dont_touch of G1972: signal is true;
	signal G1975: std_logic; attribute dont_touch of G1975: signal is true;
	signal G1978: std_logic; attribute dont_touch of G1978: signal is true;
	signal G1979: std_logic; attribute dont_touch of G1979: signal is true;
	signal G1982: std_logic; attribute dont_touch of G1982: signal is true;
	signal G1985: std_logic; attribute dont_touch of G1985: signal is true;
	signal G1988: std_logic; attribute dont_touch of G1988: signal is true;
	signal G1991: std_logic; attribute dont_touch of G1991: signal is true;
	signal G1994: std_logic; attribute dont_touch of G1994: signal is true;
	signal G1997: std_logic; attribute dont_touch of G1997: signal is true;
	signal G1998: std_logic; attribute dont_touch of G1998: signal is true;
	signal G2001: std_logic; attribute dont_touch of G2001: signal is true;
	signal G2004: std_logic; attribute dont_touch of G2004: signal is true;
	signal G2007: std_logic; attribute dont_touch of G2007: signal is true;
	signal G2008: std_logic; attribute dont_touch of G2008: signal is true;
	signal G2009: std_logic; attribute dont_touch of G2009: signal is true;
	signal G2010: std_logic; attribute dont_touch of G2010: signal is true;
	signal G2015: std_logic; attribute dont_touch of G2015: signal is true;
	signal G2018: std_logic; attribute dont_touch of G2018: signal is true;
	signal G2021: std_logic; attribute dont_touch of G2021: signal is true;
	signal G2024: std_logic; attribute dont_touch of G2024: signal is true;
	signal G2025: std_logic; attribute dont_touch of G2025: signal is true;
	signal G2026: std_logic; attribute dont_touch of G2026: signal is true;
	signal G2029: std_logic; attribute dont_touch of G2029: signal is true;
	signal G2030: std_logic; attribute dont_touch of G2030: signal is true;
	signal G2031: std_logic; attribute dont_touch of G2031: signal is true;
	signal G2032: std_logic; attribute dont_touch of G2032: signal is true;
	signal G2035: std_logic; attribute dont_touch of G2035: signal is true;
	signal G2036: std_logic; attribute dont_touch of G2036: signal is true;
	signal G2039: std_logic; attribute dont_touch of G2039: signal is true;
	signal G2040: std_logic; attribute dont_touch of G2040: signal is true;
	signal G2041: std_logic; attribute dont_touch of G2041: signal is true;
	signal G2042: std_logic; attribute dont_touch of G2042: signal is true;
	signal G2043: std_logic; attribute dont_touch of G2043: signal is true;
	signal G2044: std_logic; attribute dont_touch of G2044: signal is true;
	signal G2053: std_logic; attribute dont_touch of G2053: signal is true;
	signal G2056: std_logic; attribute dont_touch of G2056: signal is true;
	signal G2059: std_logic; attribute dont_touch of G2059: signal is true;
	signal G2060: std_logic; attribute dont_touch of G2060: signal is true;
	signal G2061: std_logic; attribute dont_touch of G2061: signal is true;
	signal G2062: std_logic; attribute dont_touch of G2062: signal is true;
	signal G2066: std_logic; attribute dont_touch of G2066: signal is true;
	signal G2067: std_logic; attribute dont_touch of G2067: signal is true;
	signal G2068: std_logic; attribute dont_touch of G2068: signal is true;
	signal G2073: std_logic; attribute dont_touch of G2073: signal is true;
	signal G2078: std_logic; attribute dont_touch of G2078: signal is true;
	signal G2079: std_logic; attribute dont_touch of G2079: signal is true;
	signal G2080: std_logic; attribute dont_touch of G2080: signal is true;
	signal G2081: std_logic; attribute dont_touch of G2081: signal is true;
	signal G2084: std_logic; attribute dont_touch of G2084: signal is true;
	signal G2085: std_logic; attribute dont_touch of G2085: signal is true;
	signal G2086: std_logic; attribute dont_touch of G2086: signal is true;
	signal G2087: std_logic; attribute dont_touch of G2087: signal is true;
	signal G2088: std_logic; attribute dont_touch of G2088: signal is true;
	signal G2089: std_logic; attribute dont_touch of G2089: signal is true;
	signal G2090: std_logic; attribute dont_touch of G2090: signal is true;
	signal G2091: std_logic; attribute dont_touch of G2091: signal is true;
	signal G2092: std_logic; attribute dont_touch of G2092: signal is true;
	signal G2095: std_logic; attribute dont_touch of G2095: signal is true;
	signal G2096: std_logic; attribute dont_touch of G2096: signal is true;
	signal G2097: std_logic; attribute dont_touch of G2097: signal is true;
	signal G2098: std_logic; attribute dont_touch of G2098: signal is true;
	signal G2099: std_logic; attribute dont_touch of G2099: signal is true;
	signal G2100: std_logic; attribute dont_touch of G2100: signal is true;
	signal G2101: std_logic; attribute dont_touch of G2101: signal is true;
	signal G2102: std_logic; attribute dont_touch of G2102: signal is true;
	signal G2103: std_logic; attribute dont_touch of G2103: signal is true;
	signal G2104: std_logic; attribute dont_touch of G2104: signal is true;
	signal G2105: std_logic; attribute dont_touch of G2105: signal is true;
	signal G2106: std_logic; attribute dont_touch of G2106: signal is true;
	signal G2107: std_logic; attribute dont_touch of G2107: signal is true;
	signal G2108: std_logic; attribute dont_touch of G2108: signal is true;
	signal G2109: std_logic; attribute dont_touch of G2109: signal is true;
	signal G2110: std_logic; attribute dont_touch of G2110: signal is true;
	signal G2111: std_logic; attribute dont_touch of G2111: signal is true;
	signal G2112: std_logic; attribute dont_touch of G2112: signal is true;
	signal G2113: std_logic; attribute dont_touch of G2113: signal is true;
	signal G2117: std_logic; attribute dont_touch of G2117: signal is true;
	signal G2118: std_logic; attribute dont_touch of G2118: signal is true;
	signal G2119: std_logic; attribute dont_touch of G2119: signal is true;
	signal G2120: std_logic; attribute dont_touch of G2120: signal is true;
	signal G2121: std_logic; attribute dont_touch of G2121: signal is true;
	signal G2125: std_logic; attribute dont_touch of G2125: signal is true;
	signal G2134: std_logic; attribute dont_touch of G2134: signal is true;
	signal G2135: std_logic; attribute dont_touch of G2135: signal is true;
	signal G2136: std_logic; attribute dont_touch of G2136: signal is true;
	signal G2137: std_logic; attribute dont_touch of G2137: signal is true;
	signal G2138: std_logic; attribute dont_touch of G2138: signal is true;
	signal G2142: std_logic; attribute dont_touch of G2142: signal is true;
	signal G2145: std_logic; attribute dont_touch of G2145: signal is true;
	signal G2154: std_logic; attribute dont_touch of G2154: signal is true;
	signal G2155: std_logic; attribute dont_touch of G2155: signal is true;
	signal G2156: std_logic; attribute dont_touch of G2156: signal is true;
	signal G2157: std_logic; attribute dont_touch of G2157: signal is true;
	signal G2158: std_logic; attribute dont_touch of G2158: signal is true;
	signal G2159: std_logic; attribute dont_touch of G2159: signal is true;
	signal G2160: std_logic; attribute dont_touch of G2160: signal is true;
	signal G2163: std_logic; attribute dont_touch of G2163: signal is true;
	signal G2164: std_logic; attribute dont_touch of G2164: signal is true;
	signal G2165: std_logic; attribute dont_touch of G2165: signal is true;
	signal G2166: std_logic; attribute dont_touch of G2166: signal is true;
	signal G2169: std_logic; attribute dont_touch of G2169: signal is true;
	signal G2170: std_logic; attribute dont_touch of G2170: signal is true;
	signal G2171: std_logic; attribute dont_touch of G2171: signal is true;
	signal G2172: std_logic; attribute dont_touch of G2172: signal is true;
	signal G2173: std_logic; attribute dont_touch of G2173: signal is true;
	signal G2174: std_logic; attribute dont_touch of G2174: signal is true;
	signal G2175: std_logic; attribute dont_touch of G2175: signal is true;
	signal G2176: std_logic; attribute dont_touch of G2176: signal is true;
	signal G2177: std_logic; attribute dont_touch of G2177: signal is true;
	signal G2178: std_logic; attribute dont_touch of G2178: signal is true;
	signal G2179: std_logic; attribute dont_touch of G2179: signal is true;
	signal G2194: std_logic; attribute dont_touch of G2194: signal is true;
	signal G2195: std_logic; attribute dont_touch of G2195: signal is true;
	signal G2196: std_logic; attribute dont_touch of G2196: signal is true;
	signal G2197: std_logic; attribute dont_touch of G2197: signal is true;
	signal G2212: std_logic; attribute dont_touch of G2212: signal is true;
	signal G2213: std_logic; attribute dont_touch of G2213: signal is true;
	signal G2214: std_logic; attribute dont_touch of G2214: signal is true;
	signal G2215: std_logic; attribute dont_touch of G2215: signal is true;
	signal G2230: std_logic; attribute dont_touch of G2230: signal is true;
	signal G2231: std_logic; attribute dont_touch of G2231: signal is true;
	signal G2232: std_logic; attribute dont_touch of G2232: signal is true;
	signal G2233: std_logic; attribute dont_touch of G2233: signal is true;
	signal G2234: std_logic; attribute dont_touch of G2234: signal is true;
	signal G2241: std_logic; attribute dont_touch of G2241: signal is true;
	signal G2242: std_logic; attribute dont_touch of G2242: signal is true;
	signal G2243: std_logic; attribute dont_touch of G2243: signal is true;
	signal G2244: std_logic; attribute dont_touch of G2244: signal is true;
	signal G2245: std_logic; attribute dont_touch of G2245: signal is true;
	signal G2252: std_logic; attribute dont_touch of G2252: signal is true;
	signal G2253: std_logic; attribute dont_touch of G2253: signal is true;
	signal G2254: std_logic; attribute dont_touch of G2254: signal is true;
	signal G2255: std_logic; attribute dont_touch of G2255: signal is true;
	signal G2256: std_logic; attribute dont_touch of G2256: signal is true;
	signal G2263: std_logic; attribute dont_touch of G2263: signal is true;
	signal G2264: std_logic; attribute dont_touch of G2264: signal is true;
	signal G2265: std_logic; attribute dont_touch of G2265: signal is true;
	signal G2266: std_logic; attribute dont_touch of G2266: signal is true;
	signal G2267: std_logic; attribute dont_touch of G2267: signal is true;
	signal G2268: std_logic; attribute dont_touch of G2268: signal is true;
	signal G2275: std_logic; attribute dont_touch of G2275: signal is true;
	signal G2276: std_logic; attribute dont_touch of G2276: signal is true;
	signal G2283: std_logic; attribute dont_touch of G2283: signal is true;
	signal G2284: std_logic; attribute dont_touch of G2284: signal is true;
	signal G2291: std_logic; attribute dont_touch of G2291: signal is true;
	signal G2292: std_logic; attribute dont_touch of G2292: signal is true;
	signal G2293: std_logic; attribute dont_touch of G2293: signal is true;
	signal G2294: std_logic; attribute dont_touch of G2294: signal is true;
	signal G2295: std_logic; attribute dont_touch of G2295: signal is true;
	signal G2296: std_logic; attribute dont_touch of G2296: signal is true;
	signal G2306: std_logic; attribute dont_touch of G2306: signal is true;
	signal G2307: std_logic; attribute dont_touch of G2307: signal is true;
	signal G2308: std_logic; attribute dont_touch of G2308: signal is true;
	signal G2311: std_logic; attribute dont_touch of G2311: signal is true;
	signal G2312: std_logic; attribute dont_touch of G2312: signal is true;
	signal G2315: std_logic; attribute dont_touch of G2315: signal is true;
	signal G2316: std_logic; attribute dont_touch of G2316: signal is true;
	signal G2317: std_logic; attribute dont_touch of G2317: signal is true;
	signal G2320: std_logic; attribute dont_touch of G2320: signal is true;
	signal G2323: std_logic; attribute dont_touch of G2323: signal is true;
	signal G2324: std_logic; attribute dont_touch of G2324: signal is true;
	signal G2327: std_logic; attribute dont_touch of G2327: signal is true;
	signal G2330: std_logic; attribute dont_touch of G2330: signal is true;
	signal G2333: std_logic; attribute dont_touch of G2333: signal is true;
	signal G2336: std_logic; attribute dont_touch of G2336: signal is true;
	signal G2339: std_logic; attribute dont_touch of G2339: signal is true;
	signal G2340: std_logic; attribute dont_touch of G2340: signal is true;
	signal G2343: std_logic; attribute dont_touch of G2343: signal is true;
	signal G2346: std_logic; attribute dont_touch of G2346: signal is true;
	signal G2347: std_logic; attribute dont_touch of G2347: signal is true;
	signal G2350: std_logic; attribute dont_touch of G2350: signal is true;
	signal G2353: std_logic; attribute dont_touch of G2353: signal is true;
	signal G2356: std_logic; attribute dont_touch of G2356: signal is true;
	signal G2357: std_logic; attribute dont_touch of G2357: signal is true;
	signal G2360: std_logic; attribute dont_touch of G2360: signal is true;
	signal G2361: std_logic; attribute dont_touch of G2361: signal is true;
	signal G2364: std_logic; attribute dont_touch of G2364: signal is true;
	signal G2367: std_logic; attribute dont_touch of G2367: signal is true;
	signal G2370: std_logic; attribute dont_touch of G2370: signal is true;
	signal G2378: std_logic; attribute dont_touch of G2378: signal is true;
	signal G2381: std_logic; attribute dont_touch of G2381: signal is true;
	signal G2390: std_logic; attribute dont_touch of G2390: signal is true;
	signal G2391: std_logic; attribute dont_touch of G2391: signal is true;
	signal G2394: std_logic; attribute dont_touch of G2394: signal is true;
	signal G2397: std_logic; attribute dont_touch of G2397: signal is true;
	signal G2405: std_logic; attribute dont_touch of G2405: signal is true;
	signal G2408: std_logic; attribute dont_touch of G2408: signal is true;
	signal G2409: std_logic; attribute dont_touch of G2409: signal is true;
	signal G2410: std_logic; attribute dont_touch of G2410: signal is true;
	signal G2413: std_logic; attribute dont_touch of G2413: signal is true;
	signal G2416: std_logic; attribute dont_touch of G2416: signal is true;
	signal G2419: std_logic; attribute dont_touch of G2419: signal is true;
	signal G2422: std_logic; attribute dont_touch of G2422: signal is true;
	signal G2430: std_logic; attribute dont_touch of G2430: signal is true;
	signal G2433: std_logic; attribute dont_touch of G2433: signal is true;
	signal G2434: std_logic; attribute dont_touch of G2434: signal is true;
	signal G2435: std_logic; attribute dont_touch of G2435: signal is true;
	signal G2436: std_logic; attribute dont_touch of G2436: signal is true;
	signal G2437: std_logic; attribute dont_touch of G2437: signal is true;
	signal G2440: std_logic; attribute dont_touch of G2440: signal is true;
	signal G2443: std_logic; attribute dont_touch of G2443: signal is true;
	signal G2446: std_logic; attribute dont_touch of G2446: signal is true;
	signal G2449: std_logic; attribute dont_touch of G2449: signal is true;
	signal G2457: std_logic; attribute dont_touch of G2457: signal is true;
	signal G2460: std_logic; attribute dont_touch of G2460: signal is true;
	signal G2461: std_logic; attribute dont_touch of G2461: signal is true;
	signal G2464: std_logic; attribute dont_touch of G2464: signal is true;
	signal G2467: std_logic; attribute dont_touch of G2467: signal is true;
	signal G2470: std_logic; attribute dont_touch of G2470: signal is true;
	signal G2473: std_logic; attribute dont_touch of G2473: signal is true;
	signal G2481: std_logic; attribute dont_touch of G2481: signal is true;
	signal G2484: std_logic; attribute dont_touch of G2484: signal is true;
	signal G2485: std_logic; attribute dont_touch of G2485: signal is true;
	signal G2488: std_logic; attribute dont_touch of G2488: signal is true;
	signal G2491: std_logic; attribute dont_touch of G2491: signal is true;
	signal G2494: std_logic; attribute dont_touch of G2494: signal is true;
	signal G2497: std_logic; attribute dont_touch of G2497: signal is true;
	signal G2505: std_logic; attribute dont_touch of G2505: signal is true;
	signal G2506: std_logic; attribute dont_touch of G2506: signal is true;
	signal G2509: std_logic; attribute dont_touch of G2509: signal is true;
	signal G2512: std_logic; attribute dont_touch of G2512: signal is true;
	signal G2515: std_logic; attribute dont_touch of G2515: signal is true;
	signal G2518: std_logic; attribute dont_touch of G2518: signal is true;
	signal G2524: std_logic; attribute dont_touch of G2524: signal is true;
	signal G2525: std_logic; attribute dont_touch of G2525: signal is true;
	signal G2535: std_logic; attribute dont_touch of G2535: signal is true;
	signal G2538: std_logic; attribute dont_touch of G2538: signal is true;
	signal G2541: std_logic; attribute dont_touch of G2541: signal is true;
	signal G2544: std_logic; attribute dont_touch of G2544: signal is true;
	signal G2550: std_logic; attribute dont_touch of G2550: signal is true;
	signal G2551: std_logic; attribute dont_touch of G2551: signal is true;
	signal G2554: std_logic; attribute dont_touch of G2554: signal is true;
	signal G2555: std_logic; attribute dont_touch of G2555: signal is true;
	signal G2565: std_logic; attribute dont_touch of G2565: signal is true;
	signal G2568: std_logic; attribute dont_touch of G2568: signal is true;
	signal G2574: std_logic; attribute dont_touch of G2574: signal is true;
	signal G2575: std_logic; attribute dont_touch of G2575: signal is true;
	signal G2576: std_logic; attribute dont_touch of G2576: signal is true;
	signal G2577: std_logic; attribute dont_touch of G2577: signal is true;
	signal G2580: std_logic; attribute dont_touch of G2580: signal is true;
	signal G2581: std_logic; attribute dont_touch of G2581: signal is true;
	signal G2582: std_logic; attribute dont_touch of G2582: signal is true;
	signal G2583: std_logic; attribute dont_touch of G2583: signal is true;
	signal G2585: std_logic; attribute dont_touch of G2585: signal is true;
	signal G2586: std_logic; attribute dont_touch of G2586: signal is true;
	signal G2587: std_logic; attribute dont_touch of G2587: signal is true;
	signal G2588: std_logic; attribute dont_touch of G2588: signal is true;
	signal G2591: std_logic; attribute dont_touch of G2591: signal is true;
	signal G2594: std_logic; attribute dont_touch of G2594: signal is true;
	signal G2598: std_logic; attribute dont_touch of G2598: signal is true;
	signal G2599: std_logic; attribute dont_touch of G2599: signal is true;
	signal G2602: std_logic; attribute dont_touch of G2602: signal is true;
	signal G2603: std_logic; attribute dont_touch of G2603: signal is true;
	signal G2604: std_logic; attribute dont_touch of G2604: signal is true;
	signal G2607: std_logic; attribute dont_touch of G2607: signal is true;
	signal G2608: std_logic; attribute dont_touch of G2608: signal is true;
	signal G2609: std_logic; attribute dont_touch of G2609: signal is true;
	signal G2612: std_logic; attribute dont_touch of G2612: signal is true;
	signal G2615: std_logic; attribute dont_touch of G2615: signal is true;
	signal G2618: std_logic; attribute dont_touch of G2618: signal is true;
	signal G2619: std_logic; attribute dont_touch of G2619: signal is true;
	signal G2622: std_logic; attribute dont_touch of G2622: signal is true;
	signal G2625: std_logic; attribute dont_touch of G2625: signal is true;
	signal G2628: std_logic; attribute dont_touch of G2628: signal is true;
	signal G2631: std_logic; attribute dont_touch of G2631: signal is true;
	signal G2634: std_logic; attribute dont_touch of G2634: signal is true;
	signal G2637: std_logic; attribute dont_touch of G2637: signal is true;
	signal G2640: std_logic; attribute dont_touch of G2640: signal is true;
	signal G2643: std_logic; attribute dont_touch of G2643: signal is true;
	signal G2644: std_logic; attribute dont_touch of G2644: signal is true;
	signal G2647: std_logic; attribute dont_touch of G2647: signal is true;
	signal G2650: std_logic; attribute dont_touch of G2650: signal is true;
	signal G2653: std_logic; attribute dont_touch of G2653: signal is true;
	signal G2656: std_logic; attribute dont_touch of G2656: signal is true;
	signal G2659: std_logic; attribute dont_touch of G2659: signal is true;
	signal G2660: std_logic; attribute dont_touch of G2660: signal is true;
	signal G2663: std_logic; attribute dont_touch of G2663: signal is true;
	signal G2664: std_logic; attribute dont_touch of G2664: signal is true;
	signal G2667: std_logic; attribute dont_touch of G2667: signal is true;
	signal G2670: std_logic; attribute dont_touch of G2670: signal is true;
	signal G2671: std_logic; attribute dont_touch of G2671: signal is true;
	signal G2672: std_logic; attribute dont_touch of G2672: signal is true;
	signal G2675: std_logic; attribute dont_touch of G2675: signal is true;
	signal G2678: std_logic; attribute dont_touch of G2678: signal is true;
	signal G2679: std_logic; attribute dont_touch of G2679: signal is true;
	signal G2682: std_logic; attribute dont_touch of G2682: signal is true;
	signal G2685: std_logic; attribute dont_touch of G2685: signal is true;
	signal G2686: std_logic; attribute dont_touch of G2686: signal is true;
	signal G2687: std_logic; attribute dont_touch of G2687: signal is true;
	signal G2688: std_logic; attribute dont_touch of G2688: signal is true;
	signal G2691: std_logic; attribute dont_touch of G2691: signal is true;
	signal G2692: std_logic; attribute dont_touch of G2692: signal is true;
	signal G2695: std_logic; attribute dont_touch of G2695: signal is true;
	signal G2698: std_logic; attribute dont_touch of G2698: signal is true;
	signal G2699: std_logic; attribute dont_touch of G2699: signal is true;
	signal G2700: std_logic; attribute dont_touch of G2700: signal is true;
	signal G2701: std_logic; attribute dont_touch of G2701: signal is true;
	signal G2705: std_logic; attribute dont_touch of G2705: signal is true;
	signal G2706: std_logic; attribute dont_touch of G2706: signal is true;
	signal G2709: std_logic; attribute dont_touch of G2709: signal is true;
	signal G2712: std_logic; attribute dont_touch of G2712: signal is true;
	signal G2713: std_logic; attribute dont_touch of G2713: signal is true;
	signal G2716: std_logic; attribute dont_touch of G2716: signal is true;
	signal G2719: std_logic; attribute dont_touch of G2719: signal is true;
	signal G2720: std_logic; attribute dont_touch of G2720: signal is true;
	signal G2721: std_logic; attribute dont_touch of G2721: signal is true;
	signal G2722: std_logic; attribute dont_touch of G2722: signal is true;
	signal G2726: std_logic; attribute dont_touch of G2726: signal is true;
	signal G2727: std_logic; attribute dont_touch of G2727: signal is true;
	signal G2728: std_logic; attribute dont_touch of G2728: signal is true;
	signal G2731: std_logic; attribute dont_touch of G2731: signal is true;
	signal G2732: std_logic; attribute dont_touch of G2732: signal is true;
	signal G2733: std_logic; attribute dont_touch of G2733: signal is true;
	signal G2734: std_logic; attribute dont_touch of G2734: signal is true;
	signal G2738: std_logic; attribute dont_touch of G2738: signal is true;
	signal G2739: std_logic; attribute dont_touch of G2739: signal is true;
	signal G2740: std_logic; attribute dont_touch of G2740: signal is true;
	signal G2743: std_logic; attribute dont_touch of G2743: signal is true;
	signal G2744: std_logic; attribute dont_touch of G2744: signal is true;
	signal G2745: std_logic; attribute dont_touch of G2745: signal is true;
	signal G2746: std_logic; attribute dont_touch of G2746: signal is true;
	signal G2747: std_logic; attribute dont_touch of G2747: signal is true;
	signal G2748: std_logic; attribute dont_touch of G2748: signal is true;
	signal G2752: std_logic; attribute dont_touch of G2752: signal is true;
	signal G2753: std_logic; attribute dont_touch of G2753: signal is true;
	signal G2754: std_logic; attribute dont_touch of G2754: signal is true;
	signal G2755: std_logic; attribute dont_touch of G2755: signal is true;
	signal G2756: std_logic; attribute dont_touch of G2756: signal is true;
	signal G2757: std_logic; attribute dont_touch of G2757: signal is true;
	signal G2758: std_logic; attribute dont_touch of G2758: signal is true;
	signal G2759: std_logic; attribute dont_touch of G2759: signal is true;
	signal G2760: std_logic; attribute dont_touch of G2760: signal is true;
	signal G2764: std_logic; attribute dont_touch of G2764: signal is true;
	signal G2765: std_logic; attribute dont_touch of G2765: signal is true;
	signal G2766: std_logic; attribute dont_touch of G2766: signal is true;
	signal G2767: std_logic; attribute dont_touch of G2767: signal is true;
	signal G2768: std_logic; attribute dont_touch of G2768: signal is true;
	signal G2769: std_logic; attribute dont_touch of G2769: signal is true;
	signal G2770: std_logic; attribute dont_touch of G2770: signal is true;
	signal G2771: std_logic; attribute dont_touch of G2771: signal is true;
	signal G2772: std_logic; attribute dont_touch of G2772: signal is true;
	signal G2776: std_logic; attribute dont_touch of G2776: signal is true;
	signal G2777: std_logic; attribute dont_touch of G2777: signal is true;
	signal G2778: std_logic; attribute dont_touch of G2778: signal is true;
	signal G2779: std_logic; attribute dont_touch of G2779: signal is true;
	signal G2780: std_logic; attribute dont_touch of G2780: signal is true;
	signal G2781: std_logic; attribute dont_touch of G2781: signal is true;
	signal G2782: std_logic; attribute dont_touch of G2782: signal is true;
	signal G2783: std_logic; attribute dont_touch of G2783: signal is true;
	signal G2787: std_logic; attribute dont_touch of G2787: signal is true;
	signal G2788: std_logic; attribute dont_touch of G2788: signal is true;
	signal G2789: std_logic; attribute dont_touch of G2789: signal is true;
	signal G2790: std_logic; attribute dont_touch of G2790: signal is true;
	signal G2791: std_logic; attribute dont_touch of G2791: signal is true;
	signal G2792: std_logic; attribute dont_touch of G2792: signal is true;
	signal G2793: std_logic; attribute dont_touch of G2793: signal is true;
	signal G2794: std_logic; attribute dont_touch of G2794: signal is true;
	signal G2795: std_logic; attribute dont_touch of G2795: signal is true;
	signal G2796: std_logic; attribute dont_touch of G2796: signal is true;
	signal G2800: std_logic; attribute dont_touch of G2800: signal is true;
	signal G2801: std_logic; attribute dont_touch of G2801: signal is true;
	signal G2802: std_logic; attribute dont_touch of G2802: signal is true;
	signal G2803: std_logic; attribute dont_touch of G2803: signal is true;
	signal G2804: std_logic; attribute dont_touch of G2804: signal is true;
	signal G2805: std_logic; attribute dont_touch of G2805: signal is true;
	signal G2806: std_logic; attribute dont_touch of G2806: signal is true;
	signal G2807: std_logic; attribute dont_touch of G2807: signal is true;
	signal G2808: std_logic; attribute dont_touch of G2808: signal is true;
	signal G2809: std_logic; attribute dont_touch of G2809: signal is true;
	signal G2813: std_logic; attribute dont_touch of G2813: signal is true;
	signal G2814: std_logic; attribute dont_touch of G2814: signal is true;
	signal G2817: std_logic; attribute dont_touch of G2817: signal is true;
	signal G2818: std_logic; attribute dont_touch of G2818: signal is true;
	signal G2819: std_logic; attribute dont_touch of G2819: signal is true;
	signal G2820: std_logic; attribute dont_touch of G2820: signal is true;
	signal G2821: std_logic; attribute dont_touch of G2821: signal is true;
	signal G2822: std_logic; attribute dont_touch of G2822: signal is true;
	signal G2826: std_logic; attribute dont_touch of G2826: signal is true;
	signal G2827: std_logic; attribute dont_touch of G2827: signal is true;
	signal G2828: std_logic; attribute dont_touch of G2828: signal is true;
	signal G2829: std_logic; attribute dont_touch of G2829: signal is true;
	signal G2830: std_logic; attribute dont_touch of G2830: signal is true;
	signal G2831: std_logic; attribute dont_touch of G2831: signal is true;
	signal G2834: std_logic; attribute dont_touch of G2834: signal is true;
	signal G2835: std_logic; attribute dont_touch of G2835: signal is true;
	signal G2836: std_logic; attribute dont_touch of G2836: signal is true;
	signal G2837: std_logic; attribute dont_touch of G2837: signal is true;
	signal G2838: std_logic; attribute dont_touch of G2838: signal is true;
	signal G2839: std_logic; attribute dont_touch of G2839: signal is true;
	signal G2840: std_logic; attribute dont_touch of G2840: signal is true;
	signal G2841: std_logic; attribute dont_touch of G2841: signal is true;
	signal G2842: std_logic; attribute dont_touch of G2842: signal is true;
	signal G2845: std_logic; attribute dont_touch of G2845: signal is true;
	signal G2846: std_logic; attribute dont_touch of G2846: signal is true;
	signal G2849: std_logic; attribute dont_touch of G2849: signal is true;
	signal G2850: std_logic; attribute dont_touch of G2850: signal is true;
	signal G2853: std_logic; attribute dont_touch of G2853: signal is true;
	signal G2856: std_logic; attribute dont_touch of G2856: signal is true;
	signal G2857: std_logic; attribute dont_touch of G2857: signal is true;
	signal G2858: std_logic; attribute dont_touch of G2858: signal is true;
	signal G2859: std_logic; attribute dont_touch of G2859: signal is true;
	signal G2860: std_logic; attribute dont_touch of G2860: signal is true;
	signal G2861: std_logic; attribute dont_touch of G2861: signal is true;
	signal G2862: std_logic; attribute dont_touch of G2862: signal is true;
	signal G2863: std_logic; attribute dont_touch of G2863: signal is true;
	signal G2864: std_logic; attribute dont_touch of G2864: signal is true;
	signal G2865: std_logic; attribute dont_touch of G2865: signal is true;
	signal G2866: std_logic; attribute dont_touch of G2866: signal is true;
	signal G2867: std_logic; attribute dont_touch of G2867: signal is true;
	signal G2868: std_logic; attribute dont_touch of G2868: signal is true;
	signal G2869: std_logic; attribute dont_touch of G2869: signal is true;
	signal G2870: std_logic; attribute dont_touch of G2870: signal is true;
	signal G2871: std_logic; attribute dont_touch of G2871: signal is true;
	signal G2872: std_logic; attribute dont_touch of G2872: signal is true;
	signal G2873: std_logic; attribute dont_touch of G2873: signal is true;
	signal G2874: std_logic; attribute dont_touch of G2874: signal is true;
	signal G2875: std_logic; attribute dont_touch of G2875: signal is true;
	signal G2876: std_logic; attribute dont_touch of G2876: signal is true;
	signal G2877: std_logic; attribute dont_touch of G2877: signal is true;
	signal G2882: std_logic; attribute dont_touch of G2882: signal is true;
	signal G2883: std_logic; attribute dont_touch of G2883: signal is true;
	signal G2884: std_logic; attribute dont_touch of G2884: signal is true;
	signal G2885: std_logic; attribute dont_touch of G2885: signal is true;
	signal G2886: std_logic; attribute dont_touch of G2886: signal is true;
	signal G2887: std_logic; attribute dont_touch of G2887: signal is true;
	signal G2888: std_logic; attribute dont_touch of G2888: signal is true;
	signal G2889: std_logic; attribute dont_touch of G2889: signal is true;
	signal G2890: std_logic; attribute dont_touch of G2890: signal is true;
	signal G2891: std_logic; attribute dont_touch of G2891: signal is true;
	signal G2892: std_logic; attribute dont_touch of G2892: signal is true;
	signal G2893: std_logic; attribute dont_touch of G2893: signal is true;
	signal G2894: std_logic; attribute dont_touch of G2894: signal is true;
	signal G2895: std_logic; attribute dont_touch of G2895: signal is true;
	signal G2896: std_logic; attribute dont_touch of G2896: signal is true;
	signal G2897: std_logic; attribute dont_touch of G2897: signal is true;
	signal G2902: std_logic; attribute dont_touch of G2902: signal is true;
	signal G2903: std_logic; attribute dont_touch of G2903: signal is true;
	signal G2904: std_logic; attribute dont_touch of G2904: signal is true;
	signal G2905: std_logic; attribute dont_touch of G2905: signal is true;
	signal G2906: std_logic; attribute dont_touch of G2906: signal is true;
	signal G2907: std_logic; attribute dont_touch of G2907: signal is true;
	signal G2908: std_logic; attribute dont_touch of G2908: signal is true;
	signal G2909: std_logic; attribute dont_touch of G2909: signal is true;
	signal G2912: std_logic; attribute dont_touch of G2912: signal is true;
	signal G2913: std_logic; attribute dont_touch of G2913: signal is true;
	signal G2914: std_logic; attribute dont_touch of G2914: signal is true;
	signal G2915: std_logic; attribute dont_touch of G2915: signal is true;
	signal G2916: std_logic; attribute dont_touch of G2916: signal is true;
	signal G2919: std_logic; attribute dont_touch of G2919: signal is true;
	signal G2920: std_logic; attribute dont_touch of G2920: signal is true;
	signal G2921: std_logic; attribute dont_touch of G2921: signal is true;
	signal G2922: std_logic; attribute dont_touch of G2922: signal is true;
	signal G2923: std_logic; attribute dont_touch of G2923: signal is true;
	signal G2924: std_logic; attribute dont_touch of G2924: signal is true;
	signal G2927: std_logic; attribute dont_touch of G2927: signal is true;
	signal G2928: std_logic; attribute dont_touch of G2928: signal is true;
	signal G2931: std_logic; attribute dont_touch of G2931: signal is true;
	signal G2932: std_logic; attribute dont_touch of G2932: signal is true;
	signal G2933: std_logic; attribute dont_touch of G2933: signal is true;
	signal G2934: std_logic; attribute dont_touch of G2934: signal is true;
	signal G2935: std_logic; attribute dont_touch of G2935: signal is true;
	signal G2936: std_logic; attribute dont_touch of G2936: signal is true;
	signal G2937: std_logic; attribute dont_touch of G2937: signal is true;
	signal G2940: std_logic; attribute dont_touch of G2940: signal is true;
	signal G2941: std_logic; attribute dont_touch of G2941: signal is true;
	signal G2944: std_logic; attribute dont_touch of G2944: signal is true;
	signal G2945: std_logic; attribute dont_touch of G2945: signal is true;
	signal G2946: std_logic; attribute dont_touch of G2946: signal is true;
	signal G2947: std_logic; attribute dont_touch of G2947: signal is true;
	signal G2948: std_logic; attribute dont_touch of G2948: signal is true;
	signal G2949: std_logic; attribute dont_touch of G2949: signal is true;
	signal G2950: std_logic; attribute dont_touch of G2950: signal is true;
	signal G2951: std_logic; attribute dont_touch of G2951: signal is true;
	signal G2952: std_logic; attribute dont_touch of G2952: signal is true;
	signal G2953: std_logic; attribute dont_touch of G2953: signal is true;
	signal G2954: std_logic; attribute dont_touch of G2954: signal is true;
	signal G2955: std_logic; attribute dont_touch of G2955: signal is true;
	signal G2956: std_logic; attribute dont_touch of G2956: signal is true;
	signal G2957: std_logic; attribute dont_touch of G2957: signal is true;
	signal G2958: std_logic; attribute dont_touch of G2958: signal is true;
	signal G2959: std_logic; attribute dont_touch of G2959: signal is true;
	signal G2960: std_logic; attribute dont_touch of G2960: signal is true;
	signal G2961: std_logic; attribute dont_touch of G2961: signal is true;
	signal G2962: std_logic; attribute dont_touch of G2962: signal is true;
	signal G2966: std_logic; attribute dont_touch of G2966: signal is true;
	signal G2967: std_logic; attribute dont_touch of G2967: signal is true;
	signal G2968: std_logic; attribute dont_touch of G2968: signal is true;
	signal G2973: std_logic; attribute dont_touch of G2973: signal is true;
	signal G2974: std_logic; attribute dont_touch of G2974: signal is true;
	signal G2975: std_logic; attribute dont_touch of G2975: signal is true;
	signal G2976: std_logic; attribute dont_touch of G2976: signal is true;
	signal G2981: std_logic; attribute dont_touch of G2981: signal is true;
	signal G2986: std_logic; attribute dont_touch of G2986: signal is true;
	signal G2995: std_logic; attribute dont_touch of G2995: signal is true;
	signal G2996: std_logic; attribute dont_touch of G2996: signal is true;
	signal G2997: std_logic; attribute dont_touch of G2997: signal is true;
	signal G2998: std_logic; attribute dont_touch of G2998: signal is true;
	signal G3001: std_logic; attribute dont_touch of G3001: signal is true;
	signal G3002: std_logic; attribute dont_touch of G3002: signal is true;
	signal G3007: std_logic; attribute dont_touch of G3007: signal is true;
	signal G3012: std_logic; attribute dont_touch of G3012: signal is true;
	signal G3013: std_logic; attribute dont_touch of G3013: signal is true;
	signal G3014: std_logic; attribute dont_touch of G3014: signal is true;
	signal G3015: std_logic; attribute dont_touch of G3015: signal is true;
	signal G3016: std_logic; attribute dont_touch of G3016: signal is true;
	signal G3019: std_logic; attribute dont_touch of G3019: signal is true;
	signal G3022: std_logic; attribute dont_touch of G3022: signal is true;
	signal G3023: std_logic; attribute dont_touch of G3023: signal is true;
	signal G3028: std_logic; attribute dont_touch of G3028: signal is true;
	signal G3029: std_logic; attribute dont_touch of G3029: signal is true;
	signal G3030: std_logic; attribute dont_touch of G3030: signal is true;
	signal G3031: std_logic; attribute dont_touch of G3031: signal is true;
	signal G3034: std_logic; attribute dont_touch of G3034: signal is true;
	signal G3037: std_logic; attribute dont_touch of G3037: signal is true;
	signal G3040: std_logic; attribute dont_touch of G3040: signal is true;
	signal G3041: std_logic; attribute dont_touch of G3041: signal is true;
	signal G3042: std_logic; attribute dont_touch of G3042: signal is true;
	signal G3043: std_logic; attribute dont_touch of G3043: signal is true;
	signal G3046: std_logic; attribute dont_touch of G3046: signal is true;
	signal G3049: std_logic; attribute dont_touch of G3049: signal is true;
	signal G3052: std_logic; attribute dont_touch of G3052: signal is true;
	signal G3053: std_logic; attribute dont_touch of G3053: signal is true;
	signal G3054: std_logic; attribute dont_touch of G3054: signal is true;
	signal G3057: std_logic; attribute dont_touch of G3057: signal is true;
	signal G3060: std_logic; attribute dont_touch of G3060: signal is true;
	signal G3063: std_logic; attribute dont_touch of G3063: signal is true;
	signal G3064: std_logic; attribute dont_touch of G3064: signal is true;
	signal G3067: std_logic; attribute dont_touch of G3067: signal is true;
	signal G3070: std_logic; attribute dont_touch of G3070: signal is true;
	signal G3073: std_logic; attribute dont_touch of G3073: signal is true;
	signal G3074: std_logic; attribute dont_touch of G3074: signal is true;
	signal G3075: std_logic; attribute dont_touch of G3075: signal is true;
	signal G3076: std_logic; attribute dont_touch of G3076: signal is true;
	signal G3079: std_logic; attribute dont_touch of G3079: signal is true;
	signal G3082: std_logic; attribute dont_touch of G3082: signal is true;
	signal G3083: std_logic; attribute dont_touch of G3083: signal is true;
	signal G3084: std_logic; attribute dont_touch of G3084: signal is true;
	signal G3085: std_logic; attribute dont_touch of G3085: signal is true;
	signal G3086: std_logic; attribute dont_touch of G3086: signal is true;
	signal G3089: std_logic; attribute dont_touch of G3089: signal is true;
	signal G3090: std_logic; attribute dont_touch of G3090: signal is true;
	signal G3093: std_logic; attribute dont_touch of G3093: signal is true;
	signal G3094: std_logic; attribute dont_touch of G3094: signal is true;
	signal G3095: std_logic; attribute dont_touch of G3095: signal is true;
	signal G3096: std_logic; attribute dont_touch of G3096: signal is true;
	signal G3099: std_logic; attribute dont_touch of G3099: signal is true;
	signal G3100: std_logic; attribute dont_touch of G3100: signal is true;
	signal G3103: std_logic; attribute dont_touch of G3103: signal is true;
	signal G3104: std_logic; attribute dont_touch of G3104: signal is true;
	signal G3108: std_logic; attribute dont_touch of G3108: signal is true;
	signal G3109: std_logic; attribute dont_touch of G3109: signal is true;
	signal G3110: std_logic; attribute dont_touch of G3110: signal is true;
	signal G3113: std_logic; attribute dont_touch of G3113: signal is true;
	signal G3114: std_logic; attribute dont_touch of G3114: signal is true;
	signal G3117: std_logic; attribute dont_touch of G3117: signal is true;
	signal G3118: std_logic; attribute dont_touch of G3118: signal is true;
	signal G3122: std_logic; attribute dont_touch of G3122: signal is true;
	signal G3123: std_logic; attribute dont_touch of G3123: signal is true;
	signal G3124: std_logic; attribute dont_touch of G3124: signal is true;
	signal G3127: std_logic; attribute dont_touch of G3127: signal is true;
	signal G3128: std_logic; attribute dont_touch of G3128: signal is true;
	signal G3132: std_logic; attribute dont_touch of G3132: signal is true;
	signal G3133: std_logic; attribute dont_touch of G3133: signal is true;
	signal G3134: std_logic; attribute dont_touch of G3134: signal is true;
	signal G3135: std_logic; attribute dont_touch of G3135: signal is true;
	signal G3136: std_logic; attribute dont_touch of G3136: signal is true;
	signal G3140: std_logic; attribute dont_touch of G3140: signal is true;
	signal G3143: std_logic; attribute dont_touch of G3143: signal is true;
	signal G3144: std_logic; attribute dont_touch of G3144: signal is true;
	signal G3145: std_logic; attribute dont_touch of G3145: signal is true;
	signal G3146: std_logic; attribute dont_touch of G3146: signal is true;
	signal G3147: std_logic; attribute dont_touch of G3147: signal is true;
	signal G3150: std_logic; attribute dont_touch of G3150: signal is true;
	signal G3154: std_logic; attribute dont_touch of G3154: signal is true;
	signal G3155: std_logic; attribute dont_touch of G3155: signal is true;
	signal G3156: std_logic; attribute dont_touch of G3156: signal is true;
	signal G3157: std_logic; attribute dont_touch of G3157: signal is true;
	signal G3158: std_logic; attribute dont_touch of G3158: signal is true;
	signal G3161: std_logic; attribute dont_touch of G3161: signal is true;
	signal G3162: std_logic; attribute dont_touch of G3162: signal is true;
	signal G3166: std_logic; attribute dont_touch of G3166: signal is true;
	signal G3167: std_logic; attribute dont_touch of G3167: signal is true;
	signal G3170: std_logic; attribute dont_touch of G3170: signal is true;
	signal G3171: std_logic; attribute dont_touch of G3171: signal is true;
	signal G3172: std_logic; attribute dont_touch of G3172: signal is true;
	signal G3173: std_logic; attribute dont_touch of G3173: signal is true;
	signal G3176: std_logic; attribute dont_touch of G3176: signal is true;
	signal G3177: std_logic; attribute dont_touch of G3177: signal is true;
	signal G3180: std_logic; attribute dont_touch of G3180: signal is true;
	signal G3181: std_logic; attribute dont_touch of G3181: signal is true;
	signal G3182: std_logic; attribute dont_touch of G3182: signal is true;
	signal G3183: std_logic; attribute dont_touch of G3183: signal is true;
	signal G3186: std_logic; attribute dont_touch of G3186: signal is true;
	signal G3187: std_logic; attribute dont_touch of G3187: signal is true;
	signal G3190: std_logic; attribute dont_touch of G3190: signal is true;
	signal G3191: std_logic; attribute dont_touch of G3191: signal is true;
	signal G3192: std_logic; attribute dont_touch of G3192: signal is true;
	signal G3195: std_logic; attribute dont_touch of G3195: signal is true;
	signal G3196: std_logic; attribute dont_touch of G3196: signal is true;
	signal G3199: std_logic; attribute dont_touch of G3199: signal is true;
	signal G3200: std_logic; attribute dont_touch of G3200: signal is true;
	signal G3203: std_logic; attribute dont_touch of G3203: signal is true;
	signal G3204: std_logic; attribute dont_touch of G3204: signal is true;
	signal G3207: std_logic; attribute dont_touch of G3207: signal is true;
	signal G3208: std_logic; attribute dont_touch of G3208: signal is true;
	signal G3209: std_logic; attribute dont_touch of G3209: signal is true;
	signal G3212: std_logic; attribute dont_touch of G3212: signal is true;
	signal G3215: std_logic; attribute dont_touch of G3215: signal is true;
	signal G3216: std_logic; attribute dont_touch of G3216: signal is true;
	signal G3219: std_logic; attribute dont_touch of G3219: signal is true;
	signal G3223: std_logic; attribute dont_touch of G3223: signal is true;
	signal G3224: std_logic; attribute dont_touch of G3224: signal is true;
	signal G3225: std_logic; attribute dont_touch of G3225: signal is true;
	signal G3226: std_logic; attribute dont_touch of G3226: signal is true;
	signal G3227: std_logic; attribute dont_touch of G3227: signal is true;
	signal G3228: std_logic; attribute dont_touch of G3228: signal is true;
	signal G3229: std_logic; attribute dont_touch of G3229: signal is true;
	signal G3230: std_logic; attribute dont_touch of G3230: signal is true;
	signal G3231: std_logic; attribute dont_touch of G3231: signal is true;
	signal G3232: std_logic; attribute dont_touch of G3232: signal is true;
	signal G3233: std_logic; attribute dont_touch of G3233: signal is true;
	signal G3234: std_logic; attribute dont_touch of G3234: signal is true;
	signal G3235: std_logic; attribute dont_touch of G3235: signal is true;
	signal G3236: std_logic; attribute dont_touch of G3236: signal is true;
	signal G3237: std_logic; attribute dont_touch of G3237: signal is true;
	signal G3238: std_logic; attribute dont_touch of G3238: signal is true;
	signal G3239: std_logic; attribute dont_touch of G3239: signal is true;
	signal G3240: std_logic; attribute dont_touch of G3240: signal is true;
	signal G3241: std_logic; attribute dont_touch of G3241: signal is true;
	signal G3242: std_logic; attribute dont_touch of G3242: signal is true;
	signal G3246: std_logic; attribute dont_touch of G3246: signal is true;
	signal G3247: std_logic; attribute dont_touch of G3247: signal is true;
	signal G3251: std_logic; attribute dont_touch of G3251: signal is true;
	signal G3258: std_logic; attribute dont_touch of G3258: signal is true;
	signal G3259: std_logic; attribute dont_touch of G3259: signal is true;
	signal G3263: std_logic; attribute dont_touch of G3263: signal is true;
	signal G3267: std_logic; attribute dont_touch of G3267: signal is true;
	signal G3271: std_logic; attribute dont_touch of G3271: signal is true;
	signal G3275: std_logic; attribute dont_touch of G3275: signal is true;
	signal G3276: std_logic; attribute dont_touch of G3276: signal is true;
	signal G3277: std_logic; attribute dont_touch of G3277: signal is true;
	signal G3278: std_logic; attribute dont_touch of G3278: signal is true;
	signal G3279: std_logic; attribute dont_touch of G3279: signal is true;
	signal G3280: std_logic; attribute dont_touch of G3280: signal is true;
	signal G3281: std_logic; attribute dont_touch of G3281: signal is true;
	signal G3282: std_logic; attribute dont_touch of G3282: signal is true;
	signal G3283: std_logic; attribute dont_touch of G3283: signal is true;
	signal G3284: std_logic; attribute dont_touch of G3284: signal is true;
	signal G3285: std_logic; attribute dont_touch of G3285: signal is true;
	signal G3286: std_logic; attribute dont_touch of G3286: signal is true;
	signal G3287: std_logic; attribute dont_touch of G3287: signal is true;
	signal G3288: std_logic; attribute dont_touch of G3288: signal is true;
	signal G3289: std_logic; attribute dont_touch of G3289: signal is true;
	signal G3290: std_logic; attribute dont_touch of G3290: signal is true;
	signal G3291: std_logic; attribute dont_touch of G3291: signal is true;
	signal G3292: std_logic; attribute dont_touch of G3292: signal is true;
	signal G3293: std_logic; attribute dont_touch of G3293: signal is true;
	signal G3294: std_logic; attribute dont_touch of G3294: signal is true;
	signal G3295: std_logic; attribute dont_touch of G3295: signal is true;
	signal G3296: std_logic; attribute dont_touch of G3296: signal is true;
	signal G3297: std_logic; attribute dont_touch of G3297: signal is true;
	signal G3298: std_logic; attribute dont_touch of G3298: signal is true;
	signal G3299: std_logic; attribute dont_touch of G3299: signal is true;
	signal G3300: std_logic; attribute dont_touch of G3300: signal is true;
	signal G3301: std_logic; attribute dont_touch of G3301: signal is true;
	signal G3302: std_logic; attribute dont_touch of G3302: signal is true;
	signal G3303: std_logic; attribute dont_touch of G3303: signal is true;
	signal G3304: std_logic; attribute dont_touch of G3304: signal is true;
	signal G3305: std_logic; attribute dont_touch of G3305: signal is true;
	signal G3306: std_logic; attribute dont_touch of G3306: signal is true;
	signal G3307: std_logic; attribute dont_touch of G3307: signal is true;
	signal G3308: std_logic; attribute dont_touch of G3308: signal is true;
	signal G3309: std_logic; attribute dont_touch of G3309: signal is true;
	signal G3310: std_logic; attribute dont_touch of G3310: signal is true;
	signal G3311: std_logic; attribute dont_touch of G3311: signal is true;
	signal G3312: std_logic; attribute dont_touch of G3312: signal is true;
	signal G3315: std_logic; attribute dont_touch of G3315: signal is true;
	signal G3316: std_logic; attribute dont_touch of G3316: signal is true;
	signal G3317: std_logic; attribute dont_touch of G3317: signal is true;
	signal G3318: std_logic; attribute dont_touch of G3318: signal is true;
	signal G3319: std_logic; attribute dont_touch of G3319: signal is true;
	signal G3320: std_logic; attribute dont_touch of G3320: signal is true;
	signal G3321: std_logic; attribute dont_touch of G3321: signal is true;
	signal G3322: std_logic; attribute dont_touch of G3322: signal is true;
	signal G3323: std_logic; attribute dont_touch of G3323: signal is true;
	signal G3324: std_logic; attribute dont_touch of G3324: signal is true;
	signal G3325: std_logic; attribute dont_touch of G3325: signal is true;
	signal G3326: std_logic; attribute dont_touch of G3326: signal is true;
	signal G3327: std_logic; attribute dont_touch of G3327: signal is true;
	signal G3328: std_logic; attribute dont_touch of G3328: signal is true;
	signal G3329: std_logic; attribute dont_touch of G3329: signal is true;
	signal G3330: std_logic; attribute dont_touch of G3330: signal is true;
	signal G3331: std_logic; attribute dont_touch of G3331: signal is true;
	signal G3332: std_logic; attribute dont_touch of G3332: signal is true;
	signal G3333: std_logic; attribute dont_touch of G3333: signal is true;
	signal G3334: std_logic; attribute dont_touch of G3334: signal is true;
	signal G3335: std_logic; attribute dont_touch of G3335: signal is true;
	signal G3336: std_logic; attribute dont_touch of G3336: signal is true;
	signal G3337: std_logic; attribute dont_touch of G3337: signal is true;
	signal G3338: std_logic; attribute dont_touch of G3338: signal is true;
	signal G3339: std_logic; attribute dont_touch of G3339: signal is true;
	signal G3340: std_logic; attribute dont_touch of G3340: signal is true;
	signal G3341: std_logic; attribute dont_touch of G3341: signal is true;
	signal G3342: std_logic; attribute dont_touch of G3342: signal is true;
	signal G3343: std_logic; attribute dont_touch of G3343: signal is true;
	signal G3344: std_logic; attribute dont_touch of G3344: signal is true;
	signal G3345: std_logic; attribute dont_touch of G3345: signal is true;
	signal G3346: std_logic; attribute dont_touch of G3346: signal is true;
	signal G3349: std_logic; attribute dont_touch of G3349: signal is true;
	signal G3350: std_logic; attribute dont_touch of G3350: signal is true;
	signal G3351: std_logic; attribute dont_touch of G3351: signal is true;
	signal G3352: std_logic; attribute dont_touch of G3352: signal is true;
	signal G3353: std_logic; attribute dont_touch of G3353: signal is true;
	signal G3354: std_logic; attribute dont_touch of G3354: signal is true;
	signal G3355: std_logic; attribute dont_touch of G3355: signal is true;
	signal G3356: std_logic; attribute dont_touch of G3356: signal is true;
	signal G3357: std_logic; attribute dont_touch of G3357: signal is true;
	signal G3358: std_logic; attribute dont_touch of G3358: signal is true;
	signal G3359: std_logic; attribute dont_touch of G3359: signal is true;
	signal G3360: std_logic; attribute dont_touch of G3360: signal is true;
	signal G3361: std_logic; attribute dont_touch of G3361: signal is true;
	signal G3362: std_logic; attribute dont_touch of G3362: signal is true;
	signal G3363: std_logic; attribute dont_touch of G3363: signal is true;
	signal G3364: std_logic; attribute dont_touch of G3364: signal is true;
	signal G3365: std_logic; attribute dont_touch of G3365: signal is true;
	signal G3366: std_logic; attribute dont_touch of G3366: signal is true;
	signal G3367: std_logic; attribute dont_touch of G3367: signal is true;
	signal G3368: std_logic; attribute dont_touch of G3368: signal is true;
	signal G3369: std_logic; attribute dont_touch of G3369: signal is true;
	signal G3370: std_logic; attribute dont_touch of G3370: signal is true;
	signal G3371: std_logic; attribute dont_touch of G3371: signal is true;
	signal G3372: std_logic; attribute dont_touch of G3372: signal is true;
	signal G3373: std_logic; attribute dont_touch of G3373: signal is true;
	signal G3374: std_logic; attribute dont_touch of G3374: signal is true;
	signal G3375: std_logic; attribute dont_touch of G3375: signal is true;
	signal G3376: std_logic; attribute dont_touch of G3376: signal is true;
	signal G3377: std_logic; attribute dont_touch of G3377: signal is true;
	signal G3378: std_logic; attribute dont_touch of G3378: signal is true;
	signal G3379: std_logic; attribute dont_touch of G3379: signal is true;
	signal G3380: std_logic; attribute dont_touch of G3380: signal is true;
	signal G3381: std_logic; attribute dont_touch of G3381: signal is true;
	signal G3382: std_logic; attribute dont_touch of G3382: signal is true;
	signal G3383: std_logic; attribute dont_touch of G3383: signal is true;
	signal G3384: std_logic; attribute dont_touch of G3384: signal is true;
	signal G3387: std_logic; attribute dont_touch of G3387: signal is true;
	signal G3388: std_logic; attribute dont_touch of G3388: signal is true;
	signal G3421: std_logic; attribute dont_touch of G3421: signal is true;
	signal G3424: std_logic; attribute dont_touch of G3424: signal is true;
	signal G3425: std_logic; attribute dont_touch of G3425: signal is true;
	signal G3433: std_logic; attribute dont_touch of G3433: signal is true;
	signal G3434: std_logic; attribute dont_touch of G3434: signal is true;
	signal G3437: std_logic; attribute dont_touch of G3437: signal is true;
	signal G3440: std_logic; attribute dont_touch of G3440: signal is true;
	signal G3441: std_logic; attribute dont_touch of G3441: signal is true;
	signal G3448: std_logic; attribute dont_touch of G3448: signal is true;
	signal G3449: std_logic; attribute dont_touch of G3449: signal is true;
	signal G3450: std_logic; attribute dont_touch of G3450: signal is true;
	signal G3451: std_logic; attribute dont_touch of G3451: signal is true;
	signal G3452: std_logic; attribute dont_touch of G3452: signal is true;
	signal G3453: std_logic; attribute dont_touch of G3453: signal is true;
	signal G3454: std_logic; attribute dont_touch of G3454: signal is true;
	signal G3455: std_logic; attribute dont_touch of G3455: signal is true;
	signal G3456: std_logic; attribute dont_touch of G3456: signal is true;
	signal G3457: std_logic; attribute dont_touch of G3457: signal is true;
	signal G3458: std_logic; attribute dont_touch of G3458: signal is true;
	signal G3459: std_logic; attribute dont_touch of G3459: signal is true;
	signal G3460: std_logic; attribute dont_touch of G3460: signal is true;
	signal G3461: std_logic; attribute dont_touch of G3461: signal is true;
	signal G3462: std_logic; attribute dont_touch of G3462: signal is true;
	signal G3463: std_logic; attribute dont_touch of G3463: signal is true;
	signal G3464: std_logic; attribute dont_touch of G3464: signal is true;
	signal G3465: std_logic; attribute dont_touch of G3465: signal is true;
	signal G3466: std_logic; attribute dont_touch of G3466: signal is true;
	signal G3477: std_logic; attribute dont_touch of G3477: signal is true;
	signal G3478: std_logic; attribute dont_touch of G3478: signal is true;
	signal G3479: std_logic; attribute dont_touch of G3479: signal is true;
	signal G3480: std_logic; attribute dont_touch of G3480: signal is true;
	signal G3481: std_logic; attribute dont_touch of G3481: signal is true;
	signal G3482: std_logic; attribute dont_touch of G3482: signal is true;
	signal G3483: std_logic; attribute dont_touch of G3483: signal is true;
	signal G3484: std_logic; attribute dont_touch of G3484: signal is true;
	signal G3485: std_logic; attribute dont_touch of G3485: signal is true;
	signal G3486: std_logic; attribute dont_touch of G3486: signal is true;
	signal G3487: std_logic; attribute dont_touch of G3487: signal is true;
	signal G3488: std_logic; attribute dont_touch of G3488: signal is true;
	signal G3489: std_logic; attribute dont_touch of G3489: signal is true;
	signal G3490: std_logic; attribute dont_touch of G3490: signal is true;
	signal G3491: std_logic; attribute dont_touch of G3491: signal is true;
	signal G3498: std_logic; attribute dont_touch of G3498: signal is true;
	signal G3499: std_logic; attribute dont_touch of G3499: signal is true;
	signal G3500: std_logic; attribute dont_touch of G3500: signal is true;
	signal G3501: std_logic; attribute dont_touch of G3501: signal is true;
	signal G3502: std_logic; attribute dont_touch of G3502: signal is true;
	signal G3503: std_logic; attribute dont_touch of G3503: signal is true;
	signal G3504: std_logic; attribute dont_touch of G3504: signal is true;
	signal G3505: std_logic; attribute dont_touch of G3505: signal is true;
	signal G3510: std_logic; attribute dont_touch of G3510: signal is true;
	signal G3511: std_logic; attribute dont_touch of G3511: signal is true;
	signal G3512: std_logic; attribute dont_touch of G3512: signal is true;
	signal G3517: std_logic; attribute dont_touch of G3517: signal is true;
	signal G3518: std_logic; attribute dont_touch of G3518: signal is true;
	signal G3519: std_logic; attribute dont_touch of G3519: signal is true;
	signal G3520: std_logic; attribute dont_touch of G3520: signal is true;
	signal G3521: std_logic; attribute dont_touch of G3521: signal is true;
	signal G3522: std_logic; attribute dont_touch of G3522: signal is true;
	signal G3525: std_logic; attribute dont_touch of G3525: signal is true;
	signal G3526: std_logic; attribute dont_touch of G3526: signal is true;
	signal G3527: std_logic; attribute dont_touch of G3527: signal is true;
	signal G3528: std_logic; attribute dont_touch of G3528: signal is true;
	signal G3529: std_logic; attribute dont_touch of G3529: signal is true;
	signal G3530: std_logic; attribute dont_touch of G3530: signal is true;
	signal G3531: std_logic; attribute dont_touch of G3531: signal is true;
	signal G3532: std_logic; attribute dont_touch of G3532: signal is true;
	signal G3533: std_logic; attribute dont_touch of G3533: signal is true;
	signal G3534: std_logic; attribute dont_touch of G3534: signal is true;
	signal G3535: std_logic; attribute dont_touch of G3535: signal is true;
	signal G3536: std_logic; attribute dont_touch of G3536: signal is true;
	signal G3537: std_logic; attribute dont_touch of G3537: signal is true;
	signal G3538: std_logic; attribute dont_touch of G3538: signal is true;
	signal G3539: std_logic; attribute dont_touch of G3539: signal is true;
	signal G3540: std_logic; attribute dont_touch of G3540: signal is true;
	signal G3541: std_logic; attribute dont_touch of G3541: signal is true;
	signal G3544: std_logic; attribute dont_touch of G3544: signal is true;
	signal G3545: std_logic; attribute dont_touch of G3545: signal is true;
	signal G3546: std_logic; attribute dont_touch of G3546: signal is true;
	signal G3551: std_logic; attribute dont_touch of G3551: signal is true;
	signal G3554: std_logic; attribute dont_touch of G3554: signal is true;
	signal G3557: std_logic; attribute dont_touch of G3557: signal is true;
	signal G3558: std_logic; attribute dont_touch of G3558: signal is true;
	signal G3559: std_logic; attribute dont_touch of G3559: signal is true;
	signal G3564: std_logic; attribute dont_touch of G3564: signal is true;
	signal G3567: std_logic; attribute dont_touch of G3567: signal is true;
	signal G3571: std_logic; attribute dont_touch of G3571: signal is true;
	signal G3575: std_logic; attribute dont_touch of G3575: signal is true;
	signal G3589: std_logic; attribute dont_touch of G3589: signal is true;
	signal G3593: std_logic; attribute dont_touch of G3593: signal is true;
	signal G3597: std_logic; attribute dont_touch of G3597: signal is true;
	signal G3598: std_logic; attribute dont_touch of G3598: signal is true;
	signal G3599: std_logic; attribute dont_touch of G3599: signal is true;
	signal G3601: std_logic; attribute dont_touch of G3601: signal is true;
	signal G3602: std_logic; attribute dont_touch of G3602: signal is true;
	signal G3603: std_logic; attribute dont_touch of G3603: signal is true;
	signal G3604: std_logic; attribute dont_touch of G3604: signal is true;
	signal G3605: std_logic; attribute dont_touch of G3605: signal is true;
	signal G3608: std_logic; attribute dont_touch of G3608: signal is true;
	signal G3609: std_logic; attribute dont_touch of G3609: signal is true;
	signal G3610: std_logic; attribute dont_touch of G3610: signal is true;
	signal G3611: std_logic; attribute dont_touch of G3611: signal is true;
	signal G3612: std_logic; attribute dont_touch of G3612: signal is true;
	signal G3613: std_logic; attribute dont_touch of G3613: signal is true;
	signal G3614: std_logic; attribute dont_touch of G3614: signal is true;
	signal G3615: std_logic; attribute dont_touch of G3615: signal is true;
	signal G3616: std_logic; attribute dont_touch of G3616: signal is true;
	signal G3617: std_logic; attribute dont_touch of G3617: signal is true;
	signal G3618: std_logic; attribute dont_touch of G3618: signal is true;
	signal G3619: std_logic; attribute dont_touch of G3619: signal is true;
	signal G3620: std_logic; attribute dont_touch of G3620: signal is true;
	signal G3621: std_logic; attribute dont_touch of G3621: signal is true;
	signal G3622: std_logic; attribute dont_touch of G3622: signal is true;
	signal G3625: std_logic; attribute dont_touch of G3625: signal is true;
	signal G3626: std_logic; attribute dont_touch of G3626: signal is true;
	signal G3627: std_logic; attribute dont_touch of G3627: signal is true;
	signal G3628: std_logic; attribute dont_touch of G3628: signal is true;
	signal G3629: std_logic; attribute dont_touch of G3629: signal is true;
	signal G3630: std_logic; attribute dont_touch of G3630: signal is true;
	signal G3631: std_logic; attribute dont_touch of G3631: signal is true;
	signal G3632: std_logic; attribute dont_touch of G3632: signal is true;
	signal G3633: std_logic; attribute dont_touch of G3633: signal is true;
	signal G3634: std_logic; attribute dont_touch of G3634: signal is true;
	signal G3635: std_logic; attribute dont_touch of G3635: signal is true;
	signal G3636: std_logic; attribute dont_touch of G3636: signal is true;
	signal G3637: std_logic; attribute dont_touch of G3637: signal is true;
	signal G3638: std_logic; attribute dont_touch of G3638: signal is true;
	signal G3641: std_logic; attribute dont_touch of G3641: signal is true;
	signal G3642: std_logic; attribute dont_touch of G3642: signal is true;
	signal G3643: std_logic; attribute dont_touch of G3643: signal is true;
	signal G3644: std_logic; attribute dont_touch of G3644: signal is true;
	signal G3645: std_logic; attribute dont_touch of G3645: signal is true;
	signal G3646: std_logic; attribute dont_touch of G3646: signal is true;
	signal G3647: std_logic; attribute dont_touch of G3647: signal is true;
	signal G3648: std_logic; attribute dont_touch of G3648: signal is true;
	signal G3649: std_logic; attribute dont_touch of G3649: signal is true;
	signal G3650: std_logic; attribute dont_touch of G3650: signal is true;
	signal G3651: std_logic; attribute dont_touch of G3651: signal is true;
	signal G3652: std_logic; attribute dont_touch of G3652: signal is true;
	signal G3653: std_logic; attribute dont_touch of G3653: signal is true;
	signal G3654: std_logic; attribute dont_touch of G3654: signal is true;
	signal G3655: std_logic; attribute dont_touch of G3655: signal is true;
	signal G3656: std_logic; attribute dont_touch of G3656: signal is true;
	signal G3657: std_logic; attribute dont_touch of G3657: signal is true;
	signal G3658: std_logic; attribute dont_touch of G3658: signal is true;
	signal G3659: std_logic; attribute dont_touch of G3659: signal is true;
	signal G3660: std_logic; attribute dont_touch of G3660: signal is true;
	signal G3661: std_logic; attribute dont_touch of G3661: signal is true;
	signal G3662: std_logic; attribute dont_touch of G3662: signal is true;
	signal G3663: std_logic; attribute dont_touch of G3663: signal is true;
	signal G3664: std_logic; attribute dont_touch of G3664: signal is true;
	signal G3665: std_logic; attribute dont_touch of G3665: signal is true;
	signal G3666: std_logic; attribute dont_touch of G3666: signal is true;
	signal G3667: std_logic; attribute dont_touch of G3667: signal is true;
	signal G3668: std_logic; attribute dont_touch of G3668: signal is true;
	signal G3669: std_logic; attribute dont_touch of G3669: signal is true;
	signal G3670: std_logic; attribute dont_touch of G3670: signal is true;
	signal G3671: std_logic; attribute dont_touch of G3671: signal is true;
	signal G3672: std_logic; attribute dont_touch of G3672: signal is true;
	signal G3673: std_logic; attribute dont_touch of G3673: signal is true;
	signal G3677: std_logic; attribute dont_touch of G3677: signal is true;
	signal G3678: std_logic; attribute dont_touch of G3678: signal is true;
	signal G3679: std_logic; attribute dont_touch of G3679: signal is true;
	signal G3680: std_logic; attribute dont_touch of G3680: signal is true;
	signal G3681: std_logic; attribute dont_touch of G3681: signal is true;
	signal G3682: std_logic; attribute dont_touch of G3682: signal is true;
	signal G3683: std_logic; attribute dont_touch of G3683: signal is true;
	signal G3684: std_logic; attribute dont_touch of G3684: signal is true;
	signal G3685: std_logic; attribute dont_touch of G3685: signal is true;
	signal G3686: std_logic; attribute dont_touch of G3686: signal is true;
	signal G3687: std_logic; attribute dont_touch of G3687: signal is true;
	signal G3688: std_logic; attribute dont_touch of G3688: signal is true;
	signal G3689: std_logic; attribute dont_touch of G3689: signal is true;
	signal G3690: std_logic; attribute dont_touch of G3690: signal is true;
	signal G3691: std_logic; attribute dont_touch of G3691: signal is true;
	signal G3692: std_logic; attribute dont_touch of G3692: signal is true;
	signal G3693: std_logic; attribute dont_touch of G3693: signal is true;
	signal G3694: std_logic; attribute dont_touch of G3694: signal is true;
	signal G3697: std_logic; attribute dont_touch of G3697: signal is true;
	signal G3698: std_logic; attribute dont_touch of G3698: signal is true;
	signal G3699: std_logic; attribute dont_touch of G3699: signal is true;
	signal G3700: std_logic; attribute dont_touch of G3700: signal is true;
	signal G3701: std_logic; attribute dont_touch of G3701: signal is true;
	signal G3702: std_logic; attribute dont_touch of G3702: signal is true;
	signal G3703: std_logic; attribute dont_touch of G3703: signal is true;
	signal G3704: std_logic; attribute dont_touch of G3704: signal is true;
	signal G3705: std_logic; attribute dont_touch of G3705: signal is true;
	signal G3709: std_logic; attribute dont_touch of G3709: signal is true;
	signal G3710: std_logic; attribute dont_touch of G3710: signal is true;
	signal G3714: std_logic; attribute dont_touch of G3714: signal is true;
	signal G3718: std_logic; attribute dont_touch of G3718: signal is true;
	signal G3719: std_logic; attribute dont_touch of G3719: signal is true;
	signal G3723: std_logic; attribute dont_touch of G3723: signal is true;
	signal G3724: std_logic; attribute dont_touch of G3724: signal is true;
	signal G3725: std_logic; attribute dont_touch of G3725: signal is true;
	signal G3726: std_logic; attribute dont_touch of G3726: signal is true;
	signal G3727: std_logic; attribute dont_touch of G3727: signal is true;
	signal G3728: std_logic; attribute dont_touch of G3728: signal is true;
	signal G3729: std_logic; attribute dont_touch of G3729: signal is true;
	signal G3730: std_logic; attribute dont_touch of G3730: signal is true;
	signal G3731: std_logic; attribute dont_touch of G3731: signal is true;
	signal G3732: std_logic; attribute dont_touch of G3732: signal is true;
	signal G3733: std_logic; attribute dont_touch of G3733: signal is true;
	signal G3739: std_logic; attribute dont_touch of G3739: signal is true;
	signal G3740: std_logic; attribute dont_touch of G3740: signal is true;
	signal G3741: std_logic; attribute dont_touch of G3741: signal is true;
	signal G3742: std_logic; attribute dont_touch of G3742: signal is true;
	signal G3743: std_logic; attribute dont_touch of G3743: signal is true;
	signal G3744: std_logic; attribute dont_touch of G3744: signal is true;
	signal G3745: std_logic; attribute dont_touch of G3745: signal is true;
	signal G3746: std_logic; attribute dont_touch of G3746: signal is true;
	signal G3747: std_logic; attribute dont_touch of G3747: signal is true;
	signal G3748: std_logic; attribute dont_touch of G3748: signal is true;
	signal G3749: std_logic; attribute dont_touch of G3749: signal is true;
	signal G3750: std_logic; attribute dont_touch of G3750: signal is true;
	signal G3751: std_logic; attribute dont_touch of G3751: signal is true;
	signal G3752: std_logic; attribute dont_touch of G3752: signal is true;
	signal G3755: std_logic; attribute dont_touch of G3755: signal is true;
	signal G3756: std_logic; attribute dont_touch of G3756: signal is true;
	signal G3757: std_logic; attribute dont_touch of G3757: signal is true;
	signal G3758: std_logic; attribute dont_touch of G3758: signal is true;
	signal G3759: std_logic; attribute dont_touch of G3759: signal is true;
	signal G3760: std_logic; attribute dont_touch of G3760: signal is true;
	signal G3761: std_logic; attribute dont_touch of G3761: signal is true;
	signal G3762: std_logic; attribute dont_touch of G3762: signal is true;
	signal G3763: std_logic; attribute dont_touch of G3763: signal is true;
	signal G3764: std_logic; attribute dont_touch of G3764: signal is true;
	signal G3765: std_logic; attribute dont_touch of G3765: signal is true;
	signal G3766: std_logic; attribute dont_touch of G3766: signal is true;
	signal G3767: std_logic; attribute dont_touch of G3767: signal is true;
	signal G3768: std_logic; attribute dont_touch of G3768: signal is true;
	signal G3769: std_logic; attribute dont_touch of G3769: signal is true;
	signal G3770: std_logic; attribute dont_touch of G3770: signal is true;
	signal G3771: std_logic; attribute dont_touch of G3771: signal is true;
	signal G3772: std_logic; attribute dont_touch of G3772: signal is true;
	signal G3773: std_logic; attribute dont_touch of G3773: signal is true;
	signal G3774: std_logic; attribute dont_touch of G3774: signal is true;
	signal G3775: std_logic; attribute dont_touch of G3775: signal is true;
	signal G3776: std_logic; attribute dont_touch of G3776: signal is true;
	signal G3777: std_logic; attribute dont_touch of G3777: signal is true;
	signal G3778: std_logic; attribute dont_touch of G3778: signal is true;
	signal G3779: std_logic; attribute dont_touch of G3779: signal is true;
	signal G3780: std_logic; attribute dont_touch of G3780: signal is true;
	signal G3781: std_logic; attribute dont_touch of G3781: signal is true;
	signal G3782: std_logic; attribute dont_touch of G3782: signal is true;
	signal G3783: std_logic; attribute dont_touch of G3783: signal is true;
	signal G3784: std_logic; attribute dont_touch of G3784: signal is true;
	signal G3785: std_logic; attribute dont_touch of G3785: signal is true;
	signal G3786: std_logic; attribute dont_touch of G3786: signal is true;
	signal G3787: std_logic; attribute dont_touch of G3787: signal is true;
	signal G3788: std_logic; attribute dont_touch of G3788: signal is true;
	signal G3789: std_logic; attribute dont_touch of G3789: signal is true;
	signal G3790: std_logic; attribute dont_touch of G3790: signal is true;
	signal G3791: std_logic; attribute dont_touch of G3791: signal is true;
	signal G3792: std_logic; attribute dont_touch of G3792: signal is true;
	signal G3793: std_logic; attribute dont_touch of G3793: signal is true;
	signal G3796: std_logic; attribute dont_touch of G3796: signal is true;
	signal G3797: std_logic; attribute dont_touch of G3797: signal is true;
	signal G3798: std_logic; attribute dont_touch of G3798: signal is true;
	signal G3799: std_logic; attribute dont_touch of G3799: signal is true;
	signal G3800: std_logic; attribute dont_touch of G3800: signal is true;
	signal G3801: std_logic; attribute dont_touch of G3801: signal is true;
	signal G3802: std_logic; attribute dont_touch of G3802: signal is true;
	signal G3803: std_logic; attribute dont_touch of G3803: signal is true;
	signal G3806: std_logic; attribute dont_touch of G3806: signal is true;
	signal G3807: std_logic; attribute dont_touch of G3807: signal is true;
	signal G3810: std_logic; attribute dont_touch of G3810: signal is true;
	signal G3813: std_logic; attribute dont_touch of G3813: signal is true;
	signal G3814: std_logic; attribute dont_touch of G3814: signal is true;
	signal G3815: std_logic; attribute dont_touch of G3815: signal is true;
	signal G3816: std_logic; attribute dont_touch of G3816: signal is true;
	signal G3819: std_logic; attribute dont_touch of G3819: signal is true;
	signal G3820: std_logic; attribute dont_touch of G3820: signal is true;
	signal G3821: std_logic; attribute dont_touch of G3821: signal is true;
	signal G3828: std_logic; attribute dont_touch of G3828: signal is true;
	signal G3829: std_logic; attribute dont_touch of G3829: signal is true;
	signal G3830: std_logic; attribute dont_touch of G3830: signal is true;
	signal G3831: std_logic; attribute dont_touch of G3831: signal is true;
	signal G3832: std_logic; attribute dont_touch of G3832: signal is true;
	signal G3833: std_logic; attribute dont_touch of G3833: signal is true;
	signal G3834: std_logic; attribute dont_touch of G3834: signal is true;
	signal G3835: std_logic; attribute dont_touch of G3835: signal is true;
	signal G3836: std_logic; attribute dont_touch of G3836: signal is true;
	signal G3837: std_logic; attribute dont_touch of G3837: signal is true;
	signal G3838: std_logic; attribute dont_touch of G3838: signal is true;
	signal G3839: std_logic; attribute dont_touch of G3839: signal is true;
	signal G3840: std_logic; attribute dont_touch of G3840: signal is true;
	signal G3841: std_logic; attribute dont_touch of G3841: signal is true;
	signal G3842: std_logic; attribute dont_touch of G3842: signal is true;
	signal G3843: std_logic; attribute dont_touch of G3843: signal is true;
	signal G3844: std_logic; attribute dont_touch of G3844: signal is true;
	signal G3845: std_logic; attribute dont_touch of G3845: signal is true;
	signal G3846: std_logic; attribute dont_touch of G3846: signal is true;
	signal G3847: std_logic; attribute dont_touch of G3847: signal is true;
	signal G3848: std_logic; attribute dont_touch of G3848: signal is true;
	signal G3849: std_logic; attribute dont_touch of G3849: signal is true;
	signal G3850: std_logic; attribute dont_touch of G3850: signal is true;
	signal G3851: std_logic; attribute dont_touch of G3851: signal is true;
	signal G3852: std_logic; attribute dont_touch of G3852: signal is true;
	signal G3853: std_logic; attribute dont_touch of G3853: signal is true;
	signal G3854: std_logic; attribute dont_touch of G3854: signal is true;
	signal G3855: std_logic; attribute dont_touch of G3855: signal is true;
	signal G3856: std_logic; attribute dont_touch of G3856: signal is true;
	signal G3857: std_logic; attribute dont_touch of G3857: signal is true;
	signal G3858: std_logic; attribute dont_touch of G3858: signal is true;
	signal G3859: std_logic; attribute dont_touch of G3859: signal is true;
	signal G3860: std_logic; attribute dont_touch of G3860: signal is true;
	signal G3861: std_logic; attribute dont_touch of G3861: signal is true;
	signal G3862: std_logic; attribute dont_touch of G3862: signal is true;
	signal G3863: std_logic; attribute dont_touch of G3863: signal is true;
	signal G3864: std_logic; attribute dont_touch of G3864: signal is true;
	signal G3865: std_logic; attribute dont_touch of G3865: signal is true;
	signal G3866: std_logic; attribute dont_touch of G3866: signal is true;
	signal G3867: std_logic; attribute dont_touch of G3867: signal is true;
	signal G3868: std_logic; attribute dont_touch of G3868: signal is true;
	signal G3869: std_logic; attribute dont_touch of G3869: signal is true;
	signal G3870: std_logic; attribute dont_touch of G3870: signal is true;
	signal G3871: std_logic; attribute dont_touch of G3871: signal is true;
	signal G3872: std_logic; attribute dont_touch of G3872: signal is true;
	signal G3873: std_logic; attribute dont_touch of G3873: signal is true;
	signal G3874: std_logic; attribute dont_touch of G3874: signal is true;
	signal G3875: std_logic; attribute dont_touch of G3875: signal is true;
	signal G3876: std_logic; attribute dont_touch of G3876: signal is true;
	signal G3877: std_logic; attribute dont_touch of G3877: signal is true;
	signal G3878: std_logic; attribute dont_touch of G3878: signal is true;
	signal G3879: std_logic; attribute dont_touch of G3879: signal is true;
	signal G3880: std_logic; attribute dont_touch of G3880: signal is true;
	signal G3881: std_logic; attribute dont_touch of G3881: signal is true;
	signal G3882: std_logic; attribute dont_touch of G3882: signal is true;
	signal G3883: std_logic; attribute dont_touch of G3883: signal is true;
	signal G3884: std_logic; attribute dont_touch of G3884: signal is true;
	signal G3885: std_logic; attribute dont_touch of G3885: signal is true;
	signal G3886: std_logic; attribute dont_touch of G3886: signal is true;
	signal G3887: std_logic; attribute dont_touch of G3887: signal is true;
	signal G3888: std_logic; attribute dont_touch of G3888: signal is true;
	signal G3889: std_logic; attribute dont_touch of G3889: signal is true;
	signal G3890: std_logic; attribute dont_touch of G3890: signal is true;
	signal G3891: std_logic; attribute dont_touch of G3891: signal is true;
	signal G3892: std_logic; attribute dont_touch of G3892: signal is true;
	signal G3893: std_logic; attribute dont_touch of G3893: signal is true;
	signal G3896: std_logic; attribute dont_touch of G3896: signal is true;
	signal G3897: std_logic; attribute dont_touch of G3897: signal is true;
	signal G3898: std_logic; attribute dont_touch of G3898: signal is true;
	signal G3899: std_logic; attribute dont_touch of G3899: signal is true;
	signal G3900: std_logic; attribute dont_touch of G3900: signal is true;
	signal G3901: std_logic; attribute dont_touch of G3901: signal is true;
	signal G3902: std_logic; attribute dont_touch of G3902: signal is true;
	signal G3903: std_logic; attribute dont_touch of G3903: signal is true;
	signal G3904: std_logic; attribute dont_touch of G3904: signal is true;
	signal G3905: std_logic; attribute dont_touch of G3905: signal is true;
	signal G3906: std_logic; attribute dont_touch of G3906: signal is true;
	signal G3907: std_logic; attribute dont_touch of G3907: signal is true;
	signal G3910: std_logic; attribute dont_touch of G3910: signal is true;
	signal G3911: std_logic; attribute dont_touch of G3911: signal is true;
	signal G3912: std_logic; attribute dont_touch of G3912: signal is true;
	signal G3913: std_logic; attribute dont_touch of G3913: signal is true;
	signal G3914: std_logic; attribute dont_touch of G3914: signal is true;
	signal G3921: std_logic; attribute dont_touch of G3921: signal is true;
	signal G3922: std_logic; attribute dont_touch of G3922: signal is true;
	signal G3923: std_logic; attribute dont_touch of G3923: signal is true;
	signal G3924: std_logic; attribute dont_touch of G3924: signal is true;
	signal G3925: std_logic; attribute dont_touch of G3925: signal is true;
	signal G3926: std_logic; attribute dont_touch of G3926: signal is true;
	signal G3927: std_logic; attribute dont_touch of G3927: signal is true;
	signal G3928: std_logic; attribute dont_touch of G3928: signal is true;
	signal G3929: std_logic; attribute dont_touch of G3929: signal is true;
	signal G3930: std_logic; attribute dont_touch of G3930: signal is true;
	signal G3931: std_logic; attribute dont_touch of G3931: signal is true;
	signal G3932: std_logic; attribute dont_touch of G3932: signal is true;
	signal G3933: std_logic; attribute dont_touch of G3933: signal is true;
	signal G3934: std_logic; attribute dont_touch of G3934: signal is true;
	signal G3935: std_logic; attribute dont_touch of G3935: signal is true;
	signal G3936: std_logic; attribute dont_touch of G3936: signal is true;
	signal G3939: std_logic; attribute dont_touch of G3939: signal is true;
	signal G3940: std_logic; attribute dont_touch of G3940: signal is true;
	signal G3941: std_logic; attribute dont_touch of G3941: signal is true;
	signal G3942: std_logic; attribute dont_touch of G3942: signal is true;
	signal G3952: std_logic; attribute dont_touch of G3952: signal is true;
	signal G3953: std_logic; attribute dont_touch of G3953: signal is true;
	signal G3954: std_logic; attribute dont_touch of G3954: signal is true;
	signal G3955: std_logic; attribute dont_touch of G3955: signal is true;
	signal G3956: std_logic; attribute dont_touch of G3956: signal is true;
	signal G3957: std_logic; attribute dont_touch of G3957: signal is true;
	signal G3958: std_logic; attribute dont_touch of G3958: signal is true;
	signal G3959: std_logic; attribute dont_touch of G3959: signal is true;
	signal G3960: std_logic; attribute dont_touch of G3960: signal is true;
	signal G3961: std_logic; attribute dont_touch of G3961: signal is true;
	signal G3962: std_logic; attribute dont_touch of G3962: signal is true;
	signal G3963: std_logic; attribute dont_touch of G3963: signal is true;
	signal G3964: std_logic; attribute dont_touch of G3964: signal is true;
	signal G3965: std_logic; attribute dont_touch of G3965: signal is true;
	signal G3966: std_logic; attribute dont_touch of G3966: signal is true;
	signal G3967: std_logic; attribute dont_touch of G3967: signal is true;
	signal G3968: std_logic; attribute dont_touch of G3968: signal is true;
	signal G3969: std_logic; attribute dont_touch of G3969: signal is true;
	signal G3970: std_logic; attribute dont_touch of G3970: signal is true;
	signal G3971: std_logic; attribute dont_touch of G3971: signal is true;
	signal G3972: std_logic; attribute dont_touch of G3972: signal is true;
	signal G3973: std_logic; attribute dont_touch of G3973: signal is true;
	signal G3974: std_logic; attribute dont_touch of G3974: signal is true;
	signal G3975: std_logic; attribute dont_touch of G3975: signal is true;
	signal G3976: std_logic; attribute dont_touch of G3976: signal is true;
	signal G3977: std_logic; attribute dont_touch of G3977: signal is true;
	signal G3978: std_logic; attribute dont_touch of G3978: signal is true;
	signal G3979: std_logic; attribute dont_touch of G3979: signal is true;
	signal G3980: std_logic; attribute dont_touch of G3980: signal is true;
	signal G3981: std_logic; attribute dont_touch of G3981: signal is true;
	signal G3982: std_logic; attribute dont_touch of G3982: signal is true;
	signal G3983: std_logic; attribute dont_touch of G3983: signal is true;
	signal G3984: std_logic; attribute dont_touch of G3984: signal is true;
	signal G3985: std_logic; attribute dont_touch of G3985: signal is true;
	signal G3986: std_logic; attribute dont_touch of G3986: signal is true;
	signal G3987: std_logic; attribute dont_touch of G3987: signal is true;
	signal G3988: std_logic; attribute dont_touch of G3988: signal is true;
	signal G3989: std_logic; attribute dont_touch of G3989: signal is true;
	signal G3990: std_logic; attribute dont_touch of G3990: signal is true;
	signal G3991: std_logic; attribute dont_touch of G3991: signal is true;
	signal G3992: std_logic; attribute dont_touch of G3992: signal is true;
	signal G3995: std_logic; attribute dont_touch of G3995: signal is true;
	signal G3996: std_logic; attribute dont_touch of G3996: signal is true;
	signal G3997: std_logic; attribute dont_touch of G3997: signal is true;
	signal G3998: std_logic; attribute dont_touch of G3998: signal is true;
	signal G3999: std_logic; attribute dont_touch of G3999: signal is true;
	signal G4000: std_logic; attribute dont_touch of G4000: signal is true;
	signal G4001: std_logic; attribute dont_touch of G4001: signal is true;
	signal G4002: std_logic; attribute dont_touch of G4002: signal is true;
	signal G4003: std_logic; attribute dont_touch of G4003: signal is true;
	signal G4004: std_logic; attribute dont_touch of G4004: signal is true;
	signal G4007: std_logic; attribute dont_touch of G4007: signal is true;
	signal G4010: std_logic; attribute dont_touch of G4010: signal is true;
	signal G4011: std_logic; attribute dont_touch of G4011: signal is true;
	signal G4014: std_logic; attribute dont_touch of G4014: signal is true;
	signal G4015: std_logic; attribute dont_touch of G4015: signal is true;
	signal G4016: std_logic; attribute dont_touch of G4016: signal is true;
	signal G4017: std_logic; attribute dont_touch of G4017: signal is true;
	signal G4020: std_logic; attribute dont_touch of G4020: signal is true;
	signal G4021: std_logic; attribute dont_touch of G4021: signal is true;
	signal G4022: std_logic; attribute dont_touch of G4022: signal is true;
	signal G4032: std_logic; attribute dont_touch of G4032: signal is true;
	signal G4033: std_logic; attribute dont_touch of G4033: signal is true;
	signal G4034: std_logic; attribute dont_touch of G4034: signal is true;
	signal G4035: std_logic; attribute dont_touch of G4035: signal is true;
	signal G4036: std_logic; attribute dont_touch of G4036: signal is true;
	signal G4037: std_logic; attribute dont_touch of G4037: signal is true;
	signal G4038: std_logic; attribute dont_touch of G4038: signal is true;
	signal G4039: std_logic; attribute dont_touch of G4039: signal is true;
	signal G4040: std_logic; attribute dont_touch of G4040: signal is true;
	signal G4041: std_logic; attribute dont_touch of G4041: signal is true;
	signal G4042: std_logic; attribute dont_touch of G4042: signal is true;
	signal G4043: std_logic; attribute dont_touch of G4043: signal is true;
	signal G4044: std_logic; attribute dont_touch of G4044: signal is true;
	signal G4045: std_logic; attribute dont_touch of G4045: signal is true;
	signal G4046: std_logic; attribute dont_touch of G4046: signal is true;
	signal G4047: std_logic; attribute dont_touch of G4047: signal is true;
	signal G4048: std_logic; attribute dont_touch of G4048: signal is true;
	signal G4049: std_logic; attribute dont_touch of G4049: signal is true;
	signal G4050: std_logic; attribute dont_touch of G4050: signal is true;
	signal G4051: std_logic; attribute dont_touch of G4051: signal is true;
	signal G4052: std_logic; attribute dont_touch of G4052: signal is true;
	signal G4053: std_logic; attribute dont_touch of G4053: signal is true;
	signal G4054: std_logic; attribute dont_touch of G4054: signal is true;
	signal G4057: std_logic; attribute dont_touch of G4057: signal is true;
	signal G4058: std_logic; attribute dont_touch of G4058: signal is true;
	signal G4059: std_logic; attribute dont_touch of G4059: signal is true;
	signal G4068: std_logic; attribute dont_touch of G4068: signal is true;
	signal G4074: std_logic; attribute dont_touch of G4074: signal is true;
	signal G4080: std_logic; attribute dont_touch of G4080: signal is true;
	signal G4086: std_logic; attribute dont_touch of G4086: signal is true;
	signal G4092: std_logic; attribute dont_touch of G4092: signal is true;
	signal G4111: std_logic; attribute dont_touch of G4111: signal is true;
	signal G4113: std_logic; attribute dont_touch of G4113: signal is true;
	signal G4114: std_logic; attribute dont_touch of G4114: signal is true;
	signal G4115: std_logic; attribute dont_touch of G4115: signal is true;
	signal G4116: std_logic; attribute dont_touch of G4116: signal is true;
	signal G4117: std_logic; attribute dont_touch of G4117: signal is true;
	signal G4118: std_logic; attribute dont_touch of G4118: signal is true;
	signal G4119: std_logic; attribute dont_touch of G4119: signal is true;
	signal G4120: std_logic; attribute dont_touch of G4120: signal is true;
	signal G4122: std_logic; attribute dont_touch of G4122: signal is true;
	signal G4123: std_logic; attribute dont_touch of G4123: signal is true;
	signal G4124: std_logic; attribute dont_touch of G4124: signal is true;
	signal G4125: std_logic; attribute dont_touch of G4125: signal is true;
	signal G4126: std_logic; attribute dont_touch of G4126: signal is true;
	signal G4127: std_logic; attribute dont_touch of G4127: signal is true;
	signal G4128: std_logic; attribute dont_touch of G4128: signal is true;
	signal G4129: std_logic; attribute dont_touch of G4129: signal is true;
	signal G4130: std_logic; attribute dont_touch of G4130: signal is true;
	signal G4131: std_logic; attribute dont_touch of G4131: signal is true;
	signal G4132: std_logic; attribute dont_touch of G4132: signal is true;
	signal G4133: std_logic; attribute dont_touch of G4133: signal is true;
	signal G4134: std_logic; attribute dont_touch of G4134: signal is true;
	signal G4135: std_logic; attribute dont_touch of G4135: signal is true;
	signal G4136: std_logic; attribute dont_touch of G4136: signal is true;
	signal G4137: std_logic; attribute dont_touch of G4137: signal is true;
	signal G4138: std_logic; attribute dont_touch of G4138: signal is true;
	signal G4139: std_logic; attribute dont_touch of G4139: signal is true;
	signal G4140: std_logic; attribute dont_touch of G4140: signal is true;
	signal G4141: std_logic; attribute dont_touch of G4141: signal is true;
	signal G4142: std_logic; attribute dont_touch of G4142: signal is true;
	signal G4143: std_logic; attribute dont_touch of G4143: signal is true;
	signal G4144: std_logic; attribute dont_touch of G4144: signal is true;
	signal G4145: std_logic; attribute dont_touch of G4145: signal is true;
	signal G4146: std_logic; attribute dont_touch of G4146: signal is true;
	signal G4147: std_logic; attribute dont_touch of G4147: signal is true;
	signal G4148: std_logic; attribute dont_touch of G4148: signal is true;
	signal G4149: std_logic; attribute dont_touch of G4149: signal is true;
	signal G4150: std_logic; attribute dont_touch of G4150: signal is true;
	signal G4151: std_logic; attribute dont_touch of G4151: signal is true;
	signal G4152: std_logic; attribute dont_touch of G4152: signal is true;
	signal G4153: std_logic; attribute dont_touch of G4153: signal is true;
	signal G4154: std_logic; attribute dont_touch of G4154: signal is true;
	signal G4155: std_logic; attribute dont_touch of G4155: signal is true;
	signal G4156: std_logic; attribute dont_touch of G4156: signal is true;
	signal G4157: std_logic; attribute dont_touch of G4157: signal is true;
	signal G4158: std_logic; attribute dont_touch of G4158: signal is true;
	signal G4159: std_logic; attribute dont_touch of G4159: signal is true;
	signal G4160: std_logic; attribute dont_touch of G4160: signal is true;
	signal G4161: std_logic; attribute dont_touch of G4161: signal is true;
	signal G4162: std_logic; attribute dont_touch of G4162: signal is true;
	signal G4163: std_logic; attribute dont_touch of G4163: signal is true;
	signal G4164: std_logic; attribute dont_touch of G4164: signal is true;
	signal G4165: std_logic; attribute dont_touch of G4165: signal is true;
	signal G4166: std_logic; attribute dont_touch of G4166: signal is true;
	signal G4167: std_logic; attribute dont_touch of G4167: signal is true;
	signal G4168: std_logic; attribute dont_touch of G4168: signal is true;
	signal G4169: std_logic; attribute dont_touch of G4169: signal is true;
	signal G4170: std_logic; attribute dont_touch of G4170: signal is true;
	signal G4171: std_logic; attribute dont_touch of G4171: signal is true;
	signal G4172: std_logic; attribute dont_touch of G4172: signal is true;
	signal G4173: std_logic; attribute dont_touch of G4173: signal is true;
	signal G4176: std_logic; attribute dont_touch of G4176: signal is true;
	signal G4177: std_logic; attribute dont_touch of G4177: signal is true;
	signal G4178: std_logic; attribute dont_touch of G4178: signal is true;
	signal G4179: std_logic; attribute dont_touch of G4179: signal is true;
	signal G4180: std_logic; attribute dont_touch of G4180: signal is true;
	signal G4181: std_logic; attribute dont_touch of G4181: signal is true;
	signal G4182: std_logic; attribute dont_touch of G4182: signal is true;
	signal G4183: std_logic; attribute dont_touch of G4183: signal is true;
	signal G4184: std_logic; attribute dont_touch of G4184: signal is true;
	signal G4185: std_logic; attribute dont_touch of G4185: signal is true;
	signal G4186: std_logic; attribute dont_touch of G4186: signal is true;
	signal G4187: std_logic; attribute dont_touch of G4187: signal is true;
	signal G4188: std_logic; attribute dont_touch of G4188: signal is true;
	signal G4189: std_logic; attribute dont_touch of G4189: signal is true;
	signal G4190: std_logic; attribute dont_touch of G4190: signal is true;
	signal G4191: std_logic; attribute dont_touch of G4191: signal is true;
	signal G4192: std_logic; attribute dont_touch of G4192: signal is true;
	signal G4193: std_logic; attribute dont_touch of G4193: signal is true;
	signal G4194: std_logic; attribute dont_touch of G4194: signal is true;
	signal G4195: std_logic; attribute dont_touch of G4195: signal is true;
	signal G4198: std_logic; attribute dont_touch of G4198: signal is true;
	signal G4199: std_logic; attribute dont_touch of G4199: signal is true;
	signal G4202: std_logic; attribute dont_touch of G4202: signal is true;
	signal G4205: std_logic; attribute dont_touch of G4205: signal is true;
	signal G4206: std_logic; attribute dont_touch of G4206: signal is true;
	signal G4209: std_logic; attribute dont_touch of G4209: signal is true;
	signal G4210: std_logic; attribute dont_touch of G4210: signal is true;
	signal G4213: std_logic; attribute dont_touch of G4213: signal is true;
	signal G4214: std_logic; attribute dont_touch of G4214: signal is true;
	signal G4215: std_logic; attribute dont_touch of G4215: signal is true;
	signal G4218: std_logic; attribute dont_touch of G4218: signal is true;
	signal G4219: std_logic; attribute dont_touch of G4219: signal is true;
	signal G4220: std_logic; attribute dont_touch of G4220: signal is true;
	signal G4221: std_logic; attribute dont_touch of G4221: signal is true;
	signal G4222: std_logic; attribute dont_touch of G4222: signal is true;
	signal G4223: std_logic; attribute dont_touch of G4223: signal is true;
	signal G4224: std_logic; attribute dont_touch of G4224: signal is true;
	signal G4225: std_logic; attribute dont_touch of G4225: signal is true;
	signal G4226: std_logic; attribute dont_touch of G4226: signal is true;
	signal G4227: std_logic; attribute dont_touch of G4227: signal is true;
	signal G4228: std_logic; attribute dont_touch of G4228: signal is true;
	signal G4229: std_logic; attribute dont_touch of G4229: signal is true;
	signal G4230: std_logic; attribute dont_touch of G4230: signal is true;
	signal G4231: std_logic; attribute dont_touch of G4231: signal is true;
	signal G4232: std_logic; attribute dont_touch of G4232: signal is true;
	signal G4233: std_logic; attribute dont_touch of G4233: signal is true;
	signal G4234: std_logic; attribute dont_touch of G4234: signal is true;
	signal G4235: std_logic; attribute dont_touch of G4235: signal is true;
	signal G4236: std_logic; attribute dont_touch of G4236: signal is true;
	signal G4237: std_logic; attribute dont_touch of G4237: signal is true;
	signal G4238: std_logic; attribute dont_touch of G4238: signal is true;
	signal G4239: std_logic; attribute dont_touch of G4239: signal is true;
	signal G4240: std_logic; attribute dont_touch of G4240: signal is true;
	signal G4241: std_logic; attribute dont_touch of G4241: signal is true;
	signal G4242: std_logic; attribute dont_touch of G4242: signal is true;
	signal G4243: std_logic; attribute dont_touch of G4243: signal is true;
	signal G4244: std_logic; attribute dont_touch of G4244: signal is true;
	signal G4245: std_logic; attribute dont_touch of G4245: signal is true;
	signal G4246: std_logic; attribute dont_touch of G4246: signal is true;
	signal G4247: std_logic; attribute dont_touch of G4247: signal is true;
	signal G4248: std_logic; attribute dont_touch of G4248: signal is true;
	signal G4249: std_logic; attribute dont_touch of G4249: signal is true;
	signal G4250: std_logic; attribute dont_touch of G4250: signal is true;
	signal G4251: std_logic; attribute dont_touch of G4251: signal is true;
	signal G4252: std_logic; attribute dont_touch of G4252: signal is true;
	signal G4253: std_logic; attribute dont_touch of G4253: signal is true;
	signal G4261: std_logic; attribute dont_touch of G4261: signal is true;
	signal G4262: std_logic; attribute dont_touch of G4262: signal is true;
	signal G4265: std_logic; attribute dont_touch of G4265: signal is true;
	signal G4266: std_logic; attribute dont_touch of G4266: signal is true;
	signal G4267: std_logic; attribute dont_touch of G4267: signal is true;
	signal G4270: std_logic; attribute dont_touch of G4270: signal is true;
	signal G4271: std_logic; attribute dont_touch of G4271: signal is true;
	signal G4272: std_logic; attribute dont_touch of G4272: signal is true;
	signal G4273: std_logic; attribute dont_touch of G4273: signal is true;
	signal G4276: std_logic; attribute dont_touch of G4276: signal is true;
	signal G4277: std_logic; attribute dont_touch of G4277: signal is true;
	signal G4280: std_logic; attribute dont_touch of G4280: signal is true;
	signal G4281: std_logic; attribute dont_touch of G4281: signal is true;
	signal G4284: std_logic; attribute dont_touch of G4284: signal is true;
	signal G4285: std_logic; attribute dont_touch of G4285: signal is true;
	signal G4286: std_logic; attribute dont_touch of G4286: signal is true;
	signal G4289: std_logic; attribute dont_touch of G4289: signal is true;
	signal G4292: std_logic; attribute dont_touch of G4292: signal is true;
	signal G4293: std_logic; attribute dont_touch of G4293: signal is true;
	signal G4296: std_logic; attribute dont_touch of G4296: signal is true;
	signal G4299: std_logic; attribute dont_touch of G4299: signal is true;
	signal G4300: std_logic; attribute dont_touch of G4300: signal is true;
	signal G4301: std_logic; attribute dont_touch of G4301: signal is true;
	signal G4302: std_logic; attribute dont_touch of G4302: signal is true;
	signal G4308: std_logic; attribute dont_touch of G4308: signal is true;
	signal G4309: std_logic; attribute dont_touch of G4309: signal is true;
	signal G4314: std_logic; attribute dont_touch of G4314: signal is true;
	signal G4319: std_logic; attribute dont_touch of G4319: signal is true;
	signal G4320: std_logic; attribute dont_touch of G4320: signal is true;
	signal G4322: std_logic; attribute dont_touch of G4322: signal is true;
	signal G4323: std_logic; attribute dont_touch of G4323: signal is true;
	signal G4328: std_logic; attribute dont_touch of G4328: signal is true;
	signal G4333: std_logic; attribute dont_touch of G4333: signal is true;
	signal G4334: std_logic; attribute dont_touch of G4334: signal is true;
	signal G4339: std_logic; attribute dont_touch of G4339: signal is true;
	signal G4340: std_logic; attribute dont_touch of G4340: signal is true;
	signal G4341: std_logic; attribute dont_touch of G4341: signal is true;
	signal G4342: std_logic; attribute dont_touch of G4342: signal is true;
	signal G4343: std_logic; attribute dont_touch of G4343: signal is true;
	signal G4344: std_logic; attribute dont_touch of G4344: signal is true;
	signal G4345: std_logic; attribute dont_touch of G4345: signal is true;
	signal G4346: std_logic; attribute dont_touch of G4346: signal is true;
	signal G4347: std_logic; attribute dont_touch of G4347: signal is true;
	signal G4348: std_logic; attribute dont_touch of G4348: signal is true;
	signal G4349: std_logic; attribute dont_touch of G4349: signal is true;
	signal G4350: std_logic; attribute dont_touch of G4350: signal is true;
	signal G4351: std_logic; attribute dont_touch of G4351: signal is true;
	signal G4352: std_logic; attribute dont_touch of G4352: signal is true;
	signal G4353: std_logic; attribute dont_touch of G4353: signal is true;
	signal G4354: std_logic; attribute dont_touch of G4354: signal is true;
	signal G4355: std_logic; attribute dont_touch of G4355: signal is true;
	signal G4356: std_logic; attribute dont_touch of G4356: signal is true;
	signal G4357: std_logic; attribute dont_touch of G4357: signal is true;
	signal G4358: std_logic; attribute dont_touch of G4358: signal is true;
	signal G4359: std_logic; attribute dont_touch of G4359: signal is true;
	signal G4360: std_logic; attribute dont_touch of G4360: signal is true;
	signal G4361: std_logic; attribute dont_touch of G4361: signal is true;
	signal G4362: std_logic; attribute dont_touch of G4362: signal is true;
	signal G4363: std_logic; attribute dont_touch of G4363: signal is true;
	signal G4364: std_logic; attribute dont_touch of G4364: signal is true;
	signal G4367: std_logic; attribute dont_touch of G4367: signal is true;
	signal G4368: std_logic; attribute dont_touch of G4368: signal is true;
	signal G4369: std_logic; attribute dont_touch of G4369: signal is true;
	signal G4370: std_logic; attribute dont_touch of G4370: signal is true;
	signal G4371: std_logic; attribute dont_touch of G4371: signal is true;
	signal G4372: std_logic; attribute dont_touch of G4372: signal is true;
	signal G4373: std_logic; attribute dont_touch of G4373: signal is true;
	signal G4374: std_logic; attribute dont_touch of G4374: signal is true;
	signal G4375: std_logic; attribute dont_touch of G4375: signal is true;
	signal G4376: std_logic; attribute dont_touch of G4376: signal is true;
	signal G4377: std_logic; attribute dont_touch of G4377: signal is true;
	signal G4378: std_logic; attribute dont_touch of G4378: signal is true;
	signal G4379: std_logic; attribute dont_touch of G4379: signal is true;
	signal G4380: std_logic; attribute dont_touch of G4380: signal is true;
	signal G4381: std_logic; attribute dont_touch of G4381: signal is true;
	signal G4382: std_logic; attribute dont_touch of G4382: signal is true;
	signal G4383: std_logic; attribute dont_touch of G4383: signal is true;
	signal G4384: std_logic; attribute dont_touch of G4384: signal is true;
	signal G4385: std_logic; attribute dont_touch of G4385: signal is true;
	signal G4386: std_logic; attribute dont_touch of G4386: signal is true;
	signal G4387: std_logic; attribute dont_touch of G4387: signal is true;
	signal G4388: std_logic; attribute dont_touch of G4388: signal is true;
	signal G4389: std_logic; attribute dont_touch of G4389: signal is true;
	signal G4390: std_logic; attribute dont_touch of G4390: signal is true;
	signal G4391: std_logic; attribute dont_touch of G4391: signal is true;
	signal G4392: std_logic; attribute dont_touch of G4392: signal is true;
	signal G4393: std_logic; attribute dont_touch of G4393: signal is true;
	signal G4394: std_logic; attribute dont_touch of G4394: signal is true;
	signal G4395: std_logic; attribute dont_touch of G4395: signal is true;
	signal G4396: std_logic; attribute dont_touch of G4396: signal is true;
	signal G4397: std_logic; attribute dont_touch of G4397: signal is true;
	signal G4398: std_logic; attribute dont_touch of G4398: signal is true;
	signal G4399: std_logic; attribute dont_touch of G4399: signal is true;
	signal G4400: std_logic; attribute dont_touch of G4400: signal is true;
	signal G4401: std_logic; attribute dont_touch of G4401: signal is true;
	signal G4402: std_logic; attribute dont_touch of G4402: signal is true;
	signal G4403: std_logic; attribute dont_touch of G4403: signal is true;
	signal G4404: std_logic; attribute dont_touch of G4404: signal is true;
	signal G4405: std_logic; attribute dont_touch of G4405: signal is true;
	signal G4406: std_logic; attribute dont_touch of G4406: signal is true;
	signal G4407: std_logic; attribute dont_touch of G4407: signal is true;
	signal G4410: std_logic; attribute dont_touch of G4410: signal is true;
	signal G4416: std_logic; attribute dont_touch of G4416: signal is true;
	signal G4423: std_logic; attribute dont_touch of G4423: signal is true;
	signal G4424: std_logic; attribute dont_touch of G4424: signal is true;
	signal G4425: std_logic; attribute dont_touch of G4425: signal is true;
	signal G4426: std_logic; attribute dont_touch of G4426: signal is true;
	signal G4427: std_logic; attribute dont_touch of G4427: signal is true;
	signal G4428: std_logic; attribute dont_touch of G4428: signal is true;
	signal G4429: std_logic; attribute dont_touch of G4429: signal is true;
	signal G4430: std_logic; attribute dont_touch of G4430: signal is true;
	signal G4431: std_logic; attribute dont_touch of G4431: signal is true;
	signal G4432: std_logic; attribute dont_touch of G4432: signal is true;
	signal G4433: std_logic; attribute dont_touch of G4433: signal is true;
	signal G4434: std_logic; attribute dont_touch of G4434: signal is true;
	signal G4435: std_logic; attribute dont_touch of G4435: signal is true;
	signal G4436: std_logic; attribute dont_touch of G4436: signal is true;
	signal G4437: std_logic; attribute dont_touch of G4437: signal is true;
	signal G4438: std_logic; attribute dont_touch of G4438: signal is true;
	signal G4439: std_logic; attribute dont_touch of G4439: signal is true;
	signal G4440: std_logic; attribute dont_touch of G4440: signal is true;
	signal G4441: std_logic; attribute dont_touch of G4441: signal is true;
	signal G4442: std_logic; attribute dont_touch of G4442: signal is true;
	signal G4443: std_logic; attribute dont_touch of G4443: signal is true;
	signal G4444: std_logic; attribute dont_touch of G4444: signal is true;
	signal G4445: std_logic; attribute dont_touch of G4445: signal is true;
	signal G4446: std_logic; attribute dont_touch of G4446: signal is true;
	signal G4447: std_logic; attribute dont_touch of G4447: signal is true;
	signal G4448: std_logic; attribute dont_touch of G4448: signal is true;
	signal G4449: std_logic; attribute dont_touch of G4449: signal is true;
	signal G4450: std_logic; attribute dont_touch of G4450: signal is true;
	signal G4451: std_logic; attribute dont_touch of G4451: signal is true;
	signal G4452: std_logic; attribute dont_touch of G4452: signal is true;
	signal G4453: std_logic; attribute dont_touch of G4453: signal is true;
	signal G4454: std_logic; attribute dont_touch of G4454: signal is true;
	signal G4455: std_logic; attribute dont_touch of G4455: signal is true;
	signal G4456: std_logic; attribute dont_touch of G4456: signal is true;
	signal G4457: std_logic; attribute dont_touch of G4457: signal is true;
	signal G4458: std_logic; attribute dont_touch of G4458: signal is true;
	signal G4459: std_logic; attribute dont_touch of G4459: signal is true;
	signal G4460: std_logic; attribute dont_touch of G4460: signal is true;
	signal G4461: std_logic; attribute dont_touch of G4461: signal is true;
	signal G4462: std_logic; attribute dont_touch of G4462: signal is true;
	signal G4463: std_logic; attribute dont_touch of G4463: signal is true;
	signal G4464: std_logic; attribute dont_touch of G4464: signal is true;
	signal G4465: std_logic; attribute dont_touch of G4465: signal is true;
	signal G4468: std_logic; attribute dont_touch of G4468: signal is true;
	signal G4471: std_logic; attribute dont_touch of G4471: signal is true;
	signal G4472: std_logic; attribute dont_touch of G4472: signal is true;
	signal G4473: std_logic; attribute dont_touch of G4473: signal is true;
	signal G4485: std_logic; attribute dont_touch of G4485: signal is true;
	signal G4486: std_logic; attribute dont_touch of G4486: signal is true;
	signal G4487: std_logic; attribute dont_touch of G4487: signal is true;
	signal G4488: std_logic; attribute dont_touch of G4488: signal is true;
	signal G4489: std_logic; attribute dont_touch of G4489: signal is true;
	signal G4490: std_logic; attribute dont_touch of G4490: signal is true;
	signal G4491: std_logic; attribute dont_touch of G4491: signal is true;
	signal G4492: std_logic; attribute dont_touch of G4492: signal is true;
	signal G4493: std_logic; attribute dont_touch of G4493: signal is true;
	signal G4494: std_logic; attribute dont_touch of G4494: signal is true;
	signal G4495: std_logic; attribute dont_touch of G4495: signal is true;
	signal G4496: std_logic; attribute dont_touch of G4496: signal is true;
	signal G4497: std_logic; attribute dont_touch of G4497: signal is true;
	signal G4498: std_logic; attribute dont_touch of G4498: signal is true;
	signal G4499: std_logic; attribute dont_touch of G4499: signal is true;
	signal G4500: std_logic; attribute dont_touch of G4500: signal is true;
	signal G4501: std_logic; attribute dont_touch of G4501: signal is true;
	signal G4502: std_logic; attribute dont_touch of G4502: signal is true;
	signal G4503: std_logic; attribute dont_touch of G4503: signal is true;
	signal G4504: std_logic; attribute dont_touch of G4504: signal is true;
	signal G4507: std_logic; attribute dont_touch of G4507: signal is true;
	signal G4508: std_logic; attribute dont_touch of G4508: signal is true;
	signal G4509: std_logic; attribute dont_touch of G4509: signal is true;
	signal G4510: std_logic; attribute dont_touch of G4510: signal is true;
	signal G4511: std_logic; attribute dont_touch of G4511: signal is true;
	signal G4512: std_logic; attribute dont_touch of G4512: signal is true;
	signal G4513: std_logic; attribute dont_touch of G4513: signal is true;
	signal G4514: std_logic; attribute dont_touch of G4514: signal is true;
	signal G4515: std_logic; attribute dont_touch of G4515: signal is true;
	signal G4516: std_logic; attribute dont_touch of G4516: signal is true;
	signal G4517: std_logic; attribute dont_touch of G4517: signal is true;
	signal G4518: std_logic; attribute dont_touch of G4518: signal is true;
	signal G4519: std_logic; attribute dont_touch of G4519: signal is true;
	signal G4520: std_logic; attribute dont_touch of G4520: signal is true;
	signal G4521: std_logic; attribute dont_touch of G4521: signal is true;
	signal G4522: std_logic; attribute dont_touch of G4522: signal is true;
	signal G4523: std_logic; attribute dont_touch of G4523: signal is true;
	signal G4524: std_logic; attribute dont_touch of G4524: signal is true;
	signal G4525: std_logic; attribute dont_touch of G4525: signal is true;
	signal G4526: std_logic; attribute dont_touch of G4526: signal is true;
	signal G4527: std_logic; attribute dont_touch of G4527: signal is true;
	signal G4528: std_logic; attribute dont_touch of G4528: signal is true;
	signal G4529: std_logic; attribute dont_touch of G4529: signal is true;
	signal G4530: std_logic; attribute dont_touch of G4530: signal is true;
	signal G4531: std_logic; attribute dont_touch of G4531: signal is true;
	signal G4532: std_logic; attribute dont_touch of G4532: signal is true;
	signal G4533: std_logic; attribute dont_touch of G4533: signal is true;
	signal G4534: std_logic; attribute dont_touch of G4534: signal is true;
	signal G4535: std_logic; attribute dont_touch of G4535: signal is true;
	signal G4536: std_logic; attribute dont_touch of G4536: signal is true;
	signal G4537: std_logic; attribute dont_touch of G4537: signal is true;
	signal G4541: std_logic; attribute dont_touch of G4541: signal is true;
	signal G4544: std_logic; attribute dont_touch of G4544: signal is true;
	signal G4545: std_logic; attribute dont_touch of G4545: signal is true;
	signal G4549: std_logic; attribute dont_touch of G4549: signal is true;
	signal G4550: std_logic; attribute dont_touch of G4550: signal is true;
	signal G4559: std_logic; attribute dont_touch of G4559: signal is true;
	signal G4560: std_logic; attribute dont_touch of G4560: signal is true;
	signal G4561: std_logic; attribute dont_touch of G4561: signal is true;
	signal G4562: std_logic; attribute dont_touch of G4562: signal is true;
	signal G4563: std_logic; attribute dont_touch of G4563: signal is true;
	signal G4564: std_logic; attribute dont_touch of G4564: signal is true;
	signal G4565: std_logic; attribute dont_touch of G4565: signal is true;
	signal G4566: std_logic; attribute dont_touch of G4566: signal is true;
	signal G4567: std_logic; attribute dont_touch of G4567: signal is true;
	signal G4568: std_logic; attribute dont_touch of G4568: signal is true;
	signal G4569: std_logic; attribute dont_touch of G4569: signal is true;
	signal G4577: std_logic; attribute dont_touch of G4577: signal is true;
	signal G4578: std_logic; attribute dont_touch of G4578: signal is true;
	signal G4579: std_logic; attribute dont_touch of G4579: signal is true;
	signal G4580: std_logic; attribute dont_touch of G4580: signal is true;
	signal G4581: std_logic; attribute dont_touch of G4581: signal is true;
	signal G4582: std_logic; attribute dont_touch of G4582: signal is true;
	signal G4583: std_logic; attribute dont_touch of G4583: signal is true;
	signal G4584: std_logic; attribute dont_touch of G4584: signal is true;
	signal G4585: std_logic; attribute dont_touch of G4585: signal is true;
	signal G4586: std_logic; attribute dont_touch of G4586: signal is true;
	signal G4587: std_logic; attribute dont_touch of G4587: signal is true;
	signal G4588: std_logic; attribute dont_touch of G4588: signal is true;
	signal G4589: std_logic; attribute dont_touch of G4589: signal is true;
	signal G4590: std_logic; attribute dont_touch of G4590: signal is true;
	signal G4591: std_logic; attribute dont_touch of G4591: signal is true;
	signal G4592: std_logic; attribute dont_touch of G4592: signal is true;
	signal G4593: std_logic; attribute dont_touch of G4593: signal is true;
	signal G4596: std_logic; attribute dont_touch of G4596: signal is true;
	signal G4597: std_logic; attribute dont_touch of G4597: signal is true;
	signal G4598: std_logic; attribute dont_touch of G4598: signal is true;
	signal G4599: std_logic; attribute dont_touch of G4599: signal is true;
	signal G4600: std_logic; attribute dont_touch of G4600: signal is true;
	signal G4601: std_logic; attribute dont_touch of G4601: signal is true;
	signal G4602: std_logic; attribute dont_touch of G4602: signal is true;
	signal G4603: std_logic; attribute dont_touch of G4603: signal is true;
	signal G4606: std_logic; attribute dont_touch of G4606: signal is true;
	signal G4607: std_logic; attribute dont_touch of G4607: signal is true;
	signal G4608: std_logic; attribute dont_touch of G4608: signal is true;
	signal G4609: std_logic; attribute dont_touch of G4609: signal is true;
	signal G4610: std_logic; attribute dont_touch of G4610: signal is true;
	signal G4611: std_logic; attribute dont_touch of G4611: signal is true;
	signal G4612: std_logic; attribute dont_touch of G4612: signal is true;
	signal G4613: std_logic; attribute dont_touch of G4613: signal is true;
	signal G4614: std_logic; attribute dont_touch of G4614: signal is true;
	signal G4615: std_logic; attribute dont_touch of G4615: signal is true;
	signal G4616: std_logic; attribute dont_touch of G4616: signal is true;
	signal G4617: std_logic; attribute dont_touch of G4617: signal is true;
	signal G4618: std_logic; attribute dont_touch of G4618: signal is true;
	signal G4619: std_logic; attribute dont_touch of G4619: signal is true;
	signal G4620: std_logic; attribute dont_touch of G4620: signal is true;
	signal G4621: std_logic; attribute dont_touch of G4621: signal is true;
	signal G4622: std_logic; attribute dont_touch of G4622: signal is true;
	signal G4623: std_logic; attribute dont_touch of G4623: signal is true;
	signal G4624: std_logic; attribute dont_touch of G4624: signal is true;
	signal G4625: std_logic; attribute dont_touch of G4625: signal is true;
	signal G4626: std_logic; attribute dont_touch of G4626: signal is true;
	signal G4627: std_logic; attribute dont_touch of G4627: signal is true;
	signal G4628: std_logic; attribute dont_touch of G4628: signal is true;
	signal G4629: std_logic; attribute dont_touch of G4629: signal is true;
	signal G4630: std_logic; attribute dont_touch of G4630: signal is true;
	signal G4631: std_logic; attribute dont_touch of G4631: signal is true;
	signal G4632: std_logic; attribute dont_touch of G4632: signal is true;
	signal G4633: std_logic; attribute dont_touch of G4633: signal is true;
	signal G4634: std_logic; attribute dont_touch of G4634: signal is true;
	signal G4635: std_logic; attribute dont_touch of G4635: signal is true;
	signal G4636: std_logic; attribute dont_touch of G4636: signal is true;
	signal G4637: std_logic; attribute dont_touch of G4637: signal is true;
	signal G4638: std_logic; attribute dont_touch of G4638: signal is true;
	signal G4639: std_logic; attribute dont_touch of G4639: signal is true;
	signal G4640: std_logic; attribute dont_touch of G4640: signal is true;
	signal G4641: std_logic; attribute dont_touch of G4641: signal is true;
	signal G4642: std_logic; attribute dont_touch of G4642: signal is true;
	signal G4643: std_logic; attribute dont_touch of G4643: signal is true;
	signal G4644: std_logic; attribute dont_touch of G4644: signal is true;
	signal G4645: std_logic; attribute dont_touch of G4645: signal is true;
	signal G4646: std_logic; attribute dont_touch of G4646: signal is true;
	signal G4647: std_logic; attribute dont_touch of G4647: signal is true;
	signal G4648: std_logic; attribute dont_touch of G4648: signal is true;
	signal G4651: std_logic; attribute dont_touch of G4651: signal is true;
	signal G4652: std_logic; attribute dont_touch of G4652: signal is true;
	signal G4653: std_logic; attribute dont_touch of G4653: signal is true;
	signal G4654: std_logic; attribute dont_touch of G4654: signal is true;
	signal G4655: std_logic; attribute dont_touch of G4655: signal is true;
	signal G4656: std_logic; attribute dont_touch of G4656: signal is true;
	signal G4657: std_logic; attribute dont_touch of G4657: signal is true;
	signal G4658: std_logic; attribute dont_touch of G4658: signal is true;
	signal G4659: std_logic; attribute dont_touch of G4659: signal is true;
	signal G4660: std_logic; attribute dont_touch of G4660: signal is true;
	signal G4661: std_logic; attribute dont_touch of G4661: signal is true;
	signal G4662: std_logic; attribute dont_touch of G4662: signal is true;
	signal G4666: std_logic; attribute dont_touch of G4666: signal is true;
	signal G4667: std_logic; attribute dont_touch of G4667: signal is true;
	signal G4668: std_logic; attribute dont_touch of G4668: signal is true;
	signal G4669: std_logic; attribute dont_touch of G4669: signal is true;
	signal G4670: std_logic; attribute dont_touch of G4670: signal is true;
	signal G4671: std_logic; attribute dont_touch of G4671: signal is true;
	signal G4672: std_logic; attribute dont_touch of G4672: signal is true;
	signal G4673: std_logic; attribute dont_touch of G4673: signal is true;
	signal G4674: std_logic; attribute dont_touch of G4674: signal is true;
	signal G4677: std_logic; attribute dont_touch of G4677: signal is true;
	signal G4678: std_logic; attribute dont_touch of G4678: signal is true;
	signal G4679: std_logic; attribute dont_touch of G4679: signal is true;
	signal G4680: std_logic; attribute dont_touch of G4680: signal is true;
	signal G4683: std_logic; attribute dont_touch of G4683: signal is true;
	signal G4684: std_logic; attribute dont_touch of G4684: signal is true;
	signal G4685: std_logic; attribute dont_touch of G4685: signal is true;
	signal G4686: std_logic; attribute dont_touch of G4686: signal is true;
	signal G4687: std_logic; attribute dont_touch of G4687: signal is true;
	signal G4688: std_logic; attribute dont_touch of G4688: signal is true;
	signal G4691: std_logic; attribute dont_touch of G4691: signal is true;
	signal G4692: std_logic; attribute dont_touch of G4692: signal is true;
	signal G4693: std_logic; attribute dont_touch of G4693: signal is true;
	signal G4694: std_logic; attribute dont_touch of G4694: signal is true;
	signal G4697: std_logic; attribute dont_touch of G4697: signal is true;
	signal G4698: std_logic; attribute dont_touch of G4698: signal is true;
	signal G4699: std_logic; attribute dont_touch of G4699: signal is true;
	signal G4700: std_logic; attribute dont_touch of G4700: signal is true;
	signal G4701: std_logic; attribute dont_touch of G4701: signal is true;
	signal G4702: std_logic; attribute dont_touch of G4702: signal is true;
	signal G4703: std_logic; attribute dont_touch of G4703: signal is true;
	signal G4704: std_logic; attribute dont_touch of G4704: signal is true;
	signal G4705: std_logic; attribute dont_touch of G4705: signal is true;
	signal G4706: std_logic; attribute dont_touch of G4706: signal is true;
	signal G4707: std_logic; attribute dont_touch of G4707: signal is true;
	signal G4708: std_logic; attribute dont_touch of G4708: signal is true;
	signal G4711: std_logic; attribute dont_touch of G4711: signal is true;
	signal G4712: std_logic; attribute dont_touch of G4712: signal is true;
	signal G4713: std_logic; attribute dont_touch of G4713: signal is true;
	signal G4714: std_logic; attribute dont_touch of G4714: signal is true;
	signal G4715: std_logic; attribute dont_touch of G4715: signal is true;
	signal G4716: std_logic; attribute dont_touch of G4716: signal is true;
	signal G4717: std_logic; attribute dont_touch of G4717: signal is true;
	signal G4718: std_logic; attribute dont_touch of G4718: signal is true;
	signal G4719: std_logic; attribute dont_touch of G4719: signal is true;
	signal G4720: std_logic; attribute dont_touch of G4720: signal is true;
	signal G4721: std_logic; attribute dont_touch of G4721: signal is true;
	signal G4722: std_logic; attribute dont_touch of G4722: signal is true;
	signal G4723: std_logic; attribute dont_touch of G4723: signal is true;
	signal G4726: std_logic; attribute dont_touch of G4726: signal is true;
	signal G4727: std_logic; attribute dont_touch of G4727: signal is true;
	signal G4730: std_logic; attribute dont_touch of G4730: signal is true;
	signal G4731: std_logic; attribute dont_touch of G4731: signal is true;
	signal G4732: std_logic; attribute dont_touch of G4732: signal is true;
	signal G4735: std_logic; attribute dont_touch of G4735: signal is true;
	signal G4736: std_logic; attribute dont_touch of G4736: signal is true;
	signal G4739: std_logic; attribute dont_touch of G4739: signal is true;
	signal G4740: std_logic; attribute dont_touch of G4740: signal is true;
	signal G4741: std_logic; attribute dont_touch of G4741: signal is true;
	signal G4744: std_logic; attribute dont_touch of G4744: signal is true;
	signal G4745: std_logic; attribute dont_touch of G4745: signal is true;
	signal G4752: std_logic; attribute dont_touch of G4752: signal is true;
	signal G4753: std_logic; attribute dont_touch of G4753: signal is true;
	signal G4756: std_logic; attribute dont_touch of G4756: signal is true;
	signal G4757: std_logic; attribute dont_touch of G4757: signal is true;
	signal G4758: std_logic; attribute dont_touch of G4758: signal is true;
	signal G4759: std_logic; attribute dont_touch of G4759: signal is true;
	signal G4760: std_logic; attribute dont_touch of G4760: signal is true;
	signal G4761: std_logic; attribute dont_touch of G4761: signal is true;
	signal G4762: std_logic; attribute dont_touch of G4762: signal is true;
	signal G4763: std_logic; attribute dont_touch of G4763: signal is true;
	signal G4764: std_logic; attribute dont_touch of G4764: signal is true;
	signal G4765: std_logic; attribute dont_touch of G4765: signal is true;
	signal G4766: std_logic; attribute dont_touch of G4766: signal is true;
	signal G4767: std_logic; attribute dont_touch of G4767: signal is true;
	signal G4768: std_logic; attribute dont_touch of G4768: signal is true;
	signal G4769: std_logic; attribute dont_touch of G4769: signal is true;
	signal G4770: std_logic; attribute dont_touch of G4770: signal is true;
	signal G4771: std_logic; attribute dont_touch of G4771: signal is true;
	signal G4772: std_logic; attribute dont_touch of G4772: signal is true;
	signal G4773: std_logic; attribute dont_touch of G4773: signal is true;
	signal G4774: std_logic; attribute dont_touch of G4774: signal is true;
	signal G4775: std_logic; attribute dont_touch of G4775: signal is true;
	signal G4776: std_logic; attribute dont_touch of G4776: signal is true;
	signal G4777: std_logic; attribute dont_touch of G4777: signal is true;
	signal G4778: std_logic; attribute dont_touch of G4778: signal is true;
	signal G4779: std_logic; attribute dont_touch of G4779: signal is true;
	signal G4780: std_logic; attribute dont_touch of G4780: signal is true;
	signal G4781: std_logic; attribute dont_touch of G4781: signal is true;
	signal G4782: std_logic; attribute dont_touch of G4782: signal is true;
	signal G4783: std_logic; attribute dont_touch of G4783: signal is true;
	signal G4784: std_logic; attribute dont_touch of G4784: signal is true;
	signal G4785: std_logic; attribute dont_touch of G4785: signal is true;
	signal G4786: std_logic; attribute dont_touch of G4786: signal is true;
	signal G4787: std_logic; attribute dont_touch of G4787: signal is true;
	signal G4788: std_logic; attribute dont_touch of G4788: signal is true;
	signal G4789: std_logic; attribute dont_touch of G4789: signal is true;
	signal G4790: std_logic; attribute dont_touch of G4790: signal is true;
	signal G4791: std_logic; attribute dont_touch of G4791: signal is true;
	signal G4792: std_logic; attribute dont_touch of G4792: signal is true;
	signal G4793: std_logic; attribute dont_touch of G4793: signal is true;
	signal G4794: std_logic; attribute dont_touch of G4794: signal is true;
	signal G4797: std_logic; attribute dont_touch of G4797: signal is true;
	signal G4798: std_logic; attribute dont_touch of G4798: signal is true;
	signal G4799: std_logic; attribute dont_touch of G4799: signal is true;
	signal G4800: std_logic; attribute dont_touch of G4800: signal is true;
	signal G4801: std_logic; attribute dont_touch of G4801: signal is true;
	signal G4802: std_logic; attribute dont_touch of G4802: signal is true;
	signal G4803: std_logic; attribute dont_touch of G4803: signal is true;
	signal G4804: std_logic; attribute dont_touch of G4804: signal is true;
	signal G4805: std_logic; attribute dont_touch of G4805: signal is true;
	signal G4806: std_logic; attribute dont_touch of G4806: signal is true;
	signal G4807: std_logic; attribute dont_touch of G4807: signal is true;
	signal G4808: std_logic; attribute dont_touch of G4808: signal is true;
	signal G4810: std_logic; attribute dont_touch of G4810: signal is true;
	signal G4811: std_logic; attribute dont_touch of G4811: signal is true;
	signal G4812: std_logic; attribute dont_touch of G4812: signal is true;
	signal G4813: std_logic; attribute dont_touch of G4813: signal is true;
	signal G4814: std_logic; attribute dont_touch of G4814: signal is true;
	signal G4815: std_logic; attribute dont_touch of G4815: signal is true;
	signal G4816: std_logic; attribute dont_touch of G4816: signal is true;
	signal G4819: std_logic; attribute dont_touch of G4819: signal is true;
	signal G4822: std_logic; attribute dont_touch of G4822: signal is true;
	signal G4823: std_logic; attribute dont_touch of G4823: signal is true;
	signal G4824: std_logic; attribute dont_touch of G4824: signal is true;
	signal G4825: std_logic; attribute dont_touch of G4825: signal is true;
	signal G4826: std_logic; attribute dont_touch of G4826: signal is true;
	signal G4827: std_logic; attribute dont_touch of G4827: signal is true;
	signal G4828: std_logic; attribute dont_touch of G4828: signal is true;
	signal G4829: std_logic; attribute dont_touch of G4829: signal is true;
	signal G4830: std_logic; attribute dont_touch of G4830: signal is true;
	signal G4831: std_logic; attribute dont_touch of G4831: signal is true;
	signal G4832: std_logic; attribute dont_touch of G4832: signal is true;
	signal G4833: std_logic; attribute dont_touch of G4833: signal is true;
	signal G4834: std_logic; attribute dont_touch of G4834: signal is true;
	signal G4835: std_logic; attribute dont_touch of G4835: signal is true;
	signal G4836: std_logic; attribute dont_touch of G4836: signal is true;
	signal G4837: std_logic; attribute dont_touch of G4837: signal is true;
	signal G4838: std_logic; attribute dont_touch of G4838: signal is true;
	signal G4839: std_logic; attribute dont_touch of G4839: signal is true;
	signal G4840: std_logic; attribute dont_touch of G4840: signal is true;
	signal G4841: std_logic; attribute dont_touch of G4841: signal is true;
	signal G4842: std_logic; attribute dont_touch of G4842: signal is true;
	signal G4843: std_logic; attribute dont_touch of G4843: signal is true;
	signal G4844: std_logic; attribute dont_touch of G4844: signal is true;
	signal G4845: std_logic; attribute dont_touch of G4845: signal is true;
	signal G4846: std_logic; attribute dont_touch of G4846: signal is true;
	signal G4847: std_logic; attribute dont_touch of G4847: signal is true;
	signal G4848: std_logic; attribute dont_touch of G4848: signal is true;
	signal G4849: std_logic; attribute dont_touch of G4849: signal is true;
	signal G4850: std_logic; attribute dont_touch of G4850: signal is true;
	signal G4851: std_logic; attribute dont_touch of G4851: signal is true;
	signal G4852: std_logic; attribute dont_touch of G4852: signal is true;
	signal G4853: std_logic; attribute dont_touch of G4853: signal is true;
	signal G4854: std_logic; attribute dont_touch of G4854: signal is true;
	signal G4855: std_logic; attribute dont_touch of G4855: signal is true;
	signal G4856: std_logic; attribute dont_touch of G4856: signal is true;
	signal G4857: std_logic; attribute dont_touch of G4857: signal is true;
	signal G4858: std_logic; attribute dont_touch of G4858: signal is true;
	signal G4859: std_logic; attribute dont_touch of G4859: signal is true;
	signal G4860: std_logic; attribute dont_touch of G4860: signal is true;
	signal G4861: std_logic; attribute dont_touch of G4861: signal is true;
	signal G4862: std_logic; attribute dont_touch of G4862: signal is true;
	signal G4863: std_logic; attribute dont_touch of G4863: signal is true;
	signal G4864: std_logic; attribute dont_touch of G4864: signal is true;
	signal G4865: std_logic; attribute dont_touch of G4865: signal is true;
	signal G4866: std_logic; attribute dont_touch of G4866: signal is true;
	signal G4867: std_logic; attribute dont_touch of G4867: signal is true;
	signal G4868: std_logic; attribute dont_touch of G4868: signal is true;
	signal G4869: std_logic; attribute dont_touch of G4869: signal is true;
	signal G4870: std_logic; attribute dont_touch of G4870: signal is true;
	signal G4871: std_logic; attribute dont_touch of G4871: signal is true;
	signal G4872: std_logic; attribute dont_touch of G4872: signal is true;
	signal G4873: std_logic; attribute dont_touch of G4873: signal is true;
	signal G4874: std_logic; attribute dont_touch of G4874: signal is true;
	signal G4877: std_logic; attribute dont_touch of G4877: signal is true;
	signal G4894: std_logic; attribute dont_touch of G4894: signal is true;
	signal G4900: std_logic; attribute dont_touch of G4900: signal is true;
	signal G4903: std_logic; attribute dont_touch of G4903: signal is true;
	signal G4904: std_logic; attribute dont_touch of G4904: signal is true;
	signal G4910: std_logic; attribute dont_touch of G4910: signal is true;
	signal G4911: std_logic; attribute dont_touch of G4911: signal is true;
	signal G4914: std_logic; attribute dont_touch of G4914: signal is true;
	signal G4915: std_logic; attribute dont_touch of G4915: signal is true;
	signal G4928: std_logic; attribute dont_touch of G4928: signal is true;
	signal G4929: std_logic; attribute dont_touch of G4929: signal is true;
	signal G4932: std_logic; attribute dont_touch of G4932: signal is true;
	signal G4933: std_logic; attribute dont_touch of G4933: signal is true;
	signal G4936: std_logic; attribute dont_touch of G4936: signal is true;
	signal G4937: std_logic; attribute dont_touch of G4937: signal is true;
	signal G4938: std_logic; attribute dont_touch of G4938: signal is true;
	signal G4941: std_logic; attribute dont_touch of G4941: signal is true;
	signal G4942: std_logic; attribute dont_touch of G4942: signal is true;
	signal G4943: std_logic; attribute dont_touch of G4943: signal is true;
	signal G4946: std_logic; attribute dont_touch of G4946: signal is true;
	signal G4947: std_logic; attribute dont_touch of G4947: signal is true;
	signal G4948: std_logic; attribute dont_touch of G4948: signal is true;
	signal G4949: std_logic; attribute dont_touch of G4949: signal is true;
	signal G4950: std_logic; attribute dont_touch of G4950: signal is true;
	signal G4967: std_logic; attribute dont_touch of G4967: signal is true;
	signal G4980: std_logic; attribute dont_touch of G4980: signal is true;
	signal G4993: std_logic; attribute dont_touch of G4993: signal is true;
	signal G5010: std_logic; attribute dont_touch of G5010: signal is true;
	signal G5011: std_logic; attribute dont_touch of G5011: signal is true;
	signal G5012: std_logic; attribute dont_touch of G5012: signal is true;
	signal G5013: std_logic; attribute dont_touch of G5013: signal is true;
	signal G5014: std_logic; attribute dont_touch of G5014: signal is true;
	signal G5015: std_logic; attribute dont_touch of G5015: signal is true;
	signal G5016: std_logic; attribute dont_touch of G5016: signal is true;
	signal G5017: std_logic; attribute dont_touch of G5017: signal is true;
	signal G5018: std_logic; attribute dont_touch of G5018: signal is true;
	signal G5019: std_logic; attribute dont_touch of G5019: signal is true;
	signal G5022: std_logic; attribute dont_touch of G5022: signal is true;
	signal G5023: std_logic; attribute dont_touch of G5023: signal is true;
	signal G5024: std_logic; attribute dont_touch of G5024: signal is true;
	signal G5025: std_logic; attribute dont_touch of G5025: signal is true;
	signal G5042: std_logic; attribute dont_touch of G5042: signal is true;
	signal G5043: std_logic; attribute dont_touch of G5043: signal is true;
	signal G5044: std_logic; attribute dont_touch of G5044: signal is true;
	signal G5045: std_logic; attribute dont_touch of G5045: signal is true;
	signal G5046: std_logic; attribute dont_touch of G5046: signal is true;
	signal G5047: std_logic; attribute dont_touch of G5047: signal is true;
	signal G5048: std_logic; attribute dont_touch of G5048: signal is true;
	signal G5049: std_logic; attribute dont_touch of G5049: signal is true;
	signal G5050: std_logic; attribute dont_touch of G5050: signal is true;
	signal G5051: std_logic; attribute dont_touch of G5051: signal is true;
	signal G5052: std_logic; attribute dont_touch of G5052: signal is true;
	signal G5053: std_logic; attribute dont_touch of G5053: signal is true;
	signal G5054: std_logic; attribute dont_touch of G5054: signal is true;
	signal G5059: std_logic; attribute dont_touch of G5059: signal is true;
	signal G5060: std_logic; attribute dont_touch of G5060: signal is true;
	signal G5061: std_logic; attribute dont_touch of G5061: signal is true;
	signal G5062: std_logic; attribute dont_touch of G5062: signal is true;
	signal G5063: std_logic; attribute dont_touch of G5063: signal is true;
	signal G5064: std_logic; attribute dont_touch of G5064: signal is true;
	signal G5065: std_logic; attribute dont_touch of G5065: signal is true;
	signal G5066: std_logic; attribute dont_touch of G5066: signal is true;
	signal G5067: std_logic; attribute dont_touch of G5067: signal is true;
	signal G5068: std_logic; attribute dont_touch of G5068: signal is true;
	signal G5069: std_logic; attribute dont_touch of G5069: signal is true;
	signal G5074: std_logic; attribute dont_touch of G5074: signal is true;
	signal G5077: std_logic; attribute dont_touch of G5077: signal is true;
	signal G5082: std_logic; attribute dont_touch of G5082: signal is true;
	signal G5083: std_logic; attribute dont_touch of G5083: signal is true;
	signal G5084: std_logic; attribute dont_touch of G5084: signal is true;
	signal G5085: std_logic; attribute dont_touch of G5085: signal is true;
	signal G5086: std_logic; attribute dont_touch of G5086: signal is true;
	signal G5087: std_logic; attribute dont_touch of G5087: signal is true;
	signal G5088: std_logic; attribute dont_touch of G5088: signal is true;
	signal G5089: std_logic; attribute dont_touch of G5089: signal is true;
	signal G5090: std_logic; attribute dont_touch of G5090: signal is true;
	signal G5091: std_logic; attribute dont_touch of G5091: signal is true;
	signal G5092: std_logic; attribute dont_touch of G5092: signal is true;
	signal G5093: std_logic; attribute dont_touch of G5093: signal is true;
	signal G5094: std_logic; attribute dont_touch of G5094: signal is true;
	signal G5095: std_logic; attribute dont_touch of G5095: signal is true;
	signal G5096: std_logic; attribute dont_touch of G5096: signal is true;
	signal G5097: std_logic; attribute dont_touch of G5097: signal is true;
	signal G5098: std_logic; attribute dont_touch of G5098: signal is true;
	signal G5099: std_logic; attribute dont_touch of G5099: signal is true;
	signal G5110: std_logic; attribute dont_touch of G5110: signal is true;
	signal G5111: std_logic; attribute dont_touch of G5111: signal is true;
	signal G5112: std_logic; attribute dont_touch of G5112: signal is true;
	signal G5113: std_logic; attribute dont_touch of G5113: signal is true;
	signal G5114: std_logic; attribute dont_touch of G5114: signal is true;
	signal G5115: std_logic; attribute dont_touch of G5115: signal is true;
	signal G5116: std_logic; attribute dont_touch of G5116: signal is true;
	signal G5117: std_logic; attribute dont_touch of G5117: signal is true;
	signal G5118: std_logic; attribute dont_touch of G5118: signal is true;
	signal G5119: std_logic; attribute dont_touch of G5119: signal is true;
	signal G5120: std_logic; attribute dont_touch of G5120: signal is true;
	signal G5121: std_logic; attribute dont_touch of G5121: signal is true;
	signal G5122: std_logic; attribute dont_touch of G5122: signal is true;
	signal G5123: std_logic; attribute dont_touch of G5123: signal is true;
	signal G5124: std_logic; attribute dont_touch of G5124: signal is true;
	signal G5135: std_logic; attribute dont_touch of G5135: signal is true;
	signal G5136: std_logic; attribute dont_touch of G5136: signal is true;
	signal G5138: std_logic; attribute dont_touch of G5138: signal is true;
	signal G5139: std_logic; attribute dont_touch of G5139: signal is true;
	signal G5140: std_logic; attribute dont_touch of G5140: signal is true;
	signal G5141: std_logic; attribute dont_touch of G5141: signal is true;
	signal G5142: std_logic; attribute dont_touch of G5142: signal is true;
	signal G5143: std_logic; attribute dont_touch of G5143: signal is true;
	signal G5144: std_logic; attribute dont_touch of G5144: signal is true;
	signal G5145: std_logic; attribute dont_touch of G5145: signal is true;
	signal G5146: std_logic; attribute dont_touch of G5146: signal is true;
	signal G5147: std_logic; attribute dont_touch of G5147: signal is true;
	signal G5148: std_logic; attribute dont_touch of G5148: signal is true;
	signal G5149: std_logic; attribute dont_touch of G5149: signal is true;
	signal G5150: std_logic; attribute dont_touch of G5150: signal is true;
	signal G5151: std_logic; attribute dont_touch of G5151: signal is true;
	signal G5152: std_logic; attribute dont_touch of G5152: signal is true;
	signal G5153: std_logic; attribute dont_touch of G5153: signal is true;
	signal G5154: std_logic; attribute dont_touch of G5154: signal is true;
	signal G5155: std_logic; attribute dont_touch of G5155: signal is true;
	signal G5156: std_logic; attribute dont_touch of G5156: signal is true;
	signal G5157: std_logic; attribute dont_touch of G5157: signal is true;
	signal G5158: std_logic; attribute dont_touch of G5158: signal is true;
	signal G5159: std_logic; attribute dont_touch of G5159: signal is true;
	signal G5160: std_logic; attribute dont_touch of G5160: signal is true;
	signal G5161: std_logic; attribute dont_touch of G5161: signal is true;
	signal G5162: std_logic; attribute dont_touch of G5162: signal is true;
	signal G5163: std_logic; attribute dont_touch of G5163: signal is true;
	signal G5164: std_logic; attribute dont_touch of G5164: signal is true;
	signal G5165: std_logic; attribute dont_touch of G5165: signal is true;
	signal G5166: std_logic; attribute dont_touch of G5166: signal is true;
	signal G5167: std_logic; attribute dont_touch of G5167: signal is true;
	signal G5168: std_logic; attribute dont_touch of G5168: signal is true;
	signal G5169: std_logic; attribute dont_touch of G5169: signal is true;
	signal G5170: std_logic; attribute dont_touch of G5170: signal is true;
	signal G5171: std_logic; attribute dont_touch of G5171: signal is true;
	signal G5172: std_logic; attribute dont_touch of G5172: signal is true;
	signal G5173: std_logic; attribute dont_touch of G5173: signal is true;
	signal G5174: std_logic; attribute dont_touch of G5174: signal is true;
	signal G5175: std_logic; attribute dont_touch of G5175: signal is true;
	signal G5176: std_logic; attribute dont_touch of G5176: signal is true;
	signal G5177: std_logic; attribute dont_touch of G5177: signal is true;
	signal G5178: std_logic; attribute dont_touch of G5178: signal is true;
	signal G5179: std_logic; attribute dont_touch of G5179: signal is true;
	signal G5180: std_logic; attribute dont_touch of G5180: signal is true;
	signal G5181: std_logic; attribute dont_touch of G5181: signal is true;
	signal G5182: std_logic; attribute dont_touch of G5182: signal is true;
	signal G5183: std_logic; attribute dont_touch of G5183: signal is true;
	signal G5184: std_logic; attribute dont_touch of G5184: signal is true;
	signal G5185: std_logic; attribute dont_touch of G5185: signal is true;
	signal G5186: std_logic; attribute dont_touch of G5186: signal is true;
	signal G5187: std_logic; attribute dont_touch of G5187: signal is true;
	signal G5188: std_logic; attribute dont_touch of G5188: signal is true;
	signal G5189: std_logic; attribute dont_touch of G5189: signal is true;
	signal G5190: std_logic; attribute dont_touch of G5190: signal is true;
	signal G5191: std_logic; attribute dont_touch of G5191: signal is true;
	signal G5192: std_logic; attribute dont_touch of G5192: signal is true;
	signal G5193: std_logic; attribute dont_touch of G5193: signal is true;
	signal G5194: std_logic; attribute dont_touch of G5194: signal is true;
	signal G5197: std_logic; attribute dont_touch of G5197: signal is true;
	signal G5198: std_logic; attribute dont_touch of G5198: signal is true;
	signal G5199: std_logic; attribute dont_touch of G5199: signal is true;
	signal G5200: std_logic; attribute dont_touch of G5200: signal is true;
	signal G5201: std_logic; attribute dont_touch of G5201: signal is true;
	signal G5202: std_logic; attribute dont_touch of G5202: signal is true;
	signal G5209: std_logic; attribute dont_touch of G5209: signal is true;
	signal G5210: std_logic; attribute dont_touch of G5210: signal is true;
	signal G5211: std_logic; attribute dont_touch of G5211: signal is true;
	signal G5212: std_logic; attribute dont_touch of G5212: signal is true;
	signal G5213: std_logic; attribute dont_touch of G5213: signal is true;
	signal G5214: std_logic; attribute dont_touch of G5214: signal is true;
	signal G5215: std_logic; attribute dont_touch of G5215: signal is true;
	signal G5216: std_logic; attribute dont_touch of G5216: signal is true;
	signal G5217: std_logic; attribute dont_touch of G5217: signal is true;
	signal G5218: std_logic; attribute dont_touch of G5218: signal is true;
	signal G5219: std_logic; attribute dont_touch of G5219: signal is true;
	signal G5220: std_logic; attribute dont_touch of G5220: signal is true;
	signal G5224: std_logic; attribute dont_touch of G5224: signal is true;
	signal G5225: std_logic; attribute dont_touch of G5225: signal is true;
	signal G5226: std_logic; attribute dont_touch of G5226: signal is true;
	signal G5227: std_logic; attribute dont_touch of G5227: signal is true;
	signal G5228: std_logic; attribute dont_touch of G5228: signal is true;
	signal G5229: std_logic; attribute dont_touch of G5229: signal is true;
	signal G5230: std_logic; attribute dont_touch of G5230: signal is true;
	signal G5231: std_logic; attribute dont_touch of G5231: signal is true;
	signal G5232: std_logic; attribute dont_touch of G5232: signal is true;
	signal G5233: std_logic; attribute dont_touch of G5233: signal is true;
	signal G5234: std_logic; attribute dont_touch of G5234: signal is true;
	signal G5235: std_logic; attribute dont_touch of G5235: signal is true;
	signal G5236: std_logic; attribute dont_touch of G5236: signal is true;
	signal G5237: std_logic; attribute dont_touch of G5237: signal is true;
	signal G5240: std_logic; attribute dont_touch of G5240: signal is true;
	signal G5241: std_logic; attribute dont_touch of G5241: signal is true;
	signal G5242: std_logic; attribute dont_touch of G5242: signal is true;
	signal G5245: std_logic; attribute dont_touch of G5245: signal is true;
	signal G5246: std_logic; attribute dont_touch of G5246: signal is true;
	signal G5247: std_logic; attribute dont_touch of G5247: signal is true;
	signal G5248: std_logic; attribute dont_touch of G5248: signal is true;
	signal G5249: std_logic; attribute dont_touch of G5249: signal is true;
	signal G5250: std_logic; attribute dont_touch of G5250: signal is true;
	signal G5251: std_logic; attribute dont_touch of G5251: signal is true;
	signal G5255: std_logic; attribute dont_touch of G5255: signal is true;
	signal G5256: std_logic; attribute dont_touch of G5256: signal is true;
	signal G5260: std_logic; attribute dont_touch of G5260: signal is true;
	signal G5261: std_logic; attribute dont_touch of G5261: signal is true;
	signal G5264: std_logic; attribute dont_touch of G5264: signal is true;
	signal G5265: std_logic; attribute dont_touch of G5265: signal is true;
	signal G5266: std_logic; attribute dont_touch of G5266: signal is true;
	signal G5269: std_logic; attribute dont_touch of G5269: signal is true;
	signal G5270: std_logic; attribute dont_touch of G5270: signal is true;
	signal G5273: std_logic; attribute dont_touch of G5273: signal is true;
	signal G5274: std_logic; attribute dont_touch of G5274: signal is true;
	signal G5277: std_logic; attribute dont_touch of G5277: signal is true;
	signal G5278: std_logic; attribute dont_touch of G5278: signal is true;
	signal G5281: std_logic; attribute dont_touch of G5281: signal is true;
	signal G5291: std_logic; attribute dont_touch of G5291: signal is true;
	signal G5292: std_logic; attribute dont_touch of G5292: signal is true;
	signal G5295: std_logic; attribute dont_touch of G5295: signal is true;
	signal G5296: std_logic; attribute dont_touch of G5296: signal is true;
	signal G5299: std_logic; attribute dont_touch of G5299: signal is true;
	signal G5300: std_logic; attribute dont_touch of G5300: signal is true;
	signal G5303: std_logic; attribute dont_touch of G5303: signal is true;
	signal G5304: std_logic; attribute dont_touch of G5304: signal is true;
	signal G5307: std_logic; attribute dont_touch of G5307: signal is true;
	signal G5308: std_logic; attribute dont_touch of G5308: signal is true;
	signal G5309: std_logic; attribute dont_touch of G5309: signal is true;
	signal G5310: std_logic; attribute dont_touch of G5310: signal is true;
	signal G5311: std_logic; attribute dont_touch of G5311: signal is true;
	signal G5314: std_logic; attribute dont_touch of G5314: signal is true;
	signal G5315: std_logic; attribute dont_touch of G5315: signal is true;
	signal G5316: std_logic; attribute dont_touch of G5316: signal is true;
	signal G5317: std_logic; attribute dont_touch of G5317: signal is true;
	signal G5318: std_logic; attribute dont_touch of G5318: signal is true;
	signal G5323: std_logic; attribute dont_touch of G5323: signal is true;
	signal G5324: std_logic; attribute dont_touch of G5324: signal is true;
	signal G5325: std_logic; attribute dont_touch of G5325: signal is true;
	signal G5326: std_logic; attribute dont_touch of G5326: signal is true;
	signal G5327: std_logic; attribute dont_touch of G5327: signal is true;
	signal G5328: std_logic; attribute dont_touch of G5328: signal is true;
	signal G5329: std_logic; attribute dont_touch of G5329: signal is true;
	signal G5330: std_logic; attribute dont_touch of G5330: signal is true;
	signal G5331: std_logic; attribute dont_touch of G5331: signal is true;
	signal G5348: std_logic; attribute dont_touch of G5348: signal is true;
	signal G5349: std_logic; attribute dont_touch of G5349: signal is true;
	signal G5350: std_logic; attribute dont_touch of G5350: signal is true;
	signal G5351: std_logic; attribute dont_touch of G5351: signal is true;
	signal G5352: std_logic; attribute dont_touch of G5352: signal is true;
	signal G5353: std_logic; attribute dont_touch of G5353: signal is true;
	signal G5354: std_logic; attribute dont_touch of G5354: signal is true;
	signal G5355: std_logic; attribute dont_touch of G5355: signal is true;
	signal G5356: std_logic; attribute dont_touch of G5356: signal is true;
	signal G5357: std_logic; attribute dont_touch of G5357: signal is true;
	signal G5358: std_logic; attribute dont_touch of G5358: signal is true;
	signal G5359: std_logic; attribute dont_touch of G5359: signal is true;
	signal G5360: std_logic; attribute dont_touch of G5360: signal is true;
	signal G5361: std_logic; attribute dont_touch of G5361: signal is true;
	signal G5362: std_logic; attribute dont_touch of G5362: signal is true;
	signal G5363: std_logic; attribute dont_touch of G5363: signal is true;
	signal G5364: std_logic; attribute dont_touch of G5364: signal is true;
	signal G5367: std_logic; attribute dont_touch of G5367: signal is true;
	signal G5368: std_logic; attribute dont_touch of G5368: signal is true;
	signal G5369: std_logic; attribute dont_touch of G5369: signal is true;
	signal G5370: std_logic; attribute dont_touch of G5370: signal is true;
	signal G5371: std_logic; attribute dont_touch of G5371: signal is true;
	signal G5372: std_logic; attribute dont_touch of G5372: signal is true;
	signal G5373: std_logic; attribute dont_touch of G5373: signal is true;
	signal G5374: std_logic; attribute dont_touch of G5374: signal is true;
	signal G5375: std_logic; attribute dont_touch of G5375: signal is true;
	signal G5376: std_logic; attribute dont_touch of G5376: signal is true;
	signal G5377: std_logic; attribute dont_touch of G5377: signal is true;
	signal G5378: std_logic; attribute dont_touch of G5378: signal is true;
	signal G5379: std_logic; attribute dont_touch of G5379: signal is true;
	signal G5380: std_logic; attribute dont_touch of G5380: signal is true;
	signal G5381: std_logic; attribute dont_touch of G5381: signal is true;
	signal G5382: std_logic; attribute dont_touch of G5382: signal is true;
	signal G5383: std_logic; attribute dont_touch of G5383: signal is true;
	signal G5384: std_logic; attribute dont_touch of G5384: signal is true;
	signal G5385: std_logic; attribute dont_touch of G5385: signal is true;
	signal G5386: std_logic; attribute dont_touch of G5386: signal is true;
	signal G5387: std_logic; attribute dont_touch of G5387: signal is true;
	signal G5388: std_logic; attribute dont_touch of G5388: signal is true;
	signal G5391: std_logic; attribute dont_touch of G5391: signal is true;
	signal G5392: std_logic; attribute dont_touch of G5392: signal is true;
	signal G5395: std_logic; attribute dont_touch of G5395: signal is true;
	signal G5398: std_logic; attribute dont_touch of G5398: signal is true;
	signal G5399: std_logic; attribute dont_touch of G5399: signal is true;
	signal G5402: std_logic; attribute dont_touch of G5402: signal is true;
	signal G5403: std_logic; attribute dont_touch of G5403: signal is true;
	signal G5406: std_logic; attribute dont_touch of G5406: signal is true;
	signal G5407: std_logic; attribute dont_touch of G5407: signal is true;
	signal G5410: std_logic; attribute dont_touch of G5410: signal is true;
	signal G5411: std_logic; attribute dont_touch of G5411: signal is true;
	signal G5414: std_logic; attribute dont_touch of G5414: signal is true;
	signal G5415: std_logic; attribute dont_touch of G5415: signal is true;
	signal G5418: std_logic; attribute dont_touch of G5418: signal is true;
	signal G5419: std_logic; attribute dont_touch of G5419: signal is true;
	signal G5420: std_logic; attribute dont_touch of G5420: signal is true;
	signal G5423: std_logic; attribute dont_touch of G5423: signal is true;
	signal G5424: std_logic; attribute dont_touch of G5424: signal is true;
	signal G5425: std_logic; attribute dont_touch of G5425: signal is true;
	signal G5428: std_logic; attribute dont_touch of G5428: signal is true;
	signal G5429: std_logic; attribute dont_touch of G5429: signal is true;
	signal G5430: std_logic; attribute dont_touch of G5430: signal is true;
	signal G5431: std_logic; attribute dont_touch of G5431: signal is true;
	signal G5432: std_logic; attribute dont_touch of G5432: signal is true;
	signal G5433: std_logic; attribute dont_touch of G5433: signal is true;
	signal G5434: std_logic; attribute dont_touch of G5434: signal is true;
	signal G5435: std_logic; attribute dont_touch of G5435: signal is true;
	signal G5436: std_logic; attribute dont_touch of G5436: signal is true;
	signal G5437: std_logic; attribute dont_touch of G5437: signal is true;
	signal G5438: std_logic; attribute dont_touch of G5438: signal is true;
	signal G5439: std_logic; attribute dont_touch of G5439: signal is true;
	signal G5440: std_logic; attribute dont_touch of G5440: signal is true;
	signal G5441: std_logic; attribute dont_touch of G5441: signal is true;
	signal G5442: std_logic; attribute dont_touch of G5442: signal is true;
	signal G5443: std_logic; attribute dont_touch of G5443: signal is true;
	signal G5444: std_logic; attribute dont_touch of G5444: signal is true;
	signal G5445: std_logic; attribute dont_touch of G5445: signal is true;
	signal G5446: std_logic; attribute dont_touch of G5446: signal is true;
	signal G5447: std_logic; attribute dont_touch of G5447: signal is true;
	signal G5448: std_logic; attribute dont_touch of G5448: signal is true;
	signal G5449: std_logic; attribute dont_touch of G5449: signal is true;
	signal G5450: std_logic; attribute dont_touch of G5450: signal is true;
	signal G5451: std_logic; attribute dont_touch of G5451: signal is true;
	signal G5452: std_logic; attribute dont_touch of G5452: signal is true;
	signal G5453: std_logic; attribute dont_touch of G5453: signal is true;
	signal G5454: std_logic; attribute dont_touch of G5454: signal is true;
	signal G5455: std_logic; attribute dont_touch of G5455: signal is true;
	signal G5456: std_logic; attribute dont_touch of G5456: signal is true;
	signal G5457: std_logic; attribute dont_touch of G5457: signal is true;
	signal G5458: std_logic; attribute dont_touch of G5458: signal is true;
	signal G5465: std_logic; attribute dont_touch of G5465: signal is true;
	signal G5466: std_logic; attribute dont_touch of G5466: signal is true;
	signal G5467: std_logic; attribute dont_touch of G5467: signal is true;
	signal G5470: std_logic; attribute dont_touch of G5470: signal is true;
	signal G5471: std_logic; attribute dont_touch of G5471: signal is true;
	signal G5472: std_logic; attribute dont_touch of G5472: signal is true;
	signal G5473: std_logic; attribute dont_touch of G5473: signal is true;
	signal G5474: std_logic; attribute dont_touch of G5474: signal is true;
	signal G5475: std_logic; attribute dont_touch of G5475: signal is true;
	signal G5476: std_logic; attribute dont_touch of G5476: signal is true;
	signal G5477: std_logic; attribute dont_touch of G5477: signal is true;
	signal G5478: std_logic; attribute dont_touch of G5478: signal is true;
	signal G5479: std_logic; attribute dont_touch of G5479: signal is true;
	signal G5480: std_logic; attribute dont_touch of G5480: signal is true;
	signal G5481: std_logic; attribute dont_touch of G5481: signal is true;
	signal G5482: std_logic; attribute dont_touch of G5482: signal is true;
	signal G5483: std_logic; attribute dont_touch of G5483: signal is true;
	signal G5484: std_logic; attribute dont_touch of G5484: signal is true;
	signal G5485: std_logic; attribute dont_touch of G5485: signal is true;
	signal G5486: std_logic; attribute dont_touch of G5486: signal is true;
	signal G5487: std_logic; attribute dont_touch of G5487: signal is true;
	signal G5488: std_logic; attribute dont_touch of G5488: signal is true;
	signal G5489: std_logic; attribute dont_touch of G5489: signal is true;
	signal G5490: std_logic; attribute dont_touch of G5490: signal is true;
	signal G5491: std_logic; attribute dont_touch of G5491: signal is true;
	signal G5492: std_logic; attribute dont_touch of G5492: signal is true;
	signal G5493: std_logic; attribute dont_touch of G5493: signal is true;
	signal G5494: std_logic; attribute dont_touch of G5494: signal is true;
	signal G5495: std_logic; attribute dont_touch of G5495: signal is true;
	signal G5496: std_logic; attribute dont_touch of G5496: signal is true;
	signal G5497: std_logic; attribute dont_touch of G5497: signal is true;
	signal G5498: std_logic; attribute dont_touch of G5498: signal is true;
	signal G5499: std_logic; attribute dont_touch of G5499: signal is true;
	signal G5500: std_logic; attribute dont_touch of G5500: signal is true;
	signal G5501: std_logic; attribute dont_touch of G5501: signal is true;
	signal G5502: std_logic; attribute dont_touch of G5502: signal is true;
	signal G5503: std_logic; attribute dont_touch of G5503: signal is true;
	signal G5504: std_logic; attribute dont_touch of G5504: signal is true;
	signal G5505: std_logic; attribute dont_touch of G5505: signal is true;
	signal G5506: std_logic; attribute dont_touch of G5506: signal is true;
	signal G5507: std_logic; attribute dont_touch of G5507: signal is true;
	signal G5508: std_logic; attribute dont_touch of G5508: signal is true;
	signal G5509: std_logic; attribute dont_touch of G5509: signal is true;
	signal G5512: std_logic; attribute dont_touch of G5512: signal is true;
	signal G5515: std_logic; attribute dont_touch of G5515: signal is true;
	signal G5518: std_logic; attribute dont_touch of G5518: signal is true;
	signal G5521: std_logic; attribute dont_touch of G5521: signal is true;
	signal G5524: std_logic; attribute dont_touch of G5524: signal is true;
	signal G5527: std_logic; attribute dont_touch of G5527: signal is true;
	signal G5530: std_logic; attribute dont_touch of G5530: signal is true;
	signal G5531: std_logic; attribute dont_touch of G5531: signal is true;
	signal G5532: std_logic; attribute dont_touch of G5532: signal is true;
	signal G5533: std_logic; attribute dont_touch of G5533: signal is true;
	signal G5534: std_logic; attribute dont_touch of G5534: signal is true;
	signal G5535: std_logic; attribute dont_touch of G5535: signal is true;
	signal G5536: std_logic; attribute dont_touch of G5536: signal is true;
	signal G5537: std_logic; attribute dont_touch of G5537: signal is true;
	signal G5538: std_logic; attribute dont_touch of G5538: signal is true;
	signal G5539: std_logic; attribute dont_touch of G5539: signal is true;
	signal G5540: std_logic; attribute dont_touch of G5540: signal is true;
	signal G5541: std_logic; attribute dont_touch of G5541: signal is true;
	signal G5542: std_logic; attribute dont_touch of G5542: signal is true;
	signal G5543: std_logic; attribute dont_touch of G5543: signal is true;
	signal G5544: std_logic; attribute dont_touch of G5544: signal is true;
	signal G5545: std_logic; attribute dont_touch of G5545: signal is true;
	signal G5546: std_logic; attribute dont_touch of G5546: signal is true;
	signal G5549: std_logic; attribute dont_touch of G5549: signal is true;
	signal G5550: std_logic; attribute dont_touch of G5550: signal is true;
	signal G5551: std_logic; attribute dont_touch of G5551: signal is true;
	signal G5552: std_logic; attribute dont_touch of G5552: signal is true;
	signal G5553: std_logic; attribute dont_touch of G5553: signal is true;
	signal G5554: std_logic; attribute dont_touch of G5554: signal is true;
	signal G5555: std_logic; attribute dont_touch of G5555: signal is true;
	signal G5556: std_logic; attribute dont_touch of G5556: signal is true;
	signal G5557: std_logic; attribute dont_touch of G5557: signal is true;
	signal G5558: std_logic; attribute dont_touch of G5558: signal is true;
	signal G5559: std_logic; attribute dont_touch of G5559: signal is true;
	signal G5560: std_logic; attribute dont_touch of G5560: signal is true;
	signal G5561: std_logic; attribute dont_touch of G5561: signal is true;
	signal G5562: std_logic; attribute dont_touch of G5562: signal is true;
	signal G5563: std_logic; attribute dont_touch of G5563: signal is true;
	signal G5564: std_logic; attribute dont_touch of G5564: signal is true;
	signal G5565: std_logic; attribute dont_touch of G5565: signal is true;
	signal G5566: std_logic; attribute dont_touch of G5566: signal is true;
	signal G5567: std_logic; attribute dont_touch of G5567: signal is true;
	signal G5568: std_logic; attribute dont_touch of G5568: signal is true;
	signal G5569: std_logic; attribute dont_touch of G5569: signal is true;
	signal G5570: std_logic; attribute dont_touch of G5570: signal is true;
	signal G5571: std_logic; attribute dont_touch of G5571: signal is true;
	signal G5572: std_logic; attribute dont_touch of G5572: signal is true;
	signal G5573: std_logic; attribute dont_touch of G5573: signal is true;
	signal G5574: std_logic; attribute dont_touch of G5574: signal is true;
	signal G5575: std_logic; attribute dont_touch of G5575: signal is true;
	signal G5576: std_logic; attribute dont_touch of G5576: signal is true;
	signal G5577: std_logic; attribute dont_touch of G5577: signal is true;
	signal G5578: std_logic; attribute dont_touch of G5578: signal is true;
	signal G5579: std_logic; attribute dont_touch of G5579: signal is true;
	signal G5580: std_logic; attribute dont_touch of G5580: signal is true;
	signal G5581: std_logic; attribute dont_touch of G5581: signal is true;
	signal G5582: std_logic; attribute dont_touch of G5582: signal is true;
	signal G5583: std_logic; attribute dont_touch of G5583: signal is true;
	signal G5584: std_logic; attribute dont_touch of G5584: signal is true;
	signal G5587: std_logic; attribute dont_touch of G5587: signal is true;
	signal G5590: std_logic; attribute dont_touch of G5590: signal is true;
	signal G5593: std_logic; attribute dont_touch of G5593: signal is true;
	signal G5596: std_logic; attribute dont_touch of G5596: signal is true;
	signal G5597: std_logic; attribute dont_touch of G5597: signal is true;
	signal G5598: std_logic; attribute dont_touch of G5598: signal is true;
	signal G5599: std_logic; attribute dont_touch of G5599: signal is true;
	signal G5600: std_logic; attribute dont_touch of G5600: signal is true;
	signal G5601: std_logic; attribute dont_touch of G5601: signal is true;
	signal G5602: std_logic; attribute dont_touch of G5602: signal is true;
	signal G5603: std_logic; attribute dont_touch of G5603: signal is true;
	signal G5604: std_logic; attribute dont_touch of G5604: signal is true;
	signal G5605: std_logic; attribute dont_touch of G5605: signal is true;
	signal G5615: std_logic; attribute dont_touch of G5615: signal is true;
	signal G5616: std_logic; attribute dont_touch of G5616: signal is true;
	signal G5617: std_logic; attribute dont_touch of G5617: signal is true;
	signal G5618: std_logic; attribute dont_touch of G5618: signal is true;
	signal G5619: std_logic; attribute dont_touch of G5619: signal is true;
	signal G5620: std_logic; attribute dont_touch of G5620: signal is true;
	signal G5621: std_logic; attribute dont_touch of G5621: signal is true;
	signal G5622: std_logic; attribute dont_touch of G5622: signal is true;
	signal G5623: std_logic; attribute dont_touch of G5623: signal is true;
	signal G5624: std_logic; attribute dont_touch of G5624: signal is true;
	signal G5625: std_logic; attribute dont_touch of G5625: signal is true;
	signal G5626: std_logic; attribute dont_touch of G5626: signal is true;
	signal G5627: std_logic; attribute dont_touch of G5627: signal is true;
	signal G5628: std_logic; attribute dont_touch of G5628: signal is true;
	signal G5629: std_logic; attribute dont_touch of G5629: signal is true;
	signal G5630: std_logic; attribute dont_touch of G5630: signal is true;
	signal G5631: std_logic; attribute dont_touch of G5631: signal is true;
	signal G5632: std_logic; attribute dont_touch of G5632: signal is true;
	signal G5633: std_logic; attribute dont_touch of G5633: signal is true;
	signal G5634: std_logic; attribute dont_touch of G5634: signal is true;
	signal G5635: std_logic; attribute dont_touch of G5635: signal is true;
	signal G5636: std_logic; attribute dont_touch of G5636: signal is true;
	signal G5637: std_logic; attribute dont_touch of G5637: signal is true;
	signal G5638: std_logic; attribute dont_touch of G5638: signal is true;
	signal G5645: std_logic; attribute dont_touch of G5645: signal is true;
	signal G5646: std_logic; attribute dont_touch of G5646: signal is true;
	signal G5647: std_logic; attribute dont_touch of G5647: signal is true;
	signal G5648: std_logic; attribute dont_touch of G5648: signal is true;
	signal G5649: std_logic; attribute dont_touch of G5649: signal is true;
	signal G5658: std_logic; attribute dont_touch of G5658: signal is true;
	signal G5659: std_logic; attribute dont_touch of G5659: signal is true;
	signal G5660: std_logic; attribute dont_touch of G5660: signal is true;
	signal G5661: std_logic; attribute dont_touch of G5661: signal is true;
	signal G5662: std_logic; attribute dont_touch of G5662: signal is true;
	signal G5663: std_logic; attribute dont_touch of G5663: signal is true;
	signal G5664: std_logic; attribute dont_touch of G5664: signal is true;
	signal G5665: std_logic; attribute dont_touch of G5665: signal is true;
	signal G5666: std_logic; attribute dont_touch of G5666: signal is true;
	signal G5667: std_logic; attribute dont_touch of G5667: signal is true;
	signal G5668: std_logic; attribute dont_touch of G5668: signal is true;
	signal G5669: std_logic; attribute dont_touch of G5669: signal is true;
	signal G5670: std_logic; attribute dont_touch of G5670: signal is true;
	signal G5671: std_logic; attribute dont_touch of G5671: signal is true;
	signal G5672: std_logic; attribute dont_touch of G5672: signal is true;
	signal G5673: std_logic; attribute dont_touch of G5673: signal is true;
	signal G5674: std_logic; attribute dont_touch of G5674: signal is true;
	signal G5675: std_logic; attribute dont_touch of G5675: signal is true;
	signal G5676: std_logic; attribute dont_touch of G5676: signal is true;
	signal G5677: std_logic; attribute dont_touch of G5677: signal is true;
	signal G5678: std_logic; attribute dont_touch of G5678: signal is true;
	signal G5679: std_logic; attribute dont_touch of G5679: signal is true;
	signal G5680: std_logic; attribute dont_touch of G5680: signal is true;
	signal G5681: std_logic; attribute dont_touch of G5681: signal is true;
	signal G5682: std_logic; attribute dont_touch of G5682: signal is true;
	signal G5683: std_logic; attribute dont_touch of G5683: signal is true;
	signal G5684: std_logic; attribute dont_touch of G5684: signal is true;
	signal G5685: std_logic; attribute dont_touch of G5685: signal is true;
	signal G5686: std_logic; attribute dont_touch of G5686: signal is true;
	signal G5687: std_logic; attribute dont_touch of G5687: signal is true;
	signal G5688: std_logic; attribute dont_touch of G5688: signal is true;
	signal G5691: std_logic; attribute dont_touch of G5691: signal is true;
	signal G5693: std_logic; attribute dont_touch of G5693: signal is true;
	signal G5694: std_logic; attribute dont_touch of G5694: signal is true;
	signal G5695: std_logic; attribute dont_touch of G5695: signal is true;
	signal G5696: std_logic; attribute dont_touch of G5696: signal is true;
	signal G5697: std_logic; attribute dont_touch of G5697: signal is true;
	signal G5698: std_logic; attribute dont_touch of G5698: signal is true;
	signal G5699: std_logic; attribute dont_touch of G5699: signal is true;
	signal G5700: std_logic; attribute dont_touch of G5700: signal is true;
	signal G5701: std_logic; attribute dont_touch of G5701: signal is true;
	signal G5702: std_logic; attribute dont_touch of G5702: signal is true;
	signal G5705: std_logic; attribute dont_touch of G5705: signal is true;
	signal G5708: std_logic; attribute dont_touch of G5708: signal is true;
	signal G5711: std_logic; attribute dont_touch of G5711: signal is true;
	signal G5714: std_logic; attribute dont_touch of G5714: signal is true;
	signal G5717: std_logic; attribute dont_touch of G5717: signal is true;
	signal G5720: std_logic; attribute dont_touch of G5720: signal is true;
	signal G5723: std_logic; attribute dont_touch of G5723: signal is true;
	signal G5726: std_logic; attribute dont_touch of G5726: signal is true;
	signal G5727: std_logic; attribute dont_touch of G5727: signal is true;
	signal G5728: std_logic; attribute dont_touch of G5728: signal is true;
	signal G5729: std_logic; attribute dont_touch of G5729: signal is true;
	signal G5730: std_logic; attribute dont_touch of G5730: signal is true;
	signal G5731: std_logic; attribute dont_touch of G5731: signal is true;
	signal G5740: std_logic; attribute dont_touch of G5740: signal is true;
	signal G5741: std_logic; attribute dont_touch of G5741: signal is true;
	signal G5742: std_logic; attribute dont_touch of G5742: signal is true;
	signal G5751: std_logic; attribute dont_touch of G5751: signal is true;
	signal G5752: std_logic; attribute dont_touch of G5752: signal is true;
	signal G5753: std_logic; attribute dont_touch of G5753: signal is true;
	signal G5770: std_logic; attribute dont_touch of G5770: signal is true;
	signal G5773: std_logic; attribute dont_touch of G5773: signal is true;
	signal G5774: std_logic; attribute dont_touch of G5774: signal is true;
	signal G5775: std_logic; attribute dont_touch of G5775: signal is true;
	signal G5776: std_logic; attribute dont_touch of G5776: signal is true;
	signal G5777: std_logic; attribute dont_touch of G5777: signal is true;
	signal G5778: std_logic; attribute dont_touch of G5778: signal is true;
	signal G5779: std_logic; attribute dont_touch of G5779: signal is true;
	signal G5780: std_logic; attribute dont_touch of G5780: signal is true;
	signal G5781: std_logic; attribute dont_touch of G5781: signal is true;
	signal G5782: std_logic; attribute dont_touch of G5782: signal is true;
	signal G5783: std_logic; attribute dont_touch of G5783: signal is true;
	signal G5784: std_logic; attribute dont_touch of G5784: signal is true;
	signal G5787: std_logic; attribute dont_touch of G5787: signal is true;
	signal G5788: std_logic; attribute dont_touch of G5788: signal is true;
	signal G5791: std_logic; attribute dont_touch of G5791: signal is true;
	signal G5794: std_logic; attribute dont_touch of G5794: signal is true;
	signal G5797: std_logic; attribute dont_touch of G5797: signal is true;
	signal G5800: std_logic; attribute dont_touch of G5800: signal is true;
	signal G5801: std_logic; attribute dont_touch of G5801: signal is true;
	signal G5804: std_logic; attribute dont_touch of G5804: signal is true;
	signal G5805: std_logic; attribute dont_touch of G5805: signal is true;
	signal G5808: std_logic; attribute dont_touch of G5808: signal is true;
	signal G5809: std_logic; attribute dont_touch of G5809: signal is true;
	signal G5812: std_logic; attribute dont_touch of G5812: signal is true;
	signal G5813: std_logic; attribute dont_touch of G5813: signal is true;
	signal G5816: std_logic; attribute dont_touch of G5816: signal is true;
	signal G5817: std_logic; attribute dont_touch of G5817: signal is true;
	signal G5818: std_logic; attribute dont_touch of G5818: signal is true;
	signal G5821: std_logic; attribute dont_touch of G5821: signal is true;
	signal G5824: std_logic; attribute dont_touch of G5824: signal is true;
	signal G5852: std_logic; attribute dont_touch of G5852: signal is true;
	signal G5853: std_logic; attribute dont_touch of G5853: signal is true;
	signal G5854: std_logic; attribute dont_touch of G5854: signal is true;
	signal G5857: std_logic; attribute dont_touch of G5857: signal is true;
	signal G5860: std_logic; attribute dont_touch of G5860: signal is true;
	signal G5861: std_logic; attribute dont_touch of G5861: signal is true;
	signal G5862: std_logic; attribute dont_touch of G5862: signal is true;
	signal G5863: std_logic; attribute dont_touch of G5863: signal is true;
	signal G5864: std_logic; attribute dont_touch of G5864: signal is true;
	signal G5865: std_logic; attribute dont_touch of G5865: signal is true;
	signal G5866: std_logic; attribute dont_touch of G5866: signal is true;
	signal G5869: std_logic; attribute dont_touch of G5869: signal is true;
	signal G5872: std_logic; attribute dont_touch of G5872: signal is true;
	signal G5873: std_logic; attribute dont_touch of G5873: signal is true;
	signal G5874: std_logic; attribute dont_touch of G5874: signal is true;
	signal G5875: std_logic; attribute dont_touch of G5875: signal is true;
	signal G5876: std_logic; attribute dont_touch of G5876: signal is true;
	signal G5877: std_logic; attribute dont_touch of G5877: signal is true;
	signal G5878: std_logic; attribute dont_touch of G5878: signal is true;
	signal G5879: std_logic; attribute dont_touch of G5879: signal is true;
	signal G5880: std_logic; attribute dont_touch of G5880: signal is true;
	signal G5883: std_logic; attribute dont_touch of G5883: signal is true;
	signal G5884: std_logic; attribute dont_touch of G5884: signal is true;
	signal G5885: std_logic; attribute dont_touch of G5885: signal is true;
	signal G5886: std_logic; attribute dont_touch of G5886: signal is true;
	signal G5887: std_logic; attribute dont_touch of G5887: signal is true;
	signal G5888: std_logic; attribute dont_touch of G5888: signal is true;
	signal G5889: std_logic; attribute dont_touch of G5889: signal is true;
	signal G5890: std_logic; attribute dont_touch of G5890: signal is true;
	signal G5891: std_logic; attribute dont_touch of G5891: signal is true;
	signal G5892: std_logic; attribute dont_touch of G5892: signal is true;
	signal G5893: std_logic; attribute dont_touch of G5893: signal is true;
	signal G5894: std_logic; attribute dont_touch of G5894: signal is true;
	signal G5895: std_logic; attribute dont_touch of G5895: signal is true;
	signal G5896: std_logic; attribute dont_touch of G5896: signal is true;
	signal G5897: std_logic; attribute dont_touch of G5897: signal is true;
	signal G5898: std_logic; attribute dont_touch of G5898: signal is true;
	signal G5899: std_logic; attribute dont_touch of G5899: signal is true;
	signal G5900: std_logic; attribute dont_touch of G5900: signal is true;
	signal G5901: std_logic; attribute dont_touch of G5901: signal is true;
	signal G5902: std_logic; attribute dont_touch of G5902: signal is true;
	signal G5903: std_logic; attribute dont_touch of G5903: signal is true;
	signal G5904: std_logic; attribute dont_touch of G5904: signal is true;
	signal G5905: std_logic; attribute dont_touch of G5905: signal is true;
	signal G5908: std_logic; attribute dont_touch of G5908: signal is true;
	signal G5909: std_logic; attribute dont_touch of G5909: signal is true;
	signal G5910: std_logic; attribute dont_touch of G5910: signal is true;
	signal G5911: std_logic; attribute dont_touch of G5911: signal is true;
	signal G5912: std_logic; attribute dont_touch of G5912: signal is true;
	signal G5915: std_logic; attribute dont_touch of G5915: signal is true;
	signal G5916: std_logic; attribute dont_touch of G5916: signal is true;
	signal G5917: std_logic; attribute dont_touch of G5917: signal is true;
	signal G5918: std_logic; attribute dont_touch of G5918: signal is true;
	signal G5919: std_logic; attribute dont_touch of G5919: signal is true;
	signal G5920: std_logic; attribute dont_touch of G5920: signal is true;
	signal G5921: std_logic; attribute dont_touch of G5921: signal is true;
	signal G5922: std_logic; attribute dont_touch of G5922: signal is true;
	signal G5923: std_logic; attribute dont_touch of G5923: signal is true;
	signal G5924: std_logic; attribute dont_touch of G5924: signal is true;
	signal G5925: std_logic; attribute dont_touch of G5925: signal is true;
	signal G5926: std_logic; attribute dont_touch of G5926: signal is true;
	signal G5935: std_logic; attribute dont_touch of G5935: signal is true;
	signal G5936: std_logic; attribute dont_touch of G5936: signal is true;
	signal G5937: std_logic; attribute dont_touch of G5937: signal is true;
	signal G5938: std_logic; attribute dont_touch of G5938: signal is true;
	signal G5939: std_logic; attribute dont_touch of G5939: signal is true;
	signal G5940: std_logic; attribute dont_touch of G5940: signal is true;
	signal G5941: std_logic; attribute dont_touch of G5941: signal is true;
	signal G5942: std_logic; attribute dont_touch of G5942: signal is true;
	signal G5943: std_logic; attribute dont_touch of G5943: signal is true;
	signal G5944: std_logic; attribute dont_touch of G5944: signal is true;
	signal G5945: std_logic; attribute dont_touch of G5945: signal is true;
	signal G5946: std_logic; attribute dont_touch of G5946: signal is true;
	signal G5947: std_logic; attribute dont_touch of G5947: signal is true;
	signal G5948: std_logic; attribute dont_touch of G5948: signal is true;
	signal G5949: std_logic; attribute dont_touch of G5949: signal is true;
	signal G5950: std_logic; attribute dont_touch of G5950: signal is true;
	signal G5951: std_logic; attribute dont_touch of G5951: signal is true;
	signal G5952: std_logic; attribute dont_touch of G5952: signal is true;
	signal G5953: std_logic; attribute dont_touch of G5953: signal is true;
	signal G5954: std_logic; attribute dont_touch of G5954: signal is true;
	signal G5955: std_logic; attribute dont_touch of G5955: signal is true;
	signal G5956: std_logic; attribute dont_touch of G5956: signal is true;
	signal G5957: std_logic; attribute dont_touch of G5957: signal is true;
	signal G5958: std_logic; attribute dont_touch of G5958: signal is true;
	signal G5975: std_logic; attribute dont_touch of G5975: signal is true;
	signal G5992: std_logic; attribute dont_touch of G5992: signal is true;
	signal G5993: std_logic; attribute dont_touch of G5993: signal is true;
	signal G5994: std_logic; attribute dont_touch of G5994: signal is true;
	signal G5995: std_logic; attribute dont_touch of G5995: signal is true;
	signal G5996: std_logic; attribute dont_touch of G5996: signal is true;
	signal G5997: std_logic; attribute dont_touch of G5997: signal is true;
	signal G6014: std_logic; attribute dont_touch of G6014: signal is true;
	signal G6015: std_logic; attribute dont_touch of G6015: signal is true;
	signal G6032: std_logic; attribute dont_touch of G6032: signal is true;
	signal G6033: std_logic; attribute dont_touch of G6033: signal is true;
	signal G6034: std_logic; attribute dont_touch of G6034: signal is true;
	signal G6035: std_logic; attribute dont_touch of G6035: signal is true;
	signal G6036: std_logic; attribute dont_touch of G6036: signal is true;
	signal G6039: std_logic; attribute dont_touch of G6039: signal is true;
	signal G6040: std_logic; attribute dont_touch of G6040: signal is true;
	signal G6043: std_logic; attribute dont_touch of G6043: signal is true;
	signal G6044: std_logic; attribute dont_touch of G6044: signal is true;
	signal G6047: std_logic; attribute dont_touch of G6047: signal is true;
	signal G6048: std_logic; attribute dont_touch of G6048: signal is true;
	signal G6051: std_logic; attribute dont_touch of G6051: signal is true;
	signal G6052: std_logic; attribute dont_touch of G6052: signal is true;
	signal G6055: std_logic; attribute dont_touch of G6055: signal is true;
	signal G6056: std_logic; attribute dont_touch of G6056: signal is true;
	signal G6057: std_logic; attribute dont_touch of G6057: signal is true;
	signal G6060: std_logic; attribute dont_touch of G6060: signal is true;
	signal G6061: std_logic; attribute dont_touch of G6061: signal is true;
	signal G6062: std_logic; attribute dont_touch of G6062: signal is true;
	signal G6065: std_logic; attribute dont_touch of G6065: signal is true;
	signal G6066: std_logic; attribute dont_touch of G6066: signal is true;
	signal G6067: std_logic; attribute dont_touch of G6067: signal is true;
	signal G6068: std_logic; attribute dont_touch of G6068: signal is true;
	signal G6069: std_logic; attribute dont_touch of G6069: signal is true;
	signal G6070: std_logic; attribute dont_touch of G6070: signal is true;
	signal G6073: std_logic; attribute dont_touch of G6073: signal is true;
	signal G6074: std_logic; attribute dont_touch of G6074: signal is true;
	signal G6075: std_logic; attribute dont_touch of G6075: signal is true;
	signal G6076: std_logic; attribute dont_touch of G6076: signal is true;
	signal G6077: std_logic; attribute dont_touch of G6077: signal is true;
	signal G6078: std_logic; attribute dont_touch of G6078: signal is true;
	signal G6079: std_logic; attribute dont_touch of G6079: signal is true;
	signal G6080: std_logic; attribute dont_touch of G6080: signal is true;
	signal G6081: std_logic; attribute dont_touch of G6081: signal is true;
	signal G6082: std_logic; attribute dont_touch of G6082: signal is true;
	signal G6083: std_logic; attribute dont_touch of G6083: signal is true;
	signal G6084: std_logic; attribute dont_touch of G6084: signal is true;
	signal G6085: std_logic; attribute dont_touch of G6085: signal is true;
	signal G6086: std_logic; attribute dont_touch of G6086: signal is true;
	signal G6087: std_logic; attribute dont_touch of G6087: signal is true;
	signal G6088: std_logic; attribute dont_touch of G6088: signal is true;
	signal G6089: std_logic; attribute dont_touch of G6089: signal is true;
	signal G6090: std_logic; attribute dont_touch of G6090: signal is true;
	signal G6091: std_logic; attribute dont_touch of G6091: signal is true;
	signal G6092: std_logic; attribute dont_touch of G6092: signal is true;
	signal G6093: std_logic; attribute dont_touch of G6093: signal is true;
	signal G6094: std_logic; attribute dont_touch of G6094: signal is true;
	signal G6095: std_logic; attribute dont_touch of G6095: signal is true;
	signal G6096: std_logic; attribute dont_touch of G6096: signal is true;
	signal G6097: std_logic; attribute dont_touch of G6097: signal is true;
	signal G6098: std_logic; attribute dont_touch of G6098: signal is true;
	signal G6099: std_logic; attribute dont_touch of G6099: signal is true;
	signal G6100: std_logic; attribute dont_touch of G6100: signal is true;
	signal G6101: std_logic; attribute dont_touch of G6101: signal is true;
	signal G6102: std_logic; attribute dont_touch of G6102: signal is true;
	signal G6103: std_logic; attribute dont_touch of G6103: signal is true;
	signal G6104: std_logic; attribute dont_touch of G6104: signal is true;
	signal G6105: std_logic; attribute dont_touch of G6105: signal is true;
	signal G6106: std_logic; attribute dont_touch of G6106: signal is true;
	signal G6107: std_logic; attribute dont_touch of G6107: signal is true;
	signal G6108: std_logic; attribute dont_touch of G6108: signal is true;
	signal G6109: std_logic; attribute dont_touch of G6109: signal is true;
	signal G6110: std_logic; attribute dont_touch of G6110: signal is true;
	signal G6113: std_logic; attribute dont_touch of G6113: signal is true;
	signal G6114: std_logic; attribute dont_touch of G6114: signal is true;
	signal G6115: std_logic; attribute dont_touch of G6115: signal is true;
	signal G6116: std_logic; attribute dont_touch of G6116: signal is true;
	signal G6117: std_logic; attribute dont_touch of G6117: signal is true;
	signal G6118: std_logic; attribute dont_touch of G6118: signal is true;
	signal G6119: std_logic; attribute dont_touch of G6119: signal is true;
	signal G6120: std_logic; attribute dont_touch of G6120: signal is true;
	signal G6121: std_logic; attribute dont_touch of G6121: signal is true;
	signal G6122: std_logic; attribute dont_touch of G6122: signal is true;
	signal G6123: std_logic; attribute dont_touch of G6123: signal is true;
	signal G6124: std_logic; attribute dont_touch of G6124: signal is true;
	signal G6125: std_logic; attribute dont_touch of G6125: signal is true;
	signal G6126: std_logic; attribute dont_touch of G6126: signal is true;
	signal G6127: std_logic; attribute dont_touch of G6127: signal is true;
	signal G6128: std_logic; attribute dont_touch of G6128: signal is true;
	signal G6129: std_logic; attribute dont_touch of G6129: signal is true;
	signal G6130: std_logic; attribute dont_touch of G6130: signal is true;
	signal G6131: std_logic; attribute dont_touch of G6131: signal is true;
	signal G6132: std_logic; attribute dont_touch of G6132: signal is true;
	signal G6133: std_logic; attribute dont_touch of G6133: signal is true;
	signal G6134: std_logic; attribute dont_touch of G6134: signal is true;
	signal G6135: std_logic; attribute dont_touch of G6135: signal is true;
	signal G6136: std_logic; attribute dont_touch of G6136: signal is true;
	signal G6137: std_logic; attribute dont_touch of G6137: signal is true;
	signal G6140: std_logic; attribute dont_touch of G6140: signal is true;
	signal G6141: std_logic; attribute dont_touch of G6141: signal is true;
	signal G6142: std_logic; attribute dont_touch of G6142: signal is true;
	signal G6143: std_logic; attribute dont_touch of G6143: signal is true;
	signal G6144: std_logic; attribute dont_touch of G6144: signal is true;
	signal G6145: std_logic; attribute dont_touch of G6145: signal is true;
	signal G6146: std_logic; attribute dont_touch of G6146: signal is true;
	signal G6147: std_logic; attribute dont_touch of G6147: signal is true;
	signal G6148: std_logic; attribute dont_touch of G6148: signal is true;
	signal G6149: std_logic; attribute dont_touch of G6149: signal is true;
	signal G6150: std_logic; attribute dont_touch of G6150: signal is true;
	signal G6151: std_logic; attribute dont_touch of G6151: signal is true;
	signal G6152: std_logic; attribute dont_touch of G6152: signal is true;
	signal G6153: std_logic; attribute dont_touch of G6153: signal is true;
	signal G6154: std_logic; attribute dont_touch of G6154: signal is true;
	signal G6155: std_logic; attribute dont_touch of G6155: signal is true;
	signal G6156: std_logic; attribute dont_touch of G6156: signal is true;
	signal G6157: std_logic; attribute dont_touch of G6157: signal is true;
	signal G6158: std_logic; attribute dont_touch of G6158: signal is true;
	signal G6159: std_logic; attribute dont_touch of G6159: signal is true;
	signal G6160: std_logic; attribute dont_touch of G6160: signal is true;
	signal G6161: std_logic; attribute dont_touch of G6161: signal is true;
	signal G6162: std_logic; attribute dont_touch of G6162: signal is true;
	signal G6163: std_logic; attribute dont_touch of G6163: signal is true;
	signal G6164: std_logic; attribute dont_touch of G6164: signal is true;
	signal G6165: std_logic; attribute dont_touch of G6165: signal is true;
	signal G6166: std_logic; attribute dont_touch of G6166: signal is true;
	signal G6167: std_logic; attribute dont_touch of G6167: signal is true;
	signal G6170: std_logic; attribute dont_touch of G6170: signal is true;
	signal G6173: std_logic; attribute dont_touch of G6173: signal is true;
	signal G6176: std_logic; attribute dont_touch of G6176: signal is true;
	signal G6179: std_logic; attribute dont_touch of G6179: signal is true;
	signal G6182: std_logic; attribute dont_touch of G6182: signal is true;
	signal G6185: std_logic; attribute dont_touch of G6185: signal is true;
	signal G6188: std_logic; attribute dont_touch of G6188: signal is true;
	signal G6189: std_logic; attribute dont_touch of G6189: signal is true;
	signal G6192: std_logic; attribute dont_touch of G6192: signal is true;
	signal G6193: std_logic; attribute dont_touch of G6193: signal is true;
	signal G6194: std_logic; attribute dont_touch of G6194: signal is true;
	signal G6211: std_logic; attribute dont_touch of G6211: signal is true;
	signal G6212: std_logic; attribute dont_touch of G6212: signal is true;
	signal G6229: std_logic; attribute dont_touch of G6229: signal is true;
	signal G6230: std_logic; attribute dont_touch of G6230: signal is true;
	signal G6231: std_logic; attribute dont_touch of G6231: signal is true;
	signal G6232: std_logic; attribute dont_touch of G6232: signal is true;
	signal G6233: std_logic; attribute dont_touch of G6233: signal is true;
	signal G6234: std_logic; attribute dont_touch of G6234: signal is true;
	signal G6235: std_logic; attribute dont_touch of G6235: signal is true;
	signal G6236: std_logic; attribute dont_touch of G6236: signal is true;
	signal G6237: std_logic; attribute dont_touch of G6237: signal is true;
	signal G6238: std_logic; attribute dont_touch of G6238: signal is true;
	signal G6239: std_logic; attribute dont_touch of G6239: signal is true;
	signal G6240: std_logic; attribute dont_touch of G6240: signal is true;
	signal G6241: std_logic; attribute dont_touch of G6241: signal is true;
	signal G6242: std_logic; attribute dont_touch of G6242: signal is true;
	signal G6243: std_logic; attribute dont_touch of G6243: signal is true;
	signal G6244: std_logic; attribute dont_touch of G6244: signal is true;
	signal G6245: std_logic; attribute dont_touch of G6245: signal is true;
	signal G6246: std_logic; attribute dont_touch of G6246: signal is true;
	signal G6247: std_logic; attribute dont_touch of G6247: signal is true;
	signal G6248: std_logic; attribute dont_touch of G6248: signal is true;
	signal G6249: std_logic; attribute dont_touch of G6249: signal is true;
	signal G6250: std_logic; attribute dont_touch of G6250: signal is true;
	signal G6251: std_logic; attribute dont_touch of G6251: signal is true;
	signal G6252: std_logic; attribute dont_touch of G6252: signal is true;
	signal G6253: std_logic; attribute dont_touch of G6253: signal is true;
	signal G6254: std_logic; attribute dont_touch of G6254: signal is true;
	signal G6255: std_logic; attribute dont_touch of G6255: signal is true;
	signal G6256: std_logic; attribute dont_touch of G6256: signal is true;
	signal G6257: std_logic; attribute dont_touch of G6257: signal is true;
	signal G6258: std_logic; attribute dont_touch of G6258: signal is true;
	signal G6259: std_logic; attribute dont_touch of G6259: signal is true;
	signal G6260: std_logic; attribute dont_touch of G6260: signal is true;
	signal G6261: std_logic; attribute dont_touch of G6261: signal is true;
	signal G6262: std_logic; attribute dont_touch of G6262: signal is true;
	signal G6263: std_logic; attribute dont_touch of G6263: signal is true;
	signal G6264: std_logic; attribute dont_touch of G6264: signal is true;
	signal G6265: std_logic; attribute dont_touch of G6265: signal is true;
	signal G6266: std_logic; attribute dont_touch of G6266: signal is true;
	signal G6267: std_logic; attribute dont_touch of G6267: signal is true;
	signal G6268: std_logic; attribute dont_touch of G6268: signal is true;
	signal G6269: std_logic; attribute dont_touch of G6269: signal is true;
	signal G6270: std_logic; attribute dont_touch of G6270: signal is true;
	signal G6271: std_logic; attribute dont_touch of G6271: signal is true;
	signal G6272: std_logic; attribute dont_touch of G6272: signal is true;
	signal G6273: std_logic; attribute dont_touch of G6273: signal is true;
	signal G6274: std_logic; attribute dont_touch of G6274: signal is true;
	signal G6275: std_logic; attribute dont_touch of G6275: signal is true;
	signal G6276: std_logic; attribute dont_touch of G6276: signal is true;
	signal G6277: std_logic; attribute dont_touch of G6277: signal is true;
	signal G6278: std_logic; attribute dont_touch of G6278: signal is true;
	signal G6279: std_logic; attribute dont_touch of G6279: signal is true;
	signal G6280: std_logic; attribute dont_touch of G6280: signal is true;
	signal G6281: std_logic; attribute dont_touch of G6281: signal is true;
	signal G6283: std_logic; attribute dont_touch of G6283: signal is true;
	signal G6285: std_logic; attribute dont_touch of G6285: signal is true;
	signal G6286: std_logic; attribute dont_touch of G6286: signal is true;
	signal G6287: std_logic; attribute dont_touch of G6287: signal is true;
	signal G6288: std_logic; attribute dont_touch of G6288: signal is true;
	signal G6289: std_logic; attribute dont_touch of G6289: signal is true;
	signal G6290: std_logic; attribute dont_touch of G6290: signal is true;
	signal G6291: std_logic; attribute dont_touch of G6291: signal is true;
	signal G6292: std_logic; attribute dont_touch of G6292: signal is true;
	signal G6293: std_logic; attribute dont_touch of G6293: signal is true;
	signal G6294: std_logic; attribute dont_touch of G6294: signal is true;
	signal G6295: std_logic; attribute dont_touch of G6295: signal is true;
	signal G6296: std_logic; attribute dont_touch of G6296: signal is true;
	signal G6297: std_logic; attribute dont_touch of G6297: signal is true;
	signal G6298: std_logic; attribute dont_touch of G6298: signal is true;
	signal G6299: std_logic; attribute dont_touch of G6299: signal is true;
	signal G6300: std_logic; attribute dont_touch of G6300: signal is true;
	signal G6301: std_logic; attribute dont_touch of G6301: signal is true;
	signal G6302: std_logic; attribute dont_touch of G6302: signal is true;
	signal G6303: std_logic; attribute dont_touch of G6303: signal is true;
	signal G6304: std_logic; attribute dont_touch of G6304: signal is true;
	signal G6305: std_logic; attribute dont_touch of G6305: signal is true;
	signal G6306: std_logic; attribute dont_touch of G6306: signal is true;
	signal G6307: std_logic; attribute dont_touch of G6307: signal is true;
	signal G6308: std_logic; attribute dont_touch of G6308: signal is true;
	signal G6309: std_logic; attribute dont_touch of G6309: signal is true;
	signal G6310: std_logic; attribute dont_touch of G6310: signal is true;
	signal G6311: std_logic; attribute dont_touch of G6311: signal is true;
	signal G6312: std_logic; attribute dont_touch of G6312: signal is true;
	signal G6313: std_logic; attribute dont_touch of G6313: signal is true;
	signal G6314: std_logic; attribute dont_touch of G6314: signal is true;
	signal G6315: std_logic; attribute dont_touch of G6315: signal is true;
	signal G6316: std_logic; attribute dont_touch of G6316: signal is true;
	signal G6317: std_logic; attribute dont_touch of G6317: signal is true;
	signal G6318: std_logic; attribute dont_touch of G6318: signal is true;
	signal G6319: std_logic; attribute dont_touch of G6319: signal is true;
	signal G6320: std_logic; attribute dont_touch of G6320: signal is true;
	signal G6321: std_logic; attribute dont_touch of G6321: signal is true;
	signal G6322: std_logic; attribute dont_touch of G6322: signal is true;
	signal G6323: std_logic; attribute dont_touch of G6323: signal is true;
	signal G6324: std_logic; attribute dont_touch of G6324: signal is true;
	signal G6325: std_logic; attribute dont_touch of G6325: signal is true;
	signal G6326: std_logic; attribute dont_touch of G6326: signal is true;
	signal G6327: std_logic; attribute dont_touch of G6327: signal is true;
	signal G6328: std_logic; attribute dont_touch of G6328: signal is true;
	signal G6329: std_logic; attribute dont_touch of G6329: signal is true;
	signal G6330: std_logic; attribute dont_touch of G6330: signal is true;
	signal G6331: std_logic; attribute dont_touch of G6331: signal is true;
	signal G6332: std_logic; attribute dont_touch of G6332: signal is true;
	signal G6333: std_logic; attribute dont_touch of G6333: signal is true;
	signal G6334: std_logic; attribute dont_touch of G6334: signal is true;
	signal G6335: std_logic; attribute dont_touch of G6335: signal is true;
	signal G6336: std_logic; attribute dont_touch of G6336: signal is true;
	signal G6337: std_logic; attribute dont_touch of G6337: signal is true;
	signal G6338: std_logic; attribute dont_touch of G6338: signal is true;
	signal G6339: std_logic; attribute dont_touch of G6339: signal is true;
	signal G6340: std_logic; attribute dont_touch of G6340: signal is true;
	signal G6341: std_logic; attribute dont_touch of G6341: signal is true;
	signal G6342: std_logic; attribute dont_touch of G6342: signal is true;
	signal G6343: std_logic; attribute dont_touch of G6343: signal is true;
	signal G6344: std_logic; attribute dont_touch of G6344: signal is true;
	signal G6345: std_logic; attribute dont_touch of G6345: signal is true;
	signal G6346: std_logic; attribute dont_touch of G6346: signal is true;
	signal G6347: std_logic; attribute dont_touch of G6347: signal is true;
	signal G6348: std_logic; attribute dont_touch of G6348: signal is true;
	signal G6351: std_logic; attribute dont_touch of G6351: signal is true;
	signal G6352: std_logic; attribute dont_touch of G6352: signal is true;
	signal G6353: std_logic; attribute dont_touch of G6353: signal is true;
	signal G6354: std_logic; attribute dont_touch of G6354: signal is true;
	signal G6357: std_logic; attribute dont_touch of G6357: signal is true;
	signal G6358: std_logic; attribute dont_touch of G6358: signal is true;
	signal G6359: std_logic; attribute dont_touch of G6359: signal is true;
	signal G6361: std_logic; attribute dont_touch of G6361: signal is true;
	signal G6363: std_logic; attribute dont_touch of G6363: signal is true;
	signal G6365: std_logic; attribute dont_touch of G6365: signal is true;
	signal G6367: std_logic; attribute dont_touch of G6367: signal is true;
	signal G6369: std_logic; attribute dont_touch of G6369: signal is true;
	signal G6371: std_logic; attribute dont_touch of G6371: signal is true;
	signal G6373: std_logic; attribute dont_touch of G6373: signal is true;
	signal G6375: std_logic; attribute dont_touch of G6375: signal is true;
	signal G6376: std_logic; attribute dont_touch of G6376: signal is true;
	signal G6385: std_logic; attribute dont_touch of G6385: signal is true;
	signal G6394: std_logic; attribute dont_touch of G6394: signal is true;
	signal G6397: std_logic; attribute dont_touch of G6397: signal is true;
	signal G6400: std_logic; attribute dont_touch of G6400: signal is true;
	signal G6401: std_logic; attribute dont_touch of G6401: signal is true;
	signal G6402: std_logic; attribute dont_touch of G6402: signal is true;
	signal G6403: std_logic; attribute dont_touch of G6403: signal is true;
	signal G6404: std_logic; attribute dont_touch of G6404: signal is true;
	signal G6405: std_logic; attribute dont_touch of G6405: signal is true;
	signal G6406: std_logic; attribute dont_touch of G6406: signal is true;
	signal G6407: std_logic; attribute dont_touch of G6407: signal is true;
	signal G6408: std_logic; attribute dont_touch of G6408: signal is true;
	signal G6409: std_logic; attribute dont_touch of G6409: signal is true;
	signal G6410: std_logic; attribute dont_touch of G6410: signal is true;
	signal G6411: std_logic; attribute dont_touch of G6411: signal is true;
	signal G6412: std_logic; attribute dont_touch of G6412: signal is true;
	signal G6413: std_logic; attribute dont_touch of G6413: signal is true;
	signal G6414: std_logic; attribute dont_touch of G6414: signal is true;
	signal G6415: std_logic; attribute dont_touch of G6415: signal is true;
	signal G6416: std_logic; attribute dont_touch of G6416: signal is true;
	signal G6417: std_logic; attribute dont_touch of G6417: signal is true;
	signal G6418: std_logic; attribute dont_touch of G6418: signal is true;
	signal G6419: std_logic; attribute dont_touch of G6419: signal is true;
	signal G6420: std_logic; attribute dont_touch of G6420: signal is true;
	signal G6421: std_logic; attribute dont_touch of G6421: signal is true;
	signal G6422: std_logic; attribute dont_touch of G6422: signal is true;
	signal G6423: std_logic; attribute dont_touch of G6423: signal is true;
	signal G6424: std_logic; attribute dont_touch of G6424: signal is true;
	signal G6425: std_logic; attribute dont_touch of G6425: signal is true;
	signal G6426: std_logic; attribute dont_touch of G6426: signal is true;
	signal G6427: std_logic; attribute dont_touch of G6427: signal is true;
	signal G6428: std_logic; attribute dont_touch of G6428: signal is true;
	signal G6429: std_logic; attribute dont_touch of G6429: signal is true;
	signal G6430: std_logic; attribute dont_touch of G6430: signal is true;
	signal G6431: std_logic; attribute dont_touch of G6431: signal is true;
	signal G6432: std_logic; attribute dont_touch of G6432: signal is true;
	signal G6433: std_logic; attribute dont_touch of G6433: signal is true;
	signal G6434: std_logic; attribute dont_touch of G6434: signal is true;
	signal G6435: std_logic; attribute dont_touch of G6435: signal is true;
	signal G6436: std_logic; attribute dont_touch of G6436: signal is true;
	signal G6437: std_logic; attribute dont_touch of G6437: signal is true;
	signal G6438: std_logic; attribute dont_touch of G6438: signal is true;
	signal G6439: std_logic; attribute dont_touch of G6439: signal is true;
	signal G6440: std_logic; attribute dont_touch of G6440: signal is true;
	signal G6441: std_logic; attribute dont_touch of G6441: signal is true;
	signal G6442: std_logic; attribute dont_touch of G6442: signal is true;
	signal G6443: std_logic; attribute dont_touch of G6443: signal is true;
	signal G6444: std_logic; attribute dont_touch of G6444: signal is true;
	signal G6445: std_logic; attribute dont_touch of G6445: signal is true;
	signal G6446: std_logic; attribute dont_touch of G6446: signal is true;
	signal G6447: std_logic; attribute dont_touch of G6447: signal is true;
	signal G6448: std_logic; attribute dont_touch of G6448: signal is true;
	signal G6449: std_logic; attribute dont_touch of G6449: signal is true;
	signal G6450: std_logic; attribute dont_touch of G6450: signal is true;
	signal G6451: std_logic; attribute dont_touch of G6451: signal is true;
	signal G6452: std_logic; attribute dont_touch of G6452: signal is true;
	signal G6453: std_logic; attribute dont_touch of G6453: signal is true;
	signal G6454: std_logic; attribute dont_touch of G6454: signal is true;
	signal G6455: std_logic; attribute dont_touch of G6455: signal is true;
	signal G6456: std_logic; attribute dont_touch of G6456: signal is true;
	signal G6457: std_logic; attribute dont_touch of G6457: signal is true;
	signal G6461: std_logic; attribute dont_touch of G6461: signal is true;
	signal G6465: std_logic; attribute dont_touch of G6465: signal is true;
	signal G6466: std_logic; attribute dont_touch of G6466: signal is true;
	signal G6467: std_logic; attribute dont_touch of G6467: signal is true;
	signal G6468: std_logic; attribute dont_touch of G6468: signal is true;
	signal G6469: std_logic; attribute dont_touch of G6469: signal is true;
	signal G6473: std_logic; attribute dont_touch of G6473: signal is true;
	signal G6474: std_logic; attribute dont_touch of G6474: signal is true;
	signal G6478: std_logic; attribute dont_touch of G6478: signal is true;
	signal G6479: std_logic; attribute dont_touch of G6479: signal is true;
	signal G6480: std_logic; attribute dont_touch of G6480: signal is true;
	signal G6481: std_logic; attribute dont_touch of G6481: signal is true;
	signal G6482: std_logic; attribute dont_touch of G6482: signal is true;
	signal G6483: std_logic; attribute dont_touch of G6483: signal is true;
	signal G6484: std_logic; attribute dont_touch of G6484: signal is true;
	signal G6485: std_logic; attribute dont_touch of G6485: signal is true;
	signal G6486: std_logic; attribute dont_touch of G6486: signal is true;
	signal G6487: std_logic; attribute dont_touch of G6487: signal is true;
	signal G6488: std_logic; attribute dont_touch of G6488: signal is true;
	signal G6489: std_logic; attribute dont_touch of G6489: signal is true;
	signal G6490: std_logic; attribute dont_touch of G6490: signal is true;
	signal G6491: std_logic; attribute dont_touch of G6491: signal is true;
	signal G6492: std_logic; attribute dont_touch of G6492: signal is true;
	signal G6493: std_logic; attribute dont_touch of G6493: signal is true;
	signal G6494: std_logic; attribute dont_touch of G6494: signal is true;
	signal G6495: std_logic; attribute dont_touch of G6495: signal is true;
	signal G6496: std_logic; attribute dont_touch of G6496: signal is true;
	signal G6497: std_logic; attribute dont_touch of G6497: signal is true;
	signal G6498: std_logic; attribute dont_touch of G6498: signal is true;
	signal G6499: std_logic; attribute dont_touch of G6499: signal is true;
	signal G6500: std_logic; attribute dont_touch of G6500: signal is true;
	signal G6501: std_logic; attribute dont_touch of G6501: signal is true;
	signal G6502: std_logic; attribute dont_touch of G6502: signal is true;
	signal G6503: std_logic; attribute dont_touch of G6503: signal is true;
	signal G6504: std_logic; attribute dont_touch of G6504: signal is true;
	signal G6505: std_logic; attribute dont_touch of G6505: signal is true;
	signal G6506: std_logic; attribute dont_touch of G6506: signal is true;
	signal G6507: std_logic; attribute dont_touch of G6507: signal is true;
	signal G6508: std_logic; attribute dont_touch of G6508: signal is true;
	signal G6509: std_logic; attribute dont_touch of G6509: signal is true;
	signal G6510: std_logic; attribute dont_touch of G6510: signal is true;
	signal G6511: std_logic; attribute dont_touch of G6511: signal is true;
	signal G6512: std_logic; attribute dont_touch of G6512: signal is true;
	signal G6513: std_logic; attribute dont_touch of G6513: signal is true;
	signal G6514: std_logic; attribute dont_touch of G6514: signal is true;
	signal G6515: std_logic; attribute dont_touch of G6515: signal is true;
	signal G6516: std_logic; attribute dont_touch of G6516: signal is true;
	signal G6517: std_logic; attribute dont_touch of G6517: signal is true;
	signal G6518: std_logic; attribute dont_touch of G6518: signal is true;
	signal G6519: std_logic; attribute dont_touch of G6519: signal is true;
	signal G6520: std_logic; attribute dont_touch of G6520: signal is true;
	signal G6521: std_logic; attribute dont_touch of G6521: signal is true;
	signal G6522: std_logic; attribute dont_touch of G6522: signal is true;
	signal G6523: std_logic; attribute dont_touch of G6523: signal is true;
	signal G6524: std_logic; attribute dont_touch of G6524: signal is true;
	signal G6525: std_logic; attribute dont_touch of G6525: signal is true;
	signal G6526: std_logic; attribute dont_touch of G6526: signal is true;
	signal G6527: std_logic; attribute dont_touch of G6527: signal is true;
	signal G6528: std_logic; attribute dont_touch of G6528: signal is true;
	signal G6529: std_logic; attribute dont_touch of G6529: signal is true;
	signal G6530: std_logic; attribute dont_touch of G6530: signal is true;
	signal G6531: std_logic; attribute dont_touch of G6531: signal is true;
	signal G6532: std_logic; attribute dont_touch of G6532: signal is true;
	signal G6533: std_logic; attribute dont_touch of G6533: signal is true;
	signal G6534: std_logic; attribute dont_touch of G6534: signal is true;
	signal G6535: std_logic; attribute dont_touch of G6535: signal is true;
	signal G6536: std_logic; attribute dont_touch of G6536: signal is true;
	signal G6537: std_logic; attribute dont_touch of G6537: signal is true;
	signal G6538: std_logic; attribute dont_touch of G6538: signal is true;
	signal G6539: std_logic; attribute dont_touch of G6539: signal is true;
	signal G6540: std_logic; attribute dont_touch of G6540: signal is true;
	signal G6541: std_logic; attribute dont_touch of G6541: signal is true;
	signal G6542: std_logic; attribute dont_touch of G6542: signal is true;
	signal G6543: std_logic; attribute dont_touch of G6543: signal is true;
	signal G6544: std_logic; attribute dont_touch of G6544: signal is true;
	signal G6545: std_logic; attribute dont_touch of G6545: signal is true;
	signal G6548: std_logic; attribute dont_touch of G6548: signal is true;
	signal G6549: std_logic; attribute dont_touch of G6549: signal is true;
	signal G6552: std_logic; attribute dont_touch of G6552: signal is true;
	signal G6553: std_logic; attribute dont_touch of G6553: signal is true;
	signal G6554: std_logic; attribute dont_touch of G6554: signal is true;
	signal G6555: std_logic; attribute dont_touch of G6555: signal is true;
	signal G6556: std_logic; attribute dont_touch of G6556: signal is true;
	signal G6557: std_logic; attribute dont_touch of G6557: signal is true;
	signal G6558: std_logic; attribute dont_touch of G6558: signal is true;
	signal G6559: std_logic; attribute dont_touch of G6559: signal is true;
	signal G6560: std_logic; attribute dont_touch of G6560: signal is true;
	signal G6561: std_logic; attribute dont_touch of G6561: signal is true;
	signal G6562: std_logic; attribute dont_touch of G6562: signal is true;
	signal G6563: std_logic; attribute dont_touch of G6563: signal is true;
	signal G6564: std_logic; attribute dont_touch of G6564: signal is true;
	signal G6565: std_logic; attribute dont_touch of G6565: signal is true;
	signal G6566: std_logic; attribute dont_touch of G6566: signal is true;
	signal G6567: std_logic; attribute dont_touch of G6567: signal is true;
	signal G6568: std_logic; attribute dont_touch of G6568: signal is true;
	signal G6569: std_logic; attribute dont_touch of G6569: signal is true;
	signal G6570: std_logic; attribute dont_touch of G6570: signal is true;
	signal G6571: std_logic; attribute dont_touch of G6571: signal is true;
	signal G6572: std_logic; attribute dont_touch of G6572: signal is true;
	signal G6573: std_logic; attribute dont_touch of G6573: signal is true;
	signal G6574: std_logic; attribute dont_touch of G6574: signal is true;
	signal G6575: std_logic; attribute dont_touch of G6575: signal is true;
	signal G6576: std_logic; attribute dont_touch of G6576: signal is true;
	signal G6577: std_logic; attribute dont_touch of G6577: signal is true;
	signal G6578: std_logic; attribute dont_touch of G6578: signal is true;
	signal G6579: std_logic; attribute dont_touch of G6579: signal is true;
	signal G6580: std_logic; attribute dont_touch of G6580: signal is true;
	signal G6581: std_logic; attribute dont_touch of G6581: signal is true;
	signal G6582: std_logic; attribute dont_touch of G6582: signal is true;
	signal G6583: std_logic; attribute dont_touch of G6583: signal is true;
	signal G6584: std_logic; attribute dont_touch of G6584: signal is true;
	signal G6585: std_logic; attribute dont_touch of G6585: signal is true;
	signal G6586: std_logic; attribute dont_touch of G6586: signal is true;
	signal G6587: std_logic; attribute dont_touch of G6587: signal is true;
	signal G6588: std_logic; attribute dont_touch of G6588: signal is true;
	signal G6589: std_logic; attribute dont_touch of G6589: signal is true;
	signal G6590: std_logic; attribute dont_touch of G6590: signal is true;
	signal G6591: std_logic; attribute dont_touch of G6591: signal is true;
	signal G6592: std_logic; attribute dont_touch of G6592: signal is true;
	signal G6593: std_logic; attribute dont_touch of G6593: signal is true;
	signal G6594: std_logic; attribute dont_touch of G6594: signal is true;
	signal G6595: std_logic; attribute dont_touch of G6595: signal is true;
	signal G6596: std_logic; attribute dont_touch of G6596: signal is true;
	signal G6597: std_logic; attribute dont_touch of G6597: signal is true;
	signal G6598: std_logic; attribute dont_touch of G6598: signal is true;
	signal G6599: std_logic; attribute dont_touch of G6599: signal is true;
	signal G6600: std_logic; attribute dont_touch of G6600: signal is true;
	signal G6601: std_logic; attribute dont_touch of G6601: signal is true;
	signal G6602: std_logic; attribute dont_touch of G6602: signal is true;
	signal G6603: std_logic; attribute dont_touch of G6603: signal is true;
	signal G6604: std_logic; attribute dont_touch of G6604: signal is true;
	signal G6605: std_logic; attribute dont_touch of G6605: signal is true;
	signal G6606: std_logic; attribute dont_touch of G6606: signal is true;
	signal G6607: std_logic; attribute dont_touch of G6607: signal is true;
	signal G6608: std_logic; attribute dont_touch of G6608: signal is true;
	signal G6609: std_logic; attribute dont_touch of G6609: signal is true;
	signal G6610: std_logic; attribute dont_touch of G6610: signal is true;
	signal G6611: std_logic; attribute dont_touch of G6611: signal is true;
	signal G6612: std_logic; attribute dont_touch of G6612: signal is true;
	signal G6613: std_logic; attribute dont_touch of G6613: signal is true;
	signal G6614: std_logic; attribute dont_touch of G6614: signal is true;
	signal G6615: std_logic; attribute dont_touch of G6615: signal is true;
	signal G6616: std_logic; attribute dont_touch of G6616: signal is true;
	signal G6617: std_logic; attribute dont_touch of G6617: signal is true;
	signal G6618: std_logic; attribute dont_touch of G6618: signal is true;
	signal G6619: std_logic; attribute dont_touch of G6619: signal is true;
	signal G6620: std_logic; attribute dont_touch of G6620: signal is true;
	signal G6621: std_logic; attribute dont_touch of G6621: signal is true;
	signal G6622: std_logic; attribute dont_touch of G6622: signal is true;
	signal G6623: std_logic; attribute dont_touch of G6623: signal is true;
	signal G6624: std_logic; attribute dont_touch of G6624: signal is true;
	signal G6625: std_logic; attribute dont_touch of G6625: signal is true;
	signal G6628: std_logic; attribute dont_touch of G6628: signal is true;
	signal G6631: std_logic; attribute dont_touch of G6631: signal is true;
	signal G6634: std_logic; attribute dont_touch of G6634: signal is true;
	signal G6637: std_logic; attribute dont_touch of G6637: signal is true;
	signal G6640: std_logic; attribute dont_touch of G6640: signal is true;
	signal G6643: std_logic; attribute dont_touch of G6643: signal is true;
	signal G6644: std_logic; attribute dont_touch of G6644: signal is true;
	signal G6645: std_logic; attribute dont_touch of G6645: signal is true;
	signal G6646: std_logic; attribute dont_touch of G6646: signal is true;
	signal G6647: std_logic; attribute dont_touch of G6647: signal is true;
	signal G6648: std_logic; attribute dont_touch of G6648: signal is true;
	signal G6649: std_logic; attribute dont_touch of G6649: signal is true;
	signal G6650: std_logic; attribute dont_touch of G6650: signal is true;
	signal G6651: std_logic; attribute dont_touch of G6651: signal is true;
	signal G6652: std_logic; attribute dont_touch of G6652: signal is true;
	signal G6653: std_logic; attribute dont_touch of G6653: signal is true;
	signal G6654: std_logic; attribute dont_touch of G6654: signal is true;
	signal G6655: std_logic; attribute dont_touch of G6655: signal is true;
	signal G6656: std_logic; attribute dont_touch of G6656: signal is true;
	signal G6657: std_logic; attribute dont_touch of G6657: signal is true;
	signal G6658: std_logic; attribute dont_touch of G6658: signal is true;
	signal G6659: std_logic; attribute dont_touch of G6659: signal is true;
	signal G6660: std_logic; attribute dont_touch of G6660: signal is true;
	signal G6661: std_logic; attribute dont_touch of G6661: signal is true;
	signal G6665: std_logic; attribute dont_touch of G6665: signal is true;
	signal G6669: std_logic; attribute dont_touch of G6669: signal is true;
	signal G6670: std_logic; attribute dont_touch of G6670: signal is true;
	signal G6673: std_logic; attribute dont_touch of G6673: signal is true;
	signal G6676: std_logic; attribute dont_touch of G6676: signal is true;
	signal G6679: std_logic; attribute dont_touch of G6679: signal is true;
	signal G6682: std_logic; attribute dont_touch of G6682: signal is true;
	signal G6683: std_logic; attribute dont_touch of G6683: signal is true;
	signal G6684: std_logic; attribute dont_touch of G6684: signal is true;
	signal G6685: std_logic; attribute dont_touch of G6685: signal is true;
	signal G6686: std_logic; attribute dont_touch of G6686: signal is true;
	signal G6687: std_logic; attribute dont_touch of G6687: signal is true;
	signal G6688: std_logic; attribute dont_touch of G6688: signal is true;
	signal G6689: std_logic; attribute dont_touch of G6689: signal is true;
	signal G6690: std_logic; attribute dont_touch of G6690: signal is true;
	signal G6691: std_logic; attribute dont_touch of G6691: signal is true;
	signal G6692: std_logic; attribute dont_touch of G6692: signal is true;
	signal G6693: std_logic; attribute dont_touch of G6693: signal is true;
	signal G6694: std_logic; attribute dont_touch of G6694: signal is true;
	signal G6695: std_logic; attribute dont_touch of G6695: signal is true;
	signal G6696: std_logic; attribute dont_touch of G6696: signal is true;
	signal G6697: std_logic; attribute dont_touch of G6697: signal is true;
	signal G6698: std_logic; attribute dont_touch of G6698: signal is true;
	signal G6699: std_logic; attribute dont_touch of G6699: signal is true;
	signal G6700: std_logic; attribute dont_touch of G6700: signal is true;
	signal G6701: std_logic; attribute dont_touch of G6701: signal is true;
	signal G6702: std_logic; attribute dont_touch of G6702: signal is true;
	signal G6703: std_logic; attribute dont_touch of G6703: signal is true;
	signal G6704: std_logic; attribute dont_touch of G6704: signal is true;
	signal G6705: std_logic; attribute dont_touch of G6705: signal is true;
	signal G6706: std_logic; attribute dont_touch of G6706: signal is true;
	signal G6707: std_logic; attribute dont_touch of G6707: signal is true;
	signal G6708: std_logic; attribute dont_touch of G6708: signal is true;
	signal G6709: std_logic; attribute dont_touch of G6709: signal is true;
	signal G6710: std_logic; attribute dont_touch of G6710: signal is true;
	signal G6711: std_logic; attribute dont_touch of G6711: signal is true;
	signal G6712: std_logic; attribute dont_touch of G6712: signal is true;
	signal G6713: std_logic; attribute dont_touch of G6713: signal is true;
	signal G6714: std_logic; attribute dont_touch of G6714: signal is true;
	signal G6715: std_logic; attribute dont_touch of G6715: signal is true;
	signal G6716: std_logic; attribute dont_touch of G6716: signal is true;
	signal G6717: std_logic; attribute dont_touch of G6717: signal is true;
	signal G6718: std_logic; attribute dont_touch of G6718: signal is true;
	signal G6719: std_logic; attribute dont_touch of G6719: signal is true;
	signal G6720: std_logic; attribute dont_touch of G6720: signal is true;
	signal G6721: std_logic; attribute dont_touch of G6721: signal is true;
	signal G6722: std_logic; attribute dont_touch of G6722: signal is true;
	signal G6723: std_logic; attribute dont_touch of G6723: signal is true;
	signal G6724: std_logic; attribute dont_touch of G6724: signal is true;
	signal G6725: std_logic; attribute dont_touch of G6725: signal is true;
	signal G6726: std_logic; attribute dont_touch of G6726: signal is true;
	signal G6727: std_logic; attribute dont_touch of G6727: signal is true;
	signal G6729: std_logic; attribute dont_touch of G6729: signal is true;
	signal G6730: std_logic; attribute dont_touch of G6730: signal is true;
	signal G6731: std_logic; attribute dont_touch of G6731: signal is true;
	signal G6732: std_logic; attribute dont_touch of G6732: signal is true;
	signal G6733: std_logic; attribute dont_touch of G6733: signal is true;
	signal G6734: std_logic; attribute dont_touch of G6734: signal is true;
	signal G6735: std_logic; attribute dont_touch of G6735: signal is true;
	signal G6736: std_logic; attribute dont_touch of G6736: signal is true;
	signal G6737: std_logic; attribute dont_touch of G6737: signal is true;
	signal G6738: std_logic; attribute dont_touch of G6738: signal is true;
	signal G6739: std_logic; attribute dont_touch of G6739: signal is true;
	signal G6740: std_logic; attribute dont_touch of G6740: signal is true;
	signal G6741: std_logic; attribute dont_touch of G6741: signal is true;
	signal G6742: std_logic; attribute dont_touch of G6742: signal is true;
	signal G6743: std_logic; attribute dont_touch of G6743: signal is true;
	signal G6744: std_logic; attribute dont_touch of G6744: signal is true;
	signal G6745: std_logic; attribute dont_touch of G6745: signal is true;
	signal G6746: std_logic; attribute dont_touch of G6746: signal is true;
	signal G6747: std_logic; attribute dont_touch of G6747: signal is true;
	signal G6748: std_logic; attribute dont_touch of G6748: signal is true;
	signal G6749: std_logic; attribute dont_touch of G6749: signal is true;
	signal G6750: std_logic; attribute dont_touch of G6750: signal is true;
	signal G6754: std_logic; attribute dont_touch of G6754: signal is true;
	signal G6758: std_logic; attribute dont_touch of G6758: signal is true;
	signal G6762: std_logic; attribute dont_touch of G6762: signal is true;
	signal G6766: std_logic; attribute dont_touch of G6766: signal is true;
	signal G6767: std_logic; attribute dont_touch of G6767: signal is true;
	signal G6768: std_logic; attribute dont_touch of G6768: signal is true;
	signal G6769: std_logic; attribute dont_touch of G6769: signal is true;
	signal G6770: std_logic; attribute dont_touch of G6770: signal is true;
	signal G6771: std_logic; attribute dont_touch of G6771: signal is true;
	signal G6772: std_logic; attribute dont_touch of G6772: signal is true;
	signal G6773: std_logic; attribute dont_touch of G6773: signal is true;
	signal G6774: std_logic; attribute dont_touch of G6774: signal is true;
	signal G6777: std_logic; attribute dont_touch of G6777: signal is true;
	signal G6778: std_logic; attribute dont_touch of G6778: signal is true;
	signal G6781: std_logic; attribute dont_touch of G6781: signal is true;
	signal G6782: std_logic; attribute dont_touch of G6782: signal is true;
	signal G6783: std_logic; attribute dont_touch of G6783: signal is true;
	signal G6784: std_logic; attribute dont_touch of G6784: signal is true;
	signal G6785: std_logic; attribute dont_touch of G6785: signal is true;
	signal G6786: std_logic; attribute dont_touch of G6786: signal is true;
	signal G6787: std_logic; attribute dont_touch of G6787: signal is true;
	signal G6788: std_logic; attribute dont_touch of G6788: signal is true;
	signal G6789: std_logic; attribute dont_touch of G6789: signal is true;
	signal G6790: std_logic; attribute dont_touch of G6790: signal is true;
	signal G6791: std_logic; attribute dont_touch of G6791: signal is true;
	signal G6792: std_logic; attribute dont_touch of G6792: signal is true;
	signal G6793: std_logic; attribute dont_touch of G6793: signal is true;
	signal G6794: std_logic; attribute dont_touch of G6794: signal is true;
	signal G6795: std_logic; attribute dont_touch of G6795: signal is true;
	signal G6796: std_logic; attribute dont_touch of G6796: signal is true;
	signal G6797: std_logic; attribute dont_touch of G6797: signal is true;
	signal G6798: std_logic; attribute dont_touch of G6798: signal is true;
	signal G6799: std_logic; attribute dont_touch of G6799: signal is true;
	signal G6800: std_logic; attribute dont_touch of G6800: signal is true;
	signal G6801: std_logic; attribute dont_touch of G6801: signal is true;
	signal G6802: std_logic; attribute dont_touch of G6802: signal is true;
	signal G6803: std_logic; attribute dont_touch of G6803: signal is true;
	signal G6806: std_logic; attribute dont_touch of G6806: signal is true;
	signal G6809: std_logic; attribute dont_touch of G6809: signal is true;
	signal G6812: std_logic; attribute dont_touch of G6812: signal is true;
	signal G6816: std_logic; attribute dont_touch of G6816: signal is true;
	signal G6817: std_logic; attribute dont_touch of G6817: signal is true;
	signal G6818: std_logic; attribute dont_touch of G6818: signal is true;
	signal G6819: std_logic; attribute dont_touch of G6819: signal is true;
	signal G6820: std_logic; attribute dont_touch of G6820: signal is true;
	signal G6821: std_logic; attribute dont_touch of G6821: signal is true;
	signal G6822: std_logic; attribute dont_touch of G6822: signal is true;
	signal G6823: std_logic; attribute dont_touch of G6823: signal is true;
	signal G6824: std_logic; attribute dont_touch of G6824: signal is true;
	signal G6825: std_logic; attribute dont_touch of G6825: signal is true;
	signal G6826: std_logic; attribute dont_touch of G6826: signal is true;
	signal G6827: std_logic; attribute dont_touch of G6827: signal is true;
	signal G6828: std_logic; attribute dont_touch of G6828: signal is true;
	signal G6829: std_logic; attribute dont_touch of G6829: signal is true;
	signal G6830: std_logic; attribute dont_touch of G6830: signal is true;
	signal G6831: std_logic; attribute dont_touch of G6831: signal is true;
	signal G6832: std_logic; attribute dont_touch of G6832: signal is true;
	signal G6833: std_logic; attribute dont_touch of G6833: signal is true;
	signal G6834: std_logic; attribute dont_touch of G6834: signal is true;
	signal G6835: std_logic; attribute dont_touch of G6835: signal is true;
	signal G6836: std_logic; attribute dont_touch of G6836: signal is true;
	signal G6837: std_logic; attribute dont_touch of G6837: signal is true;
	signal G6838: std_logic; attribute dont_touch of G6838: signal is true;
	signal G6839: std_logic; attribute dont_touch of G6839: signal is true;
	signal G6840: std_logic; attribute dont_touch of G6840: signal is true;
	signal G6841: std_logic; attribute dont_touch of G6841: signal is true;
	signal G6842: std_logic; attribute dont_touch of G6842: signal is true;
	signal G6843: std_logic; attribute dont_touch of G6843: signal is true;
	signal G6844: std_logic; attribute dont_touch of G6844: signal is true;
	signal G6845: std_logic; attribute dont_touch of G6845: signal is true;
	signal G6846: std_logic; attribute dont_touch of G6846: signal is true;
	signal G6847: std_logic; attribute dont_touch of G6847: signal is true;
	signal G6848: std_logic; attribute dont_touch of G6848: signal is true;
	signal G6849: std_logic; attribute dont_touch of G6849: signal is true;
	signal G6850: std_logic; attribute dont_touch of G6850: signal is true;
	signal G6851: std_logic; attribute dont_touch of G6851: signal is true;
	signal G6852: std_logic; attribute dont_touch of G6852: signal is true;
	signal G6853: std_logic; attribute dont_touch of G6853: signal is true;
	signal G6854: std_logic; attribute dont_touch of G6854: signal is true;
	signal G6855: std_logic; attribute dont_touch of G6855: signal is true;
	signal G6864: std_logic; attribute dont_touch of G6864: signal is true;
	signal G6873: std_logic; attribute dont_touch of G6873: signal is true;
	signal G6874: std_logic; attribute dont_touch of G6874: signal is true;
	signal G6875: std_logic; attribute dont_touch of G6875: signal is true;
	signal G6876: std_logic; attribute dont_touch of G6876: signal is true;
	signal G6877: std_logic; attribute dont_touch of G6877: signal is true;
	signal G6878: std_logic; attribute dont_touch of G6878: signal is true;
	signal G6879: std_logic; attribute dont_touch of G6879: signal is true;
	signal G6880: std_logic; attribute dont_touch of G6880: signal is true;
	signal G6881: std_logic; attribute dont_touch of G6881: signal is true;
	signal G6882: std_logic; attribute dont_touch of G6882: signal is true;
	signal G6883: std_logic; attribute dont_touch of G6883: signal is true;
	signal G6884: std_logic; attribute dont_touch of G6884: signal is true;
	signal G6885: std_logic; attribute dont_touch of G6885: signal is true;
	signal G6886: std_logic; attribute dont_touch of G6886: signal is true;
	signal G6887: std_logic; attribute dont_touch of G6887: signal is true;
	signal G6888: std_logic; attribute dont_touch of G6888: signal is true;
	signal G6889: std_logic; attribute dont_touch of G6889: signal is true;
	signal G6890: std_logic; attribute dont_touch of G6890: signal is true;
	signal G6891: std_logic; attribute dont_touch of G6891: signal is true;
	signal G6892: std_logic; attribute dont_touch of G6892: signal is true;
	signal G6893: std_logic; attribute dont_touch of G6893: signal is true;
	signal G6894: std_logic; attribute dont_touch of G6894: signal is true;
	signal G6895: std_logic; attribute dont_touch of G6895: signal is true;
	signal G6896: std_logic; attribute dont_touch of G6896: signal is true;
	signal G6897: std_logic; attribute dont_touch of G6897: signal is true;
	signal G6898: std_logic; attribute dont_touch of G6898: signal is true;
	signal G6899: std_logic; attribute dont_touch of G6899: signal is true;
	signal G6900: std_logic; attribute dont_touch of G6900: signal is true;
	signal G6901: std_logic; attribute dont_touch of G6901: signal is true;
	signal G6902: std_logic; attribute dont_touch of G6902: signal is true;
	signal G6903: std_logic; attribute dont_touch of G6903: signal is true;
	signal G6904: std_logic; attribute dont_touch of G6904: signal is true;
	signal G6905: std_logic; attribute dont_touch of G6905: signal is true;
	signal G6906: std_logic; attribute dont_touch of G6906: signal is true;
	signal G6907: std_logic; attribute dont_touch of G6907: signal is true;
	signal G6908: std_logic; attribute dont_touch of G6908: signal is true;
	signal G6909: std_logic; attribute dont_touch of G6909: signal is true;
	signal G6910: std_logic; attribute dont_touch of G6910: signal is true;
	signal G6911: std_logic; attribute dont_touch of G6911: signal is true;
	signal G6912: std_logic; attribute dont_touch of G6912: signal is true;
	signal G6913: std_logic; attribute dont_touch of G6913: signal is true;
	signal G6914: std_logic; attribute dont_touch of G6914: signal is true;
	signal G6915: std_logic; attribute dont_touch of G6915: signal is true;
	signal G6916: std_logic; attribute dont_touch of G6916: signal is true;
	signal G6917: std_logic; attribute dont_touch of G6917: signal is true;
	signal G6918: std_logic; attribute dont_touch of G6918: signal is true;
	signal G6919: std_logic; attribute dont_touch of G6919: signal is true;
	signal G6920: std_logic; attribute dont_touch of G6920: signal is true;
	signal G6921: std_logic; attribute dont_touch of G6921: signal is true;
	signal G6922: std_logic; attribute dont_touch of G6922: signal is true;
	signal G6923: std_logic; attribute dont_touch of G6923: signal is true;
	signal G6924: std_logic; attribute dont_touch of G6924: signal is true;
	signal G6925: std_logic; attribute dont_touch of G6925: signal is true;
	signal G6926: std_logic; attribute dont_touch of G6926: signal is true;
	signal G6927: std_logic; attribute dont_touch of G6927: signal is true;
	signal G6928: std_logic; attribute dont_touch of G6928: signal is true;
	signal G6929: std_logic; attribute dont_touch of G6929: signal is true;
	signal G6930: std_logic; attribute dont_touch of G6930: signal is true;
	signal G6931: std_logic; attribute dont_touch of G6931: signal is true;
	signal G6932: std_logic; attribute dont_touch of G6932: signal is true;
	signal G6933: std_logic; attribute dont_touch of G6933: signal is true;
	signal G6934: std_logic; attribute dont_touch of G6934: signal is true;
	signal G6935: std_logic; attribute dont_touch of G6935: signal is true;
	signal G6936: std_logic; attribute dont_touch of G6936: signal is true;
	signal G6937: std_logic; attribute dont_touch of G6937: signal is true;
	signal G6938: std_logic; attribute dont_touch of G6938: signal is true;
	signal G6939: std_logic; attribute dont_touch of G6939: signal is true;
	signal G6940: std_logic; attribute dont_touch of G6940: signal is true;
	signal G6941: std_logic; attribute dont_touch of G6941: signal is true;
	signal I1825: std_logic; attribute dont_touch of I1825: signal is true;
	signal I1832: std_logic; attribute dont_touch of I1832: signal is true;
	signal I1835: std_logic; attribute dont_touch of I1835: signal is true;
	signal I1838: std_logic; attribute dont_touch of I1838: signal is true;
	signal I1841: std_logic; attribute dont_touch of I1841: signal is true;
	signal I1844: std_logic; attribute dont_touch of I1844: signal is true;
	signal I1847: std_logic; attribute dont_touch of I1847: signal is true;
	signal I1850: std_logic; attribute dont_touch of I1850: signal is true;
	signal I1853: std_logic; attribute dont_touch of I1853: signal is true;
	signal I1856: std_logic; attribute dont_touch of I1856: signal is true;
	signal I1859: std_logic; attribute dont_touch of I1859: signal is true;
	signal I1862: std_logic; attribute dont_touch of I1862: signal is true;
	signal I1865: std_logic; attribute dont_touch of I1865: signal is true;
	signal I1868: std_logic; attribute dont_touch of I1868: signal is true;
	signal I1871: std_logic; attribute dont_touch of I1871: signal is true;
	signal I1874: std_logic; attribute dont_touch of I1874: signal is true;
	signal I1877: std_logic; attribute dont_touch of I1877: signal is true;
	signal I1880: std_logic; attribute dont_touch of I1880: signal is true;
	signal I1917: std_logic; attribute dont_touch of I1917: signal is true;
	signal I1924: std_logic; attribute dont_touch of I1924: signal is true;
	signal I1927: std_logic; attribute dont_touch of I1927: signal is true;
	signal I1932: std_logic; attribute dont_touch of I1932: signal is true;
	signal I1935: std_logic; attribute dont_touch of I1935: signal is true;
	signal I1938: std_logic; attribute dont_touch of I1938: signal is true;
	signal I1942: std_logic; attribute dont_touch of I1942: signal is true;
	signal I1947: std_logic; attribute dont_touch of I1947: signal is true;
	signal I1951: std_logic; attribute dont_touch of I1951: signal is true;
	signal I1952: std_logic; attribute dont_touch of I1952: signal is true;
	signal I1953: std_logic; attribute dont_touch of I1953: signal is true;
	signal I1958: std_logic; attribute dont_touch of I1958: signal is true;
	signal I1961: std_logic; attribute dont_touch of I1961: signal is true;
	signal I1962: std_logic; attribute dont_touch of I1962: signal is true;
	signal I1963: std_logic; attribute dont_touch of I1963: signal is true;
	signal I1969: std_logic; attribute dont_touch of I1969: signal is true;
	signal I1970: std_logic; attribute dont_touch of I1970: signal is true;
	signal I1971: std_logic; attribute dont_touch of I1971: signal is true;
	signal I1978: std_logic; attribute dont_touch of I1978: signal is true;
	signal I1979: std_logic; attribute dont_touch of I1979: signal is true;
	signal I1980: std_logic; attribute dont_touch of I1980: signal is true;
	signal I1986: std_logic; attribute dont_touch of I1986: signal is true;
	signal I1987: std_logic; attribute dont_touch of I1987: signal is true;
	signal I1988: std_logic; attribute dont_touch of I1988: signal is true;
	signal I1994: std_logic; attribute dont_touch of I1994: signal is true;
	signal I1995: std_logic; attribute dont_touch of I1995: signal is true;
	signal I1996: std_logic; attribute dont_touch of I1996: signal is true;
	signal I2003: std_logic; attribute dont_touch of I2003: signal is true;
	signal I2004: std_logic; attribute dont_touch of I2004: signal is true;
	signal I2005: std_logic; attribute dont_touch of I2005: signal is true;
	signal I2013: std_logic; attribute dont_touch of I2013: signal is true;
	signal I2014: std_logic; attribute dont_touch of I2014: signal is true;
	signal I2015: std_logic; attribute dont_touch of I2015: signal is true;
	signal I2021: std_logic; attribute dont_touch of I2021: signal is true;
	signal I2022: std_logic; attribute dont_touch of I2022: signal is true;
	signal I2023: std_logic; attribute dont_touch of I2023: signal is true;
	signal I2029: std_logic; attribute dont_touch of I2029: signal is true;
	signal I2033: std_logic; attribute dont_touch of I2033: signal is true;
	signal I2037: std_logic; attribute dont_touch of I2037: signal is true;
	signal I2041: std_logic; attribute dont_touch of I2041: signal is true;
	signal I2044: std_logic; attribute dont_touch of I2044: signal is true;
	signal I2047: std_logic; attribute dont_touch of I2047: signal is true;
	signal I2050: std_logic; attribute dont_touch of I2050: signal is true;
	signal I2053: std_logic; attribute dont_touch of I2053: signal is true;
	signal I2057: std_logic; attribute dont_touch of I2057: signal is true;
	signal I2060: std_logic; attribute dont_touch of I2060: signal is true;
	signal I2061: std_logic; attribute dont_touch of I2061: signal is true;
	signal I2062: std_logic; attribute dont_touch of I2062: signal is true;
	signal I2067: std_logic; attribute dont_touch of I2067: signal is true;
	signal I2072: std_logic; attribute dont_touch of I2072: signal is true;
	signal I2073: std_logic; attribute dont_touch of I2073: signal is true;
	signal I2074: std_logic; attribute dont_touch of I2074: signal is true;
	signal I2080: std_logic; attribute dont_touch of I2080: signal is true;
	signal I2081: std_logic; attribute dont_touch of I2081: signal is true;
	signal I2082: std_logic; attribute dont_touch of I2082: signal is true;
	signal I2089: std_logic; attribute dont_touch of I2089: signal is true;
	signal I2090: std_logic; attribute dont_touch of I2090: signal is true;
	signal I2091: std_logic; attribute dont_touch of I2091: signal is true;
	signal I2108: std_logic; attribute dont_touch of I2108: signal is true;
	signal I2109: std_logic; attribute dont_touch of I2109: signal is true;
	signal I2110: std_logic; attribute dont_touch of I2110: signal is true;
	signal I2115: std_logic; attribute dont_touch of I2115: signal is true;
	signal I2119: std_logic; attribute dont_touch of I2119: signal is true;
	signal I2122: std_logic; attribute dont_touch of I2122: signal is true;
	signal I2125: std_logic; attribute dont_touch of I2125: signal is true;
	signal I2128: std_logic; attribute dont_touch of I2128: signal is true;
	signal I2131: std_logic; attribute dont_touch of I2131: signal is true;
	signal I2134: std_logic; attribute dont_touch of I2134: signal is true;
	signal I2137: std_logic; attribute dont_touch of I2137: signal is true;
	signal I2140: std_logic; attribute dont_touch of I2140: signal is true;
	signal I2143: std_logic; attribute dont_touch of I2143: signal is true;
	signal I2147: std_logic; attribute dont_touch of I2147: signal is true;
	signal I2150: std_logic; attribute dont_touch of I2150: signal is true;
	signal I2154: std_logic; attribute dont_touch of I2154: signal is true;
	signal I2159: std_logic; attribute dont_touch of I2159: signal is true;
	signal I2162: std_logic; attribute dont_touch of I2162: signal is true;
	signal I2165: std_logic; attribute dont_touch of I2165: signal is true;
	signal I2169: std_logic; attribute dont_touch of I2169: signal is true;
	signal I2172: std_logic; attribute dont_touch of I2172: signal is true;
	signal I2175: std_logic; attribute dont_touch of I2175: signal is true;
	signal I2179: std_logic; attribute dont_touch of I2179: signal is true;
	signal I2182: std_logic; attribute dont_touch of I2182: signal is true;
	signal I2185: std_logic; attribute dont_touch of I2185: signal is true;
	signal I2190: std_logic; attribute dont_touch of I2190: signal is true;
	signal I2193: std_logic; attribute dont_touch of I2193: signal is true;
	signal I2196: std_logic; attribute dont_touch of I2196: signal is true;
	signal I2199: std_logic; attribute dont_touch of I2199: signal is true;
	signal I2204: std_logic; attribute dont_touch of I2204: signal is true;
	signal I2207: std_logic; attribute dont_touch of I2207: signal is true;
	signal I2212: std_logic; attribute dont_touch of I2212: signal is true;
	signal I2215: std_logic; attribute dont_touch of I2215: signal is true;
	signal I2218: std_logic; attribute dont_touch of I2218: signal is true;
	signal I2221: std_logic; attribute dont_touch of I2221: signal is true;
	signal I2225: std_logic; attribute dont_touch of I2225: signal is true;
	signal I2228: std_logic; attribute dont_touch of I2228: signal is true;
	signal I2231: std_logic; attribute dont_touch of I2231: signal is true;
	signal I2234: std_logic; attribute dont_touch of I2234: signal is true;
	signal I2237: std_logic; attribute dont_touch of I2237: signal is true;
	signal I2240: std_logic; attribute dont_touch of I2240: signal is true;
	signal I2244: std_logic; attribute dont_touch of I2244: signal is true;
	signal I2245: std_logic; attribute dont_touch of I2245: signal is true;
	signal I2246: std_logic; attribute dont_touch of I2246: signal is true;
	signal I2269: std_logic; attribute dont_touch of I2269: signal is true;
	signal I2272: std_logic; attribute dont_touch of I2272: signal is true;
	signal I2275: std_logic; attribute dont_touch of I2275: signal is true;
	signal I2278: std_logic; attribute dont_touch of I2278: signal is true;
	signal I2281: std_logic; attribute dont_touch of I2281: signal is true;
	signal I2284: std_logic; attribute dont_touch of I2284: signal is true;
	signal I2287: std_logic; attribute dont_touch of I2287: signal is true;
	signal I2290: std_logic; attribute dont_touch of I2290: signal is true;
	signal I2293: std_logic; attribute dont_touch of I2293: signal is true;
	signal I2296: std_logic; attribute dont_touch of I2296: signal is true;
	signal I2299: std_logic; attribute dont_touch of I2299: signal is true;
	signal I2300: std_logic; attribute dont_touch of I2300: signal is true;
	signal I2301: std_logic; attribute dont_touch of I2301: signal is true;
	signal I2306: std_logic; attribute dont_touch of I2306: signal is true;
	signal I2309: std_logic; attribute dont_touch of I2309: signal is true;
	signal I2312: std_logic; attribute dont_touch of I2312: signal is true;
	signal I2315: std_logic; attribute dont_touch of I2315: signal is true;
	signal I2318: std_logic; attribute dont_touch of I2318: signal is true;
	signal I2321: std_logic; attribute dont_touch of I2321: signal is true;
	signal I2324: std_logic; attribute dont_touch of I2324: signal is true;
	signal I2327: std_logic; attribute dont_touch of I2327: signal is true;
	signal I2330: std_logic; attribute dont_touch of I2330: signal is true;
	signal I2334: std_logic; attribute dont_touch of I2334: signal is true;
	signal I2337: std_logic; attribute dont_touch of I2337: signal is true;
	signal I2340: std_logic; attribute dont_touch of I2340: signal is true;
	signal I2343: std_logic; attribute dont_touch of I2343: signal is true;
	signal I2346: std_logic; attribute dont_touch of I2346: signal is true;
	signal I2349: std_logic; attribute dont_touch of I2349: signal is true;
	signal I2352: std_logic; attribute dont_touch of I2352: signal is true;
	signal I2355: std_logic; attribute dont_touch of I2355: signal is true;
	signal I2358: std_logic; attribute dont_touch of I2358: signal is true;
	signal I2361: std_logic; attribute dont_touch of I2361: signal is true;
	signal I2364: std_logic; attribute dont_touch of I2364: signal is true;
	signal I2367: std_logic; attribute dont_touch of I2367: signal is true;
	signal I2370: std_logic; attribute dont_touch of I2370: signal is true;
	signal I2373: std_logic; attribute dont_touch of I2373: signal is true;
	signal I2376: std_logic; attribute dont_touch of I2376: signal is true;
	signal I2379: std_logic; attribute dont_touch of I2379: signal is true;
	signal I2382: std_logic; attribute dont_touch of I2382: signal is true;
	signal I2385: std_logic; attribute dont_touch of I2385: signal is true;
	signal I2388: std_logic; attribute dont_touch of I2388: signal is true;
	signal I2391: std_logic; attribute dont_touch of I2391: signal is true;
	signal I2394: std_logic; attribute dont_touch of I2394: signal is true;
	signal I2399: std_logic; attribute dont_touch of I2399: signal is true;
	signal I2402: std_logic; attribute dont_touch of I2402: signal is true;
	signal I2405: std_logic; attribute dont_touch of I2405: signal is true;
	signal I2408: std_logic; attribute dont_touch of I2408: signal is true;
	signal I2411: std_logic; attribute dont_touch of I2411: signal is true;
	signal I2414: std_logic; attribute dont_touch of I2414: signal is true;
	signal I2417: std_logic; attribute dont_touch of I2417: signal is true;
	signal I2420: std_logic; attribute dont_touch of I2420: signal is true;
	signal I2424: std_logic; attribute dont_touch of I2424: signal is true;
	signal I2428: std_logic; attribute dont_touch of I2428: signal is true;
	signal I2442: std_logic; attribute dont_touch of I2442: signal is true;
	signal I2445: std_logic; attribute dont_touch of I2445: signal is true;
	signal I2449: std_logic; attribute dont_touch of I2449: signal is true;
	signal I2453: std_logic; attribute dont_touch of I2453: signal is true;
	signal I2457: std_logic; attribute dont_touch of I2457: signal is true;
	signal I2460: std_logic; attribute dont_touch of I2460: signal is true;
	signal I2464: std_logic; attribute dont_touch of I2464: signal is true;
	signal I2473: std_logic; attribute dont_touch of I2473: signal is true;
	signal I2476: std_logic; attribute dont_touch of I2476: signal is true;
	signal I2479: std_logic; attribute dont_touch of I2479: signal is true;
	signal I2485: std_logic; attribute dont_touch of I2485: signal is true;
	signal I2491: std_logic; attribute dont_touch of I2491: signal is true;
	signal I2497: std_logic; attribute dont_touch of I2497: signal is true;
	signal I2498: std_logic; attribute dont_touch of I2498: signal is true;
	signal I2499: std_logic; attribute dont_touch of I2499: signal is true;
	signal I2506: std_logic; attribute dont_touch of I2506: signal is true;
	signal I2507: std_logic; attribute dont_touch of I2507: signal is true;
	signal I2508: std_logic; attribute dont_touch of I2508: signal is true;
	signal I2521: std_logic; attribute dont_touch of I2521: signal is true;
	signal I2526: std_logic; attribute dont_touch of I2526: signal is true;
	signal I2527: std_logic; attribute dont_touch of I2527: signal is true;
	signal I2528: std_logic; attribute dont_touch of I2528: signal is true;
	signal I2537: std_logic; attribute dont_touch of I2537: signal is true;
	signal I2542: std_logic; attribute dont_touch of I2542: signal is true;
	signal I2543: std_logic; attribute dont_touch of I2543: signal is true;
	signal I2544: std_logic; attribute dont_touch of I2544: signal is true;
	signal I2552: std_logic; attribute dont_touch of I2552: signal is true;
	signal I2566: std_logic; attribute dont_touch of I2566: signal is true;
	signal I2570: std_logic; attribute dont_touch of I2570: signal is true;
	signal I2574: std_logic; attribute dont_touch of I2574: signal is true;
	signal I2578: std_logic; attribute dont_touch of I2578: signal is true;
	signal I2581: std_logic; attribute dont_touch of I2581: signal is true;
	signal I2584: std_logic; attribute dont_touch of I2584: signal is true;
	signal I2588: std_logic; attribute dont_touch of I2588: signal is true;
	signal I2593: std_logic; attribute dont_touch of I2593: signal is true;
	signal I2596: std_logic; attribute dont_touch of I2596: signal is true;
	signal I2601: std_logic; attribute dont_touch of I2601: signal is true;
	signal I2604: std_logic; attribute dont_touch of I2604: signal is true;
	signal I2608: std_logic; attribute dont_touch of I2608: signal is true;
	signal I2611: std_logic; attribute dont_touch of I2611: signal is true;
	signal I2614: std_logic; attribute dont_touch of I2614: signal is true;
	signal I2617: std_logic; attribute dont_touch of I2617: signal is true;
	signal I2620: std_logic; attribute dont_touch of I2620: signal is true;
	signal I2623: std_logic; attribute dont_touch of I2623: signal is true;
	signal I2627: std_logic; attribute dont_touch of I2627: signal is true;
	signal I2630: std_logic; attribute dont_touch of I2630: signal is true;
	signal I2635: std_logic; attribute dont_touch of I2635: signal is true;
	signal I2638: std_logic; attribute dont_touch of I2638: signal is true;
	signal I2643: std_logic; attribute dont_touch of I2643: signal is true;
	signal I2648: std_logic; attribute dont_touch of I2648: signal is true;
	signal I2653: std_logic; attribute dont_touch of I2653: signal is true;
	signal I2658: std_logic; attribute dont_touch of I2658: signal is true;
	signal I2663: std_logic; attribute dont_touch of I2663: signal is true;
	signal I2668: std_logic; attribute dont_touch of I2668: signal is true;
	signal I2671: std_logic; attribute dont_touch of I2671: signal is true;
	signal I2674: std_logic; attribute dont_touch of I2674: signal is true;
	signal I2675: std_logic; attribute dont_touch of I2675: signal is true;
	signal I2676: std_logic; attribute dont_touch of I2676: signal is true;
	signal I2681: std_logic; attribute dont_touch of I2681: signal is true;
	signal I2682: std_logic; attribute dont_touch of I2682: signal is true;
	signal I2683: std_logic; attribute dont_touch of I2683: signal is true;
	signal I2688: std_logic; attribute dont_touch of I2688: signal is true;
	signal I2692: std_logic; attribute dont_touch of I2692: signal is true;
	signal I2696: std_logic; attribute dont_touch of I2696: signal is true;
	signal I2700: std_logic; attribute dont_touch of I2700: signal is true;
	signal I2703: std_logic; attribute dont_touch of I2703: signal is true;
	signal I2707: std_logic; attribute dont_touch of I2707: signal is true;
	signal I2712: std_logic; attribute dont_touch of I2712: signal is true;
	signal I2716: std_logic; attribute dont_touch of I2716: signal is true;
	signal I2721: std_logic; attribute dont_touch of I2721: signal is true;
	signal I2724: std_logic; attribute dont_touch of I2724: signal is true;
	signal I2728: std_logic; attribute dont_touch of I2728: signal is true;
	signal I2731: std_logic; attribute dont_touch of I2731: signal is true;
	signal I2735: std_logic; attribute dont_touch of I2735: signal is true;
	signal I2738: std_logic; attribute dont_touch of I2738: signal is true;
	signal I2741: std_logic; attribute dont_touch of I2741: signal is true;
	signal I2745: std_logic; attribute dont_touch of I2745: signal is true;
	signal I2749: std_logic; attribute dont_touch of I2749: signal is true;
	signal I2753: std_logic; attribute dont_touch of I2753: signal is true;
	signal I2756: std_logic; attribute dont_touch of I2756: signal is true;
	signal I2760: std_logic; attribute dont_touch of I2760: signal is true;
	signal I2763: std_logic; attribute dont_touch of I2763: signal is true;
	signal I2766: std_logic; attribute dont_touch of I2766: signal is true;
	signal I2767: std_logic; attribute dont_touch of I2767: signal is true;
	signal I2768: std_logic; attribute dont_touch of I2768: signal is true;
	signal I2773: std_logic; attribute dont_touch of I2773: signal is true;
	signal I2776: std_logic; attribute dont_touch of I2776: signal is true;
	signal I2779: std_logic; attribute dont_touch of I2779: signal is true;
	signal I2782: std_logic; attribute dont_touch of I2782: signal is true;
	signal I2785: std_logic; attribute dont_touch of I2785: signal is true;
	signal I2788: std_logic; attribute dont_touch of I2788: signal is true;
	signal I2791: std_logic; attribute dont_touch of I2791: signal is true;
	signal I2795: std_logic; attribute dont_touch of I2795: signal is true;
	signal I2796: std_logic; attribute dont_touch of I2796: signal is true;
	signal I2797: std_logic; attribute dont_touch of I2797: signal is true;
	signal I2802: std_logic; attribute dont_touch of I2802: signal is true;
	signal I2805: std_logic; attribute dont_touch of I2805: signal is true;
	signal I2808: std_logic; attribute dont_touch of I2808: signal is true;
	signal I2811: std_logic; attribute dont_touch of I2811: signal is true;
	signal I2814: std_logic; attribute dont_touch of I2814: signal is true;
	signal I2817: std_logic; attribute dont_touch of I2817: signal is true;
	signal I2821: std_logic; attribute dont_touch of I2821: signal is true;
	signal I2825: std_logic; attribute dont_touch of I2825: signal is true;
	signal I2828: std_logic; attribute dont_touch of I2828: signal is true;
	signal I2831: std_logic; attribute dont_touch of I2831: signal is true;
	signal I2835: std_logic; attribute dont_touch of I2835: signal is true;
	signal I2839: std_logic; attribute dont_touch of I2839: signal is true;
	signal I2842: std_logic; attribute dont_touch of I2842: signal is true;
	signal I2845: std_logic; attribute dont_touch of I2845: signal is true;
	signal I2848: std_logic; attribute dont_touch of I2848: signal is true;
	signal I2854: std_logic; attribute dont_touch of I2854: signal is true;
	signal I2857: std_logic; attribute dont_touch of I2857: signal is true;
	signal I2860: std_logic; attribute dont_touch of I2860: signal is true;
	signal I2864: std_logic; attribute dont_touch of I2864: signal is true;
	signal I2867: std_logic; attribute dont_touch of I2867: signal is true;
	signal I2870: std_logic; attribute dont_touch of I2870: signal is true;
	signal I2873: std_logic; attribute dont_touch of I2873: signal is true;
	signal I2877: std_logic; attribute dont_touch of I2877: signal is true;
	signal I2880: std_logic; attribute dont_touch of I2880: signal is true;
	signal I2883: std_logic; attribute dont_touch of I2883: signal is true;
	signal I2887: std_logic; attribute dont_touch of I2887: signal is true;
	signal I2890: std_logic; attribute dont_touch of I2890: signal is true;
	signal I2893: std_logic; attribute dont_touch of I2893: signal is true;
	signal I2897: std_logic; attribute dont_touch of I2897: signal is true;
	signal I2898: std_logic; attribute dont_touch of I2898: signal is true;
	signal I2899: std_logic; attribute dont_touch of I2899: signal is true;
	signal I2904: std_logic; attribute dont_touch of I2904: signal is true;
	signal I2907: std_logic; attribute dont_touch of I2907: signal is true;
	signal I2910: std_logic; attribute dont_touch of I2910: signal is true;
	signal I2913: std_logic; attribute dont_touch of I2913: signal is true;
	signal I2916: std_logic; attribute dont_touch of I2916: signal is true;
	signal I2919: std_logic; attribute dont_touch of I2919: signal is true;
	signal I2922: std_logic; attribute dont_touch of I2922: signal is true;
	signal I2925: std_logic; attribute dont_touch of I2925: signal is true;
	signal I2929: std_logic; attribute dont_touch of I2929: signal is true;
	signal I2933: std_logic; attribute dont_touch of I2933: signal is true;
	signal I2934: std_logic; attribute dont_touch of I2934: signal is true;
	signal I2935: std_logic; attribute dont_touch of I2935: signal is true;
	signal I2940: std_logic; attribute dont_touch of I2940: signal is true;
	signal I2943: std_logic; attribute dont_touch of I2943: signal is true;
	signal I2946: std_logic; attribute dont_touch of I2946: signal is true;
	signal I2949: std_logic; attribute dont_touch of I2949: signal is true;
	signal I2952: std_logic; attribute dont_touch of I2952: signal is true;
	signal I2955: std_logic; attribute dont_touch of I2955: signal is true;
	signal I2958: std_logic; attribute dont_touch of I2958: signal is true;
	signal I2961: std_logic; attribute dont_touch of I2961: signal is true;
	signal I2964: std_logic; attribute dont_touch of I2964: signal is true;
	signal I2967: std_logic; attribute dont_touch of I2967: signal is true;
	signal I2970: std_logic; attribute dont_touch of I2970: signal is true;
	signal I2973: std_logic; attribute dont_touch of I2973: signal is true;
	signal I2979: std_logic; attribute dont_touch of I2979: signal is true;
	signal I2982: std_logic; attribute dont_touch of I2982: signal is true;
	signal I2986: std_logic; attribute dont_touch of I2986: signal is true;
	signal I2989: std_logic; attribute dont_touch of I2989: signal is true;
	signal I2992: std_logic; attribute dont_touch of I2992: signal is true;
	signal I2995: std_logic; attribute dont_touch of I2995: signal is true;
	signal I2998: std_logic; attribute dont_touch of I2998: signal is true;
	signal I3001: std_logic; attribute dont_touch of I3001: signal is true;
	signal I3004: std_logic; attribute dont_touch of I3004: signal is true;
	signal I3007: std_logic; attribute dont_touch of I3007: signal is true;
	signal I3010: std_logic; attribute dont_touch of I3010: signal is true;
	signal I3013: std_logic; attribute dont_touch of I3013: signal is true;
	signal I3016: std_logic; attribute dont_touch of I3016: signal is true;
	signal I3019: std_logic; attribute dont_touch of I3019: signal is true;
	signal I3022: std_logic; attribute dont_touch of I3022: signal is true;
	signal I3025: std_logic; attribute dont_touch of I3025: signal is true;
	signal I3028: std_logic; attribute dont_touch of I3028: signal is true;
	signal I3031: std_logic; attribute dont_touch of I3031: signal is true;
	signal I3034: std_logic; attribute dont_touch of I3034: signal is true;
	signal I3037: std_logic; attribute dont_touch of I3037: signal is true;
	signal I3040: std_logic; attribute dont_touch of I3040: signal is true;
	signal I3044: std_logic; attribute dont_touch of I3044: signal is true;
	signal I3047: std_logic; attribute dont_touch of I3047: signal is true;
	signal I3050: std_logic; attribute dont_touch of I3050: signal is true;
	signal I3053: std_logic; attribute dont_touch of I3053: signal is true;
	signal I3056: std_logic; attribute dont_touch of I3056: signal is true;
	signal I3059: std_logic; attribute dont_touch of I3059: signal is true;
	signal I3062: std_logic; attribute dont_touch of I3062: signal is true;
	signal I3065: std_logic; attribute dont_touch of I3065: signal is true;
	signal I3068: std_logic; attribute dont_touch of I3068: signal is true;
	signal I3071: std_logic; attribute dont_touch of I3071: signal is true;
	signal I3074: std_logic; attribute dont_touch of I3074: signal is true;
	signal I3077: std_logic; attribute dont_touch of I3077: signal is true;
	signal I3080: std_logic; attribute dont_touch of I3080: signal is true;
	signal I3083: std_logic; attribute dont_touch of I3083: signal is true;
	signal I3086: std_logic; attribute dont_touch of I3086: signal is true;
	signal I3090: std_logic; attribute dont_touch of I3090: signal is true;
	signal I3093: std_logic; attribute dont_touch of I3093: signal is true;
	signal I3096: std_logic; attribute dont_touch of I3096: signal is true;
	signal I3099: std_logic; attribute dont_touch of I3099: signal is true;
	signal I3102: std_logic; attribute dont_touch of I3102: signal is true;
	signal I3105: std_logic; attribute dont_touch of I3105: signal is true;
	signal I3109: std_logic; attribute dont_touch of I3109: signal is true;
	signal I3112: std_logic; attribute dont_touch of I3112: signal is true;
	signal I3115: std_logic; attribute dont_touch of I3115: signal is true;
	signal I3125: std_logic; attribute dont_touch of I3125: signal is true;
	signal I3126: std_logic; attribute dont_touch of I3126: signal is true;
	signal I3127: std_logic; attribute dont_touch of I3127: signal is true;
	signal I3134: std_logic; attribute dont_touch of I3134: signal is true;
	signal I3137: std_logic; attribute dont_touch of I3137: signal is true;
	signal I3140: std_logic; attribute dont_touch of I3140: signal is true;
	signal I3144: std_logic; attribute dont_touch of I3144: signal is true;
	signal I3148: std_logic; attribute dont_touch of I3148: signal is true;
	signal I3152: std_logic; attribute dont_touch of I3152: signal is true;
	signal I3155: std_logic; attribute dont_touch of I3155: signal is true;
	signal I3158: std_logic; attribute dont_touch of I3158: signal is true;
	signal I3161: std_logic; attribute dont_touch of I3161: signal is true;
	signal I3168: std_logic; attribute dont_touch of I3168: signal is true;
	signal I3169: std_logic; attribute dont_touch of I3169: signal is true;
	signal I3170: std_logic; attribute dont_touch of I3170: signal is true;
	signal I3177: std_logic; attribute dont_touch of I3177: signal is true;
	signal I3178: std_logic; attribute dont_touch of I3178: signal is true;
	signal I3179: std_logic; attribute dont_touch of I3179: signal is true;
	signal I3188: std_logic; attribute dont_touch of I3188: signal is true;
	signal I3189: std_logic; attribute dont_touch of I3189: signal is true;
	signal I3190: std_logic; attribute dont_touch of I3190: signal is true;
	signal I3198: std_logic; attribute dont_touch of I3198: signal is true;
	signal I3202: std_logic; attribute dont_touch of I3202: signal is true;
	signal I3206: std_logic; attribute dont_touch of I3206: signal is true;
	signal I3212: std_logic; attribute dont_touch of I3212: signal is true;
	signal I3215: std_logic; attribute dont_touch of I3215: signal is true;
	signal I3222: std_logic; attribute dont_touch of I3222: signal is true;
	signal I3225: std_logic; attribute dont_touch of I3225: signal is true;
	signal I3232: std_logic; attribute dont_touch of I3232: signal is true;
	signal I3235: std_logic; attribute dont_touch of I3235: signal is true;
	signal I3240: std_logic; attribute dont_touch of I3240: signal is true;
	signal I3244: std_logic; attribute dont_touch of I3244: signal is true;
	signal I3247: std_logic; attribute dont_touch of I3247: signal is true;
	signal I3251: std_logic; attribute dont_touch of I3251: signal is true;
	signal I3255: std_logic; attribute dont_touch of I3255: signal is true;
	signal I3258: std_logic; attribute dont_touch of I3258: signal is true;
	signal I3261: std_logic; attribute dont_touch of I3261: signal is true;
	signal I3268: std_logic; attribute dont_touch of I3268: signal is true;
	signal I3271: std_logic; attribute dont_touch of I3271: signal is true;
	signal I3274: std_logic; attribute dont_touch of I3274: signal is true;
	signal I3278: std_logic; attribute dont_touch of I3278: signal is true;
	signal I3281: std_logic; attribute dont_touch of I3281: signal is true;
	signal I3284: std_logic; attribute dont_touch of I3284: signal is true;
	signal I3288: std_logic; attribute dont_touch of I3288: signal is true;
	signal I3291: std_logic; attribute dont_touch of I3291: signal is true;
	signal I3294: std_logic; attribute dont_touch of I3294: signal is true;
	signal I3298: std_logic; attribute dont_touch of I3298: signal is true;
	signal I3301: std_logic; attribute dont_touch of I3301: signal is true;
	signal I3304: std_logic; attribute dont_touch of I3304: signal is true;
	signal I3307: std_logic; attribute dont_touch of I3307: signal is true;
	signal I3310: std_logic; attribute dont_touch of I3310: signal is true;
	signal I3313: std_logic; attribute dont_touch of I3313: signal is true;
	signal I3316: std_logic; attribute dont_touch of I3316: signal is true;
	signal I3319: std_logic; attribute dont_touch of I3319: signal is true;
	signal I3322: std_logic; attribute dont_touch of I3322: signal is true;
	signal I3325: std_logic; attribute dont_touch of I3325: signal is true;
	signal I3328: std_logic; attribute dont_touch of I3328: signal is true;
	signal I3331: std_logic; attribute dont_touch of I3331: signal is true;
	signal I3334: std_logic; attribute dont_touch of I3334: signal is true;
	signal I3337: std_logic; attribute dont_touch of I3337: signal is true;
	signal I3340: std_logic; attribute dont_touch of I3340: signal is true;
	signal I3343: std_logic; attribute dont_touch of I3343: signal is true;
	signal I3346: std_logic; attribute dont_touch of I3346: signal is true;
	signal I3349: std_logic; attribute dont_touch of I3349: signal is true;
	signal I3352: std_logic; attribute dont_touch of I3352: signal is true;
	signal I3355: std_logic; attribute dont_touch of I3355: signal is true;
	signal I3358: std_logic; attribute dont_touch of I3358: signal is true;
	signal I3361: std_logic; attribute dont_touch of I3361: signal is true;
	signal I3364: std_logic; attribute dont_touch of I3364: signal is true;
	signal I3367: std_logic; attribute dont_touch of I3367: signal is true;
	signal I3370: std_logic; attribute dont_touch of I3370: signal is true;
	signal I3373: std_logic; attribute dont_touch of I3373: signal is true;
	signal I3376: std_logic; attribute dont_touch of I3376: signal is true;
	signal I3379: std_logic; attribute dont_touch of I3379: signal is true;
	signal I3382: std_logic; attribute dont_touch of I3382: signal is true;
	signal I3385: std_logic; attribute dont_touch of I3385: signal is true;
	signal I3388: std_logic; attribute dont_touch of I3388: signal is true;
	signal I3391: std_logic; attribute dont_touch of I3391: signal is true;
	signal I3395: std_logic; attribute dont_touch of I3395: signal is true;
	signal I3398: std_logic; attribute dont_touch of I3398: signal is true;
	signal I3399: std_logic; attribute dont_touch of I3399: signal is true;
	signal I3400: std_logic; attribute dont_touch of I3400: signal is true;
	signal I3405: std_logic; attribute dont_touch of I3405: signal is true;
	signal I3408: std_logic; attribute dont_touch of I3408: signal is true;
	signal I3411: std_logic; attribute dont_touch of I3411: signal is true;
	signal I3412: std_logic; attribute dont_touch of I3412: signal is true;
	signal I3413: std_logic; attribute dont_touch of I3413: signal is true;
	signal I3419: std_logic; attribute dont_touch of I3419: signal is true;
	signal I3422: std_logic; attribute dont_touch of I3422: signal is true;
	signal I3425: std_logic; attribute dont_touch of I3425: signal is true;
	signal I3428: std_logic; attribute dont_touch of I3428: signal is true;
	signal I3431: std_logic; attribute dont_touch of I3431: signal is true;
	signal I3434: std_logic; attribute dont_touch of I3434: signal is true;
	signal I3441: std_logic; attribute dont_touch of I3441: signal is true;
	signal I3445: std_logic; attribute dont_touch of I3445: signal is true;
	signal I3446: std_logic; attribute dont_touch of I3446: signal is true;
	signal I3447: std_logic; attribute dont_touch of I3447: signal is true;
	signal I3452: std_logic; attribute dont_touch of I3452: signal is true;
	signal I3455: std_logic; attribute dont_touch of I3455: signal is true;
	signal I3456: std_logic; attribute dont_touch of I3456: signal is true;
	signal I3457: std_logic; attribute dont_touch of I3457: signal is true;
	signal I3462: std_logic; attribute dont_touch of I3462: signal is true;
	signal I3465: std_logic; attribute dont_touch of I3465: signal is true;
	signal I3468: std_logic; attribute dont_touch of I3468: signal is true;
	signal I3471: std_logic; attribute dont_touch of I3471: signal is true;
	signal I3474: std_logic; attribute dont_touch of I3474: signal is true;
	signal I3478: std_logic; attribute dont_touch of I3478: signal is true;
	signal I3481: std_logic; attribute dont_touch of I3481: signal is true;
	signal I3485: std_logic; attribute dont_touch of I3485: signal is true;
	signal I3488: std_logic; attribute dont_touch of I3488: signal is true;
	signal I3493: std_logic; attribute dont_touch of I3493: signal is true;
	signal I3496: std_logic; attribute dont_touch of I3496: signal is true;
	signal I3499: std_logic; attribute dont_touch of I3499: signal is true;
	signal I3502: std_logic; attribute dont_touch of I3502: signal is true;
	signal I3505: std_logic; attribute dont_touch of I3505: signal is true;
	signal I3509: std_logic; attribute dont_touch of I3509: signal is true;
	signal I3513: std_logic; attribute dont_touch of I3513: signal is true;
	signal I3516: std_logic; attribute dont_touch of I3516: signal is true;
	signal I3519: std_logic; attribute dont_touch of I3519: signal is true;
	signal I3522: std_logic; attribute dont_touch of I3522: signal is true;
	signal I3525: std_logic; attribute dont_touch of I3525: signal is true;
	signal I3528: std_logic; attribute dont_touch of I3528: signal is true;
	signal I3531: std_logic; attribute dont_touch of I3531: signal is true;
	signal I3534: std_logic; attribute dont_touch of I3534: signal is true;
	signal I3537: std_logic; attribute dont_touch of I3537: signal is true;
	signal I3540: std_logic; attribute dont_touch of I3540: signal is true;
	signal I3543: std_logic; attribute dont_touch of I3543: signal is true;
	signal I3546: std_logic; attribute dont_touch of I3546: signal is true;
	signal I3550: std_logic; attribute dont_touch of I3550: signal is true;
	signal I3553: std_logic; attribute dont_touch of I3553: signal is true;
	signal I3556: std_logic; attribute dont_touch of I3556: signal is true;
	signal I3560: std_logic; attribute dont_touch of I3560: signal is true;
	signal I3563: std_logic; attribute dont_touch of I3563: signal is true;
	signal I3569: std_logic; attribute dont_touch of I3569: signal is true;
	signal I3572: std_logic; attribute dont_touch of I3572: signal is true;
	signal I3575: std_logic; attribute dont_touch of I3575: signal is true;
	signal I3578: std_logic; attribute dont_touch of I3578: signal is true;
	signal I3581: std_logic; attribute dont_touch of I3581: signal is true;
	signal I3584: std_logic; attribute dont_touch of I3584: signal is true;
	signal I3587: std_logic; attribute dont_touch of I3587: signal is true;
	signal I3590: std_logic; attribute dont_touch of I3590: signal is true;
	signal I3593: std_logic; attribute dont_touch of I3593: signal is true;
	signal I3596: std_logic; attribute dont_touch of I3596: signal is true;
	signal I3599: std_logic; attribute dont_touch of I3599: signal is true;
	signal I3602: std_logic; attribute dont_touch of I3602: signal is true;
	signal I3605: std_logic; attribute dont_touch of I3605: signal is true;
	signal I3608: std_logic; attribute dont_touch of I3608: signal is true;
	signal I3611: std_logic; attribute dont_touch of I3611: signal is true;
	signal I3614: std_logic; attribute dont_touch of I3614: signal is true;
	signal I3617: std_logic; attribute dont_touch of I3617: signal is true;
	signal I3620: std_logic; attribute dont_touch of I3620: signal is true;
	signal I3623: std_logic; attribute dont_touch of I3623: signal is true;
	signal I3626: std_logic; attribute dont_touch of I3626: signal is true;
	signal I3629: std_logic; attribute dont_touch of I3629: signal is true;
	signal I3632: std_logic; attribute dont_touch of I3632: signal is true;
	signal I3635: std_logic; attribute dont_touch of I3635: signal is true;
	signal I3638: std_logic; attribute dont_touch of I3638: signal is true;
	signal I3641: std_logic; attribute dont_touch of I3641: signal is true;
	signal I3644: std_logic; attribute dont_touch of I3644: signal is true;
	signal I3647: std_logic; attribute dont_touch of I3647: signal is true;
	signal I3650: std_logic; attribute dont_touch of I3650: signal is true;
	signal I3653: std_logic; attribute dont_touch of I3653: signal is true;
	signal I3656: std_logic; attribute dont_touch of I3656: signal is true;
	signal I3659: std_logic; attribute dont_touch of I3659: signal is true;
	signal I3662: std_logic; attribute dont_touch of I3662: signal is true;
	signal I3665: std_logic; attribute dont_touch of I3665: signal is true;
	signal I3669: std_logic; attribute dont_touch of I3669: signal is true;
	signal I3672: std_logic; attribute dont_touch of I3672: signal is true;
	signal I3675: std_logic; attribute dont_touch of I3675: signal is true;
	signal I3678: std_logic; attribute dont_touch of I3678: signal is true;
	signal I3681: std_logic; attribute dont_touch of I3681: signal is true;
	signal I3684: std_logic; attribute dont_touch of I3684: signal is true;
	signal I3687: std_logic; attribute dont_touch of I3687: signal is true;
	signal I3691: std_logic; attribute dont_touch of I3691: signal is true;
	signal I3694: std_logic; attribute dont_touch of I3694: signal is true;
	signal I3697: std_logic; attribute dont_touch of I3697: signal is true;
	signal I3698: std_logic; attribute dont_touch of I3698: signal is true;
	signal I3699: std_logic; attribute dont_touch of I3699: signal is true;
	signal I3705: std_logic; attribute dont_touch of I3705: signal is true;
	signal I3708: std_logic; attribute dont_touch of I3708: signal is true;
	signal I3711: std_logic; attribute dont_touch of I3711: signal is true;
	signal I3714: std_logic; attribute dont_touch of I3714: signal is true;
	signal I3717: std_logic; attribute dont_touch of I3717: signal is true;
	signal I3720: std_logic; attribute dont_touch of I3720: signal is true;
	signal I3723: std_logic; attribute dont_touch of I3723: signal is true;
	signal I3726: std_logic; attribute dont_touch of I3726: signal is true;
	signal I3729: std_logic; attribute dont_touch of I3729: signal is true;
	signal I3733: std_logic; attribute dont_touch of I3733: signal is true;
	signal I3736: std_logic; attribute dont_touch of I3736: signal is true;
	signal I3739: std_logic; attribute dont_touch of I3739: signal is true;
	signal I3740: std_logic; attribute dont_touch of I3740: signal is true;
	signal I3741: std_logic; attribute dont_touch of I3741: signal is true;
	signal I3746: std_logic; attribute dont_touch of I3746: signal is true;
	signal I3749: std_logic; attribute dont_touch of I3749: signal is true;
	signal I3752: std_logic; attribute dont_touch of I3752: signal is true;
	signal I3755: std_logic; attribute dont_touch of I3755: signal is true;
	signal I3758: std_logic; attribute dont_touch of I3758: signal is true;
	signal I3761: std_logic; attribute dont_touch of I3761: signal is true;
	signal I3764: std_logic; attribute dont_touch of I3764: signal is true;
	signal I3767: std_logic; attribute dont_touch of I3767: signal is true;
	signal I3770: std_logic; attribute dont_touch of I3770: signal is true;
	signal I3773: std_logic; attribute dont_touch of I3773: signal is true;
	signal I3776: std_logic; attribute dont_touch of I3776: signal is true;
	signal I3779: std_logic; attribute dont_touch of I3779: signal is true;
	signal I3782: std_logic; attribute dont_touch of I3782: signal is true;
	signal I3785: std_logic; attribute dont_touch of I3785: signal is true;
	signal I3788: std_logic; attribute dont_touch of I3788: signal is true;
	signal I3791: std_logic; attribute dont_touch of I3791: signal is true;
	signal I3794: std_logic; attribute dont_touch of I3794: signal is true;
	signal I3797: std_logic; attribute dont_touch of I3797: signal is true;
	signal I3800: std_logic; attribute dont_touch of I3800: signal is true;
	signal I3804: std_logic; attribute dont_touch of I3804: signal is true;
	signal I3808: std_logic; attribute dont_touch of I3808: signal is true;
	signal I3811: std_logic; attribute dont_touch of I3811: signal is true;
	signal I3816: std_logic; attribute dont_touch of I3816: signal is true;
	signal I3819: std_logic; attribute dont_touch of I3819: signal is true;
	signal I3823: std_logic; attribute dont_touch of I3823: signal is true;
	signal I3826: std_logic; attribute dont_touch of I3826: signal is true;
	signal I3830: std_logic; attribute dont_touch of I3830: signal is true;
	signal I3833: std_logic; attribute dont_touch of I3833: signal is true;
	signal I3836: std_logic; attribute dont_touch of I3836: signal is true;
	signal I3840: std_logic; attribute dont_touch of I3840: signal is true;
	signal I3843: std_logic; attribute dont_touch of I3843: signal is true;
	signal I3846: std_logic; attribute dont_touch of I3846: signal is true;
	signal I3847: std_logic; attribute dont_touch of I3847: signal is true;
	signal I3848: std_logic; attribute dont_touch of I3848: signal is true;
	signal I3855: std_logic; attribute dont_touch of I3855: signal is true;
	signal I3858: std_logic; attribute dont_touch of I3858: signal is true;
	signal I3861: std_logic; attribute dont_touch of I3861: signal is true;
	signal I3864: std_logic; attribute dont_touch of I3864: signal is true;
	signal I3868: std_logic; attribute dont_touch of I3868: signal is true;
	signal I3871: std_logic; attribute dont_touch of I3871: signal is true;
	signal I3874: std_logic; attribute dont_touch of I3874: signal is true;
	signal I3875: std_logic; attribute dont_touch of I3875: signal is true;
	signal I3876: std_logic; attribute dont_touch of I3876: signal is true;
	signal I3883: std_logic; attribute dont_touch of I3883: signal is true;
	signal I3886: std_logic; attribute dont_touch of I3886: signal is true;
	signal I3890: std_logic; attribute dont_touch of I3890: signal is true;
	signal I3893: std_logic; attribute dont_touch of I3893: signal is true;
	signal I3894: std_logic; attribute dont_touch of I3894: signal is true;
	signal I3895: std_logic; attribute dont_touch of I3895: signal is true;
	signal I3902: std_logic; attribute dont_touch of I3902: signal is true;
	signal I3906: std_logic; attribute dont_touch of I3906: signal is true;
	signal I3909: std_logic; attribute dont_touch of I3909: signal is true;
	signal I3914: std_logic; attribute dont_touch of I3914: signal is true;
	signal I3915: std_logic; attribute dont_touch of I3915: signal is true;
	signal I3916: std_logic; attribute dont_touch of I3916: signal is true;
	signal I3923: std_logic; attribute dont_touch of I3923: signal is true;
	signal I3927: std_logic; attribute dont_touch of I3927: signal is true;
	signal I3933: std_logic; attribute dont_touch of I3933: signal is true;
	signal I3934: std_logic; attribute dont_touch of I3934: signal is true;
	signal I3935: std_logic; attribute dont_touch of I3935: signal is true;
	signal I3942: std_logic; attribute dont_touch of I3942: signal is true;
	signal I3946: std_logic; attribute dont_touch of I3946: signal is true;
	signal I3952: std_logic; attribute dont_touch of I3952: signal is true;
	signal I3953: std_logic; attribute dont_touch of I3953: signal is true;
	signal I3954: std_logic; attribute dont_touch of I3954: signal is true;
	signal I3961: std_logic; attribute dont_touch of I3961: signal is true;
	signal I3965: std_logic; attribute dont_touch of I3965: signal is true;
	signal I3970: std_logic; attribute dont_touch of I3970: signal is true;
	signal I3971: std_logic; attribute dont_touch of I3971: signal is true;
	signal I3972: std_logic; attribute dont_touch of I3972: signal is true;
	signal I3979: std_logic; attribute dont_touch of I3979: signal is true;
	signal I3983: std_logic; attribute dont_touch of I3983: signal is true;
	signal I3988: std_logic; attribute dont_touch of I3988: signal is true;
	signal I3989: std_logic; attribute dont_touch of I3989: signal is true;
	signal I3990: std_logic; attribute dont_touch of I3990: signal is true;
	signal I3999: std_logic; attribute dont_touch of I3999: signal is true;
	signal I4003: std_logic; attribute dont_touch of I4003: signal is true;
	signal I4008: std_logic; attribute dont_touch of I4008: signal is true;
	signal I4009: std_logic; attribute dont_touch of I4009: signal is true;
	signal I4010: std_logic; attribute dont_touch of I4010: signal is true;
	signal I4019: std_logic; attribute dont_touch of I4019: signal is true;
	signal I4023: std_logic; attribute dont_touch of I4023: signal is true;
	signal I4031: std_logic; attribute dont_touch of I4031: signal is true;
	signal I4040: std_logic; attribute dont_touch of I4040: signal is true;
	signal I4050: std_logic; attribute dont_touch of I4050: signal is true;
	signal I4059: std_logic; attribute dont_touch of I4059: signal is true;
	signal I4066: std_logic; attribute dont_touch of I4066: signal is true;
	signal I4123: std_logic; attribute dont_touch of I4123: signal is true;
	signal I4133: std_logic; attribute dont_touch of I4133: signal is true;
	signal I4150: std_logic; attribute dont_touch of I4150: signal is true;
	signal I4151: std_logic; attribute dont_touch of I4151: signal is true;
	signal I4152: std_logic; attribute dont_touch of I4152: signal is true;
	signal I4159: std_logic; attribute dont_touch of I4159: signal is true;
	signal I4160: std_logic; attribute dont_touch of I4160: signal is true;
	signal I4161: std_logic; attribute dont_touch of I4161: signal is true;
	signal I4166: std_logic; attribute dont_touch of I4166: signal is true;
	signal I4170: std_logic; attribute dont_touch of I4170: signal is true;
	signal I4173: std_logic; attribute dont_touch of I4173: signal is true;
	signal I4176: std_logic; attribute dont_touch of I4176: signal is true;
	signal I4182: std_logic; attribute dont_touch of I4182: signal is true;
	signal I4183: std_logic; attribute dont_touch of I4183: signal is true;
	signal I4184: std_logic; attribute dont_touch of I4184: signal is true;
	signal I4189: std_logic; attribute dont_touch of I4189: signal is true;
	signal I4192: std_logic; attribute dont_touch of I4192: signal is true;
	signal I4195: std_logic; attribute dont_touch of I4195: signal is true;
	signal I4198: std_logic; attribute dont_touch of I4198: signal is true;
	signal I4203: std_logic; attribute dont_touch of I4203: signal is true;
	signal I4204: std_logic; attribute dont_touch of I4204: signal is true;
	signal I4205: std_logic; attribute dont_touch of I4205: signal is true;
	signal I4210: std_logic; attribute dont_touch of I4210: signal is true;
	signal I4211: std_logic; attribute dont_touch of I4211: signal is true;
	signal I4212: std_logic; attribute dont_touch of I4212: signal is true;
	signal I4217: std_logic; attribute dont_touch of I4217: signal is true;
	signal I4220: std_logic; attribute dont_touch of I4220: signal is true;
	signal I4223: std_logic; attribute dont_touch of I4223: signal is true;
	signal I4226: std_logic; attribute dont_touch of I4226: signal is true;
	signal I4229: std_logic; attribute dont_touch of I4229: signal is true;
	signal I4233: std_logic; attribute dont_touch of I4233: signal is true;
	signal I4234: std_logic; attribute dont_touch of I4234: signal is true;
	signal I4235: std_logic; attribute dont_touch of I4235: signal is true;
	signal I4240: std_logic; attribute dont_touch of I4240: signal is true;
	signal I4243: std_logic; attribute dont_touch of I4243: signal is true;
	signal I4246: std_logic; attribute dont_touch of I4246: signal is true;
	signal I4249: std_logic; attribute dont_touch of I4249: signal is true;
	signal I4252: std_logic; attribute dont_touch of I4252: signal is true;
	signal I4255: std_logic; attribute dont_touch of I4255: signal is true;
	signal I4258: std_logic; attribute dont_touch of I4258: signal is true;
	signal I4261: std_logic; attribute dont_touch of I4261: signal is true;
	signal I4264: std_logic; attribute dont_touch of I4264: signal is true;
	signal I4267: std_logic; attribute dont_touch of I4267: signal is true;
	signal I4270: std_logic; attribute dont_touch of I4270: signal is true;
	signal I4273: std_logic; attribute dont_touch of I4273: signal is true;
	signal I4276: std_logic; attribute dont_touch of I4276: signal is true;
	signal I4279: std_logic; attribute dont_touch of I4279: signal is true;
	signal I4282: std_logic; attribute dont_touch of I4282: signal is true;
	signal I4285: std_logic; attribute dont_touch of I4285: signal is true;
	signal I4288: std_logic; attribute dont_touch of I4288: signal is true;
	signal I4291: std_logic; attribute dont_touch of I4291: signal is true;
	signal I4294: std_logic; attribute dont_touch of I4294: signal is true;
	signal I4297: std_logic; attribute dont_touch of I4297: signal is true;
	signal I4300: std_logic; attribute dont_touch of I4300: signal is true;
	signal I4303: std_logic; attribute dont_touch of I4303: signal is true;
	signal I4306: std_logic; attribute dont_touch of I4306: signal is true;
	signal I4309: std_logic; attribute dont_touch of I4309: signal is true;
	signal I4312: std_logic; attribute dont_touch of I4312: signal is true;
	signal I4315: std_logic; attribute dont_touch of I4315: signal is true;
	signal I4318: std_logic; attribute dont_touch of I4318: signal is true;
	signal I4321: std_logic; attribute dont_touch of I4321: signal is true;
	signal I4324: std_logic; attribute dont_touch of I4324: signal is true;
	signal I4327: std_logic; attribute dont_touch of I4327: signal is true;
	signal I4331: std_logic; attribute dont_touch of I4331: signal is true;
	signal I4334: std_logic; attribute dont_touch of I4334: signal is true;
	signal I4337: std_logic; attribute dont_touch of I4337: signal is true;
	signal I4340: std_logic; attribute dont_touch of I4340: signal is true;
	signal I4343: std_logic; attribute dont_touch of I4343: signal is true;
	signal I4347: std_logic; attribute dont_touch of I4347: signal is true;
	signal I4351: std_logic; attribute dont_touch of I4351: signal is true;
	signal I4354: std_logic; attribute dont_touch of I4354: signal is true;
	signal I4358: std_logic; attribute dont_touch of I4358: signal is true;
	signal I4362: std_logic; attribute dont_touch of I4362: signal is true;
	signal I4366: std_logic; attribute dont_touch of I4366: signal is true;
	signal I4371: std_logic; attribute dont_touch of I4371: signal is true;
	signal I4375: std_logic; attribute dont_touch of I4375: signal is true;
	signal I4382: std_logic; attribute dont_touch of I4382: signal is true;
	signal I4391: std_logic; attribute dont_touch of I4391: signal is true;
	signal I4398: std_logic; attribute dont_touch of I4398: signal is true;
	signal I4402: std_logic; attribute dont_touch of I4402: signal is true;
	signal I4410: std_logic; attribute dont_touch of I4410: signal is true;
	signal I4414: std_logic; attribute dont_touch of I4414: signal is true;
	signal I4420: std_logic; attribute dont_touch of I4420: signal is true;
	signal I4424: std_logic; attribute dont_touch of I4424: signal is true;
	signal I4429: std_logic; attribute dont_touch of I4429: signal is true;
	signal I4433: std_logic; attribute dont_touch of I4433: signal is true;
	signal I4437: std_logic; attribute dont_touch of I4437: signal is true;
	signal I4441: std_logic; attribute dont_touch of I4441: signal is true;
	signal I4444: std_logic; attribute dont_touch of I4444: signal is true;
	signal I4445: std_logic; attribute dont_touch of I4445: signal is true;
	signal I4446: std_logic; attribute dont_touch of I4446: signal is true;
	signal I4452: std_logic; attribute dont_touch of I4452: signal is true;
	signal I4455: std_logic; attribute dont_touch of I4455: signal is true;
	signal I4459: std_logic; attribute dont_touch of I4459: signal is true;
	signal I4462: std_logic; attribute dont_touch of I4462: signal is true;
	signal I4465: std_logic; attribute dont_touch of I4465: signal is true;
	signal I4468: std_logic; attribute dont_touch of I4468: signal is true;
	signal I4471: std_logic; attribute dont_touch of I4471: signal is true;
	signal I4474: std_logic; attribute dont_touch of I4474: signal is true;
	signal I4477: std_logic; attribute dont_touch of I4477: signal is true;
	signal I4480: std_logic; attribute dont_touch of I4480: signal is true;
	signal I4483: std_logic; attribute dont_touch of I4483: signal is true;
	signal I4486: std_logic; attribute dont_touch of I4486: signal is true;
	signal I4489: std_logic; attribute dont_touch of I4489: signal is true;
	signal I4492: std_logic; attribute dont_touch of I4492: signal is true;
	signal I4495: std_logic; attribute dont_touch of I4495: signal is true;
	signal I4498: std_logic; attribute dont_touch of I4498: signal is true;
	signal I4501: std_logic; attribute dont_touch of I4501: signal is true;
	signal I4504: std_logic; attribute dont_touch of I4504: signal is true;
	signal I4507: std_logic; attribute dont_touch of I4507: signal is true;
	signal I4510: std_logic; attribute dont_touch of I4510: signal is true;
	signal I4513: std_logic; attribute dont_touch of I4513: signal is true;
	signal I4516: std_logic; attribute dont_touch of I4516: signal is true;
	signal I4519: std_logic; attribute dont_touch of I4519: signal is true;
	signal I4522: std_logic; attribute dont_touch of I4522: signal is true;
	signal I4526: std_logic; attribute dont_touch of I4526: signal is true;
	signal I4527: std_logic; attribute dont_touch of I4527: signal is true;
	signal I4528: std_logic; attribute dont_touch of I4528: signal is true;
	signal I4534: std_logic; attribute dont_touch of I4534: signal is true;
	signal I4537: std_logic; attribute dont_touch of I4537: signal is true;
	signal I4545: std_logic; attribute dont_touch of I4545: signal is true;
	signal I4546: std_logic; attribute dont_touch of I4546: signal is true;
	signal I4547: std_logic; attribute dont_touch of I4547: signal is true;
	signal I4587: std_logic; attribute dont_touch of I4587: signal is true;
	signal I4593: std_logic; attribute dont_touch of I4593: signal is true;
	signal I4623: std_logic; attribute dont_touch of I4623: signal is true;
	signal I4646: std_logic; attribute dont_touch of I4646: signal is true;
	signal I4664: std_logic; attribute dont_touch of I4664: signal is true;
	signal I4667: std_logic; attribute dont_touch of I4667: signal is true;
	signal I4671: std_logic; attribute dont_touch of I4671: signal is true;
	signal I4678: std_logic; attribute dont_touch of I4678: signal is true;
	signal I4681: std_logic; attribute dont_touch of I4681: signal is true;
	signal I4684: std_logic; attribute dont_touch of I4684: signal is true;
	signal I4688: std_logic; attribute dont_touch of I4688: signal is true;
	signal I4706: std_logic; attribute dont_touch of I4706: signal is true;
	signal I4743: std_logic; attribute dont_touch of I4743: signal is true;
	signal I4752: std_logic; attribute dont_touch of I4752: signal is true;
	signal I4757: std_logic; attribute dont_touch of I4757: signal is true;
	signal I4762: std_logic; attribute dont_touch of I4762: signal is true;
	signal I4777: std_logic; attribute dont_touch of I4777: signal is true;
	signal I4782: std_logic; attribute dont_touch of I4782: signal is true;
	signal I4783: std_logic; attribute dont_touch of I4783: signal is true;
	signal I4784: std_logic; attribute dont_touch of I4784: signal is true;
	signal I4791: std_logic; attribute dont_touch of I4791: signal is true;
	signal I4794: std_logic; attribute dont_touch of I4794: signal is true;
	signal I4799: std_logic; attribute dont_touch of I4799: signal is true;
	signal I4802: std_logic; attribute dont_touch of I4802: signal is true;
	signal I4809: std_logic; attribute dont_touch of I4809: signal is true;
	signal I4821: std_logic; attribute dont_touch of I4821: signal is true;
	signal I4903: std_logic; attribute dont_touch of I4903: signal is true;
	signal I4919: std_logic; attribute dont_touch of I4919: signal is true;
	signal I4920: std_logic; attribute dont_touch of I4920: signal is true;
	signal I4921: std_logic; attribute dont_touch of I4921: signal is true;
	signal I4935: std_logic; attribute dont_touch of I4935: signal is true;
	signal I4939: std_logic; attribute dont_touch of I4939: signal is true;
	signal I4940: std_logic; attribute dont_touch of I4940: signal is true;
	signal I4941: std_logic; attribute dont_touch of I4941: signal is true;
	signal I4955: std_logic; attribute dont_touch of I4955: signal is true;
	signal I4961: std_logic; attribute dont_touch of I4961: signal is true;
	signal I4964: std_logic; attribute dont_touch of I4964: signal is true;
	signal I4976: std_logic; attribute dont_touch of I4976: signal is true;
	signal I4980: std_logic; attribute dont_touch of I4980: signal is true;
	signal I4986: std_logic; attribute dont_touch of I4986: signal is true;
	signal I5002: std_logic; attribute dont_touch of I5002: signal is true;
	signal I5006: std_logic; attribute dont_touch of I5006: signal is true;
	signal I5019: std_logic; attribute dont_touch of I5019: signal is true;
	signal I5023: std_logic; attribute dont_touch of I5023: signal is true;
	signal I5027: std_logic; attribute dont_touch of I5027: signal is true;
	signal I5030: std_logic; attribute dont_touch of I5030: signal is true;
	signal I5033: std_logic; attribute dont_touch of I5033: signal is true;
	signal I5037: std_logic; attribute dont_touch of I5037: signal is true;
	signal I5040: std_logic; attribute dont_touch of I5040: signal is true;
	signal I5043: std_logic; attribute dont_touch of I5043: signal is true;
	signal I5050: std_logic; attribute dont_touch of I5050: signal is true;
	signal I5053: std_logic; attribute dont_touch of I5053: signal is true;
	signal I5056: std_logic; attribute dont_touch of I5056: signal is true;
	signal I5059: std_logic; attribute dont_touch of I5059: signal is true;
	signal I5065: std_logic; attribute dont_touch of I5065: signal is true;
	signal I5068: std_logic; attribute dont_touch of I5068: signal is true;
	signal I5071: std_logic; attribute dont_touch of I5071: signal is true;
	signal I5078: std_logic; attribute dont_touch of I5078: signal is true;
	signal I5081: std_logic; attribute dont_touch of I5081: signal is true;
	signal I5084: std_logic; attribute dont_touch of I5084: signal is true;
	signal I5091: std_logic; attribute dont_touch of I5091: signal is true;
	signal I5094: std_logic; attribute dont_touch of I5094: signal is true;
	signal I5103: std_logic; attribute dont_touch of I5103: signal is true;
	signal I5106: std_logic; attribute dont_touch of I5106: signal is true;
	signal I5109: std_logic; attribute dont_touch of I5109: signal is true;
	signal I5116: std_logic; attribute dont_touch of I5116: signal is true;
	signal I5119: std_logic; attribute dont_touch of I5119: signal is true;
	signal I5124: std_logic; attribute dont_touch of I5124: signal is true;
	signal I5148: std_logic; attribute dont_touch of I5148: signal is true;
	signal I5153: std_logic; attribute dont_touch of I5153: signal is true;
	signal I5157: std_logic; attribute dont_touch of I5157: signal is true;
	signal I5169: std_logic; attribute dont_touch of I5169: signal is true;
	signal I5177: std_logic; attribute dont_touch of I5177: signal is true;
	signal I5182: std_logic; attribute dont_touch of I5182: signal is true;
	signal I5187: std_logic; attribute dont_touch of I5187: signal is true;
	signal I5188: std_logic; attribute dont_touch of I5188: signal is true;
	signal I5189: std_logic; attribute dont_touch of I5189: signal is true;
	signal I5195: std_logic; attribute dont_touch of I5195: signal is true;
	signal I5196: std_logic; attribute dont_touch of I5196: signal is true;
	signal I5197: std_logic; attribute dont_touch of I5197: signal is true;
	signal I5204: std_logic; attribute dont_touch of I5204: signal is true;
	signal I5207: std_logic; attribute dont_touch of I5207: signal is true;
	signal I5208: std_logic; attribute dont_touch of I5208: signal is true;
	signal I5209: std_logic; attribute dont_touch of I5209: signal is true;
	signal I5214: std_logic; attribute dont_touch of I5214: signal is true;
	signal I5217: std_logic; attribute dont_touch of I5217: signal is true;
	signal I5223: std_logic; attribute dont_touch of I5223: signal is true;
	signal I5226: std_logic; attribute dont_touch of I5226: signal is true;
	signal I5227: std_logic; attribute dont_touch of I5227: signal is true;
	signal I5228: std_logic; attribute dont_touch of I5228: signal is true;
	signal I5233: std_logic; attribute dont_touch of I5233: signal is true;
	signal I5236: std_logic; attribute dont_touch of I5236: signal is true;
	signal I5242: std_logic; attribute dont_touch of I5242: signal is true;
	signal I5243: std_logic; attribute dont_touch of I5243: signal is true;
	signal I5244: std_logic; attribute dont_touch of I5244: signal is true;
	signal I5249: std_logic; attribute dont_touch of I5249: signal is true;
	signal I5252: std_logic; attribute dont_touch of I5252: signal is true;
	signal I5257: std_logic; attribute dont_touch of I5257: signal is true;
	signal I5258: std_logic; attribute dont_touch of I5258: signal is true;
	signal I5259: std_logic; attribute dont_touch of I5259: signal is true;
	signal I5264: std_logic; attribute dont_touch of I5264: signal is true;
	signal I5269: std_logic; attribute dont_touch of I5269: signal is true;
	signal I5270: std_logic; attribute dont_touch of I5270: signal is true;
	signal I5271: std_logic; attribute dont_touch of I5271: signal is true;
	signal I5292: std_logic; attribute dont_touch of I5292: signal is true;
	signal I5293: std_logic; attribute dont_touch of I5293: signal is true;
	signal I5294: std_logic; attribute dont_touch of I5294: signal is true;
	signal I5300: std_logic; attribute dont_touch of I5300: signal is true;
	signal I5301: std_logic; attribute dont_touch of I5301: signal is true;
	signal I5302: std_logic; attribute dont_touch of I5302: signal is true;
	signal I5307: std_logic; attribute dont_touch of I5307: signal is true;
	signal I5308: std_logic; attribute dont_touch of I5308: signal is true;
	signal I5309: std_logic; attribute dont_touch of I5309: signal is true;
	signal I5316: std_logic; attribute dont_touch of I5316: signal is true;
	signal I5320: std_logic; attribute dont_touch of I5320: signal is true;
	signal I5324: std_logic; attribute dont_touch of I5324: signal is true;
	signal I5328: std_logic; attribute dont_touch of I5328: signal is true;
	signal I5333: std_logic; attribute dont_touch of I5333: signal is true;
	signal I5337: std_logic; attribute dont_touch of I5337: signal is true;
	signal I5343: std_logic; attribute dont_touch of I5343: signal is true;
	signal I5351: std_logic; attribute dont_touch of I5351: signal is true;
	signal I5352: std_logic; attribute dont_touch of I5352: signal is true;
	signal I5359: std_logic; attribute dont_touch of I5359: signal is true;
	signal I5360: std_logic; attribute dont_touch of I5360: signal is true;
	signal I5376: std_logic; attribute dont_touch of I5376: signal is true;
	signal I5379: std_logic; attribute dont_touch of I5379: signal is true;
	signal I5382: std_logic; attribute dont_touch of I5382: signal is true;
	signal I5385: std_logic; attribute dont_touch of I5385: signal is true;
	signal I5388: std_logic; attribute dont_touch of I5388: signal is true;
	signal I5391: std_logic; attribute dont_touch of I5391: signal is true;
	signal I5394: std_logic; attribute dont_touch of I5394: signal is true;
	signal I5397: std_logic; attribute dont_touch of I5397: signal is true;
	signal I5400: std_logic; attribute dont_touch of I5400: signal is true;
	signal I5403: std_logic; attribute dont_touch of I5403: signal is true;
	signal I5406: std_logic; attribute dont_touch of I5406: signal is true;
	signal I5409: std_logic; attribute dont_touch of I5409: signal is true;
	signal I5412: std_logic; attribute dont_touch of I5412: signal is true;
	signal I5415: std_logic; attribute dont_touch of I5415: signal is true;
	signal I5418: std_logic; attribute dont_touch of I5418: signal is true;
	signal I5421: std_logic; attribute dont_touch of I5421: signal is true;
	signal I5424: std_logic; attribute dont_touch of I5424: signal is true;
	signal I5427: std_logic; attribute dont_touch of I5427: signal is true;
	signal I5430: std_logic; attribute dont_touch of I5430: signal is true;
	signal I5433: std_logic; attribute dont_touch of I5433: signal is true;
	signal I5436: std_logic; attribute dont_touch of I5436: signal is true;
	signal I5439: std_logic; attribute dont_touch of I5439: signal is true;
	signal I5442: std_logic; attribute dont_touch of I5442: signal is true;
	signal I5445: std_logic; attribute dont_touch of I5445: signal is true;
	signal I5448: std_logic; attribute dont_touch of I5448: signal is true;
	signal I5451: std_logic; attribute dont_touch of I5451: signal is true;
	signal I5454: std_logic; attribute dont_touch of I5454: signal is true;
	signal I5457: std_logic; attribute dont_touch of I5457: signal is true;
	signal I5460: std_logic; attribute dont_touch of I5460: signal is true;
	signal I5463: std_logic; attribute dont_touch of I5463: signal is true;
	signal I5466: std_logic; attribute dont_touch of I5466: signal is true;
	signal I5469: std_logic; attribute dont_touch of I5469: signal is true;
	signal I5472: std_logic; attribute dont_touch of I5472: signal is true;
	signal I5475: std_logic; attribute dont_touch of I5475: signal is true;
	signal I5478: std_logic; attribute dont_touch of I5478: signal is true;
	signal I5481: std_logic; attribute dont_touch of I5481: signal is true;
	signal I5484: std_logic; attribute dont_touch of I5484: signal is true;
	signal I5487: std_logic; attribute dont_touch of I5487: signal is true;
	signal I5490: std_logic; attribute dont_touch of I5490: signal is true;
	signal I5493: std_logic; attribute dont_touch of I5493: signal is true;
	signal I5496: std_logic; attribute dont_touch of I5496: signal is true;
	signal I5499: std_logic; attribute dont_touch of I5499: signal is true;
	signal I5502: std_logic; attribute dont_touch of I5502: signal is true;
	signal I5505: std_logic; attribute dont_touch of I5505: signal is true;
	signal I5508: std_logic; attribute dont_touch of I5508: signal is true;
	signal I5511: std_logic; attribute dont_touch of I5511: signal is true;
	signal I5514: std_logic; attribute dont_touch of I5514: signal is true;
	signal I5517: std_logic; attribute dont_touch of I5517: signal is true;
	signal I5520: std_logic; attribute dont_touch of I5520: signal is true;
	signal I5523: std_logic; attribute dont_touch of I5523: signal is true;
	signal I5526: std_logic; attribute dont_touch of I5526: signal is true;
	signal I5529: std_logic; attribute dont_touch of I5529: signal is true;
	signal I5532: std_logic; attribute dont_touch of I5532: signal is true;
	signal I5535: std_logic; attribute dont_touch of I5535: signal is true;
	signal I5536: std_logic; attribute dont_touch of I5536: signal is true;
	signal I5537: std_logic; attribute dont_touch of I5537: signal is true;
	signal I5542: std_logic; attribute dont_touch of I5542: signal is true;
	signal I5545: std_logic; attribute dont_touch of I5545: signal is true;
	signal I5548: std_logic; attribute dont_touch of I5548: signal is true;
	signal I5551: std_logic; attribute dont_touch of I5551: signal is true;
	signal I5556: std_logic; attribute dont_touch of I5556: signal is true;
	signal I5562: std_logic; attribute dont_touch of I5562: signal is true;
	signal I5568: std_logic; attribute dont_touch of I5568: signal is true;
	signal I5577: std_logic; attribute dont_touch of I5577: signal is true;
	signal I5591: std_logic; attribute dont_touch of I5591: signal is true;
	signal I5594: std_logic; attribute dont_touch of I5594: signal is true;
	signal I5597: std_logic; attribute dont_touch of I5597: signal is true;
	signal I5600: std_logic; attribute dont_touch of I5600: signal is true;
	signal I5603: std_logic; attribute dont_touch of I5603: signal is true;
	signal I5606: std_logic; attribute dont_touch of I5606: signal is true;
	signal I5609: std_logic; attribute dont_touch of I5609: signal is true;
	signal I5612: std_logic; attribute dont_touch of I5612: signal is true;
	signal I5615: std_logic; attribute dont_touch of I5615: signal is true;
	signal I5618: std_logic; attribute dont_touch of I5618: signal is true;
	signal I5622: std_logic; attribute dont_touch of I5622: signal is true;
	signal I5626: std_logic; attribute dont_touch of I5626: signal is true;
	signal I5630: std_logic; attribute dont_touch of I5630: signal is true;
	signal I5633: std_logic; attribute dont_touch of I5633: signal is true;
	signal I5637: std_logic; attribute dont_touch of I5637: signal is true;
	signal I5640: std_logic; attribute dont_touch of I5640: signal is true;
	signal I5644: std_logic; attribute dont_touch of I5644: signal is true;
	signal I5647: std_logic; attribute dont_touch of I5647: signal is true;
	signal I5648: std_logic; attribute dont_touch of I5648: signal is true;
	signal I5649: std_logic; attribute dont_touch of I5649: signal is true;
	signal I5654: std_logic; attribute dont_touch of I5654: signal is true;
	signal I5657: std_logic; attribute dont_touch of I5657: signal is true;
	signal I5658: std_logic; attribute dont_touch of I5658: signal is true;
	signal I5659: std_logic; attribute dont_touch of I5659: signal is true;
	signal I5668: std_logic; attribute dont_touch of I5668: signal is true;
	signal I5674: std_logic; attribute dont_touch of I5674: signal is true;
	signal I5686: std_logic; attribute dont_touch of I5686: signal is true;
	signal I5692: std_logic; attribute dont_touch of I5692: signal is true;
	signal I5696: std_logic; attribute dont_touch of I5696: signal is true;
	signal I5699: std_logic; attribute dont_touch of I5699: signal is true;
	signal I5702: std_logic; attribute dont_touch of I5702: signal is true;
	signal I5705: std_logic; attribute dont_touch of I5705: signal is true;
	signal I5708: std_logic; attribute dont_touch of I5708: signal is true;
	signal I5713: std_logic; attribute dont_touch of I5713: signal is true;
	signal I5716: std_logic; attribute dont_touch of I5716: signal is true;
	signal I5720: std_logic; attribute dont_touch of I5720: signal is true;
	signal I5723: std_logic; attribute dont_touch of I5723: signal is true;
	signal I5728: std_logic; attribute dont_touch of I5728: signal is true;
	signal I5731: std_logic; attribute dont_touch of I5731: signal is true;
	signal I5736: std_logic; attribute dont_touch of I5736: signal is true;
	signal I5739: std_logic; attribute dont_touch of I5739: signal is true;
	signal I5743: std_logic; attribute dont_touch of I5743: signal is true;
	signal I5746: std_logic; attribute dont_touch of I5746: signal is true;
	signal I5750: std_logic; attribute dont_touch of I5750: signal is true;
	signal I5753: std_logic; attribute dont_touch of I5753: signal is true;
	signal I5756: std_logic; attribute dont_touch of I5756: signal is true;
	signal I5759: std_logic; attribute dont_touch of I5759: signal is true;
	signal I5760: std_logic; attribute dont_touch of I5760: signal is true;
	signal I5761: std_logic; attribute dont_touch of I5761: signal is true;
	signal I5766: std_logic; attribute dont_touch of I5766: signal is true;
	signal I5767: std_logic; attribute dont_touch of I5767: signal is true;
	signal I5768: std_logic; attribute dont_touch of I5768: signal is true;
	signal I5774: std_logic; attribute dont_touch of I5774: signal is true;
	signal I5777: std_logic; attribute dont_touch of I5777: signal is true;
	signal I5782: std_logic; attribute dont_touch of I5782: signal is true;
	signal I5783: std_logic; attribute dont_touch of I5783: signal is true;
	signal I5784: std_logic; attribute dont_touch of I5784: signal is true;
	signal I5790: std_logic; attribute dont_touch of I5790: signal is true;
	signal I5793: std_logic; attribute dont_touch of I5793: signal is true;
	signal I5825: std_logic; attribute dont_touch of I5825: signal is true;
	signal I5831: std_logic; attribute dont_touch of I5831: signal is true;
	signal I5837: std_logic; attribute dont_touch of I5837: signal is true;
	signal I5840: std_logic; attribute dont_touch of I5840: signal is true;
	signal I5843: std_logic; attribute dont_touch of I5843: signal is true;
	signal I5848: std_logic; attribute dont_touch of I5848: signal is true;
	signal I5851: std_logic; attribute dont_touch of I5851: signal is true;
	signal I5854: std_logic; attribute dont_touch of I5854: signal is true;
	signal I5857: std_logic; attribute dont_touch of I5857: signal is true;
	signal I5862: std_logic; attribute dont_touch of I5862: signal is true;
	signal I5865: std_logic; attribute dont_touch of I5865: signal is true;
	signal I5868: std_logic; attribute dont_touch of I5868: signal is true;
	signal I5871: std_logic; attribute dont_touch of I5871: signal is true;
	signal I5876: std_logic; attribute dont_touch of I5876: signal is true;
	signal I5879: std_logic; attribute dont_touch of I5879: signal is true;
	signal I5882: std_logic; attribute dont_touch of I5882: signal is true;
	signal I5885: std_logic; attribute dont_touch of I5885: signal is true;
	signal I5890: std_logic; attribute dont_touch of I5890: signal is true;
	signal I5893: std_logic; attribute dont_touch of I5893: signal is true;
	signal I5896: std_logic; attribute dont_touch of I5896: signal is true;
	signal I5899: std_logic; attribute dont_touch of I5899: signal is true;
	signal I5904: std_logic; attribute dont_touch of I5904: signal is true;
	signal I5907: std_logic; attribute dont_touch of I5907: signal is true;
	signal I5910: std_logic; attribute dont_touch of I5910: signal is true;
	signal I5913: std_logic; attribute dont_touch of I5913: signal is true;
	signal I5920: std_logic; attribute dont_touch of I5920: signal is true;
	signal I5923: std_logic; attribute dont_touch of I5923: signal is true;
	signal I5926: std_logic; attribute dont_touch of I5926: signal is true;
	signal I5929: std_logic; attribute dont_touch of I5929: signal is true;
	signal I5933: std_logic; attribute dont_touch of I5933: signal is true;
	signal I5938: std_logic; attribute dont_touch of I5938: signal is true;
	signal I5944: std_logic; attribute dont_touch of I5944: signal is true;
	signal I5948: std_logic; attribute dont_touch of I5948: signal is true;
	signal I5952: std_logic; attribute dont_touch of I5952: signal is true;
	signal I5977: std_logic; attribute dont_touch of I5977: signal is true;
	signal I5987: std_logic; attribute dont_touch of I5987: signal is true;
	signal I5991: std_logic; attribute dont_touch of I5991: signal is true;
	signal I5998: std_logic; attribute dont_touch of I5998: signal is true;
	signal I6001: std_logic; attribute dont_touch of I6001: signal is true;
	signal I6004: std_logic; attribute dont_touch of I6004: signal is true;
	signal I6008: std_logic; attribute dont_touch of I6008: signal is true;
	signal I6012: std_logic; attribute dont_touch of I6012: signal is true;
	signal I6015: std_logic; attribute dont_touch of I6015: signal is true;
	signal I6020: std_logic; attribute dont_touch of I6020: signal is true;
	signal I6023: std_logic; attribute dont_touch of I6023: signal is true;
	signal I6026: std_logic; attribute dont_touch of I6026: signal is true;
	signal I6027: std_logic; attribute dont_touch of I6027: signal is true;
	signal I6028: std_logic; attribute dont_touch of I6028: signal is true;
	signal I6033: std_logic; attribute dont_touch of I6033: signal is true;
	signal I6036: std_logic; attribute dont_touch of I6036: signal is true;
	signal I6039: std_logic; attribute dont_touch of I6039: signal is true;
	signal I6042: std_logic; attribute dont_touch of I6042: signal is true;
	signal I6045: std_logic; attribute dont_touch of I6045: signal is true;
	signal I6048: std_logic; attribute dont_touch of I6048: signal is true;
	signal I6051: std_logic; attribute dont_touch of I6051: signal is true;
	signal I6054: std_logic; attribute dont_touch of I6054: signal is true;
	signal I6057: std_logic; attribute dont_touch of I6057: signal is true;
	signal I6060: std_logic; attribute dont_touch of I6060: signal is true;
	signal I6063: std_logic; attribute dont_touch of I6063: signal is true;
	signal I6066: std_logic; attribute dont_touch of I6066: signal is true;
	signal I6069: std_logic; attribute dont_touch of I6069: signal is true;
	signal I6072: std_logic; attribute dont_touch of I6072: signal is true;
	signal I6075: std_logic; attribute dont_touch of I6075: signal is true;
	signal I6078: std_logic; attribute dont_touch of I6078: signal is true;
	signal I6081: std_logic; attribute dont_touch of I6081: signal is true;
	signal I6084: std_logic; attribute dont_touch of I6084: signal is true;
	signal I6087: std_logic; attribute dont_touch of I6087: signal is true;
	signal I6090: std_logic; attribute dont_touch of I6090: signal is true;
	signal I6093: std_logic; attribute dont_touch of I6093: signal is true;
	signal I6096: std_logic; attribute dont_touch of I6096: signal is true;
	signal I6099: std_logic; attribute dont_touch of I6099: signal is true;
	signal I6102: std_logic; attribute dont_touch of I6102: signal is true;
	signal I6105: std_logic; attribute dont_touch of I6105: signal is true;
	signal I6108: std_logic; attribute dont_touch of I6108: signal is true;
	signal I6111: std_logic; attribute dont_touch of I6111: signal is true;
	signal I6114: std_logic; attribute dont_touch of I6114: signal is true;
	signal I6118: std_logic; attribute dont_touch of I6118: signal is true;
	signal I6126: std_logic; attribute dont_touch of I6126: signal is true;
	signal I6132: std_logic; attribute dont_touch of I6132: signal is true;
	signal I6139: std_logic; attribute dont_touch of I6139: signal is true;
	signal I6143: std_logic; attribute dont_touch of I6143: signal is true;
	signal I6170: std_logic; attribute dont_touch of I6170: signal is true;
	signal I6175: std_logic; attribute dont_touch of I6175: signal is true;
	signal I6176: std_logic; attribute dont_touch of I6176: signal is true;
	signal I6177: std_logic; attribute dont_touch of I6177: signal is true;
	signal I6182: std_logic; attribute dont_touch of I6182: signal is true;
	signal I6185: std_logic; attribute dont_touch of I6185: signal is true;
	signal I6186: std_logic; attribute dont_touch of I6186: signal is true;
	signal I6187: std_logic; attribute dont_touch of I6187: signal is true;
	signal I6194: std_logic; attribute dont_touch of I6194: signal is true;
	signal I6195: std_logic; attribute dont_touch of I6195: signal is true;
	signal I6196: std_logic; attribute dont_touch of I6196: signal is true;
	signal I6231: std_logic; attribute dont_touch of I6231: signal is true;
	signal I6244: std_logic; attribute dont_touch of I6244: signal is true;
	signal I6247: std_logic; attribute dont_touch of I6247: signal is true;
	signal I6250: std_logic; attribute dont_touch of I6250: signal is true;
	signal I6253: std_logic; attribute dont_touch of I6253: signal is true;
	signal I6269: std_logic; attribute dont_touch of I6269: signal is true;
	signal I6280: std_logic; attribute dont_touch of I6280: signal is true;
	signal I6283: std_logic; attribute dont_touch of I6283: signal is true;
	signal I6289: std_logic; attribute dont_touch of I6289: signal is true;
	signal I6292: std_logic; attribute dont_touch of I6292: signal is true;
	signal I6296: std_logic; attribute dont_touch of I6296: signal is true;
	signal I6299: std_logic; attribute dont_touch of I6299: signal is true;
	signal I6302: std_logic; attribute dont_touch of I6302: signal is true;
	signal I6305: std_logic; attribute dont_touch of I6305: signal is true;
	signal I6308: std_logic; attribute dont_touch of I6308: signal is true;
	signal I6311: std_logic; attribute dont_touch of I6311: signal is true;
	signal I6315: std_logic; attribute dont_touch of I6315: signal is true;
	signal I6318: std_logic; attribute dont_touch of I6318: signal is true;
	signal I6321: std_logic; attribute dont_touch of I6321: signal is true;
	signal I6324: std_logic; attribute dont_touch of I6324: signal is true;
	signal I6327: std_logic; attribute dont_touch of I6327: signal is true;
	signal I6330: std_logic; attribute dont_touch of I6330: signal is true;
	signal I6334: std_logic; attribute dont_touch of I6334: signal is true;
	signal I6337: std_logic; attribute dont_touch of I6337: signal is true;
	signal I6340: std_logic; attribute dont_touch of I6340: signal is true;
	signal I6343: std_logic; attribute dont_touch of I6343: signal is true;
	signal I6346: std_logic; attribute dont_touch of I6346: signal is true;
	signal I6349: std_logic; attribute dont_touch of I6349: signal is true;
	signal I6352: std_logic; attribute dont_touch of I6352: signal is true;
	signal I6355: std_logic; attribute dont_touch of I6355: signal is true;
	signal I6359: std_logic; attribute dont_touch of I6359: signal is true;
	signal I6362: std_logic; attribute dont_touch of I6362: signal is true;
	signal I6366: std_logic; attribute dont_touch of I6366: signal is true;
	signal I6371: std_logic; attribute dont_touch of I6371: signal is true;
	signal I6377: std_logic; attribute dont_touch of I6377: signal is true;
	signal I6382: std_logic; attribute dont_touch of I6382: signal is true;
	signal I6386: std_logic; attribute dont_touch of I6386: signal is true;
	signal I6390: std_logic; attribute dont_touch of I6390: signal is true;
	signal I6391: std_logic; attribute dont_touch of I6391: signal is true;
	signal I6392: std_logic; attribute dont_touch of I6392: signal is true;
	signal I6397: std_logic; attribute dont_touch of I6397: signal is true;
	signal I6400: std_logic; attribute dont_touch of I6400: signal is true;
	signal I6403: std_logic; attribute dont_touch of I6403: signal is true;
	signal I6406: std_logic; attribute dont_touch of I6406: signal is true;
	signal I6410: std_logic; attribute dont_touch of I6410: signal is true;
	signal I6414: std_logic; attribute dont_touch of I6414: signal is true;
	signal I6417: std_logic; attribute dont_touch of I6417: signal is true;
	signal I6420: std_logic; attribute dont_touch of I6420: signal is true;
	signal I6425: std_logic; attribute dont_touch of I6425: signal is true;
	signal I6430: std_logic; attribute dont_touch of I6430: signal is true;
	signal I6434: std_logic; attribute dont_touch of I6434: signal is true;
	signal I6437: std_logic; attribute dont_touch of I6437: signal is true;
	signal I6441: std_logic; attribute dont_touch of I6441: signal is true;
	signal I6444: std_logic; attribute dont_touch of I6444: signal is true;
	signal I6448: std_logic; attribute dont_touch of I6448: signal is true;
	signal I6452: std_logic; attribute dont_touch of I6452: signal is true;
	signal I6456: std_logic; attribute dont_touch of I6456: signal is true;
	signal I6464: std_logic; attribute dont_touch of I6464: signal is true;
	signal I6470: std_logic; attribute dont_touch of I6470: signal is true;
	signal I6473: std_logic; attribute dont_touch of I6473: signal is true;
	signal I6474: std_logic; attribute dont_touch of I6474: signal is true;
	signal I6475: std_logic; attribute dont_touch of I6475: signal is true;
	signal I6485: std_logic; attribute dont_touch of I6485: signal is true;
	signal I6488: std_logic; attribute dont_touch of I6488: signal is true;
	signal I6495: std_logic; attribute dont_touch of I6495: signal is true;
	signal I6499: std_logic; attribute dont_touch of I6499: signal is true;
	signal I6500: std_logic; attribute dont_touch of I6500: signal is true;
	signal I6501: std_logic; attribute dont_touch of I6501: signal is true;
	signal I6507: std_logic; attribute dont_touch of I6507: signal is true;
	signal I6525: std_logic; attribute dont_touch of I6525: signal is true;
	signal I6528: std_logic; attribute dont_touch of I6528: signal is true;
	signal I6531: std_logic; attribute dont_touch of I6531: signal is true;
	signal I6534: std_logic; attribute dont_touch of I6534: signal is true;
	signal I6537: std_logic; attribute dont_touch of I6537: signal is true;
	signal I6540: std_logic; attribute dont_touch of I6540: signal is true;
	signal I6543: std_logic; attribute dont_touch of I6543: signal is true;
	signal I6546: std_logic; attribute dont_touch of I6546: signal is true;
	signal I6549: std_logic; attribute dont_touch of I6549: signal is true;
	signal I6552: std_logic; attribute dont_touch of I6552: signal is true;
	signal I6555: std_logic; attribute dont_touch of I6555: signal is true;
	signal I6558: std_logic; attribute dont_touch of I6558: signal is true;
	signal I6561: std_logic; attribute dont_touch of I6561: signal is true;
	signal I6564: std_logic; attribute dont_touch of I6564: signal is true;
	signal I6567: std_logic; attribute dont_touch of I6567: signal is true;
	signal I6570: std_logic; attribute dont_touch of I6570: signal is true;
	signal I6573: std_logic; attribute dont_touch of I6573: signal is true;
	signal I6576: std_logic; attribute dont_touch of I6576: signal is true;
	signal I6579: std_logic; attribute dont_touch of I6579: signal is true;
	signal I6582: std_logic; attribute dont_touch of I6582: signal is true;
	signal I6587: std_logic; attribute dont_touch of I6587: signal is true;
	signal I6599: std_logic; attribute dont_touch of I6599: signal is true;
	signal I6607: std_logic; attribute dont_touch of I6607: signal is true;
	signal I6612: std_logic; attribute dont_touch of I6612: signal is true;
	signal I6615: std_logic; attribute dont_touch of I6615: signal is true;
	signal I6621: std_logic; attribute dont_touch of I6621: signal is true;
	signal I6625: std_logic; attribute dont_touch of I6625: signal is true;
	signal I6630: std_logic; attribute dont_touch of I6630: signal is true;
	signal I6635: std_logic; attribute dont_touch of I6635: signal is true;
	signal I6646: std_logic; attribute dont_touch of I6646: signal is true;
	signal I6649: std_logic; attribute dont_touch of I6649: signal is true;
	signal I6659: std_logic; attribute dont_touch of I6659: signal is true;
	signal I6660: std_logic; attribute dont_touch of I6660: signal is true;
	signal I6661: std_logic; attribute dont_touch of I6661: signal is true;
	signal I6666: std_logic; attribute dont_touch of I6666: signal is true;
	signal I6672: std_logic; attribute dont_touch of I6672: signal is true;
	signal I6677: std_logic; attribute dont_touch of I6677: signal is true;
	signal I6680: std_logic; attribute dont_touch of I6680: signal is true;
	signal I6685: std_logic; attribute dont_touch of I6685: signal is true;
	signal I6689: std_logic; attribute dont_touch of I6689: signal is true;
	signal I6692: std_logic; attribute dont_touch of I6692: signal is true;
	signal I6697: std_logic; attribute dont_touch of I6697: signal is true;
	signal I6701: std_logic; attribute dont_touch of I6701: signal is true;
	signal I6706: std_logic; attribute dont_touch of I6706: signal is true;
	signal I6723: std_logic; attribute dont_touch of I6723: signal is true;
	signal I6733: std_logic; attribute dont_touch of I6733: signal is true;
	signal I6737: std_logic; attribute dont_touch of I6737: signal is true;
	signal I6740: std_logic; attribute dont_touch of I6740: signal is true;
	signal I6743: std_logic; attribute dont_touch of I6743: signal is true;
	signal I6744: std_logic; attribute dont_touch of I6744: signal is true;
	signal I6745: std_logic; attribute dont_touch of I6745: signal is true;
	signal I6750: std_logic; attribute dont_touch of I6750: signal is true;
	signal I6753: std_logic; attribute dont_touch of I6753: signal is true;
	signal I6756: std_logic; attribute dont_touch of I6756: signal is true;
	signal I6759: std_logic; attribute dont_touch of I6759: signal is true;
	signal I6763: std_logic; attribute dont_touch of I6763: signal is true;
	signal I6766: std_logic; attribute dont_touch of I6766: signal is true;
	signal I6769: std_logic; attribute dont_touch of I6769: signal is true;
	signal I6772: std_logic; attribute dont_touch of I6772: signal is true;
	signal I6775: std_logic; attribute dont_touch of I6775: signal is true;
	signal I6780: std_logic; attribute dont_touch of I6780: signal is true;
	signal I6783: std_logic; attribute dont_touch of I6783: signal is true;
	signal I6786: std_logic; attribute dont_touch of I6786: signal is true;
	signal I6789: std_logic; attribute dont_touch of I6789: signal is true;
	signal I6792: std_logic; attribute dont_touch of I6792: signal is true;
	signal I6795: std_logic; attribute dont_touch of I6795: signal is true;
	signal I6798: std_logic; attribute dont_touch of I6798: signal is true;
	signal I6801: std_logic; attribute dont_touch of I6801: signal is true;
	signal I6809: std_logic; attribute dont_touch of I6809: signal is true;
	signal I6812: std_logic; attribute dont_touch of I6812: signal is true;
	signal I6816: std_logic; attribute dont_touch of I6816: signal is true;
	signal I6819: std_logic; attribute dont_touch of I6819: signal is true;
	signal I6867: std_logic; attribute dont_touch of I6867: signal is true;
	signal I6874: std_logic; attribute dont_touch of I6874: signal is true;
	signal I6885: std_logic; attribute dont_touch of I6885: signal is true;
	signal I6895: std_logic; attribute dont_touch of I6895: signal is true;
	signal I6918: std_logic; attribute dont_touch of I6918: signal is true;
	signal I6923: std_logic; attribute dont_touch of I6923: signal is true;
	signal I6927: std_logic; attribute dont_touch of I6927: signal is true;
	signal I6930: std_logic; attribute dont_touch of I6930: signal is true;
	signal I6933: std_logic; attribute dont_touch of I6933: signal is true;
	signal I6937: std_logic; attribute dont_touch of I6937: signal is true;
	signal I6942: std_logic; attribute dont_touch of I6942: signal is true;
	signal I6946: std_logic; attribute dont_touch of I6946: signal is true;
	signal I6949: std_logic; attribute dont_touch of I6949: signal is true;
	signal I6952: std_logic; attribute dont_touch of I6952: signal is true;
	signal I6956: std_logic; attribute dont_touch of I6956: signal is true;
	signal I6959: std_logic; attribute dont_touch of I6959: signal is true;
	signal I6962: std_logic; attribute dont_touch of I6962: signal is true;
	signal I6963: std_logic; attribute dont_touch of I6963: signal is true;
	signal I6964: std_logic; attribute dont_touch of I6964: signal is true;
	signal I6972: std_logic; attribute dont_touch of I6972: signal is true;
	signal I6976: std_logic; attribute dont_touch of I6976: signal is true;
	signal I6986: std_logic; attribute dont_touch of I6986: signal is true;
	signal I6989: std_logic; attribute dont_touch of I6989: signal is true;
	signal I6992: std_logic; attribute dont_touch of I6992: signal is true;
	signal I6995: std_logic; attribute dont_touch of I6995: signal is true;
	signal I7002: std_logic; attribute dont_touch of I7002: signal is true;
	signal I7007: std_logic; attribute dont_touch of I7007: signal is true;
	signal I7012: std_logic; attribute dont_touch of I7012: signal is true;
	signal I7029: std_logic; attribute dont_touch of I7029: signal is true;
	signal I7035: std_logic; attribute dont_touch of I7035: signal is true;
	signal I7039: std_logic; attribute dont_touch of I7039: signal is true;
	signal I7042: std_logic; attribute dont_touch of I7042: signal is true;
	signal I7045: std_logic; attribute dont_touch of I7045: signal is true;
	signal I7051: std_logic; attribute dont_touch of I7051: signal is true;
	signal I7055: std_logic; attribute dont_touch of I7055: signal is true;
	signal I7058: std_logic; attribute dont_touch of I7058: signal is true;
	signal I7061: std_logic; attribute dont_touch of I7061: signal is true;
	signal I7065: std_logic; attribute dont_touch of I7065: signal is true;
	signal I7069: std_logic; attribute dont_touch of I7069: signal is true;
	signal I7073: std_logic; attribute dont_touch of I7073: signal is true;
	signal I7077: std_logic; attribute dont_touch of I7077: signal is true;
	signal I7081: std_logic; attribute dont_touch of I7081: signal is true;
	signal I7086: std_logic; attribute dont_touch of I7086: signal is true;
	signal I7091: std_logic; attribute dont_touch of I7091: signal is true;
	signal I7097: std_logic; attribute dont_touch of I7097: signal is true;
	signal I7098: std_logic; attribute dont_touch of I7098: signal is true;
	signal I7099: std_logic; attribute dont_touch of I7099: signal is true;
	signal I7104: std_logic; attribute dont_touch of I7104: signal is true;
	signal I7107: std_logic; attribute dont_touch of I7107: signal is true;
	signal I7110: std_logic; attribute dont_touch of I7110: signal is true;
	signal I7113: std_logic; attribute dont_touch of I7113: signal is true;
	signal I7116: std_logic; attribute dont_touch of I7116: signal is true;
	signal I7119: std_logic; attribute dont_touch of I7119: signal is true;
	signal I7143: std_logic; attribute dont_touch of I7143: signal is true;
	signal I7146: std_logic; attribute dont_touch of I7146: signal is true;
	signal I7150: std_logic; attribute dont_touch of I7150: signal is true;
	signal I7153: std_logic; attribute dont_touch of I7153: signal is true;
	signal I7161: std_logic; attribute dont_touch of I7161: signal is true;
	signal I7164: std_logic; attribute dont_touch of I7164: signal is true;
	signal I7167: std_logic; attribute dont_touch of I7167: signal is true;
	signal I7170: std_logic; attribute dont_touch of I7170: signal is true;
	signal I7173: std_logic; attribute dont_touch of I7173: signal is true;
	signal I7176: std_logic; attribute dont_touch of I7176: signal is true;
	signal I7187: std_logic; attribute dont_touch of I7187: signal is true;
	signal I7190: std_logic; attribute dont_touch of I7190: signal is true;
	signal I7193: std_logic; attribute dont_touch of I7193: signal is true;
	signal I7197: std_logic; attribute dont_touch of I7197: signal is true;
	signal I7208: std_logic; attribute dont_touch of I7208: signal is true;
	signal I7209: std_logic; attribute dont_touch of I7209: signal is true;
	signal I7210: std_logic; attribute dont_touch of I7210: signal is true;
	signal I7216: std_logic; attribute dont_touch of I7216: signal is true;
	signal I7217: std_logic; attribute dont_touch of I7217: signal is true;
	signal I7218: std_logic; attribute dont_touch of I7218: signal is true;
	signal I7223: std_logic; attribute dont_touch of I7223: signal is true;
	signal I7224: std_logic; attribute dont_touch of I7224: signal is true;
	signal I7225: std_logic; attribute dont_touch of I7225: signal is true;
	signal I7230: std_logic; attribute dont_touch of I7230: signal is true;
	signal I7231: std_logic; attribute dont_touch of I7231: signal is true;
	signal I7232: std_logic; attribute dont_touch of I7232: signal is true;
	signal I7237: std_logic; attribute dont_touch of I7237: signal is true;
	signal I7238: std_logic; attribute dont_touch of I7238: signal is true;
	signal I7239: std_logic; attribute dont_touch of I7239: signal is true;
	signal I7244: std_logic; attribute dont_touch of I7244: signal is true;
	signal I7245: std_logic; attribute dont_touch of I7245: signal is true;
	signal I7246: std_logic; attribute dont_touch of I7246: signal is true;
	signal I7251: std_logic; attribute dont_touch of I7251: signal is true;
	signal I7254: std_logic; attribute dont_touch of I7254: signal is true;
	signal I7258: std_logic; attribute dont_touch of I7258: signal is true;
	signal I7261: std_logic; attribute dont_touch of I7261: signal is true;
	signal I7264: std_logic; attribute dont_touch of I7264: signal is true;
	signal I7267: std_logic; attribute dont_touch of I7267: signal is true;
	signal I7270: std_logic; attribute dont_touch of I7270: signal is true;
	signal I7276: std_logic; attribute dont_touch of I7276: signal is true;
	signal I7284: std_logic; attribute dont_touch of I7284: signal is true;
	signal I7295: std_logic; attribute dont_touch of I7295: signal is true;
	signal I7311: std_logic; attribute dont_touch of I7311: signal is true;
	signal I7312: std_logic; attribute dont_touch of I7312: signal is true;
	signal I7313: std_logic; attribute dont_touch of I7313: signal is true;
	signal I7318: std_logic; attribute dont_touch of I7318: signal is true;
	signal I7333: std_logic; attribute dont_touch of I7333: signal is true;
	signal I7336: std_logic; attribute dont_touch of I7336: signal is true;
	signal I7339: std_logic; attribute dont_touch of I7339: signal is true;
	signal I7342: std_logic; attribute dont_touch of I7342: signal is true;
	signal I7346: std_logic; attribute dont_touch of I7346: signal is true;
	signal I7349: std_logic; attribute dont_touch of I7349: signal is true;
	signal I7352: std_logic; attribute dont_touch of I7352: signal is true;
	signal I7355: std_logic; attribute dont_touch of I7355: signal is true;
	signal I7358: std_logic; attribute dont_touch of I7358: signal is true;
	signal I7361: std_logic; attribute dont_touch of I7361: signal is true;
	signal I7372: std_logic; attribute dont_touch of I7372: signal is true;
	signal I7397: std_logic; attribute dont_touch of I7397: signal is true;
	signal I7404: std_logic; attribute dont_touch of I7404: signal is true;
	signal I7432: std_logic; attribute dont_touch of I7432: signal is true;
	signal I7433: std_logic; attribute dont_touch of I7433: signal is true;
	signal I7434: std_logic; attribute dont_touch of I7434: signal is true;
	signal I7439: std_logic; attribute dont_touch of I7439: signal is true;
	signal I7440: std_logic; attribute dont_touch of I7440: signal is true;
	signal I7441: std_logic; attribute dont_touch of I7441: signal is true;
	signal I7451: std_logic; attribute dont_touch of I7451: signal is true;
	signal I7463: std_logic; attribute dont_touch of I7463: signal is true;
	signal I7466: std_logic; attribute dont_touch of I7466: signal is true;
	signal I7469: std_logic; attribute dont_touch of I7469: signal is true;
	signal I7472: std_logic; attribute dont_touch of I7472: signal is true;
	signal I7475: std_logic; attribute dont_touch of I7475: signal is true;
	signal I7478: std_logic; attribute dont_touch of I7478: signal is true;
	signal I7481: std_logic; attribute dont_touch of I7481: signal is true;
	signal I7484: std_logic; attribute dont_touch of I7484: signal is true;
	signal I7487: std_logic; attribute dont_touch of I7487: signal is true;
	signal I7490: std_logic; attribute dont_touch of I7490: signal is true;
	signal I7494: std_logic; attribute dont_touch of I7494: signal is true;
	signal I7497: std_logic; attribute dont_touch of I7497: signal is true;
	signal I7501: std_logic; attribute dont_touch of I7501: signal is true;
	signal I7506: std_logic; attribute dont_touch of I7506: signal is true;
	signal I7509: std_logic; attribute dont_touch of I7509: signal is true;
	signal I7514: std_logic; attribute dont_touch of I7514: signal is true;
	signal I7517: std_logic; attribute dont_touch of I7517: signal is true;
	signal I7520: std_logic; attribute dont_touch of I7520: signal is true;
	signal I7521: std_logic; attribute dont_touch of I7521: signal is true;
	signal I7522: std_logic; attribute dont_touch of I7522: signal is true;
	signal I7527: std_logic; attribute dont_touch of I7527: signal is true;
	signal I7528: std_logic; attribute dont_touch of I7528: signal is true;
	signal I7529: std_logic; attribute dont_touch of I7529: signal is true;
	signal I7534: std_logic; attribute dont_touch of I7534: signal is true;
	signal I7535: std_logic; attribute dont_touch of I7535: signal is true;
	signal I7536: std_logic; attribute dont_touch of I7536: signal is true;
	signal I7541: std_logic; attribute dont_touch of I7541: signal is true;
	signal I7542: std_logic; attribute dont_touch of I7542: signal is true;
	signal I7543: std_logic; attribute dont_touch of I7543: signal is true;
	signal I7548: std_logic; attribute dont_touch of I7548: signal is true;
	signal I7549: std_logic; attribute dont_touch of I7549: signal is true;
	signal I7550: std_logic; attribute dont_touch of I7550: signal is true;
	signal I7555: std_logic; attribute dont_touch of I7555: signal is true;
	signal I7556: std_logic; attribute dont_touch of I7556: signal is true;
	signal I7557: std_logic; attribute dont_touch of I7557: signal is true;
	signal I7562: std_logic; attribute dont_touch of I7562: signal is true;
	signal I7563: std_logic; attribute dont_touch of I7563: signal is true;
	signal I7564: std_logic; attribute dont_touch of I7564: signal is true;
	signal I7569: std_logic; attribute dont_touch of I7569: signal is true;
	signal I7570: std_logic; attribute dont_touch of I7570: signal is true;
	signal I7571: std_logic; attribute dont_touch of I7571: signal is true;
	signal I7576: std_logic; attribute dont_touch of I7576: signal is true;
	signal I7577: std_logic; attribute dont_touch of I7577: signal is true;
	signal I7578: std_logic; attribute dont_touch of I7578: signal is true;
	signal I7583: std_logic; attribute dont_touch of I7583: signal is true;
	signal I7587: std_logic; attribute dont_touch of I7587: signal is true;
	signal I7590: std_logic; attribute dont_touch of I7590: signal is true;
	signal I7593: std_logic; attribute dont_touch of I7593: signal is true;
	signal I7596: std_logic; attribute dont_touch of I7596: signal is true;
	signal I7600: std_logic; attribute dont_touch of I7600: signal is true;
	signal I7604: std_logic; attribute dont_touch of I7604: signal is true;
	signal I7608: std_logic; attribute dont_touch of I7608: signal is true;
	signal I7612: std_logic; attribute dont_touch of I7612: signal is true;
	signal I7634: std_logic; attribute dont_touch of I7634: signal is true;
	signal I7637: std_logic; attribute dont_touch of I7637: signal is true;
	signal I7640: std_logic; attribute dont_touch of I7640: signal is true;
	signal I7643: std_logic; attribute dont_touch of I7643: signal is true;
	signal I7646: std_logic; attribute dont_touch of I7646: signal is true;
	signal I7679: std_logic; attribute dont_touch of I7679: signal is true;
	signal I7683: std_logic; attribute dont_touch of I7683: signal is true;
	signal I7686: std_logic; attribute dont_touch of I7686: signal is true;
	signal I7689: std_logic; attribute dont_touch of I7689: signal is true;
	signal I7692: std_logic; attribute dont_touch of I7692: signal is true;
	signal I7695: std_logic; attribute dont_touch of I7695: signal is true;
	signal I7698: std_logic; attribute dont_touch of I7698: signal is true;
	signal I7701: std_logic; attribute dont_touch of I7701: signal is true;
	signal I7704: std_logic; attribute dont_touch of I7704: signal is true;
	signal I7707: std_logic; attribute dont_touch of I7707: signal is true;
	signal I7796: std_logic; attribute dont_touch of I7796: signal is true;
	signal I7799: std_logic; attribute dont_touch of I7799: signal is true;
	signal I7802: std_logic; attribute dont_touch of I7802: signal is true;
	signal I7805: std_logic; attribute dont_touch of I7805: signal is true;
	signal I7808: std_logic; attribute dont_touch of I7808: signal is true;
	signal I7811: std_logic; attribute dont_touch of I7811: signal is true;
	signal I7814: std_logic; attribute dont_touch of I7814: signal is true;
	signal I7817: std_logic; attribute dont_touch of I7817: signal is true;
	signal I7829: std_logic; attribute dont_touch of I7829: signal is true;
	signal I7832: std_logic; attribute dont_touch of I7832: signal is true;
	signal I7835: std_logic; attribute dont_touch of I7835: signal is true;
	signal I7838: std_logic; attribute dont_touch of I7838: signal is true;
	signal I7852: std_logic; attribute dont_touch of I7852: signal is true;
	signal I7856: std_logic; attribute dont_touch of I7856: signal is true;
	signal I7859: std_logic; attribute dont_touch of I7859: signal is true;
	signal I7865: std_logic; attribute dont_touch of I7865: signal is true;
	signal I7871: std_logic; attribute dont_touch of I7871: signal is true;
	signal I7892: std_logic; attribute dont_touch of I7892: signal is true;
	signal I7906: std_logic; attribute dont_touch of I7906: signal is true;
	signal I7910: std_logic; attribute dont_touch of I7910: signal is true;
	signal I7960: std_logic; attribute dont_touch of I7960: signal is true;
	signal I7963: std_logic; attribute dont_touch of I7963: signal is true;
	signal I7966: std_logic; attribute dont_touch of I7966: signal is true;
	signal I7969: std_logic; attribute dont_touch of I7969: signal is true;
	signal I7970: std_logic; attribute dont_touch of I7970: signal is true;
	signal I7971: std_logic; attribute dont_touch of I7971: signal is true;
	signal I7972: std_logic; attribute dont_touch of I7972: signal is true;
	signal I7978: std_logic; attribute dont_touch of I7978: signal is true;
	signal I7979: std_logic; attribute dont_touch of I7979: signal is true;
	signal I7980: std_logic; attribute dont_touch of I7980: signal is true;
	signal I7981: std_logic; attribute dont_touch of I7981: signal is true;
	signal I7987: std_logic; attribute dont_touch of I7987: signal is true;
	signal I7988: std_logic; attribute dont_touch of I7988: signal is true;
	signal I7989: std_logic; attribute dont_touch of I7989: signal is true;
	signal I7990: std_logic; attribute dont_touch of I7990: signal is true;
	signal I7996: std_logic; attribute dont_touch of I7996: signal is true;
	signal I7999: std_logic; attribute dont_touch of I7999: signal is true;
	signal I8002: std_logic; attribute dont_touch of I8002: signal is true;
	signal I8005: std_logic; attribute dont_touch of I8005: signal is true;
	signal I8027: std_logic; attribute dont_touch of I8027: signal is true;
	signal I8030: std_logic; attribute dont_touch of I8030: signal is true;
	signal I8034: std_logic; attribute dont_touch of I8034: signal is true;
	signal I8040: std_logic; attribute dont_touch of I8040: signal is true;
	signal I8044: std_logic; attribute dont_touch of I8044: signal is true;
	signal I8051: std_logic; attribute dont_touch of I8051: signal is true;
	signal I8056: std_logic; attribute dont_touch of I8056: signal is true;
	signal I8061: std_logic; attribute dont_touch of I8061: signal is true;
	signal I8066: std_logic; attribute dont_touch of I8066: signal is true;
	signal I8070: std_logic; attribute dont_touch of I8070: signal is true;
	signal I8074: std_logic; attribute dont_touch of I8074: signal is true;
	signal I8079: std_logic; attribute dont_touch of I8079: signal is true;
	signal I8080: std_logic; attribute dont_touch of I8080: signal is true;
	signal I8081: std_logic; attribute dont_touch of I8081: signal is true;
	signal I8082: std_logic; attribute dont_touch of I8082: signal is true;
	signal I8089: std_logic; attribute dont_touch of I8089: signal is true;
	signal I8093: std_logic; attribute dont_touch of I8093: signal is true;
	signal I8103: std_logic; attribute dont_touch of I8103: signal is true;
	signal I8107: std_logic; attribute dont_touch of I8107: signal is true;
	signal I8110: std_logic; attribute dont_touch of I8110: signal is true;
	signal I8113: std_logic; attribute dont_touch of I8113: signal is true;
	signal I8117: std_logic; attribute dont_touch of I8117: signal is true;
	signal I8118: std_logic; attribute dont_touch of I8118: signal is true;
	signal I8119: std_logic; attribute dont_touch of I8119: signal is true;
	signal I8120: std_logic; attribute dont_touch of I8120: signal is true;
	signal I8126: std_logic; attribute dont_touch of I8126: signal is true;
	signal I8127: std_logic; attribute dont_touch of I8127: signal is true;
	signal I8128: std_logic; attribute dont_touch of I8128: signal is true;
	signal I8129: std_logic; attribute dont_touch of I8129: signal is true;
	signal I8135: std_logic; attribute dont_touch of I8135: signal is true;
	signal I8136: std_logic; attribute dont_touch of I8136: signal is true;
	signal I8137: std_logic; attribute dont_touch of I8137: signal is true;
	signal I8138: std_logic; attribute dont_touch of I8138: signal is true;
	signal I8144: std_logic; attribute dont_touch of I8144: signal is true;
	signal I8147: std_logic; attribute dont_touch of I8147: signal is true;
	signal I8150: std_logic; attribute dont_touch of I8150: signal is true;
	signal I8153: std_logic; attribute dont_touch of I8153: signal is true;
	signal I8156: std_logic; attribute dont_touch of I8156: signal is true;
	signal I8159: std_logic; attribute dont_touch of I8159: signal is true;
	signal I8162: std_logic; attribute dont_touch of I8162: signal is true;
	signal I8165: std_logic; attribute dont_touch of I8165: signal is true;
	signal I8168: std_logic; attribute dont_touch of I8168: signal is true;
	signal I8171: std_logic; attribute dont_touch of I8171: signal is true;
	signal I8174: std_logic; attribute dont_touch of I8174: signal is true;
	signal I8177: std_logic; attribute dont_touch of I8177: signal is true;
	signal I8180: std_logic; attribute dont_touch of I8180: signal is true;
	signal I8183: std_logic; attribute dont_touch of I8183: signal is true;
	signal I8186: std_logic; attribute dont_touch of I8186: signal is true;
	signal I8189: std_logic; attribute dont_touch of I8189: signal is true;
	signal I8194: std_logic; attribute dont_touch of I8194: signal is true;
	signal I8195: std_logic; attribute dont_touch of I8195: signal is true;
	signal I8196: std_logic; attribute dont_touch of I8196: signal is true;
	signal I8201: std_logic; attribute dont_touch of I8201: signal is true;
	signal I8202: std_logic; attribute dont_touch of I8202: signal is true;
	signal I8203: std_logic; attribute dont_touch of I8203: signal is true;
	signal I8208: std_logic; attribute dont_touch of I8208: signal is true;
	signal I8209: std_logic; attribute dont_touch of I8209: signal is true;
	signal I8210: std_logic; attribute dont_touch of I8210: signal is true;
	signal I8211: std_logic; attribute dont_touch of I8211: signal is true;
	signal I8217: std_logic; attribute dont_touch of I8217: signal is true;
	signal I8220: std_logic; attribute dont_touch of I8220: signal is true;
	signal I8223: std_logic; attribute dont_touch of I8223: signal is true;
	signal I8226: std_logic; attribute dont_touch of I8226: signal is true;
	signal I8229: std_logic; attribute dont_touch of I8229: signal is true;
	signal I8232: std_logic; attribute dont_touch of I8232: signal is true;
	signal I8235: std_logic; attribute dont_touch of I8235: signal is true;
	signal I8240: std_logic; attribute dont_touch of I8240: signal is true;
	signal I8243: std_logic; attribute dont_touch of I8243: signal is true;
	signal I8246: std_logic; attribute dont_touch of I8246: signal is true;
	signal I8249: std_logic; attribute dont_touch of I8249: signal is true;
	signal I8252: std_logic; attribute dont_touch of I8252: signal is true;
	signal I8255: std_logic; attribute dont_touch of I8255: signal is true;
	signal I8258: std_logic; attribute dont_touch of I8258: signal is true;
	signal I8261: std_logic; attribute dont_touch of I8261: signal is true;
	signal I8264: std_logic; attribute dont_touch of I8264: signal is true;
	signal I8267: std_logic; attribute dont_touch of I8267: signal is true;
	signal I8270: std_logic; attribute dont_touch of I8270: signal is true;
	signal I8273: std_logic; attribute dont_touch of I8273: signal is true;
	signal I8276: std_logic; attribute dont_touch of I8276: signal is true;
	signal I8279: std_logic; attribute dont_touch of I8279: signal is true;
	signal I8282: std_logic; attribute dont_touch of I8282: signal is true;
	signal I8285: std_logic; attribute dont_touch of I8285: signal is true;
	signal I8290: std_logic; attribute dont_touch of I8290: signal is true;
	signal I8295: std_logic; attribute dont_touch of I8295: signal is true;
	signal I8300: std_logic; attribute dont_touch of I8300: signal is true;
	signal I8309: std_logic; attribute dont_touch of I8309: signal is true;
	signal I8329: std_logic; attribute dont_touch of I8329: signal is true;
	signal I8332: std_logic; attribute dont_touch of I8332: signal is true;
	signal I8335: std_logic; attribute dont_touch of I8335: signal is true;
	signal I8342: std_logic; attribute dont_touch of I8342: signal is true;
	signal I8345: std_logic; attribute dont_touch of I8345: signal is true;
	signal I8346: std_logic; attribute dont_touch of I8346: signal is true;
	signal I8347: std_logic; attribute dont_touch of I8347: signal is true;
	signal I8348: std_logic; attribute dont_touch of I8348: signal is true;
	signal I8349: std_logic; attribute dont_touch of I8349: signal is true;
	signal I8356: std_logic; attribute dont_touch of I8356: signal is true;
	signal I8357: std_logic; attribute dont_touch of I8357: signal is true;
	signal I8358: std_logic; attribute dont_touch of I8358: signal is true;
	signal I8359: std_logic; attribute dont_touch of I8359: signal is true;
	signal I8360: std_logic; attribute dont_touch of I8360: signal is true;
	signal I8367: std_logic; attribute dont_touch of I8367: signal is true;
	signal I8368: std_logic; attribute dont_touch of I8368: signal is true;
	signal I8369: std_logic; attribute dont_touch of I8369: signal is true;
	signal I8370: std_logic; attribute dont_touch of I8370: signal is true;
	signal I8376: std_logic; attribute dont_touch of I8376: signal is true;
	signal I8377: std_logic; attribute dont_touch of I8377: signal is true;
	signal I8378: std_logic; attribute dont_touch of I8378: signal is true;
	signal I8379: std_logic; attribute dont_touch of I8379: signal is true;
	signal I8385: std_logic; attribute dont_touch of I8385: signal is true;
	signal I8386: std_logic; attribute dont_touch of I8386: signal is true;
	signal I8387: std_logic; attribute dont_touch of I8387: signal is true;
	signal I8393: std_logic; attribute dont_touch of I8393: signal is true;
	signal I8394: std_logic; attribute dont_touch of I8394: signal is true;
	signal I8395: std_logic; attribute dont_touch of I8395: signal is true;
	signal I8411: std_logic; attribute dont_touch of I8411: signal is true;
	signal I8414: std_logic; attribute dont_touch of I8414: signal is true;
	signal I8417: std_logic; attribute dont_touch of I8417: signal is true;
	signal I8420: std_logic; attribute dont_touch of I8420: signal is true;
	signal I8423: std_logic; attribute dont_touch of I8423: signal is true;
	signal I8426: std_logic; attribute dont_touch of I8426: signal is true;
	signal I8429: std_logic; attribute dont_touch of I8429: signal is true;
	signal I8432: std_logic; attribute dont_touch of I8432: signal is true;
	signal I8435: std_logic; attribute dont_touch of I8435: signal is true;
	signal I8438: std_logic; attribute dont_touch of I8438: signal is true;
	signal I8441: std_logic; attribute dont_touch of I8441: signal is true;
	signal I8444: std_logic; attribute dont_touch of I8444: signal is true;
	signal I8447: std_logic; attribute dont_touch of I8447: signal is true;
	signal I8450: std_logic; attribute dont_touch of I8450: signal is true;
	signal I8453: std_logic; attribute dont_touch of I8453: signal is true;
	signal I8456: std_logic; attribute dont_touch of I8456: signal is true;
	signal I8459: std_logic; attribute dont_touch of I8459: signal is true;
	signal I8462: std_logic; attribute dont_touch of I8462: signal is true;
	signal I8467: std_logic; attribute dont_touch of I8467: signal is true;
	signal I8470: std_logic; attribute dont_touch of I8470: signal is true;
	signal I8473: std_logic; attribute dont_touch of I8473: signal is true;
	signal I8476: std_logic; attribute dont_touch of I8476: signal is true;
	signal I8479: std_logic; attribute dont_touch of I8479: signal is true;
	signal I8482: std_logic; attribute dont_touch of I8482: signal is true;
	signal I8485: std_logic; attribute dont_touch of I8485: signal is true;
	signal I8488: std_logic; attribute dont_touch of I8488: signal is true;
	signal I8491: std_logic; attribute dont_touch of I8491: signal is true;
	signal I8494: std_logic; attribute dont_touch of I8494: signal is true;
	signal I8497: std_logic; attribute dont_touch of I8497: signal is true;
	signal I8500: std_logic; attribute dont_touch of I8500: signal is true;
	signal I8503: std_logic; attribute dont_touch of I8503: signal is true;
	signal I8506: std_logic; attribute dont_touch of I8506: signal is true;
	signal I8509: std_logic; attribute dont_touch of I8509: signal is true;
	signal I8512: std_logic; attribute dont_touch of I8512: signal is true;
	signal I8515: std_logic; attribute dont_touch of I8515: signal is true;
	signal I8518: std_logic; attribute dont_touch of I8518: signal is true;
	signal I8521: std_logic; attribute dont_touch of I8521: signal is true;
	signal I8524: std_logic; attribute dont_touch of I8524: signal is true;
	signal I8527: std_logic; attribute dont_touch of I8527: signal is true;
	signal I8531: std_logic; attribute dont_touch of I8531: signal is true;
	signal I8535: std_logic; attribute dont_touch of I8535: signal is true;
	signal I8538: std_logic; attribute dont_touch of I8538: signal is true;
	signal I8541: std_logic; attribute dont_touch of I8541: signal is true;
	signal I8544: std_logic; attribute dont_touch of I8544: signal is true;
	signal I8548: std_logic; attribute dont_touch of I8548: signal is true;
	signal I8552: std_logic; attribute dont_touch of I8552: signal is true;
	signal I8555: std_logic; attribute dont_touch of I8555: signal is true;
	signal I8564: std_logic; attribute dont_touch of I8564: signal is true;
	signal I8567: std_logic; attribute dont_touch of I8567: signal is true;
	signal I8570: std_logic; attribute dont_touch of I8570: signal is true;
	signal I8573: std_logic; attribute dont_touch of I8573: signal is true;
	signal I8576: std_logic; attribute dont_touch of I8576: signal is true;
	signal I8579: std_logic; attribute dont_touch of I8579: signal is true;
	signal I8582: std_logic; attribute dont_touch of I8582: signal is true;
	signal I8585: std_logic; attribute dont_touch of I8585: signal is true;
	signal I8588: std_logic; attribute dont_touch of I8588: signal is true;
	signal I8591: std_logic; attribute dont_touch of I8591: signal is true;
	signal I8594: std_logic; attribute dont_touch of I8594: signal is true;
	signal I8597: std_logic; attribute dont_touch of I8597: signal is true;
	signal I8600: std_logic; attribute dont_touch of I8600: signal is true;
	signal I8603: std_logic; attribute dont_touch of I8603: signal is true;
	signal I8614: std_logic; attribute dont_touch of I8614: signal is true;
	signal I8617: std_logic; attribute dont_touch of I8617: signal is true;
	signal I8620: std_logic; attribute dont_touch of I8620: signal is true;
	signal I8623: std_logic; attribute dont_touch of I8623: signal is true;
	signal I8626: std_logic; attribute dont_touch of I8626: signal is true;
	signal I8629: std_logic; attribute dont_touch of I8629: signal is true;
	signal I8632: std_logic; attribute dont_touch of I8632: signal is true;
	signal I8635: std_logic; attribute dont_touch of I8635: signal is true;
	signal I8638: std_logic; attribute dont_touch of I8638: signal is true;
	signal I8641: std_logic; attribute dont_touch of I8641: signal is true;
	signal I8644: std_logic; attribute dont_touch of I8644: signal is true;
	signal I8647: std_logic; attribute dont_touch of I8647: signal is true;
	signal I8650: std_logic; attribute dont_touch of I8650: signal is true;
	signal I8653: std_logic; attribute dont_touch of I8653: signal is true;
	signal I8656: std_logic; attribute dont_touch of I8656: signal is true;
	signal I8659: std_logic; attribute dont_touch of I8659: signal is true;
	signal I8662: std_logic; attribute dont_touch of I8662: signal is true;
	signal I8665: std_logic; attribute dont_touch of I8665: signal is true;
	signal I8668: std_logic; attribute dont_touch of I8668: signal is true;
	signal I8671: std_logic; attribute dont_touch of I8671: signal is true;
	signal I8674: std_logic; attribute dont_touch of I8674: signal is true;
	signal I8678: std_logic; attribute dont_touch of I8678: signal is true;
	signal I8681: std_logic; attribute dont_touch of I8681: signal is true;
	signal I8684: std_logic; attribute dont_touch of I8684: signal is true;
	signal I8687: std_logic; attribute dont_touch of I8687: signal is true;
	signal I8690: std_logic; attribute dont_touch of I8690: signal is true;
	signal I8693: std_logic; attribute dont_touch of I8693: signal is true;
	signal I8696: std_logic; attribute dont_touch of I8696: signal is true;
	signal I8699: std_logic; attribute dont_touch of I8699: signal is true;
	signal I8702: std_logic; attribute dont_touch of I8702: signal is true;
	signal I8707: std_logic; attribute dont_touch of I8707: signal is true;
	signal I8710: std_logic; attribute dont_touch of I8710: signal is true;
	signal I8713: std_logic; attribute dont_touch of I8713: signal is true;
	signal I8716: std_logic; attribute dont_touch of I8716: signal is true;
	signal I8721: std_logic; attribute dont_touch of I8721: signal is true;
	signal I8724: std_logic; attribute dont_touch of I8724: signal is true;
	signal I8727: std_logic; attribute dont_touch of I8727: signal is true;
	signal I8730: std_logic; attribute dont_touch of I8730: signal is true;
	signal I8745: std_logic; attribute dont_touch of I8745: signal is true;
	signal I8749: std_logic; attribute dont_touch of I8749: signal is true;
	signal I8752: std_logic; attribute dont_touch of I8752: signal is true;
	signal I8755: std_logic; attribute dont_touch of I8755: signal is true;
	signal I8758: std_logic; attribute dont_touch of I8758: signal is true;
	signal I8761: std_logic; attribute dont_touch of I8761: signal is true;
	signal I8764: std_logic; attribute dont_touch of I8764: signal is true;
	signal I8767: std_logic; attribute dont_touch of I8767: signal is true;
	signal I8773: std_logic; attribute dont_touch of I8773: signal is true;
	signal I8774: std_logic; attribute dont_touch of I8774: signal is true;
	signal I8778: std_logic; attribute dont_touch of I8778: signal is true;
	signal I8779: std_logic; attribute dont_touch of I8779: signal is true;
	signal I8800: std_logic; attribute dont_touch of I8800: signal is true;
	signal I8803: std_logic; attribute dont_touch of I8803: signal is true;
	signal I8806: std_logic; attribute dont_touch of I8806: signal is true;
	signal I8809: std_logic; attribute dont_touch of I8809: signal is true;
	signal I8812: std_logic; attribute dont_touch of I8812: signal is true;
	signal I8815: std_logic; attribute dont_touch of I8815: signal is true;
	signal I8818: std_logic; attribute dont_touch of I8818: signal is true;
	signal I8821: std_logic; attribute dont_touch of I8821: signal is true;
	signal I8828: std_logic; attribute dont_touch of I8828: signal is true;
	signal I8831: std_logic; attribute dont_touch of I8831: signal is true;
	signal I8834: std_logic; attribute dont_touch of I8834: signal is true;
	signal I8837: std_logic; attribute dont_touch of I8837: signal is true;
	signal I8840: std_logic; attribute dont_touch of I8840: signal is true;
	signal I8843: std_logic; attribute dont_touch of I8843: signal is true;
	signal I8854: std_logic; attribute dont_touch of I8854: signal is true;
	signal I8857: std_logic; attribute dont_touch of I8857: signal is true;
	signal I8860: std_logic; attribute dont_touch of I8860: signal is true;
	signal I8863: std_logic; attribute dont_touch of I8863: signal is true;
	signal I8866: std_logic; attribute dont_touch of I8866: signal is true;
	signal I8869: std_logic; attribute dont_touch of I8869: signal is true;
	signal I8872: std_logic; attribute dont_touch of I8872: signal is true;
	signal I8875: std_logic; attribute dont_touch of I8875: signal is true;
	signal I8878: std_logic; attribute dont_touch of I8878: signal is true;
	signal I8881: std_logic; attribute dont_touch of I8881: signal is true;
	signal I8884: std_logic; attribute dont_touch of I8884: signal is true;
	signal I8888: std_logic; attribute dont_touch of I8888: signal is true;
	signal I8891: std_logic; attribute dont_touch of I8891: signal is true;
	signal I8894: std_logic; attribute dont_touch of I8894: signal is true;
	signal I8897: std_logic; attribute dont_touch of I8897: signal is true;
	signal I8907: std_logic; attribute dont_touch of I8907: signal is true;
	signal I8910: std_logic; attribute dont_touch of I8910: signal is true;
	signal I8913: std_logic; attribute dont_touch of I8913: signal is true;
	signal I8916: std_logic; attribute dont_touch of I8916: signal is true;
	signal I8940: std_logic; attribute dont_touch of I8940: signal is true;
	signal I8943: std_logic; attribute dont_touch of I8943: signal is true;
	signal I8946: std_logic; attribute dont_touch of I8946: signal is true;
	signal I8958: std_logic; attribute dont_touch of I8958: signal is true;
	signal I8961: std_logic; attribute dont_touch of I8961: signal is true;
	signal I8966: std_logic; attribute dont_touch of I8966: signal is true;
	signal I8969: std_logic; attribute dont_touch of I8969: signal is true;
	signal I8972: std_logic; attribute dont_touch of I8972: signal is true;
	signal I8975: std_logic; attribute dont_touch of I8975: signal is true;
	signal I8978: std_logic; attribute dont_touch of I8978: signal is true;
	signal I8981: std_logic; attribute dont_touch of I8981: signal is true;
	signal I8984: std_logic; attribute dont_touch of I8984: signal is true;
	signal I8988: std_logic; attribute dont_touch of I8988: signal is true;
	signal I8991: std_logic; attribute dont_touch of I8991: signal is true;
	signal I8994: std_logic; attribute dont_touch of I8994: signal is true;
	signal I8997: std_logic; attribute dont_touch of I8997: signal is true;
	signal I9002: std_logic; attribute dont_touch of I9002: signal is true;
	signal I9005: std_logic; attribute dont_touch of I9005: signal is true;
	signal I9008: std_logic; attribute dont_touch of I9008: signal is true;
	signal I9011: std_logic; attribute dont_touch of I9011: signal is true;
	signal I9014: std_logic; attribute dont_touch of I9014: signal is true;
	signal I9021: std_logic; attribute dont_touch of I9021: signal is true;
	signal I9024: std_logic; attribute dont_touch of I9024: signal is true;
	signal I9028: std_logic; attribute dont_touch of I9028: signal is true;
	signal I9031: std_logic; attribute dont_touch of I9031: signal is true;
	signal I9035: std_logic; attribute dont_touch of I9035: signal is true;
	signal I9038: std_logic; attribute dont_touch of I9038: signal is true;
	signal I9041: std_logic; attribute dont_touch of I9041: signal is true;
	signal I9044: std_logic; attribute dont_touch of I9044: signal is true;
	signal I9047: std_logic; attribute dont_touch of I9047: signal is true;
	signal I9050: std_logic; attribute dont_touch of I9050: signal is true;
	signal I9051: std_logic; attribute dont_touch of I9051: signal is true;
	signal I9052: std_logic; attribute dont_touch of I9052: signal is true;
	signal I9057: std_logic; attribute dont_touch of I9057: signal is true;
	signal I9058: std_logic; attribute dont_touch of I9058: signal is true;
	signal I9059: std_logic; attribute dont_touch of I9059: signal is true;
	signal I9064: std_logic; attribute dont_touch of I9064: signal is true;
	signal I9065: std_logic; attribute dont_touch of I9065: signal is true;
	signal I9066: std_logic; attribute dont_touch of I9066: signal is true;
	signal I9074: std_logic; attribute dont_touch of I9074: signal is true;
	signal I9077: std_logic; attribute dont_touch of I9077: signal is true;
	signal I9082: std_logic; attribute dont_touch of I9082: signal is true;
	signal I9085: std_logic; attribute dont_touch of I9085: signal is true;
	signal I9092: std_logic; attribute dont_touch of I9092: signal is true;
	signal I9095: std_logic; attribute dont_touch of I9095: signal is true;
	signal I9098: std_logic; attribute dont_touch of I9098: signal is true;
	signal I9101: std_logic; attribute dont_touch of I9101: signal is true;
	signal I9104: std_logic; attribute dont_touch of I9104: signal is true;
	signal I9107: std_logic; attribute dont_touch of I9107: signal is true;
	signal I9110: std_logic; attribute dont_touch of I9110: signal is true;
	signal I9113: std_logic; attribute dont_touch of I9113: signal is true;
	signal I9116: std_logic; attribute dont_touch of I9116: signal is true;
	signal I9119: std_logic; attribute dont_touch of I9119: signal is true;
	signal I9122: std_logic; attribute dont_touch of I9122: signal is true;
	signal I9125: std_logic; attribute dont_touch of I9125: signal is true;
	signal I9128: std_logic; attribute dont_touch of I9128: signal is true;
	signal I9131: std_logic; attribute dont_touch of I9131: signal is true;
	signal I9134: std_logic; attribute dont_touch of I9134: signal is true;
	signal I9137: std_logic; attribute dont_touch of I9137: signal is true;
	signal I9140: std_logic; attribute dont_touch of I9140: signal is true;
	signal I9143: std_logic; attribute dont_touch of I9143: signal is true;
	signal I9146: std_logic; attribute dont_touch of I9146: signal is true;
	signal I9149: std_logic; attribute dont_touch of I9149: signal is true;
	signal I9152: std_logic; attribute dont_touch of I9152: signal is true;
	signal I9155: std_logic; attribute dont_touch of I9155: signal is true;
	signal I9158: std_logic; attribute dont_touch of I9158: signal is true;
	signal I9161: std_logic; attribute dont_touch of I9161: signal is true;
	signal I9164: std_logic; attribute dont_touch of I9164: signal is true;
	signal I9167: std_logic; attribute dont_touch of I9167: signal is true;
	signal I9170: std_logic; attribute dont_touch of I9170: signal is true;
	signal I9173: std_logic; attribute dont_touch of I9173: signal is true;
	signal I9176: std_logic; attribute dont_touch of I9176: signal is true;
	signal I9179: std_logic; attribute dont_touch of I9179: signal is true;
	signal I9182: std_logic; attribute dont_touch of I9182: signal is true;
	signal I9185: std_logic; attribute dont_touch of I9185: signal is true;
	signal I9203: std_logic; attribute dont_touch of I9203: signal is true;
	signal I9208: std_logic; attribute dont_touch of I9208: signal is true;
	signal I9217: std_logic; attribute dont_touch of I9217: signal is true;
	signal I9220: std_logic; attribute dont_touch of I9220: signal is true;
	signal I9227: std_logic; attribute dont_touch of I9227: signal is true;
	signal I9230: std_logic; attribute dont_touch of I9230: signal is true;
	signal I9233: std_logic; attribute dont_touch of I9233: signal is true;
	signal I9236: std_logic; attribute dont_touch of I9236: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			G1<=G6720;
			G2<=G6721;
			G3<=G6597;
			G6<=G6722;
			G7<=G6598;
			G10<=G6723;
			G11<=G6599;
			G14<=G6724;
			G15<=G6602;
			G18<=G6725;
			G19<=G6600;
			G24<=G6726;
			G25<=G6601;
			G28<=G6727;
			G29<=G6853;
			G33<=G6854;
			G43<=G6407;
			G48<=G6729;
			G49<=G6583;
			G54<=G6584;
			G59<=G6585;
			G64<=G6586;
			G69<=G6587;
			G74<=G6588;
			G79<=G6589;
			G84<=G6590;
			G111<=G6277;
			G114<=G4116;
			G117<=G4839;
			G118<=G4113;
			G119<=G4114;
			G122<=G4115;
			G123<=G6940;
			G127<=G6941;
			G128<=G5138;
			G131<=G5139;
			G135<=G5140;
			G139<=G5141;
			G143<=G6401;
			G148<=G5874;
			G152<=G6402;
			G157<=G5470;
			G161<=G6403;
			G166<=G5471;
			G170<=G6404;
			G175<=G5472;
			G179<=G6405;
			G184<=G5473;
			G188<=G6406;
			G193<=G5474;
			G197<=G6509;
			G204<=G5875;
			G205<=G6100;
			G206<=G6101;
			G207<=G6102;
			G208<=G5876;
			G209<=G6103;
			G210<=G6839;
			G211<=G6840;
			G212<=G3233;
			G218<=G3234;
			G224<=G3235;
			G230<=G3236;
			G236<=G3237;
			G242<=G3238;
			G248<=G3239;
			G254<=G3240;
			G260<=G3241;
			G266<=G4659;
			G269<=G6510;
			G276<=G5877;
			G277<=G6104;
			G278<=G6105;
			G279<=G6106;
			G280<=G5878;
			G281<=G6107;
			G282<=G6841;
			G283<=G6842;
			G284<=G3224;
			G285<=G3225;
			G286<=G3226;
			G287<=G3227;
			G288<=G3228;
			G289<=G3229;
			G290<=G3230;
			G291<=G3231;
			G292<=G3232;
			G293<=G6511;
			G297<=G6512;
			G323<=G4120;
			G326<=G4840;
			G327<=G4117;
			G328<=G4118;
			G331<=G4119;
			G332<=G6823;
			G336<=G6925;
			G337<=G2585;
			G338<=G5475;
			G341<=G5476;
			G345<=G5477;
			G349<=G5478;
			G353<=G5479;
			G357<=G5480;
			G361<=G6582;
			G366<=G6278;
			G370<=G5693;
			G374<=G5694;
			G378<=G5695;
			G382<=G5696;
			G386<=G5697;
			G390<=G5698;
			G394<=G5699;
			G398<=G5700;
			G402<=G4849;
			G406<=G4850;
			G410<=G4851;
			G414<=G4852;
			G418<=G4853;
			G422<=G4854;
			G426<=G4855;
			G430<=G4856;
			G434<=G4848;
			G437<=G4847;
			G441<=G4846;
			G445<=G4845;
			G449<=G4844;
			G453<=G4843;
			G457<=G4842;
			G461<=G4841;
			G465<=G6507;
			G471<=G1291;
			G478<=G1292;
			G485<=G6801;
			G486<=G2586;
			G489<=G2587;
			G492<=G6744;
			G496<=G6745;
			G500<=G6497;
			G504<=G6498;
			G508<=G6499;
			G512<=G6500;
			G516<=G6501;
			G520<=G6502;
			G524<=G6503;
			G528<=G6504;
			G532<=G6508;
			G536<=G6506;
			G541<=G6505;
			G545<=G6824;
			G548<=G6825;
			G551<=G6826;
			G554<=G6827;
			G571<=G5580;
			G574<=G6591;
			G578<=G6592;
			G582<=G6593;
			G586<=G6594;
			G590<=G6595;
			G594<=G6596;
			G598<=G4122;
			G602<=G4123;
			G606<=G4857;
			G610<=G4124;
			G613<=G4423;
			G616<=G4657;
			G619<=G4858;
			G622<=G5147;
			G625<=G5328;
			G628<=G5489;
			G631<=G5581;
			G634<=G4424;
			G638<=G1289;
			G642<=G4658;
			G646<=G5148;
			G650<=G5329;
			G654<=G5490;
			G658<=G4425;
			G662<=G1831;
			G663<=G4125;
			G664<=G1288;
			G665<=G4126;
			G666<=G4128;
			G667<=G4127;
			G668<=G6800;
			G669<=G5582;
			G672<=G5491;
			G675<=G1294;
			G676<=G5330;
			G677<=G4129;
			G678<=G4130;
			G679<=G4131;
			G680<=G4132;
			G681<=G4133;
			G682<=G4134;
			G683<=G4135;
			G684<=G4136;
			G685<=G4137;
			G686<=G4138;
			G687<=G4139;
			G688<=G4140;
			G689<=G4141;
			G690<=G4142;
			G691<=G4143;
			G692<=G4144;
			G693<=G4145;
			G694<=G4146;
			G695<=G4147;
			G696<=G4148;
			G697<=G4149;
			G698<=G4150;
			G699<=G4426;
		end if;
	end process;
	G706<= not I1825;
	G709<= not G114;
	G710<= not G128;
	G714<= not G131;
	G715<= not G135;
	G716<= not I1832;
	G719<= not I1835;
	G729<= not I1838;
	G736<= not I1841;
	G743<= not I1844;
	G749<= not I1847;
	G754<= not I1850;
	G760<= not I1853;
	G766<= not I1856;
	G774<= not I1859;
	G784<= not I1862;
	G791<= not I1865;
	G798<= not I1868;
	G804<= not I1871;
	G809<= not I1874;
	G815<= not I1877;
	G821<= not I1880;
	G829<= not G323;
	G830<= not G338;
	G834<= not G341;
	G835<= not G345;
	G836<= not G349;
	G837<= not G353;
	G838<= not G564;
	G839<= not G567;
	G842<= not G571;
	G843<= not G574;
	G844<= not G578;
	G845<= not G582;
	G846<= not G586;
	G847<= not G590;
	G848<= not G594;
	G849<= not G598;
	G850<= not G602;
	G851<= not G606;
	G852<= not G634;
	G853<= not G642;
	G854<= not G646;
	G855<= not G650;
	G856<= not G654;
	G857<= not G170;
	G858<= not G301;
	G861<= not G179;
	G862<= not G319;
	G865<= not G188;
	G866<= not G314;
	G872<= not G143;
	G873<= not G306;
	G878<= not G639;
	G889<= not G310;
	G893<= not G23;
	G894<= not I1917;
	G895<= not G139;
	G896<= not G22;
	G897<= not G41;
	G898<= not G47;
	G899<= not I1924;
	G900<= not I1927;
	G908<= not I1932;
	G909<= not I1935;
	G910<= not I1938;
	G913<= not G658;
	G917<= not I1942;
	G921<= not G111;
	G922<= not I1947;
	G923<= not G332;
	G927<= not I1958;
	G929<= not G49;
	G931<= not G54;
	G932<= not G337;
	G938<= not G59;
	G940<= not G64;
	G942<= not G69;
	G943<= not G496;
	G945<= not G536;
	G946<= not G361;
	G947<= not G74;
	G949<= not G79;
	G951<= not G84;
	G952<= not I2029;
	G964<= not G357;
	G965<= not I2033;
	G971<= not G658;
	G980<= not I2037;
	G985<= not G638;
	G996<= not I2041;
	G1001<= not I2044;
	G1006<= not I2047;
	G1011<= not I2050;
	G1017<= not I2053;
	G1030<= not I2057;
	G1037<= not I2067;
	G1038<= not G127;
	G1039<= not G662;
	G1043<= not G486;
	G1045<= not G699;
	G1046<= not G489;
	G1048<= not G492;
	G1049<= not G266;
	G1052<= not G668;
	G1053<= not G197;
	G1054<= not G485;
	G1055<= not G269;
	G1056<= not G89;
	G1059<= not G702;
	G1060<= not G107;
	G1063<= not G675;
	G1064<= not G102;
	G1070<= not G94;
	G1076<= not I2115;
	G1084<= not G98;
	G1088<= not I2119;
	G1094<= not I2122;
	G1101<= not I2125;
	G1106<= not I2128;
	G1107<= not I2131;
	G1108<= not I2134;
	G1109<= not I2137;
	G1110<= not I2140;
	G1111<= not I2143;
	G1112<= not G336;
	G1113<= not I2147;
	G1114<= not I2150;
	G1115<= not G40;
	G1116<= not I2154;
	G1117<= not G32;
	G1118<= not G36;
	G1119<= not I2159;
	G1122<= not I2162;
	G1123<= not I2165;
	G1142<= not I2169;
	G1143<= not I2172;
	G1156<= not I2175;
	G1160<= not I2179;
	G1161<= not I2182;
	G1173<= not I2185;
	G1174<= not G37;
	G1175<= not G42;
	G1176<= not I2190;
	G1177<= not I2193;
	G1189<= not I2196;
	G1190<= not I2199;
	G1191<= not G38;
	G1192<= not G44;
	G1193<= not I2204;
	G1203<= not I2207;
	G1204<= not G39;
	G1205<= not G45;
	G1206<= not I2212;
	G1209<= not I2215;
	G1219<= not I2218;
	G1220<= not I2221;
	G1221<= not G46;
	G1222<= not I2225;
	G1232<= not I2228;
	G1233<= not I2231;
	G1236<= not I2234;
	G1246<= not I2237;
	G1249<= not I2240;
	G1250<= not G123;
	G1254<= not G152;
	G1255<= not G161;
	G1256<= not G838;
	G1257<= not G845;
	G1263<= not G846;
	G1267<= not G843;
	G1270<= not G844;
	G1273<= not G839;
	G1274<= not G856;
	G1275<= not G842;
	G1276<= not G847;
	G1279<= not G848;
	G1282<= not G849;
	G1283<= not G853;
	G1284<= not G851;
	G1285<= not G852;
	G1286<= not G854;
	G1287<= not G855;
	G1288<= not I2269;
	G1289<= not I2272;
	G1290<= not I2275;
	G1291<= not I2278;
	G1292<= not I2281;
	G1293<= not I2284;
	G1294<= not I2287;
	G1295<= not I2290;
	G1305<= not I2293;
	G1315<= not I2296;
	G1317<= not I2306;
	G1318<= not I2309;
	G1319<= not I2312;
	G1320<= not I2315;
	G1321<= not I2318;
	G1322<= not I2321;
	G1323<= not I2324;
	G1324<= not I2327;
	G1325<= not I2330;
	G1326<= not G894;
	G1327<= not I2334;
	G1328<= not I2337;
	G1329<= not I2340;
	G1330<= not I2343;
	G1331<= not I2346;
	G1332<= not I2349;
	G1333<= not I2352;
	G1334<= not I2355;
	G1335<= not I2358;
	G1336<= not I2361;
	G1337<= not I2364;
	G1338<= not I2367;
	G1339<= not I2370;
	G1340<= not I2373;
	G1341<= not I2376;
	G1344<= not I2379;
	G1345<= not I2382;
	G1348<= not I2385;
	G1351<= not I2388;
	G1352<= not I2391;
	G1355<= not I2394;
	G1358<= not G1119;
	G1363<= not I2399;
	G1366<= not I2402;
	G1369<= not I2405;
	G1372<= not I2408;
	G1375<= not I2411;
	G1378<= not I2414;
	G1381<= not I2417;
	G1384<= not I2420;
	G1391<= not I2424;
	G1394<= not G1206;
	G1395<= not I2428;
	G1410<= not G1233;
	G1415<= not G1246;
	G1423<= not I2442;
	G1426<= not I2445;
	G1439<= not I2449;
	G1450<= not I2453;
	G1460<= not I2457;
	G1461<= not I2460;
	G1471<= not I2464;
	G1472<= not G952;
	G1477<= not G952;
	G1480<= not G985;
	G1484<= not I2473;
	G1491<= not I2476;
	G1498<= not I2479;
	G1502<= not G709;
	G1503<= not G878;
	G1504<= not I2485;
	G1513<= not G878;
	G1519<= not I2491;
	G1528<= not G878;
	G1529<= not G1076;
	G1533<= not G878;
	G1535<= not G1088;
	G1539<= not G878;
	G1541<= not G1094;
	G1542<= not G878;
	G1543<= not G1006;
	G1546<= not G1101;
	G1549<= not G878;
	G1550<= not G996;
	G1551<= not G1011;
	G1552<= not G1030;
	G1555<= not I2521;
	G1556<= not G878;
	G1557<= not G1017;
	G1559<= not G965;
	G1563<= not G1006;
	G1564<= not G1030;
	G1567<= not I2537;
	G1577<= not G1001;
	G1578<= not I2552;
	G1581<= not G910;
	G1583<= not G1001;
	G1584<= not G743;
	G1586<= not G1052;
	G1587<= not G1123;
	G1588<= not G798;
	G1593<= not G1054;
	G1594<= not G1143;
	G1608<= not I2570;
	G1623<= not I2578;
	G1624<= not I2581;
	G1627<= not I2584;
	G1631<= not I2588;
	G1632<= not G760;
	G1636<= not I2593;
	G1637<= not I2596;
	G1638<= not G754;
	G1639<= not G815;
	G1640<= not I2601;
	G1641<= not I2604;
	G1642<= not G809;
	G1643<= not I2608;
	G1644<= not I2611;
	G1645<= not I2614;
	G1646<= not I2617;
	G1647<= not I2620;
	G1648<= not I2623;
	G1649<= not G985;
	G1650<= not I2627;
	G1653<= not I2630;
	G1654<= not G878;
	G1655<= not G985;
	G1656<= not I2635;
	G1659<= not I2638;
	G1660<= not G985;
	G1661<= not G1076;
	G1664<= not I2643;
	G1665<= not G985;
	G1666<= not G1088;
	G1670<= not I2648;
	G1671<= not G985;
	G1672<= not G1094;
	G1673<= not I2653;
	G1674<= not G985;
	G1675<= not G1101;
	G1678<= not I2658;
	G1679<= not G985;
	G1680<= not G1011;
	G1681<= not I2663;
	G1682<= not G829;
	G1683<= not G1017;
	G1684<= not I2668;
	G1685<= not I2671;
	G1688<= not I2688;
	G1690<= not I2692;
	G1692<= not I2696;
	G1695<= not G1106;
	G1696<= not I2700;
	G1699<= not I2703;
	G1702<= not G1107;
	G1703<= not I2707;
	G1710<= not G1109;
	G1711<= not I2712;
	G1714<= not G1110;
	G1715<= not I2716;
	G1720<= not G1111;
	G1721<= not I2721;
	G1724<= not I2724;
	G1725<= not G1113;
	G1726<= not I2728;
	G1729<= not I2731;
	G1730<= not G1114;
	G1731<= not I2735;
	G1732<= not I2738;
	G1733<= not I2741;
	G1734<= not G952;
	G1735<= not I2745;
	G1738<= not G1108;
	G1739<= not I2749;
	G1740<= not G1116;
	G1741<= not I2753;
	G1742<= not I2756;
	G1747<= not I2760;
	G1748<= not I2763;
	G1754<= not I2773;
	G1755<= not I2776;
	G1756<= not I2779;
	G1759<= not I2782;
	G1760<= not I2785;
	G1761<= not I2788;
	G1762<= not I2791;
	G1769<= not I2802;
	G1770<= not I2805;
	G1771<= not I2808;
	G1772<= not I2811;
	G1773<= not I2814;
	G1774<= not I2817;
	G1775<= not G952;
	G1776<= not I2821;
	G1781<= not I2825;
	G1782<= not I2828;
	G1783<= not I2831;
	G1787<= not I2835;
	G1788<= not G985;
	G1789<= not I2839;
	G1790<= not I2842;
	G1791<= not I2845;
	G1792<= not I2848;
	G1805<= not I2854;
	G1806<= not I2857;
	G1807<= not I2860;
	G1811<= not I2864;
	G1812<= not I2867;
	G1813<= not I2870;
	G1814<= not I2873;
	G1819<= not I2877;
	G1820<= not I2880;
	G1821<= not I2883;
	G1823<= not I2887;
	G1824<= not I2890;
	G1825<= not I2893;
	G1830<= not I2904;
	G1831<= not I2907;
	G1832<= not I2910;
	G1833<= not I2913;
	G1834<= not I2916;
	G1835<= not I2919;
	G1836<= not I2922;
	G1837<= not I2925;
	G1838<= not G1595;
	G1841<= not I2929;
	G1842<= not G1612;
	G1846<= not I2940;
	G1847<= not I2943;
	G1848<= not I2946;
	G1849<= not I2949;
	G1852<= not I2952;
	G1853<= not I2955;
	G1854<= not I2958;
	G1857<= not I2961;
	G1858<= not I2964;
	G1861<= not I2967;
	G1875<= not I2970;
	G1878<= not I2973;
	G1880<= not G1603;
	G1883<= not G1797;
	G1884<= not I2979;
	G1887<= not I2982;
	G1890<= not G1359;
	G1891<= not I2986;
	G1894<= not I2989;
	G1897<= not I2992;
	G1898<= not I2995;
	G1899<= not I2998;
	G1902<= not I3001;
	G1905<= not I3004;
	G1908<= not I3007;
	G1911<= not I3010;
	G1914<= not I3013;
	G1917<= not I3016;
	G1918<= not I3019;
	G1919<= not I3022;
	G1922<= not I3025;
	G1925<= not I3028;
	G1928<= not I3031;
	G1931<= not I3034;
	G1934<= not I3037;
	G1935<= not I3040;
	G1936<= not G1756;
	G1937<= not I3044;
	G1940<= not I3047;
	G1943<= not I3050;
	G1946<= not I3053;
	G1947<= not I3056;
	G1950<= not I3059;
	G1953<= not I3062;
	G1954<= not I3065;
	G1957<= not I3068;
	G1960<= not I3071;
	G1963<= not I3074;
	G1966<= not I3077;
	G1969<= not I3080;
	G1972<= not I3083;
	G1975<= not I3086;
	G1978<= not G1387;
	G1979<= not I3090;
	G1982<= not I3093;
	G1985<= not I3096;
	G1988<= not I3099;
	G1991<= not I3102;
	G1994<= not I3105;
	G1997<= not G1398;
	G1998<= not I3109;
	G2001<= not I3112;
	G2004<= not I3115;
	G2007<= not G1411;
	G2025<= not G1276;
	G2029<= not I3134;
	G2030<= not I3137;
	G2031<= not I3140;
	G2032<= not G1749;
	G2035<= not I3144;
	G2036<= not G1764;
	G2039<= not I3148;
	G2040<= not G1738;
	G2041<= not I3152;
	G2042<= not I3155;
	G2043<= not I3158;
	G2044<= not I3161;
	G2059<= not G1402;
	G2060<= not G1369;
	G2066<= not G1341;
	G2078<= not G1345;
	G2079<= not G1348;
	G2086<= not I3198;
	G2087<= not G1352;
	G2088<= not I3202;
	G2090<= not I3206;
	G2091<= not G1355;
	G2096<= not I3212;
	G2097<= not I3215;
	G2098<= not G1363;
	G2099<= not G1366;
	G2102<= not I3222;
	G2103<= not I3225;
	G2104<= not G1372;
	G2105<= not G1375;
	G2106<= not G1378;
	G2108<= not I3232;
	G2109<= not I3235;
	G2110<= not G1381;
	G2111<= not G1384;
	G2112<= not I3240;
	G2117<= not I3244;
	G2118<= not I3247;
	G2119<= not G1391;
	G2120<= not I3251;
	G2125<= not I3255;
	G2134<= not I3258;
	G2135<= not I3261;
	G2136<= not G1395;
	G2145<= not I3268;
	G2154<= not I3271;
	G2155<= not I3274;
	G2157<= not I3278;
	G2158<= not I3281;
	G2159<= not I3284;
	G2163<= not I3288;
	G2164<= not I3291;
	G2165<= not I3294;
	G2169<= not I3298;
	G2170<= not I3301;
	G2171<= not I3304;
	G2172<= not I3307;
	G2173<= not I3310;
	G2174<= not I3313;
	G2175<= not I3316;
	G2176<= not I3319;
	G2177<= not I3322;
	G2178<= not I3325;
	G2179<= not I3328;
	G2194<= not I3331;
	G2195<= not I3334;
	G2196<= not I3337;
	G2197<= not I3340;
	G2212<= not I3343;
	G2213<= not I3346;
	G2214<= not I3349;
	G2215<= not I3352;
	G2230<= not I3355;
	G2231<= not I3358;
	G2232<= not I3361;
	G2233<= not I3364;
	G2234<= not I3367;
	G2241<= not I3370;
	G2242<= not I3373;
	G2243<= not I3376;
	G2244<= not I3379;
	G2245<= not I3382;
	G2252<= not I3385;
	G2253<= not I3388;
	G2254<= not I3391;
	G2256<= not I3395;
	G2264<= not I3405;
	G2265<= not I3408;
	G2268<= not I3419;
	G2275<= not I3422;
	G2276<= not I3425;
	G2283<= not I3428;
	G2284<= not I3431;
	G2291<= not I3434;
	G2293<= not G1567;
	G2295<= not G1578;
	G2296<= not I3441;
	G2306<= not G1743;
	G2308<= not I3452;
	G2312<= not I3462;
	G2315<= not I3465;
	G2316<= not I3468;
	G2317<= not I3471;
	G2320<= not I3474;
	G2324<= not I3478;
	G2327<= not I3481;
	G2330<= not G1777;
	G2333<= not I3485;
	G2336<= not I3488;
	G2343<= not I3493;
	G2346<= not I3496;
	G2347<= not I3499;
	G2350<= not I3502;
	G2353<= not I3505;
	G2357<= not I3509;
	G2360<= not G1793;
	G2361<= not I3513;
	G2364<= not I3516;
	G2367<= not I3519;
	G2370<= not I3522;
	G2378<= not I3525;
	G2381<= not I3528;
	G2390<= not I3531;
	G2391<= not I3534;
	G2394<= not I3537;
	G2397<= not I3540;
	G2405<= not I3543;
	G2408<= not I3546;
	G2409<= not G1815;
	G2410<= not I3550;
	G2413<= not I3553;
	G2416<= not I3556;
	G2422<= not I3560;
	G2430<= not I3563;
	G2436<= not I3569;
	G2437<= not I3572;
	G2440<= not I3575;
	G2443<= not I3578;
	G2446<= not I3581;
	G2449<= not I3584;
	G2457<= not I3587;
	G2460<= not I3590;
	G2461<= not I3593;
	G2464<= not I3596;
	G2467<= not I3599;
	G2470<= not I3602;
	G2473<= not I3605;
	G2481<= not I3608;
	G2484<= not I3611;
	G2485<= not I3614;
	G2488<= not I3617;
	G2491<= not I3620;
	G2494<= not I3623;
	G2497<= not I3626;
	G2505<= not I3629;
	G2506<= not I3632;
	G2509<= not I3635;
	G2512<= not I3638;
	G2515<= not I3641;
	G2518<= not I3644;
	G2524<= not I3647;
	G2525<= not I3650;
	G2535<= not I3653;
	G2538<= not I3656;
	G2541<= not I3659;
	G2544<= not I3662;
	G2550<= not I3665;
	G2554<= not I3669;
	G2555<= not I3672;
	G2565<= not I3675;
	G2568<= not I3678;
	G2574<= not I3681;
	G2575<= not I3684;
	G2576<= not I3687;
	G2580<= not I3691;
	G2581<= not I3694;
	G2583<= not G1830;
	G2584<= not I3705;
	G2585<= not I3708;
	G2586<= not I3711;
	G2587<= not I3714;
	G2588<= not I3717;
	G2591<= not I3720;
	G2594<= not I3723;
	G2598<= not I3726;
	G2599<= not I3729;
	G2602<= not G2061;
	G2603<= not I3733;
	G2604<= not I3736;
	G2608<= not I3746;
	G2609<= not I3749;
	G2612<= not I3752;
	G2615<= not I3755;
	G2618<= not I3758;
	G2619<= not I3761;
	G2622<= not I3764;
	G2625<= not I3767;
	G2628<= not I3770;
	G2631<= not I3773;
	G2634<= not I3776;
	G2637<= not I3779;
	G2640<= not I3782;
	G2643<= not I3785;
	G2644<= not I3788;
	G2647<= not I3791;
	G2650<= not I3794;
	G2653<= not I3797;
	G2656<= not I3800;
	G2660<= not I3804;
	G2663<= not G2308;
	G2664<= not I3808;
	G2667<= not I3811;
	G2672<= not I3816;
	G2675<= not I3819;
	G2678<= not G2312;
	G2679<= not I3823;
	G2682<= not I3826;
	G2686<= not I3830;
	G2687<= not I3833;
	G2688<= not I3836;
	G2691<= not G2317;
	G2692<= not I3840;
	G2695<= not I3843;
	G2701<= not I3855;
	G2705<= not I3858;
	G2706<= not I3861;
	G2709<= not I3864;
	G2712<= not G2320;
	G2713<= not I3868;
	G2716<= not I3871;
	G2722<= not I3883;
	G2726<= not I3886;
	G2727<= not G2324;
	G2728<= not I3890;
	G2734<= not I3902;
	G2738<= not G2327;
	G2739<= not I3906;
	G2740<= not I3909;
	G2743<= not G2333;
	G2744<= not G2336;
	G2748<= not I3923;
	G2752<= not G2343;
	G2753<= not I3927;
	G2754<= not G2347;
	G2755<= not G2350;
	G2756<= not G2353;
	G2760<= not I3942;
	G2764<= not G2357;
	G2765<= not I3946;
	G2766<= not G2361;
	G2767<= not G2364;
	G2768<= not G2367;
	G2772<= not I3961;
	G2776<= not G2378;
	G2777<= not I3965;
	G2778<= not G2391;
	G2779<= not G2394;
	G2783<= not I3979;
	G2787<= not G2405;
	G2788<= not I3983;
	G2789<= not G2410;
	G2790<= not G2413;
	G2792<= not G2416;
	G2796<= not I3999;
	G2800<= not G2430;
	G2801<= not I4003;
	G2802<= not G2437;
	G2803<= not G2440;
	G2805<= not G2443;
	G2806<= not G2446;
	G2809<= not I4019;
	G2813<= not G2457;
	G2814<= not I4023;
	G2817<= not G2461;
	G2818<= not G2464;
	G2819<= not G2467;
	G2820<= not G2470;
	G2822<= not I4031;
	G2826<= not G2481;
	G2827<= not G2485;
	G2828<= not G2488;
	G2829<= not G2491;
	G2830<= not G2494;
	G2835<= not G2506;
	G2836<= not G2509;
	G2837<= not G2512;
	G2838<= not G2515;
	G2839<= not G2535;
	G2840<= not G2538;
	G2841<= not G2541;
	G2842<= not I4050;
	G2845<= not G2565;
	G2849<= not G2577;
	G2856<= not G2010;
	G2857<= not I4059;
	G2862<= not I4066;
	G2863<= not G2296;
	G2864<= not G1887;
	G2865<= not G2296;
	G2866<= not G1905;
	G2867<= not G1908;
	G2869<= not G2433;
	G2870<= not G2296;
	G2871<= not G1919;
	G2872<= not G1922;
	G2874<= not G1849;
	G2875<= not G1940;
	G2876<= not G1943;
	G2877<= not G2434;
	G2882<= not G1854;
	G2883<= not G1954;
	G2884<= not G1957;
	G2885<= not G1963;
	G2886<= not G1966;
	G2887<= not G1858;
	G2888<= not G1972;
	G2889<= not G1975;
	G2890<= not G1875;
	G2891<= not G1884;
	G2892<= not G1982;
	G2893<= not G1985;
	G2894<= not G1891;
	G2895<= not G1894;
	G2902<= not G1899;
	G2903<= not G1902;
	G2904<= not G1991;
	G2905<= not G1994;
	G2906<= not G1911;
	G2907<= not G1914;
	G2912<= not G2001;
	G2913<= not G1925;
	G2914<= not G1928;
	G2915<= not G1931;
	G2919<= not G1937;
	G2920<= not G1947;
	G2921<= not G1950;
	G2922<= not G1960;
	G2923<= not G1969;
	G2927<= not G1979;
	G2931<= not G1988;
	G2932<= not G1998;
	G2933<= not I4123;
	G2934<= not G2004;
	G2936<= not G2026;
	G2945<= not I4133;
	G2946<= not G2296;
	G2952<= not G2381;
	G2954<= not G2381;
	G2956<= not G1861;
	G2957<= not G1861;
	G2958<= not G1861;
	G2959<= not G1861;
	G2961<= not G1861;
	G2962<= not G2008;
	G2967<= not I4166;
	G2968<= not G2179;
	G2973<= not I4170;
	G2974<= not I4173;
	G2975<= not I4176;
	G2976<= not G2197;
	G2981<= not G2179;
	G2986<= not G2010;
	G2996<= not I4189;
	G2997<= not I4192;
	G2998<= not I4195;
	G3001<= not I4198;
	G3002<= not G2215;
	G3007<= not G2197;
	G3014<= not I4217;
	G3015<= not I4220;
	G3016<= not I4223;
	G3019<= not I4226;
	G3022<= not I4229;
	G3023<= not G2215;
	G3029<= not I4240;
	G3030<= not I4243;
	G3031<= not I4246;
	G3034<= not I4249;
	G3037<= not I4252;
	G3040<= not I4255;
	G3041<= not I4258;
	G3042<= not I4261;
	G3043<= not I4264;
	G3046<= not I4267;
	G3049<= not I4270;
	G3052<= not I4273;
	G3053<= not I4276;
	G3054<= not I4279;
	G3057<= not I4282;
	G3060<= not I4285;
	G3063<= not I4288;
	G3064<= not I4291;
	G3067<= not I4294;
	G3070<= not I4297;
	G3073<= not I4300;
	G3074<= not I4303;
	G3075<= not I4306;
	G3076<= not I4309;
	G3079<= not I4312;
	G3082<= not I4315;
	G3083<= not I4318;
	G3084<= not I4321;
	G3085<= not I4324;
	G3086<= not I4327;
	G3090<= not I4331;
	G3093<= not I4334;
	G3094<= not I4337;
	G3095<= not I4340;
	G3096<= not I4343;
	G3100<= not I4347;
	G3104<= not I4351;
	G3108<= not I4354;
	G3110<= not I4358;
	G3114<= not I4362;
	G3118<= not I4366;
	G3124<= not I4371;
	G3128<= not I4375;
	G3136<= not I4382;
	G3150<= not I4391;
	G3158<= not I4398;
	G3162<= not I4402;
	G3173<= not I4410;
	G3177<= not I4414;
	G3183<= not I4420;
	G3187<= not I4424;
	G3192<= not I4429;
	G3196<= not I4433;
	G3199<= not G1861;
	G3200<= not I4437;
	G3204<= not I4441;
	G3209<= not I4452;
	G3212<= not I4455;
	G3216<= not I4459;
	G3219<= not I4462;
	G3222<= not I4465;
	G3223<= not I4468;
	G3224<= not I4471;
	G3225<= not I4474;
	G3226<= not I4477;
	G3227<= not I4480;
	G3228<= not I4483;
	G3229<= not I4486;
	G3230<= not I4489;
	G3231<= not I4492;
	G3232<= not I4495;
	G3233<= not I4498;
	G3234<= not I4501;
	G3235<= not I4504;
	G3236<= not I4507;
	G3237<= not I4510;
	G3238<= not I4513;
	G3239<= not I4516;
	G3240<= not I4519;
	G3241<= not I4522;
	G3242<= not G3083;
	G3247<= not G2973;
	G3251<= not I4534;
	G3258<= not I4537;
	G3259<= not G2996;
	G3263<= not G3015;
	G3267<= not G3030;
	G3271<= not G3042;
	G3284<= not G3019;
	G3289<= not G3034;
	G3291<= not G3037;
	G3297<= not G3046;
	G3299<= not G3049;
	G3306<= not G3057;
	G3308<= not G3060;
	G3312<= not I4587;
	G3318<= not I4593;
	G3320<= not G3067;
	G3322<= not G3070;
	G3331<= not G3076;
	G3332<= not G3079;
	G3342<= not G3086;
	G3343<= not G3090;
	G3346<= not I4623;
	G3354<= not G3096;
	G3355<= not G3100;
	G3363<= not G3110;
	G3364<= not G3114;
	G3369<= not I4646;
	G3370<= not G3124;
	G3380<= not G2831;
	G3384<= not G2834;
	G3387<= not I4664;
	G3388<= not I4667;
	G3424<= not I4671;
	G3440<= not I4678;
	G3441<= not I4681;
	G3448<= not I4684;
	G3450<= not I4688;
	G3451<= not G2615;
	G3452<= not G2625;
	G3453<= not G2628;
	G3455<= not G2637;
	G3456<= not G2640;
	G3457<= not G2653;
	G3458<= not G2656;
	G3459<= not G2664;
	G3460<= not G2667;
	G3461<= not G2986;
	G3462<= not G2679;
	G3463<= not G2682;
	G3465<= not G2986;
	G3466<= not I4706;
	G3477<= not G2692;
	G3478<= not G2695;
	G3480<= not G2986;
	G3481<= not G2612;
	G3482<= not G2713;
	G3483<= not G2716;
	G3485<= not G2986;
	G3486<= not G2869;
	G3487<= not G2622;
	G3488<= not G2728;
	G3491<= not G2608;
	G3498<= not G2634;
	G3500<= not G2647;
	G3501<= not G2650;
	G3504<= not G2675;
	G3510<= not G2709;
	G3519<= not G2740;
	G3527<= not I4743;
	G3534<= not I4752;
	G3537<= not I4757;
	G3540<= not I4762;
	G3541<= not G2643;
	G3545<= not G3085;
	G3546<= not G3095;
	G3557<= not G2598;
	G3559<= not G2603;
	G3564<= not G2618;
	G3567<= not G3074;
	G3571<= not G3084;
	G3575<= not I4777;
	G3589<= not G3094;
	G3593<= not G2997;
	G3600<= not I4791;
	G3601<= not I4794;
	G3604<= not I4799;
	G3605<= not I4802;
	G3612<= not I4809;
	G3622<= not I4821;
	G3638<= not G3108;
	G3673<= not G3075;
	G3677<= not G3140;
	G3705<= not G3014;
	G3710<= not G3029;
	G3714<= not G3041;
	G3719<= not G3053;
	G3723<= not I4903;
	G3752<= not I4935;
	G3761<= not G3605;
	G3766<= not I4955;
	G3769<= not G3622;
	G3770<= not I4961;
	G3771<= not I4964;
	G3772<= not G3466;
	G3773<= not G3466;
	G3775<= not G3388;
	G3776<= not G3466;
	G3777<= not G3388;
	G3778<= not G3388;
	G3779<= not G3466;
	G3781<= not I4976;
	G3782<= not G3388;
	G3783<= not I4980;
	G3785<= not G3466;
	G3786<= not G3388;
	G3787<= not I4986;
	G3788<= not G3466;
	G3789<= not G3388;
	G3790<= not G3388;
	G3791<= not G3388;
	G3792<= not G3388;
	G3793<= not G3491;
	G3796<= not G3388;
	G3797<= not G3388;
	G3798<= not G3388;
	G3799<= not G3388;
	G3800<= not G3388;
	G3801<= not G3388;
	G3802<= not G3388;
	G3803<= not I5002;
	G3807<= not I5006;
	G3813<= not G3258;
	G3830<= not I5019;
	G3832<= not I5023;
	G3834<= not I5027;
	G3835<= not I5030;
	G3836<= not I5033;
	G3838<= not I5037;
	G3839<= not I5040;
	G3840<= not I5043;
	G3845<= not I5050;
	G3846<= not I5053;
	G3847<= not I5056;
	G3848<= not I5059;
	G3852<= not I5065;
	G3853<= not I5068;
	G3854<= not I5071;
	G3859<= not I5078;
	G3860<= not I5081;
	G3861<= not I5084;
	G3866<= not I5091;
	G3867<= not I5094;
	G3868<= not G3491;
	G3872<= not G3312;
	G3874<= not I5103;
	G3875<= not I5106;
	G3876<= not I5109;
	G3881<= not I5116;
	G3882<= not I5119;
	G3885<= not I5124;
	G3886<= not G3346;
	G3889<= not G3575;
	G3890<= not G3575;
	G3892<= not G3575;
	G3897<= not G3251;
	G3898<= not G3575;
	G3900<= not G3575;
	G3901<= not G3575;
	G3902<= not G3575;
	G3904<= not G3575;
	G3906<= not G3575;
	G3911<= not I5148;
	G3912<= not G3505;
	G3914<= not I5153;
	G3921<= not G3512;
	G3922<= not I5157;
	G3932<= not I5169;
	G3940<= not I5177;
	G3952<= not I5182;
	G3960<= not I5204;
	G3962<= not I5214;
	G3963<= not I5217;
	G3967<= not I5223;
	G3969<= not I5233;
	G3970<= not I5236;
	G3975<= not I5249;
	G3976<= not I5252;
	G3980<= not I5264;
	G3984<= not G3564;
	G4003<= not G3441;
	G4010<= not G3601;
	G4011<= not G3486;
	G4014<= not I5316;
	G4016<= not I5320;
	G4020<= not I5324;
	G4022<= not I5328;
	G4034<= not I5333;
	G4036<= not I5337;
	G4040<= not I5343;
	G4098<= not I5376;
	G4099<= not I5379;
	G4100<= not I5382;
	G4101<= not I5385;
	G4102<= not I5388;
	G4103<= not I5391;
	G4104<= not I5394;
	G4105<= not I5397;
	G4106<= not I5400;
	G4107<= not I5403;
	G4108<= not I5406;
	G4109<= not I5409;
	G4110<= not I5412;
	G4111<= not I5415;
	G4112<= not I5418;
	G4113<= not I5421;
	G4114<= not I5424;
	G4115<= not I5427;
	G4116<= not I5430;
	G4117<= not I5433;
	G4118<= not I5436;
	G4119<= not I5439;
	G4120<= not I5442;
	G4121<= not I5445;
	G4122<= not I5448;
	G4123<= not I5451;
	G4124<= not I5454;
	G4125<= not I5457;
	G4126<= not I5460;
	G4127<= not I5463;
	G4128<= not I5466;
	G4129<= not I5469;
	G4130<= not I5472;
	G4131<= not I5475;
	G4132<= not I5478;
	G4133<= not I5481;
	G4134<= not I5484;
	G4135<= not I5487;
	G4136<= not I5490;
	G4137<= not I5493;
	G4138<= not I5496;
	G4139<= not I5499;
	G4140<= not I5502;
	G4141<= not I5505;
	G4142<= not I5508;
	G4143<= not I5511;
	G4144<= not I5514;
	G4145<= not I5517;
	G4146<= not I5520;
	G4147<= not I5523;
	G4148<= not I5526;
	G4149<= not I5529;
	G4150<= not I5532;
	G4152<= not I5542;
	G4153<= not I5545;
	G4154<= not I5548;
	G4155<= not I5551;
	G4158<= not I5556;
	G4162<= not I5562;
	G4166<= not I5568;
	G4173<= not I5577;
	G4187<= not I5591;
	G4188<= not I5594;
	G4189<= not I5597;
	G4190<= not I5600;
	G4191<= not I5603;
	G4192<= not I5606;
	G4193<= not I5609;
	G4194<= not I5612;
	G4195<= not I5615;
	G4198<= not I5618;
	G4202<= not I5622;
	G4206<= not I5626;
	G4210<= not I5630;
	G4213<= not I5633;
	G4215<= not I5637;
	G4218<= not I5640;
	G4220<= not I5644;
	G4222<= not I5654;
	G4224<= not G4046;
	G4225<= not G4059;
	G4226<= not G4050;
	G4227<= not G4059;
	G4228<= not I5668;
	G4229<= not G4059;
	G4232<= not I5674;
	G4242<= not I5686;
	G4246<= not I5692;
	G4248<= not I5696;
	G4249<= not I5699;
	G4250<= not I5702;
	G4251<= not I5705;
	G4252<= not I5708;
	G4262<= not I5713;
	G4265<= not I5716;
	G4267<= not I5720;
	G4270<= not I5723;
	G4273<= not I5728;
	G4276<= not I5731;
	G4281<= not I5736;
	G4284<= not I5739;
	G4286<= not I5743;
	G4289<= not I5746;
	G4292<= not G4059;
	G4293<= not I5750;
	G4296<= not I5753;
	G4299<= not I5756;
	G4302<= not G4068;
	G4307<= not I5774;
	G4308<= not I5777;
	G4309<= not G4074;
	G4314<= not G4080;
	G4320<= not G4011;
	G4321<= not I5790;
	G4322<= not I5793;
	G4323<= not G4086;
	G4328<= not G4092;
	G4334<= not G3733;
	G4343<= not G4011;
	G4350<= not G4010;
	G4364<= not I5825;
	G4370<= not I5831;
	G4374<= not I5837;
	G4375<= not I5840;
	G4376<= not I5843;
	G4379<= not I5848;
	G4380<= not I5851;
	G4381<= not I5854;
	G4382<= not I5857;
	G4385<= not I5862;
	G4386<= not I5865;
	G4387<= not I5868;
	G4388<= not I5871;
	G4391<= not I5876;
	G4392<= not I5879;
	G4393<= not I5882;
	G4394<= not I5885;
	G4397<= not I5890;
	G4398<= not I5893;
	G4399<= not I5896;
	G4400<= not I5899;
	G4402<= not G4017;
	G4403<= not I5904;
	G4404<= not I5907;
	G4405<= not I5910;
	G4406<= not I5913;
	G4422<= not G4111;
	G4423<= not I5920;
	G4424<= not I5923;
	G4425<= not I5926;
	G4426<= not I5929;
	G4428<= not I5933;
	G4431<= not I5938;
	G4435<= not I5944;
	G4437<= not I5948;
	G4439<= not I5952;
	G4462<= not I5977;
	G4463<= not G4364;
	G4485<= not I5987;
	G4487<= not I5991;
	G4492<= not I5998;
	G4493<= not I6001;
	G4494<= not I6004;
	G4496<= not I6008;
	G4498<= not I6012;
	G4499<= not I6015;
	G4502<= not I6020;
	G4503<= not I6023;
	G4507<= not I6033;
	G4508<= not I6036;
	G4509<= not I6039;
	G4510<= not I6042;
	G4511<= not I6045;
	G4512<= not I6048;
	G4513<= not I6051;
	G4514<= not I6054;
	G4515<= not I6057;
	G4516<= not I6060;
	G4517<= not I6063;
	G4518<= not I6066;
	G4519<= not I6069;
	G4520<= not I6072;
	G4521<= not I6075;
	G4522<= not I6078;
	G4523<= not I6081;
	G4524<= not I6084;
	G4525<= not I6087;
	G4526<= not I6090;
	G4527<= not I6093;
	G4528<= not I6096;
	G4529<= not I6099;
	G4530<= not I6102;
	G4531<= not I6105;
	G4532<= not I6108;
	G4533<= not I6111;
	G4534<= not I6114;
	G4535<= not G4173;
	G4536<= not I6118;
	G4537<= not G4410;
	G4545<= not G4416;
	G4550<= not I6126;
	G4559<= not G4187;
	G4560<= not G4188;
	G4561<= not G4189;
	G4562<= not I6132;
	G4563<= not G4190;
	G4564<= not G4192;
	G4565<= not G4195;
	G4566<= not G4198;
	G4567<= not I6139;
	G4569<= not I6143;
	G4577<= not G4202;
	G4579<= not G4206;
	G4582<= not G4210;
	G4587<= not G4215;
	G4601<= not G4191;
	G4603<= not I6170;
	G4606<= not G4193;
	G4609<= not I6182;
	G4612<= not G4320;
	G4614<= not G4308;
	G4615<= not G4322;
	G4617<= not G4242;
	G4618<= not G4246;
	G4619<= not G4248;
	G4620<= not G4251;
	G4622<= not G4252;
	G4623<= not G4262;
	G4624<= not G4265;
	G4625<= not G4267;
	G4626<= not G4270;
	G4628<= not G4273;
	G4629<= not G4276;
	G4632<= not G4281;
	G4633<= not G4284;
	G4636<= not G4286;
	G4639<= not G4289;
	G4643<= not G4293;
	G4644<= not I6231;
	G4647<= not G4296;
	G4657<= not I6244;
	G4658<= not I6247;
	G4659<= not I6250;
	G4660<= not I6253;
	G4662<= not G4640;
	G4679<= not I6269;
	G4692<= not I6280;
	G4693<= not I6283;
	G4699<= not I6289;
	G4700<= not I6292;
	G4702<= not I6296;
	G4703<= not I6299;
	G4704<= not I6302;
	G4705<= not I6305;
	G4706<= not I6308;
	G4707<= not I6311;
	G4711<= not I6315;
	G4712<= not I6318;
	G4713<= not I6321;
	G4714<= not I6324;
	G4715<= not I6327;
	G4716<= not I6330;
	G4717<= not G4465;
	G4718<= not I6334;
	G4719<= not I6337;
	G4720<= not I6340;
	G4721<= not I6343;
	G4722<= not I6346;
	G4723<= not I6349;
	G4726<= not I6352;
	G4727<= not I6355;
	G4731<= not I6359;
	G4732<= not I6362;
	G4736<= not I6366;
	G4741<= not I6371;
	G4753<= not I6377;
	G4758<= not I6382;
	G4760<= not I6386;
	G4763<= not I6397;
	G4764<= not I6400;
	G4765<= not I6403;
	G4766<= not I6406;
	G4767<= not G4601;
	G4768<= not I6410;
	G4769<= not G4606;
	G4770<= not I6414;
	G4771<= not I6417;
	G4772<= not I6420;
	G4775<= not I6425;
	G4778<= not I6430;
	G4780<= not I6434;
	G4781<= not I6437;
	G4783<= not I6441;
	G4784<= not I6444;
	G4786<= not I6448;
	G4788<= not I6452;
	G4790<= not I6456;
	G4798<= not I6464;
	G4799<= not G4485;
	G4801<= not G4487;
	G4802<= not I6470;
	G4804<= not G4473;
	G4805<= not G4473;
	G4806<= not G4473;
	G4807<= not G4473;
	G4808<= not G4473;
	G4809<= not I6485;
	G4810<= not I6488;
	G4815<= not I6495;
	G4822<= not G4614;
	G4823<= not I6507;
	G4824<= not G4615;
	G4837<= not G4473;
	G4839<= not I6525;
	G4840<= not I6528;
	G4841<= not I6531;
	G4842<= not I6534;
	G4843<= not I6537;
	G4844<= not I6540;
	G4845<= not I6543;
	G4846<= not I6546;
	G4847<= not I6549;
	G4848<= not I6552;
	G4849<= not I6555;
	G4850<= not I6558;
	G4851<= not I6561;
	G4852<= not I6564;
	G4853<= not I6567;
	G4854<= not I6570;
	G4855<= not I6573;
	G4856<= not I6576;
	G4857<= not I6579;
	G4858<= not I6582;
	G4861<= not I6587;
	G4869<= not G4662;
	G4871<= not I6599;
	G4894<= not G4813;
	G4900<= not I6607;
	G4904<= not G4812;
	G4910<= not I6612;
	G4911<= not I6615;
	G4914<= not G4816;
	G4915<= not G4669;
	G4929<= not I6621;
	G4933<= not I6625;
	G4938<= not I6630;
	G4943<= not I6635;
	G4980<= not G4678;
	G5010<= not I6646;
	G5011<= not I6649;
	G5022<= not I6666;
	G5025<= not G4814;
	G5042<= not I6672;
	G5045<= not I6677;
	G5046<= not I6680;
	G5049<= not I6685;
	G5051<= not I6689;
	G5052<= not I6692;
	G5054<= not G4816;
	G5059<= not I6697;
	G5061<= not I6701;
	G5063<= not G4799;
	G5064<= not I6706;
	G5067<= not G4801;
	G5082<= not G4723;
	G5084<= not G4727;
	G5086<= not G4732;
	G5087<= not G4736;
	G5089<= not I6723;
	G5090<= not G4741;
	G5092<= not G4753;
	G5097<= not I6733;
	G5099<= not I6737;
	G5110<= not I6740;
	G5112<= not I6750;
	G5113<= not I6753;
	G5114<= not I6756;
	G5115<= not I6759;
	G5116<= not G4810;
	G5117<= not I6763;
	G5118<= not I6766;
	G5119<= not I6769;
	G5120<= not I6772;
	G5121<= not I6775;
	G5124<= not I6780;
	G5135<= not I6783;
	G5136<= not I6786;
	G5137<= not I6789;
	G5138<= not I6792;
	G5139<= not I6795;
	G5140<= not I6798;
	G5141<= not I6801;
	G5147<= not I6809;
	G5148<= not I6812;
	G5150<= not I6816;
	G5151<= not I6819;
	G5155<= not G5099;
	G5160<= not G5099;
	G5168<= not G5099;
	G5174<= not G5099;
	G5179<= not G5099;
	G5199<= not I6867;
	G5210<= not I6874;
	G5219<= not I6885;
	G5220<= not G4903;
	G5230<= not I6895;
	G5237<= not G5083;
	G5242<= not G5085;
	G5247<= not G4900;
	G5248<= not G4911;
	G5250<= not G4929;
	G5251<= not G5069;
	G5255<= not G4933;
	G5256<= not G5077;
	G5260<= not G4938;
	G5261<= not I6918;
	G5264<= not G4943;
	G5266<= not I6923;
	G5270<= not I6927;
	G5273<= not I6930;
	G5274<= not I6933;
	G5278<= not I6937;
	G5292<= not I6942;
	G5296<= not I6946;
	G5299<= not I6949;
	G5300<= not I6952;
	G5304<= not I6956;
	G5307<= not I6959;
	G5309<= not G5063;
	G5310<= not G5067;
	G5314<= not I6972;
	G5315<= not G5116;
	G5316<= not I6976;
	G5328<= not I6986;
	G5329<= not I6989;
	G5330<= not I6992;
	G5331<= not I6995;
	G5352<= not I7002;
	G5355<= not I7007;
	G5358<= not I7012;
	G5375<= not I7029;
	G5379<= not I7035;
	G5381<= not I7039;
	G5382<= not I7042;
	G5383<= not I7045;
	G5384<= not G5220;
	G5387<= not I7051;
	G5391<= not I7055;
	G5392<= not I7058;
	G5395<= not I7061;
	G5399<= not I7065;
	G5403<= not I7069;
	G5407<= not I7073;
	G5411<= not I7077;
	G5415<= not I7081;
	G5420<= not I7086;
	G5425<= not I7091;
	G5432<= not I7104;
	G5433<= not I7107;
	G5434<= not I7110;
	G5435<= not I7113;
	G5436<= not I7116;
	G5437<= not I7119;
	G5439<= not G5261;
	G5440<= not G5266;
	G5442<= not G5270;
	G5445<= not G5274;
	G5448<= not G5278;
	G5450<= not G5292;
	G5453<= not G5296;
	G5456<= not G5300;
	G5457<= not G5304;
	G5465<= not I7143;
	G5466<= not I7146;
	G5468<= not I7150;
	G5469<= not I7153;
	G5475<= not I7161;
	G5476<= not I7164;
	G5477<= not I7167;
	G5478<= not I7170;
	G5479<= not I7173;
	G5480<= not I7176;
	G5489<= not I7187;
	G5490<= not I7190;
	G5491<= not I7193;
	G5493<= not I7197;
	G5509<= not I7251;
	G5512<= not I7254;
	G5518<= not I7258;
	G5521<= not I7261;
	G5524<= not I7264;
	G5527<= not I7267;
	G5530<= not I7270;
	G5534<= not I7276;
	G5536<= not G5467;
	G5537<= not G5385;
	G5538<= not G5331;
	G5539<= not G5331;
	G5540<= not I7284;
	G5542<= not G5331;
	G5543<= not G5331;
	G5544<= not G5331;
	G5545<= not G5331;
	G5546<= not G5388;
	G5549<= not G5331;
	G5550<= not G5331;
	G5551<= not I7295;
	G5554<= not G5455;
	G5563<= not G5381;
	G5564<= not G5382;
	G5566<= not I7318;
	G5567<= not G5418;
	G5568<= not G5423;
	G5570<= not G5392;
	G5571<= not G5395;
	G5572<= not G5399;
	G5573<= not G5403;
	G5574<= not G5407;
	G5575<= not G5411;
	G5576<= not G5415;
	G5577<= not G5420;
	G5578<= not G5425;
	G5579<= not I7333;
	G5580<= not I7336;
	G5581<= not I7339;
	G5582<= not I7342;
	G5584<= not I7346;
	G5587<= not I7349;
	G5590<= not I7352;
	G5593<= not I7355;
	G5596<= not I7358;
	G5597<= not I7361;
	G5615<= not I7372;
	G5631<= not G5536;
	G5638<= not I7397;
	G5645<= not G5537;
	G5647<= not G5509;
	G5649<= not I7404;
	G5658<= not G5512;
	G5661<= not G5518;
	G5664<= not G5521;
	G5667<= not G5524;
	G5670<= not G5527;
	G5685<= not G5552;
	G5687<= not G5567;
	G5691<= not G5568;
	G5692<= not I7451;
	G5702<= not I7463;
	G5705<= not I7466;
	G5708<= not I7469;
	G5711<= not I7472;
	G5714<= not I7475;
	G5717<= not I7478;
	G5720<= not I7481;
	G5723<= not I7484;
	G5726<= not I7487;
	G5727<= not I7490;
	G5729<= not I7494;
	G5730<= not I7497;
	G5740<= not I7501;
	G5741<= not G5602;
	G5742<= not G5686;
	G5751<= not I7506;
	G5752<= not I7509;
	G5770<= not G5645;
	G5773<= not I7514;
	G5774<= not I7517;
	G5784<= not I7583;
	G5787<= not G5685;
	G5788<= not I7587;
	G5791<= not I7590;
	G5794<= not I7593;
	G5797<= not I7596;
	G5801<= not I7600;
	G5805<= not I7604;
	G5809<= not I7608;
	G5813<= not I7612;
	G5824<= not G5631;
	G5860<= not G5634;
	G5861<= not G5636;
	G5874<= not I7634;
	G5875<= not I7637;
	G5876<= not I7640;
	G5877<= not I7643;
	G5878<= not I7646;
	G5879<= not G5770;
	G5880<= not G5824;
	G5884<= not G5864;
	G5885<= not G5865;
	G5886<= not G5753;
	G5887<= not G5742;
	G5888<= not G5731;
	G5889<= not G5742;
	G5890<= not G5753;
	G5891<= not G5731;
	G5892<= not G5742;
	G5893<= not G5753;
	G5894<= not G5731;
	G5895<= not G5742;
	G5896<= not G5753;
	G5897<= not G5731;
	G5899<= not G5753;
	G5901<= not G5753;
	G5903<= not G5753;
	G5905<= not G5852;
	G5908<= not G5753;
	G5912<= not G5853;
	G5915<= not I7679;
	G5917<= not I7683;
	G5918<= not I7686;
	G5919<= not I7689;
	G5920<= not I7692;
	G5921<= not I7695;
	G5922<= not I7698;
	G5923<= not I7701;
	G5924<= not I7704;
	G5925<= not I7707;
	G5946<= not G5729;
	G5950<= not G5730;
	G5957<= not G5866;
	G5958<= not G5818;
	G5975<= not G5821;
	G5992<= not G5869;
	G5993<= not G5872;
	G5994<= not G5873;
	G5995<= not G5824;
	G5996<= not G5824;
	G5997<= not G5854;
	G6014<= not G5824;
	G6015<= not G5857;
	G6032<= not G5770;
	G6033<= not G5824;
	G6034<= not G5824;
	G6035<= not G5824;
	G6036<= not G5824;
	G6039<= not G5824;
	G6040<= not G5824;
	G6043<= not G5824;
	G6044<= not G5824;
	G6048<= not G5824;
	G6051<= not G5824;
	G6052<= not G5824;
	G6057<= not G5824;
	G6062<= not G5824;
	G6065<= not G5784;
	G6067<= not G5788;
	G6069<= not G5791;
	G6070<= not G5824;
	G6074<= not G5794;
	G6076<= not G5797;
	G6078<= not G5801;
	G6080<= not G5805;
	G6083<= not G5809;
	G6087<= not G5813;
	G6100<= not I7796;
	G6101<= not I7799;
	G6102<= not I7802;
	G6103<= not I7805;
	G6104<= not I7808;
	G6105<= not I7811;
	G6106<= not I7814;
	G6107<= not I7817;
	G6115<= not G5879;
	G6117<= not G5880;
	G6119<= not I7829;
	G6120<= not I7832;
	G6121<= not I7835;
	G6122<= not I7838;
	G6134<= not I7852;
	G6136<= not I7856;
	G6137<= not I7859;
	G6143<= not I7865;
	G6147<= not I7871;
	G6160<= not G5926;
	G6161<= not G5926;
	G6162<= not G5926;
	G6163<= not G5926;
	G6164<= not G5926;
	G6165<= not G5926;
	G6166<= not I7892;
	G6188<= not G5950;
	G6192<= not G5946;
	G6193<= not G5957;
	G6194<= not I7906;
	G6211<= not G5992;
	G6212<= not I7910;
	G6229<= not G6036;
	G6230<= not G6040;
	G6231<= not G6044;
	G6232<= not G6048;
	G6233<= not G6052;
	G6234<= not G6057;
	G6235<= not G6062;
	G6236<= not G6070;
	G6276<= not I7960;
	G6277<= not I7963;
	G6278<= not I7966;
	G6282<= not I7996;
	G6283<= not I7999;
	G6284<= not I8002;
	G6285<= not I8005;
	G6305<= not I8027;
	G6306<= not I8030;
	G6308<= not I8034;
	G6312<= not I8040;
	G6314<= not I8044;
	G6319<= not I8051;
	G6322<= not I8056;
	G6325<= not I8061;
	G6328<= not I8066;
	G6330<= not I8070;
	G6332<= not I8074;
	G6337<= not I8089;
	G6339<= not I8093;
	G6347<= not I8103;
	G6351<= not I8107;
	G6352<= not I8110;
	G6353<= not I8113;
	G6360<= not I8144;
	G6361<= not I8147;
	G6362<= not I8150;
	G6363<= not I8153;
	G6364<= not I8156;
	G6365<= not I8159;
	G6366<= not I8162;
	G6367<= not I8165;
	G6368<= not I8168;
	G6369<= not I8171;
	G6370<= not I8174;
	G6371<= not I8177;
	G6372<= not I8180;
	G6373<= not I8183;
	G6374<= not I8186;
	G6375<= not I8189;
	G6376<= not G6267;
	G6385<= not G6271;
	G6401<= not I8217;
	G6402<= not I8220;
	G6403<= not I8223;
	G6404<= not I8226;
	G6405<= not I8229;
	G6406<= not I8232;
	G6407<= not I8235;
	G6408<= not G6283;
	G6409<= not G6285;
	G6410<= not I8240;
	G6411<= not I8243;
	G6412<= not I8246;
	G6413<= not I8249;
	G6414<= not I8252;
	G6415<= not I8255;
	G6416<= not I8258;
	G6417<= not I8261;
	G6418<= not I8264;
	G6419<= not I8267;
	G6420<= not I8270;
	G6421<= not I8273;
	G6422<= not I8276;
	G6423<= not I8279;
	G6424<= not I8282;
	G6425<= not I8285;
	G6428<= not I8290;
	G6431<= not I8295;
	G6434<= not I8300;
	G6441<= not I8309;
	G6465<= not I8329;
	G6466<= not I8332;
	G6467<= not I8335;
	G6478<= not I8342;
	G6484<= not G6361;
	G6486<= not G6363;
	G6487<= not G6365;
	G6488<= not G6367;
	G6489<= not G6369;
	G6490<= not G6371;
	G6491<= not G6373;
	G6493<= not G6375;
	G6497<= not I8411;
	G6498<= not I8414;
	G6499<= not I8417;
	G6500<= not I8420;
	G6501<= not I8423;
	G6502<= not I8426;
	G6503<= not I8429;
	G6504<= not I8432;
	G6505<= not I8435;
	G6506<= not I8438;
	G6507<= not I8441;
	G6508<= not I8444;
	G6509<= not I8447;
	G6510<= not I8450;
	G6511<= not I8453;
	G6512<= not I8456;
	G6513<= not I8459;
	G6514<= not I8462;
	G6515<= not G6408;
	G6516<= not G6409;
	G6517<= not I8467;
	G6518<= not I8470;
	G6519<= not I8473;
	G6520<= not I8476;
	G6521<= not I8479;
	G6522<= not I8482;
	G6523<= not I8485;
	G6524<= not I8488;
	G6525<= not I8491;
	G6526<= not I8494;
	G6527<= not I8497;
	G6528<= not I8500;
	G6529<= not I8503;
	G6530<= not I8506;
	G6531<= not I8509;
	G6532<= not I8512;
	G6533<= not I8515;
	G6534<= not I8518;
	G6535<= not I8521;
	G6536<= not I8524;
	G6537<= not I8527;
	G6538<= not G6469;
	G6539<= not I8531;
	G6540<= not G6474;
	G6541<= not I8535;
	G6542<= not I8538;
	G6543<= not I8541;
	G6544<= not I8544;
	G6548<= not I8548;
	G6552<= not I8552;
	G6553<= not I8555;
	G6560<= not I8564;
	G6561<= not I8567;
	G6562<= not I8570;
	G6563<= not I8573;
	G6564<= not I8576;
	G6565<= not I8579;
	G6566<= not I8582;
	G6567<= not I8585;
	G6568<= not I8588;
	G6569<= not I8591;
	G6570<= not I8594;
	G6571<= not I8597;
	G6572<= not I8600;
	G6573<= not I8603;
	G6574<= not G6484;
	G6575<= not G6486;
	G6576<= not G6487;
	G6577<= not G6488;
	G6578<= not G6489;
	G6579<= not G6490;
	G6580<= not G6491;
	G6581<= not G6493;
	G6582<= not I8614;
	G6583<= not I8617;
	G6584<= not I8620;
	G6585<= not I8623;
	G6586<= not I8626;
	G6587<= not I8629;
	G6588<= not I8632;
	G6589<= not I8635;
	G6590<= not I8638;
	G6591<= not I8641;
	G6592<= not I8644;
	G6593<= not I8647;
	G6594<= not I8650;
	G6595<= not I8653;
	G6596<= not I8656;
	G6597<= not I8659;
	G6598<= not I8662;
	G6599<= not I8665;
	G6600<= not I8668;
	G6601<= not I8671;
	G6602<= not I8674;
	G6604<= not I8678;
	G6605<= not I8681;
	G6606<= not I8684;
	G6607<= not I8687;
	G6608<= not I8690;
	G6609<= not I8693;
	G6610<= not I8696;
	G6611<= not I8699;
	G6612<= not I8702;
	G6615<= not I8707;
	G6616<= not I8710;
	G6617<= not I8713;
	G6618<= not I8716;
	G6621<= not I8721;
	G6622<= not I8724;
	G6623<= not I8727;
	G6624<= not I8730;
	G6649<= not I8745;
	G6651<= not I8749;
	G6652<= not I8752;
	G6653<= not I8755;
	G6654<= not I8758;
	G6655<= not I8761;
	G6656<= not I8764;
	G6657<= not I8767;
	G6694<= not I8800;
	G6695<= not I8803;
	G6696<= not I8806;
	G6697<= not I8809;
	G6698<= not I8812;
	G6699<= not I8815;
	G6700<= not I8818;
	G6701<= not I8821;
	G6706<= not I8828;
	G6707<= not I8831;
	G6708<= not I8834;
	G6709<= not I8837;
	G6710<= not I8840;
	G6711<= not I8843;
	G6712<= not G6676;
	G6713<= not G6679;
	G6714<= not G6670;
	G6715<= not G6673;
	G6720<= not I8854;
	G6721<= not I8857;
	G6722<= not I8860;
	G6723<= not I8863;
	G6724<= not I8866;
	G6725<= not I8869;
	G6726<= not I8872;
	G6727<= not I8875;
	G6728<= not I8878;
	G6729<= not I8881;
	G6730<= not I8884;
	G6732<= not I8888;
	G6733<= not I8891;
	G6734<= not I8894;
	G6735<= not I8897;
	G6743<= not I8907;
	G6744<= not I8910;
	G6745<= not I8913;
	G6746<= not I8916;
	G6784<= not I8940;
	G6785<= not I8943;
	G6786<= not I8946;
	G6796<= not I8958;
	G6797<= not I8961;
	G6800<= not I8966;
	G6801<= not I8969;
	G6802<= not I8972;
	G6803<= not I8975;
	G6806<= not I8978;
	G6809<= not I8981;
	G6812<= not I8984;
	G6817<= not I8988;
	G6818<= not I8991;
	G6819<= not I8994;
	G6820<= not I8997;
	G6821<= not G6785;
	G6822<= not G6786;
	G6823<= not I9002;
	G6824<= not I9005;
	G6825<= not I9008;
	G6826<= not I9011;
	G6827<= not I9014;
	G6832<= not I9021;
	G6833<= not I9024;
	G6834<= not G6821;
	G6835<= not I9028;
	G6836<= not I9031;
	G6837<= not G6822;
	G6838<= not I9035;
	G6839<= not I9038;
	G6840<= not I9041;
	G6841<= not I9044;
	G6842<= not I9047;
	G6849<= not I9074;
	G6850<= not I9077;
	G6853<= not I9082;
	G6854<= not I9085;
	G6875<= not I9092;
	G6876<= not I9095;
	G6877<= not I9098;
	G6878<= not I9101;
	G6879<= not I9104;
	G6880<= not I9107;
	G6881<= not I9110;
	G6882<= not I9113;
	G6883<= not I9116;
	G6884<= not I9119;
	G6885<= not I9122;
	G6886<= not I9125;
	G6887<= not I9128;
	G6888<= not I9131;
	G6889<= not I9134;
	G6890<= not I9137;
	G6891<= not I9140;
	G6892<= not I9143;
	G6893<= not I9146;
	G6894<= not I9149;
	G6895<= not I9152;
	G6896<= not I9155;
	G6897<= not I9158;
	G6898<= not I9161;
	G6899<= not I9164;
	G6900<= not I9167;
	G6901<= not I9170;
	G6902<= not I9173;
	G6903<= not I9176;
	G6904<= not I9179;
	G6905<= not I9182;
	G6906<= not I9185;
	G6922<= not I9203;
	G6925<= not I9208;
	G6932<= not I9217;
	G6933<= not I9220;
	G6938<= not I9227;
	G6939<= not I9230;
	G6940<= not I9233;
	G6941<= not I9236;
	I1825<= not G361;
	I1832<= not G143;
	I1835<= not G205;
	I1838<= not G206;
	I1841<= not G207;
	I1844<= not G208;
	I1847<= not G209;
	I1850<= not G210;
	I1853<= not G211;
	I1856<= not G204;
	I1859<= not G277;
	I1862<= not G278;
	I1865<= not G279;
	I1868<= not G280;
	I1871<= not G281;
	I1874<= not G282;
	I1877<= not G283;
	I1880<= not G276;
	I1917<= not G48;
	I1924<= not G663;
	I1927<= not G665;
	I1932<= not G667;
	I1935<= not G666;
	I1938<= not G332;
	I1942<= not G664;
	I1947<= not G699;
	I1958<= not G702;
	I2029<= not G677;
	I2033<= not G678;
	I2037<= not G679;
	I2041<= not G680;
	I2044<= not G681;
	I2047<= not G682;
	I2050<= not G683;
	I2053<= not G684;
	I2057<= not G685;
	I2067<= not G686;
	I2115<= not G687;
	I2119<= not G688;
	I2122<= not G689;
	I2125<= not G698;
	I2128<= not G18;
	I2131<= not G24;
	I2134<= not G705;
	I2137<= not G1;
	I2140<= not G28;
	I2143<= not G2;
	I2147<= not G6;
	I2150<= not G10;
	I2154<= not G14;
	I2159<= not G465;
	I2162<= not G197;
	I2165<= not G690;
	I2169<= not G269;
	I2172<= not G691;
	I2175<= not G25;
	I2179<= not G293;
	I2182<= not G692;
	I2185<= not G29;
	I2190<= not G297;
	I2193<= not G693;
	I2196<= not G3;
	I2199<= not G33;
	I2204<= not G694;
	I2207<= not G7;
	I2212<= not G123;
	I2215<= not G695;
	I2218<= not G11;
	I2221<= not G43;
	I2225<= not G696;
	I2228<= not G15;
	I2231<= not G465;
	I2234<= not G697;
	I2237<= not G465;
	I2240<= not G19;
	I2269<= not G899;
	I2272<= not G908;
	I2275<= not G909;
	I2278<= not G917;
	I2281<= not G900;
	I2284<= not G922;
	I2287<= not G927;
	I2290<= not G971;
	I2293<= not G971;
	I2296<= not G893;
	I2306<= not G896;
	I2309<= not G1236;
	I2312<= not G897;
	I2315<= not G1222;
	I2318<= not G1236;
	I2321<= not G898;
	I2324<= not G1209;
	I2327<= not G1222;
	I2330<= not G1122;
	I2334<= not G1193;
	I2337<= not G1209;
	I2340<= not G1142;
	I2343<= not G1177;
	I2346<= not G1193;
	I2349<= not G1160;
	I2352<= not G1161;
	I2355<= not G1177;
	I2358<= not G1176;
	I2361<= not G1075;
	I2364<= not G1143;
	I2367<= not G1161;
	I2370<= not G1123;
	I2373<= not G1143;
	I2376<= not G729;
	I2379<= not G1123;
	I2382<= not G719;
	I2385<= not G784;
	I2388<= not G878;
	I2391<= not G774;
	I2394<= not G719;
	I2399<= not G729;
	I2402<= not G774;
	I2405<= not G1112;
	I2408<= not G719;
	I2411<= not G736;
	I2414<= not G784;
	I2417<= not G774;
	I2420<= not G791;
	I2424<= not G719;
	I2428<= not G774;
	I2442<= not G872;
	I2445<= not G971;
	I2449<= not G971;
	I2453<= not G952;
	I2457<= not G1253;
	I2460<= not G952;
	I2464<= not G850;
	I2473<= not G971;
	I2476<= not G971;
	I2479<= not G1049;
	I2485<= not G766;
	I2491<= not G821;
	I2521<= not G1063;
	I2537<= not G971;
	I2552<= not G971;
	I2570<= not G1222;
	I2578<= not G1209;
	I2581<= not G946;
	I2584<= not G839;
	I2588<= not G1193;
	I2593<= not G1177;
	I2596<= not G985;
	I2601<= not G1161;
	I2604<= not G1222;
	I2608<= not G1143;
	I2611<= not G1209;
	I2614<= not G1123;
	I2617<= not G1193;
	I2620<= not G1177;
	I2623<= not G1161;
	I2627<= not G1053;
	I2630<= not G1143;
	I2635<= not G1055;
	I2638<= not G1123;
	I2643<= not G965;
	I2648<= not G980;
	I2653<= not G996;
	I2658<= not G1001;
	I2663<= not G1006;
	I2668<= not G1011;
	I2671<= not G1017;
	I2688<= not G1030;
	I2692<= not G1037;
	I2696<= not G1156;
	I2700<= not G1173;
	I2703<= not G1189;
	I2707<= not G1190;
	I2712<= not G1203;
	I2716<= not G1115;
	I2721<= not G1219;
	I2724<= not G1220;
	I2728<= not G1232;
	I2731<= not G1117;
	I2735<= not G1118;
	I2738<= not G1236;
	I2741<= not G1222;
	I2745<= not G1249;
	I2749<= not G1209;
	I2753<= not G1174;
	I2756<= not G1175;
	I2760<= not G1193;
	I2763<= not G1236;
	I2773<= not G1191;
	I2776<= not G1192;
	I2779<= not G1038;
	I2782<= not G1177;
	I2785<= not G1222;
	I2788<= not G1236;
	I2791<= not G1236;
	I2802<= not G1204;
	I2805<= not G1205;
	I2808<= not G1161;
	I2811<= not G1209;
	I2814<= not G1222;
	I2817<= not G1222;
	I2821<= not G1221;
	I2825<= not G1143;
	I2828<= not G1193;
	I2831<= not G1209;
	I2835<= not G1209;
	I2839<= not G1123;
	I2842<= not G1177;
	I2845<= not G1193;
	I2848<= not G1193;
	I2854<= not G1236;
	I2857<= not G1161;
	I2860<= not G1177;
	I2864<= not G1177;
	I2867<= not G1143;
	I2870<= not G1161;
	I2873<= not G1161;
	I2877<= not G1123;
	I2880<= not G1143;
	I2883<= not G1143;
	I2887<= not G1123;
	I2890<= not G1123;
	I2893<= not G1236;
	I2904<= not G1256;
	I2907<= not G1498;
	I2910<= not G1645;
	I2913<= not G1792;
	I2916<= not G1643;
	I2919<= not G1787;
	I2922<= not G1774;
	I2925<= not G1762;
	I2929<= not G1659;
	I2940<= not G1653;
	I2943<= not G1715;
	I2946<= not G1587;
	I2949<= not G1263;
	I2952<= not G1594;
	I2955<= not G1729;
	I2958<= not G1257;
	I2961<= not G1731;
	I2964<= not G1257;
	I2967<= not G1682;
	I2970<= not G1504;
	I2973<= not G1687;
	I2979<= not G1263;
	I2982<= not G1426;
	I2986<= not G1504;
	I2989<= not G1519;
	I2992<= not G1741;
	I2995<= not G1742;
	I2998<= not G1257;
	I3001<= not G1267;
	I3004<= not G1426;
	I3007<= not G1439;
	I3010<= not G1504;
	I3013<= not G1519;
	I3016<= not G1754;
	I3019<= not G1755;
	I3022<= not G1426;
	I3025<= not G1439;
	I3028<= not G1504;
	I3031<= not G1504;
	I3034<= not G1519;
	I3037<= not G1769;
	I3040<= not G1770;
	I3044<= not G1257;
	I3047<= not G1426;
	I3050<= not G1439;
	I3053<= not G1407;
	I3056<= not G1519;
	I3059<= not G1519;
	I3062<= not G1776;
	I3065<= not G1426;
	I3068<= not G1439;
	I3071<= not G1504;
	I3074<= not G1426;
	I3077<= not G1439;
	I3080<= not G1519;
	I3083<= not G1426;
	I3086<= not G1439;
	I3090<= not G1504;
	I3093<= not G1426;
	I3096<= not G1439;
	I3099<= not G1519;
	I3102<= not G1426;
	I3105<= not G1439;
	I3109<= not G1504;
	I3112<= not G1439;
	I3115<= not G1519;
	I3134<= not G1336;
	I3137<= not G1315;
	I3140<= not G1317;
	I3144<= not G1319;
	I3148<= not G1595;
	I3152<= not G1322;
	I3155<= not G1612;
	I3158<= not G1829;
	I3161<= not G1270;
	I3198<= not G1819;
	I3202<= not G1812;
	I3206<= not G1823;
	I3212<= not G1806;
	I3215<= not G1820;
	I3222<= not G1790;
	I3225<= not G1813;
	I3232<= not G1782;
	I3235<= not G1807;
	I3240<= not G1460;
	I3244<= not G1772;
	I3247<= not G1791;
	I3251<= not G1471;
	I3255<= not G1650;
	I3258<= not G1760;
	I3261<= not G1783;
	I3268<= not G1656;
	I3271<= not G1748;
	I3274<= not G1773;
	I3278<= not G1695;
	I3281<= not G1761;
	I3284<= not G1702;
	I3288<= not G1710;
	I3291<= not G1714;
	I3294<= not G1720;
	I3298<= not G1725;
	I3301<= not G1730;
	I3304<= not G1740;
	I3307<= not G1339;
	I3310<= not G1640;
	I3313<= not G1337;
	I3316<= not G1344;
	I3319<= not G1636;
	I3322<= not G1333;
	I3325<= not G1340;
	I3328<= not G1273;
	I3331<= not G1631;
	I3334<= not G1330;
	I3337<= not G1338;
	I3340<= not G1282;
	I3343<= not G1623;
	I3346<= not G1327;
	I3349<= not G1334;
	I3352<= not G1285;
	I3355<= not G1608;
	I3358<= not G1323;
	I3361<= not G1331;
	I3364<= not G1648;
	I3367<= not G1283;
	I3370<= not G1805;
	I3373<= not G1320;
	I3376<= not G1328;
	I3379<= not G1647;
	I3382<= not G1284;
	I3385<= not G1318;
	I3388<= not G1324;
	I3391<= not G1646;
	I3395<= not G1286;
	I3405<= not G1321;
	I3408<= not G1644;
	I3419<= not G1287;
	I3422<= not G1641;
	I3425<= not G1274;
	I3428<= not G1825;
	I3431<= not G1275;
	I3434<= not G1627;
	I3441<= not G1502;
	I3452<= not G1450;
	I3462<= not G1450;
	I3465<= not G1724;
	I3468<= not G1802;
	I3471<= not G1450;
	I3474<= not G1450;
	I3478<= not G1450;
	I3481<= not G1461;
	I3485<= not G1450;
	I3488<= not G1295;
	I3493<= not G1461;
	I3496<= not G1326;
	I3499<= not G1450;
	I3502<= not G1295;
	I3505<= not G1305;
	I3509<= not G1461;
	I3513<= not G1450;
	I3516<= not G1295;
	I3519<= not G1305;
	I3522<= not G1664;
	I3525<= not G1461;
	I3528<= not G1422;
	I3531<= not G1593;
	I3534<= not G1295;
	I3537<= not G1305;
	I3540<= not G1670;
	I3543<= not G1461;
	I3546<= not G1586;
	I3550<= not G1295;
	I3553<= not G1305;
	I3556<= not G1484;
	I3560<= not G1673;
	I3563<= not G1461;
	I3569<= not G1789;
	I3572<= not G1295;
	I3575<= not G1305;
	I3578<= not G1484;
	I3581<= not G1491;
	I3584<= not G1678;
	I3587<= not G1461;
	I3590<= not G1781;
	I3593<= not G1295;
	I3596<= not G1305;
	I3599<= not G1484;
	I3602<= not G1491;
	I3605<= not G1681;
	I3608<= not G1461;
	I3611<= not G1771;
	I3614<= not G1295;
	I3617<= not G1305;
	I3620<= not G1484;
	I3623<= not G1491;
	I3626<= not G1684;
	I3629<= not G1759;
	I3632<= not G1295;
	I3635<= not G1305;
	I3638<= not G1484;
	I3641<= not G1491;
	I3644<= not G1685;
	I3647<= not G1747;
	I3650<= not G1650;
	I3653<= not G1305;
	I3656<= not G1484;
	I3659<= not G1491;
	I3662<= not G1688;
	I3665<= not G1824;
	I3669<= not G1739;
	I3672<= not G1656;
	I3675<= not G1491;
	I3678<= not G1690;
	I3681<= not G1821;
	I3684<= not G1733;
	I3687<= not G1814;
	I3691<= not G1732;
	I3694<= not G1811;
	I3705<= not G2316;
	I3708<= not G1946;
	I3711<= not G1848;
	I3714<= not G1852;
	I3717<= not G2154;
	I3720<= not G2155;
	I3723<= not G2158;
	I3726<= not G2030;
	I3729<= not G2436;
	I3733<= not G2031;
	I3736<= not G2460;
	I3746<= not G2035;
	I3749<= not G2484;
	I3752<= not G2044;
	I3755<= not G2125;
	I3758<= not G2041;
	I3761<= not G2505;
	I3764<= not G2044;
	I3767<= not G2125;
	I3770<= not G2145;
	I3773<= not G2524;
	I3776<= not G2044;
	I3779<= not G2125;
	I3782<= not G2145;
	I3785<= not G2346;
	I3788<= not G2554;
	I3791<= not G2044;
	I3794<= not G2044;
	I3797<= not G2125;
	I3800<= not G2145;
	I3804<= not G2575;
	I3808<= not G2125;
	I3811<= not G2145;
	I3816<= not G2580;
	I3819<= not G2044;
	I3823<= not G2125;
	I3826<= not G2145;
	I3830<= not G2179;
	I3833<= not G2266;
	I3836<= not G1832;
	I3840<= not G2125;
	I3843<= not G2145;
	I3855<= not G2550;
	I3858<= not G2197;
	I3861<= not G1834;
	I3864<= not G2044;
	I3868<= not G2125;
	I3871<= not G2145;
	I3883<= not G2574;
	I3886<= not G2215;
	I3890<= not G2145;
	I3902<= not G2576;
	I3906<= not G2234;
	I3909<= not G2044;
	I3923<= not G2581;
	I3927<= not G2245;
	I3942<= not G1833;
	I3946<= not G2256;
	I3961<= not G1835;
	I3965<= not G2268;
	I3979<= not G1836;
	I3983<= not G2276;
	I3999<= not G1837;
	I4003<= not G2284;
	I4019<= not G1841;
	I4023<= not G2315;
	I4031<= not G1846;
	I4050<= not G2059;
	I4059<= not G1878;
	I4066<= not G2582;
	I4123<= not G2043;
	I4133<= not G2040;
	I4166<= not G2390;
	I4170<= not G2157;
	I4173<= not G2408;
	I4176<= not G2268;
	I4189<= not G2159;
	I4192<= not G1847;
	I4195<= not G2173;
	I4198<= not G2276;
	I4217<= not G2163;
	I4220<= not G2164;
	I4223<= not G2176;
	I4226<= not G2525;
	I4229<= not G2284;
	I4240<= not G2165;
	I4243<= not G1853;
	I4246<= not G2194;
	I4249<= not G2525;
	I4252<= not G2555;
	I4255<= not G2179;
	I4258<= not G2169;
	I4261<= not G1857;
	I4264<= not G2212;
	I4267<= not G2525;
	I4270<= not G2555;
	I4273<= not G2197;
	I4276<= not G2170;
	I4279<= not G2230;
	I4282<= not G2525;
	I4285<= not G2555;
	I4288<= not G2215;
	I4291<= not G2241;
	I4294<= not G2525;
	I4297<= not G2555;
	I4300<= not G2234;
	I4303<= not G1897;
	I4306<= not G1898;
	I4309<= not G2525;
	I4312<= not G2555;
	I4315<= not G2245;
	I4318<= not G2171;
	I4321<= not G1917;
	I4324<= not G1918;
	I4327<= not G2525;
	I4331<= not G2555;
	I4334<= not G2256;
	I4337<= not G1934;
	I4340<= not G1935;
	I4343<= not G2525;
	I4347<= not G2555;
	I4351<= not G2233;
	I4354<= not G1953;
	I4358<= not G2525;
	I4362<= not G2555;
	I4366<= not G2244;
	I4371<= not G2555;
	I4375<= not G2254;
	I4382<= not G2265;
	I4391<= not G2275;
	I4398<= not G2086;
	I4402<= not G2283;
	I4410<= not G2088;
	I4414<= not G2090;
	I4420<= not G2096;
	I4424<= not G2097;
	I4429<= not G2102;
	I4433<= not G2103;
	I4437<= not G2108;
	I4441<= not G2109;
	I4452<= not G2117;
	I4455<= not G2118;
	I4459<= not G2134;
	I4462<= not G2135;
	I4465<= not G2945;
	I4468<= not G2583;
	I4471<= not G3040;
	I4474<= not G3052;
	I4477<= not G3063;
	I4480<= not G3073;
	I4483<= not G3082;
	I4486<= not G3093;
	I4489<= not G2975;
	I4492<= not G3001;
	I4495<= not G3022;
	I4498<= not G2686;
	I4501<= not G2705;
	I4504<= not G2726;
	I4507<= not G2739;
	I4510<= not G2753;
	I4513<= not G2765;
	I4516<= not G2777;
	I4519<= not G2788;
	I4522<= not G2801;
	I4534<= not G2858;
	I4537<= not G2877;
	I4587<= not G2962;
	I4593<= not G2966;
	I4623<= not G2962;
	I4646<= not G2602;
	I4664<= not G2924;
	I4667<= not G2908;
	I4671<= not G2928;
	I4678<= not G2670;
	I4681<= not G2947;
	I4684<= not G2687;
	I4688<= not G3207;
	I4706<= not G2877;
	I4743<= not G2594;
	I4752<= not G2859;
	I4757<= not G2861;
	I4762<= not G2862;
	I4777<= not G2962;
	I4791<= not G2814;
	I4794<= not G2814;
	I4799<= not G2967;
	I4802<= not G2877;
	I4809<= not G2974;
	I4821<= not G2877;
	I4903<= not G3223;
	I4935<= not G3369;
	I4955<= not G3673;
	I4961<= not G3597;
	I4964<= not G3673;
	I4976<= not G3575;
	I4980<= not G3546;
	I4986<= not G3638;
	I5002<= not G3612;
	I5006<= not G3604;
	I5019<= not G3318;
	I5023<= not G3263;
	I5027<= not G3267;
	I5030<= not G3242;
	I5033<= not G3527;
	I5037<= not G3705;
	I5040<= not G3271;
	I5043<= not G3247;
	I5050<= not G3246;
	I5053<= not G3710;
	I5056<= not G3567;
	I5059<= not G3259;
	I5065<= not G3714;
	I5068<= not G3571;
	I5071<= not G3263;
	I5078<= not G3719;
	I5081<= not G3589;
	I5084<= not G3593;
	I5091<= not G3242;
	I5094<= not G3705;
	I5103<= not G3440;
	I5106<= not G3247;
	I5109<= not G3710;
	I5116<= not G3259;
	I5119<= not G3714;
	I5124<= not G3719;
	I5148<= not G3450;
	I5153<= not G3330;
	I5157<= not G3454;
	I5169<= not G3593;
	I5177<= not G3267;
	I5182<= not G3271;
	I5204<= not G3534;
	I5214<= not G3567;
	I5217<= not G3673;
	I5223<= not G3537;
	I5233<= not G3571;
	I5236<= not G3545;
	I5249<= not G3589;
	I5252<= not G3546;
	I5264<= not G3638;
	I5316<= not G3557;
	I5320<= not G3559;
	I5324<= not G3466;
	I5328<= not G3502;
	I5333<= not G3491;
	I5337<= not G3564;
	I5343<= not G3599;
	I5376<= not G4014;
	I5379<= not G3940;
	I5382<= not G3952;
	I5385<= not G3962;
	I5388<= not G3969;
	I5391<= not G3975;
	I5394<= not G4016;
	I5397<= not G3932;
	I5400<= not G3963;
	I5403<= not G3970;
	I5406<= not G3976;
	I5409<= not G3980;
	I5412<= not G4034;
	I5415<= not G3723;
	I5418<= not G4036;
	I5421<= not G3724;
	I5424<= not G3725;
	I5427<= not G3726;
	I5430<= not G3727;
	I5433<= not G3728;
	I5436<= not G3729;
	I5439<= not G3730;
	I5442<= not G3731;
	I5445<= not G4040;
	I5448<= not G3960;
	I5451<= not G3967;
	I5454<= not G3874;
	I5457<= not G3766;
	I5460<= not G3771;
	I5463<= not G3783;
	I5466<= not G3787;
	I5469<= not G3838;
	I5472<= not G3846;
	I5475<= not G3852;
	I5478<= not G3859;
	I5481<= not G3866;
	I5484<= not G3875;
	I5487<= not G3881;
	I5490<= not G3832;
	I5493<= not G3834;
	I5496<= not G3839;
	I5499<= not G3847;
	I5502<= not G3853;
	I5505<= not G3860;
	I5508<= not G3867;
	I5511<= not G3876;
	I5514<= not G3882;
	I5517<= not G3885;
	I5520<= not G3835;
	I5523<= not G3840;
	I5526<= not G3848;
	I5529<= not G3854;
	I5532<= not G3861;
	I5542<= not G3984;
	I5545<= not G3814;
	I5548<= not G4059;
	I5551<= not G4059;
	I5556<= not G4059;
	I5562<= not G4002;
	I5568<= not G3897;
	I5577<= not G4022;
	I5591<= not G3821;
	I5594<= not G3821;
	I5597<= not G3821;
	I5600<= not G3821;
	I5603<= not G3893;
	I5606<= not G3821;
	I5609<= not G3893;
	I5612<= not G3910;
	I5615<= not G3914;
	I5618<= not G3821;
	I5622<= not G3914;
	I5626<= not G3914;
	I5630<= not G3914;
	I5633<= not G3768;
	I5637<= not G3914;
	I5640<= not G3770;
	I5644<= not G4059;
	I5654<= not G3742;
	I5668<= not G3828;
	I5674<= not G4003;
	I5686<= not G3942;
	I5692<= not G3942;
	I5696<= not G3942;
	I5699<= not G3844;
	I5702<= not G3845;
	I5705<= not G3942;
	I5708<= not G3942;
	I5713<= not G4022;
	I5716<= not G3942;
	I5720<= not G4022;
	I5723<= not G3942;
	I5728<= not G4022;
	I5731<= not G3942;
	I5736<= not G4022;
	I5739<= not G3942;
	I5743<= not G4022;
	I5746<= not G4022;
	I5750<= not G4022;
	I5753<= not G4022;
	I5756<= not G3922;
	I5774<= not G3807;
	I5777<= not G3807;
	I5790<= not G3803;
	I5793<= not G3803;
	I5825<= not G3914;
	I5831<= not G3842;
	I5837<= not G3850;
	I5840<= not G3732;
	I5843<= not G3851;
	I5848<= not G3856;
	I5851<= not G3739;
	I5854<= not G3857;
	I5857<= not G3740;
	I5862<= not G3863;
	I5865<= not G3743;
	I5868<= not G3864;
	I5871<= not G3744;
	I5876<= not G3870;
	I5879<= not G3745;
	I5882<= not G3871;
	I5885<= not G3746;
	I5890<= not G3878;
	I5893<= not G3747;
	I5896<= not G3879;
	I5899<= not G3748;
	I5904<= not G3749;
	I5907<= not G3883;
	I5910<= not G3750;
	I5913<= not G3751;
	I5920<= not G4228;
	I5923<= not G4299;
	I5926<= not G4153;
	I5929<= not G4152;
	I5933<= not G4346;
	I5938<= not G4351;
	I5944<= not G4356;
	I5948<= not G4360;
	I5952<= not G4367;
	I5977<= not G4319;
	I5987<= not G4224;
	I5991<= not G4226;
	I5998<= not G4157;
	I6001<= not G4162;
	I6004<= not G4159;
	I6008<= not G4163;
	I6012<= not G4167;
	I6015<= not G4170;
	I6020<= not G4176;
	I6023<= not G4151;
	I6033<= not G4179;
	I6036<= not G4370;
	I6039<= not G4182;
	I6042<= not G4374;
	I6045<= not G4375;
	I6048<= not G4376;
	I6051<= not G4185;
	I6054<= not G4194;
	I6057<= not G4379;
	I6060<= not G4380;
	I6063<= not G4381;
	I6066<= not G4382;
	I6069<= not G4213;
	I6072<= not G4385;
	I6075<= not G4386;
	I6078<= not G4387;
	I6081<= not G4388;
	I6084<= not G4391;
	I6087<= not G4392;
	I6090<= not G4393;
	I6093<= not G4394;
	I6096<= not G4397;
	I6099<= not G4398;
	I6102<= not G4399;
	I6105<= not G4400;
	I6108<= not G4403;
	I6111<= not G4404;
	I6114<= not G4405;
	I6118<= not G4406;
	I6126<= not G4240;
	I6132<= not G4219;
	I6139<= not G4222;
	I6143<= not G4237;
	I6170<= not G4343;
	I6182<= not G4249;
	I6231<= not G4350;
	I6244<= not G4519;
	I6247<= not G4609;
	I6250<= not G4514;
	I6253<= not G4608;
	I6269<= not G4655;
	I6280<= not G4430;
	I6283<= not G4613;
	I6289<= not G4433;
	I6292<= not G4434;
	I6296<= not G4436;
	I6299<= not G4438;
	I6302<= not G4440;
	I6305<= not G4441;
	I6308<= not G4443;
	I6311<= not G4444;
	I6315<= not G4446;
	I6318<= not G4447;
	I6321<= not G4559;
	I6324<= not G4450;
	I6327<= not G4451;
	I6330<= not G4560;
	I6334<= not G4454;
	I6337<= not G4455;
	I6340<= not G4561;
	I6343<= not G4458;
	I6346<= not G4563;
	I6349<= not G4569;
	I6352<= not G4564;
	I6355<= not G4569;
	I6359<= not G4566;
	I6362<= not G4569;
	I6366<= not G4569;
	I6371<= not G4569;
	I6377<= not G4569;
	I6382<= not G4460;
	I6386<= not G4462;
	I6397<= not G4473;
	I6400<= not G4473;
	I6403<= not G4492;
	I6406<= not G4473;
	I6410<= not G4473;
	I6414<= not G4497;
	I6417<= not G4617;
	I6420<= not G4618;
	I6425<= not G4619;
	I6430<= not G4620;
	I6434<= not G4622;
	I6437<= not G4501;
	I6441<= not G4624;
	I6444<= not G4503;
	I6448<= not G4626;
	I6452<= not G4629;
	I6456<= not G4633;
	I6464<= not G4562;
	I6470<= not G4473;
	I6485<= not G4603;
	I6488<= not G4603;
	I6495<= not G4607;
	I6507<= not G4644;
	I6525<= not G4770;
	I6528<= not G4815;
	I6531<= not G4704;
	I6534<= not G4706;
	I6537<= not G4711;
	I6540<= not G4714;
	I6543<= not G4718;
	I6546<= not G4692;
	I6549<= not G4699;
	I6552<= not G4702;
	I6555<= not G4703;
	I6558<= not G4705;
	I6561<= not G4707;
	I6564<= not G4712;
	I6567<= not G4715;
	I6570<= not G4719;
	I6573<= not G4721;
	I6576<= not G4700;
	I6579<= not G4798;
	I6582<= not G4765;
	I6587<= not G4803;
	I6599<= not G4823;
	I6607<= not G4745;
	I6612<= not G4660;
	I6615<= not G4745;
	I6621<= not G4745;
	I6625<= not G4745;
	I6630<= not G4745;
	I6635<= not G4745;
	I6646<= not G4687;
	I6649<= not G4693;
	I6666<= not G4740;
	I6672<= not G4752;
	I6677<= not G4757;
	I6680<= not G4713;
	I6685<= not G4716;
	I6689<= not G4758;
	I6692<= not G4720;
	I6697<= not G4722;
	I6701<= not G4726;
	I6706<= not G4731;
	I6723<= not G4761;
	I6733<= not G4773;
	I6737<= not G4662;
	I6740<= not G4781;
	I6750<= not G4771;
	I6753<= not G4772;
	I6756<= not G4775;
	I6759<= not G4778;
	I6763<= not G4780;
	I6766<= not G4783;
	I6769<= not G4786;
	I6772<= not G4788;
	I6775<= not G4790;
	I6780<= not G4825;
	I6783<= not G4822;
	I6786<= not G4824;
	I6789<= not G4871;
	I6792<= not G5097;
	I6795<= not G5022;
	I6798<= not G5042;
	I6801<= not G5045;
	I6809<= not G5051;
	I6812<= not G5110;
	I6816<= not G5111;
	I6819<= not G5019;
	I6867<= not G5082;
	I6874<= not G4861;
	I6885<= not G4872;
	I6895<= not G5010;
	I6918<= not G5124;
	I6923<= not G5124;
	I6927<= not G5124;
	I6930<= not G5017;
	I6933<= not G5124;
	I6937<= not G5124;
	I6942<= not G5124;
	I6946<= not G5124;
	I6949<= not G5050;
	I6952<= not G5124;
	I6956<= not G5124;
	I6959<= not G5089;
	I6972<= not G5135;
	I6976<= not G5136;
	I6986<= not G5230;
	I6989<= not G5307;
	I6992<= not G5151;
	I6995<= not G5220;
	I7002<= not G5308;
	I7007<= not G5314;
	I7012<= not G5316;
	I7029<= not G5149;
	I7035<= not G5150;
	I7039<= not G5309;
	I7042<= not G5310;
	I7045<= not G5167;
	I7051<= not G5219;
	I7055<= not G5318;
	I7058<= not G5281;
	I7061<= not G5281;
	I7065<= not G5281;
	I7069<= not G5281;
	I7073<= not G5281;
	I7077<= not G5281;
	I7081<= not G5281;
	I7086<= not G5281;
	I7091<= not G5281;
	I7104<= not G5273;
	I7107<= not G5277;
	I7110<= not G5291;
	I7113<= not G5295;
	I7116<= not G5299;
	I7119<= not G5303;
	I7143<= not G5323;
	I7146<= not G5231;
	I7150<= not G5355;
	I7153<= not G5358;
	I7161<= not G5465;
	I7164<= not G5433;
	I7167<= not G5434;
	I7170<= not G5435;
	I7173<= not G5436;
	I7176<= not G5437;
	I7187<= not G5387;
	I7190<= not G5432;
	I7193<= not G5466;
	I7197<= not G5431;
	I7251<= not G5458;
	I7254<= not G5458;
	I7258<= not G5458;
	I7261<= not G5458;
	I7264<= not G5458;
	I7267<= not G5458;
	I7270<= not G5352;
	I7276<= not G5375;
	I7284<= not G5383;
	I7295<= not G5439;
	I7318<= not G5452;
	I7333<= not G5386;
	I7336<= not G5534;
	I7339<= not G5540;
	I7342<= not G5579;
	I7346<= not G5531;
	I7349<= not G5532;
	I7352<= not G5533;
	I7355<= not G5535;
	I7358<= not G5565;
	I7361<= not G5566;
	I7372<= not G5493;
	I7397<= not G5561;
	I7404<= not G5541;
	I7451<= not G5597;
	I7463<= not G5622;
	I7466<= not G5624;
	I7469<= not G5625;
	I7472<= not G5626;
	I7475<= not G5627;
	I7478<= not G5628;
	I7481<= not G5629;
	I7484<= not G5630;
	I7487<= not G5684;
	I7490<= not G5583;
	I7494<= not G5691;
	I7497<= not G5687;
	I7501<= not G5596;
	I7506<= not G5584;
	I7509<= not G5587;
	I7514<= not G5590;
	I7517<= not G5593;
	I7583<= not G5605;
	I7587<= not G5605;
	I7590<= not G5605;
	I7593<= not G5605;
	I7596<= not G5605;
	I7600<= not G5605;
	I7604<= not G5605;
	I7608<= not G5605;
	I7612<= not G5605;
	I7634<= not G5727;
	I7637<= not G5751;
	I7640<= not G5773;
	I7643<= not G5752;
	I7646<= not G5774;
	I7679<= not G5726;
	I7683<= not G5702;
	I7686<= not G5705;
	I7689<= not G5708;
	I7692<= not G5711;
	I7695<= not G5714;
	I7698<= not G5717;
	I7701<= not G5720;
	I7704<= not G5723;
	I7707<= not G5701;
	I7796<= not G5917;
	I7799<= not G5918;
	I7802<= not G5920;
	I7805<= not G5923;
	I7808<= not G5919;
	I7811<= not G5921;
	I7814<= not G5922;
	I7817<= not G5924;
	I7829<= not G5926;
	I7832<= not G5943;
	I7835<= not G5926;
	I7838<= not G5947;
	I7852<= not G5993;
	I7856<= not G5994;
	I7859<= not G6032;
	I7865<= not G6095;
	I7871<= not G6097;
	I7892<= not G5916;
	I7906<= not G5912;
	I7910<= not G5905;
	I7960<= not G5925;
	I7963<= not G6276;
	I7966<= not G6166;
	I7996<= not G6137;
	I7999<= not G6137;
	I8002<= not G6110;
	I8005<= not G6110;
	I8027<= not G6237;
	I8030<= not G6239;
	I8034<= not G6242;
	I8040<= not G6142;
	I8044<= not G6252;
	I8051<= not G6108;
	I8056<= not G6109;
	I8061<= not G6113;
	I8066<= not G6114;
	I8070<= not G6116;
	I8074<= not G6118;
	I8089<= not G6120;
	I8093<= not G6122;
	I8103<= not G6134;
	I8107<= not G6136;
	I8110<= not G6143;
	I8113<= not G6147;
	I8144<= not G6182;
	I8147<= not G6182;
	I8150<= not G6185;
	I8153<= not G6185;
	I8156<= not G6167;
	I8159<= not G6167;
	I8162<= not G6189;
	I8165<= not G6189;
	I8168<= not G6170;
	I8171<= not G6170;
	I8174<= not G6173;
	I8177<= not G6173;
	I8180<= not G6176;
	I8183<= not G6176;
	I8186<= not G6179;
	I8189<= not G6179;
	I8217<= not G6319;
	I8220<= not G6322;
	I8223<= not G6325;
	I8226<= not G6328;
	I8229<= not G6330;
	I8232<= not G6332;
	I8235<= not G6312;
	I8240<= not G6287;
	I8243<= not G6286;
	I8246<= not G6290;
	I8249<= not G6289;
	I8252<= not G6294;
	I8255<= not G6292;
	I8258<= not G6293;
	I8261<= not G6298;
	I8264<= not G6296;
	I8267<= not G6297;
	I8270<= not G6300;
	I8273<= not G6301;
	I8276<= not G6303;
	I8279<= not G6307;
	I8282<= not G6309;
	I8285<= not G6310;
	I8290<= not G6291;
	I8295<= not G6295;
	I8300<= not G6299;
	I8309<= not G6304;
	I8329<= not G6305;
	I8332<= not G6306;
	I8335<= not G6308;
	I8342<= not G6314;
	I8411<= not G6415;
	I8414<= not G6418;
	I8417<= not G6420;
	I8420<= not G6422;
	I8423<= not G6423;
	I8426<= not G6424;
	I8429<= not G6425;
	I8432<= not G6411;
	I8435<= not G6413;
	I8438<= not G6416;
	I8441<= not G6419;
	I8444<= not G6421;
	I8447<= not G6410;
	I8450<= not G6412;
	I8453<= not G6414;
	I8456<= not G6417;
	I8459<= not G6427;
	I8462<= not G6430;
	I8467<= not G6457;
	I8470<= not G6461;
	I8473<= not G6485;
	I8476<= not G6457;
	I8479<= not G6482;
	I8482<= not G6461;
	I8485<= not G6479;
	I8488<= not G6426;
	I8491<= not G6480;
	I8494<= not G6428;
	I8497<= not G6481;
	I8500<= not G6431;
	I8503<= not G6434;
	I8506<= not G6483;
	I8509<= not G6437;
	I8512<= not G6441;
	I8515<= not G6492;
	I8518<= not G6494;
	I8521<= not G6495;
	I8524<= not G6496;
	I8527<= not G6440;
	I8531<= not G6444;
	I8535<= not G6447;
	I8538<= not G6450;
	I8541<= not G6452;
	I8544<= not G6453;
	I8548<= not G6454;
	I8552<= not G6455;
	I8555<= not G6456;
	I8564<= not G6429;
	I8567<= not G6432;
	I8570<= not G6433;
	I8573<= not G6435;
	I8576<= not G6436;
	I8579<= not G6438;
	I8582<= not G6439;
	I8585<= not G6442;
	I8588<= not G6443;
	I8591<= not G6448;
	I8594<= not G6446;
	I8597<= not G6445;
	I8600<= not G6451;
	I8603<= not G6449;
	I8614<= not G6537;
	I8617<= not G6539;
	I8620<= not G6541;
	I8623<= not G6542;
	I8626<= not G6543;
	I8629<= not G6544;
	I8632<= not G6548;
	I8635<= not G6552;
	I8638<= not G6553;
	I8641<= not G6524;
	I8644<= not G6526;
	I8647<= not G6528;
	I8650<= not G6529;
	I8653<= not G6531;
	I8656<= not G6532;
	I8659<= not G6523;
	I8662<= not G6525;
	I8665<= not G6527;
	I8668<= not G6530;
	I8671<= not G6519;
	I8674<= not G6521;
	I8678<= not G6565;
	I8681<= not G6566;
	I8684<= not G6567;
	I8687<= not G6568;
	I8690<= not G6571;
	I8693<= not G6570;
	I8696<= not G6569;
	I8699<= not G6573;
	I8702<= not G6572;
	I8707<= not G6520;
	I8710<= not G6517;
	I8713<= not G6522;
	I8716<= not G6518;
	I8721<= not G6534;
	I8724<= not G6533;
	I8727<= not G6536;
	I8730<= not G6535;
	I8745<= not G6513;
	I8749<= not G6560;
	I8752<= not G6514;
	I8755<= not G6561;
	I8758<= not G6562;
	I8761<= not G6563;
	I8764<= not G6564;
	I8767<= not G6619;
	I8800<= not G6684;
	I8803<= not G6685;
	I8806<= not G6686;
	I8809<= not G6687;
	I8812<= not G6688;
	I8815<= not G6689;
	I8818<= not G6690;
	I8821<= not G6691;
	I8828<= not G6661;
	I8831<= not G6665;
	I8834<= not G6661;
	I8837<= not G6665;
	I8840<= not G6657;
	I8843<= not G6658;
	I8854<= not G6696;
	I8857<= not G6698;
	I8860<= not G6699;
	I8863<= not G6700;
	I8866<= not G6701;
	I8869<= not G6694;
	I8872<= not G6695;
	I8875<= not G6697;
	I8878<= not G6710;
	I8881<= not G6711;
	I8884<= not G6704;
	I8888<= not G6708;
	I8891<= not G6706;
	I8894<= not G6709;
	I8897<= not G6707;
	I8907<= not G6702;
	I8910<= not G6730;
	I8913<= not G6743;
	I8916<= not G6742;
	I8940<= not G6783;
	I8943<= not G6774;
	I8946<= not G6778;
	I8958<= not G6774;
	I8961<= not G6778;
	I8966<= not G6796;
	I8969<= not G6797;
	I8972<= not G6795;
	I8975<= not G6791;
	I8978<= not G6792;
	I8981<= not G6793;
	I8984<= not G6794;
	I8988<= not G6787;
	I8991<= not G6788;
	I8994<= not G6789;
	I8997<= not G6790;
	I9002<= not G6802;
	I9005<= not G6817;
	I9008<= not G6818;
	I9011<= not G6819;
	I9014<= not G6820;
	I9021<= not G6812;
	I9024<= not G6803;
	I9028<= not G6806;
	I9031<= not G6809;
	I9035<= not G6812;
	I9038<= not G6833;
	I9041<= not G6835;
	I9044<= not G6836;
	I9047<= not G6838;
	I9074<= not G6844;
	I9077<= not G6845;
	I9082<= not G6849;
	I9085<= not G6850;
	I9092<= not G6855;
	I9095<= not G6855;
	I9098<= not G6864;
	I9101<= not G6855;
	I9104<= not G6864;
	I9107<= not G6855;
	I9110<= not G6864;
	I9113<= not G6855;
	I9116<= not G6864;
	I9119<= not G6855;
	I9122<= not G6864;
	I9125<= not G6855;
	I9128<= not G6864;
	I9131<= not G6855;
	I9134<= not G6864;
	I9137<= not G6864;
	I9140<= not G6888;
	I9143<= not G6886;
	I9146<= not G6890;
	I9149<= not G6884;
	I9152<= not G6889;
	I9155<= not G6882;
	I9158<= not G6887;
	I9161<= not G6880;
	I9164<= not G6885;
	I9167<= not G6878;
	I9170<= not G6883;
	I9173<= not G6876;
	I9176<= not G6881;
	I9179<= not G6875;
	I9182<= not G6879;
	I9185<= not G6877;
	I9203<= not G6921;
	I9208<= not G6922;
	I9217<= not G6931;
	I9220<= not G6930;
	I9227<= not G6937;
	I9230<= not G6936;
	I9233<= not G6938;
	I9236<= not G6939;
	G918<=G610 and G602;
	G1027<=G598 and G567;
	G1407<=G301 and G866;
	G1416<=G913 and G266;
	G1419<=G613 and G918;
	G1436<=G834 and G830;
	G1499<=G1101 and G1094;
	G1514<=G1017 and G1011;
	G1570<=G634 and G1027;
	G1575<=G980 and G965;
	G1576<=G1101 and G1094;
	G1585<=G1017 and G1011;
	G1595<=G729 and G719 and G766 and I2566;
	G1609<=G760 and G754;
	G1612<=G784 and G774 and G821 and I2574;
	G1620<=G1056 and G1084;
	G1628<=G815 and G809;
	G1633<=G716 and G152;
	G1689<=G766 and G719;
	G1691<=G821 and G774;
	G1706<=G766 and G719 and G729;
	G1716<=G821 and G774 and G784;
	G1763<=G478 and G1119;
	G1784<=G858 and G889;
	G1802<=G89 and G1064;
	G1808<=G706 and G49;
	G1826<=G714 and G710;
	G2015<=G616 and G1419;
	G2018<=G1423 and G1254;
	G2021<=G835 and G1436;
	G2026<=G1359 and G1402 and G1398 and G901;
	G2053<=G1094 and G1675;
	G2056<=G1672 and G1675;
	G2062<=G1499 and G1666;
	G2068<=G1541 and G1546;
	G2073<=G1088 and G1499;
	G2081<=G1094 and G1546;
	G2084<=G1577 and G1563;
	G2085<=G1123 and G1567;
	G2089<=G1123 and G1578;
	G2092<=G642 and G1570;
	G2101<=G1001 and G1543;
	G2107<=G1583 and G1543;
	G2113<=G1576 and G1535;
	G2121<=G1632 and G754;
	G2137<=G760 and G1638;
	G2138<=G1639 and G809;
	G2142<=G1793 and G1777;
	G2156<=G815 and G1642;
	G2160<=G1624 and G929;
	G2166<=G1633 and G161;
	G2255<=G1706 and G736;
	G2267<=G1716 and G791;
	G2292<=G1706 and G736 and G743;
	G2294<=G1716 and G791 and G798;
	G2323<=G471 and G1358;
	G2339<=G1603 and G197;
	G2340<=G1398 and G1387;
	G2356<=G1603 and G269;
	G2419<=G1808 and G54;
	G2551<=G715 and G1826;
	G2577<=G1743 and G1797 and G1793 and G1138;
	G2659<=G1686 and G2296;
	G2670<=G2029 and G1503;
	G2671<=G2263 and G2296;
	G2685<=G2370 and G1887;
	G2699<=G2397 and G1905;
	G2700<=G2370 and G1908;
	G2720<=G2422 and G1919;
	G2721<=G2397 and G1922;
	G2732<=G2449 and G1940;
	G2733<=G2422 and G1943;
	G2746<=G2473 and G1954;
	G2747<=G2449 and G1957;
	G2758<=G2497 and G1963;
	G2759<=G2473 and G1966;
	G2770<=G2518 and G1972;
	G2771<=G2497 and G1975;
	G2781<=G2544 and G1982;
	G2782<=G2518 and G1985;
	G2793<=G2568 and G1991;
	G2794<=G2544 and G1994;
	G2807<=G2568 and G2001;
	G2808<=G2009 and G1581;
	G2821<=G1890 and G910;
	G2834<=G1263 and G1257 and G1270 and I4040;
	G2846<=G619 and G2015;
	G2850<=G2018 and G1255;
	G2853<=G836 and G2021;
	G2859<=G2112 and G1649;
	G2860<=G710 and G2296;
	G2861<=G2120 and G1654;
	G2868<=G1316 and G1861;
	G2873<=G1845 and G1861;
	G2897<=G1030 and G2062;
	G2909<=G606 and G2092;
	G2916<=G1030 and G2113;
	G2935<=G2291 and G1788;
	G2937<=G2160 and G931;
	G2941<=G2166 and G170;
	G2948<=G2137 and G1595;
	G2949<=G830 and G1861;
	G2950<=G2156 and G1612;
	G2953<=G2381 and G293;
	G2955<=G2381 and G297;
	G3089<=G212 and G2336;
	G3099<=G218 and G2350;
	G3103<=G212 and G2353;
	G3113<=G224 and G2364;
	G3117<=G218 and G2367;
	G3122<=G2435 and G1394;
	G3123<=G230 and G2391;
	G3127<=G224 and G2394;
	G3132<=G2306 and G1206;
	G3133<=G236 and G2410;
	G3134<=G230 and G2413;
	G3135<=G2370 and G2416;
	G3143<=G242 and G2437;
	G3144<=G236 and G2440;
	G3145<=G2397 and G2443;
	G3146<=G2370 and G2446;
	G3147<=G2419 and G59;
	G3154<=G2039 and G1410;
	G3155<=G248 and G2461;
	G3156<=G242 and G2464;
	G3157<=G2422 and G2467;
	G3161<=G2397 and G2470;
	G3166<=G2042 and G1233;
	G3167<=G1883 and G921;
	G3170<=G254 and G2485;
	G3171<=G248 and G2488;
	G3172<=G2449 and G2491;
	G3176<=G2422 and G2494;
	G3180<=G260 and G2506;
	G3181<=G254 and G2509;
	G3182<=G2473 and G2512;
	G3186<=G2449 and G2515;
	G3190<=G260 and G2535;
	G3191<=G2497 and G2538;
	G3195<=G2473 and G2541;
	G3203<=G2497 and G2565;
	G3208<=G895 and G2551;
	G3275<=G2172 and G2615;
	G3277<=G2174 and G2625;
	G3278<=G2175 and G2628;
	G3279<=G2599 and G2612;
	G3280<=G2177 and G2637;
	G3281<=G2178 and G2640;
	G3282<=G131 and G2863;
	G3283<=G2609 and G2622;
	G3285<=G2195 and G2653;
	G3286<=G2196 and G2656;
	G3287<=G135 and G2865;
	G3288<=G2631 and G2634;
	G3290<=G2213 and G2664;
	G3292<=G2214 and G2667;
	G3293<=G212 and G2864;
	G3294<=G139 and G2870;
	G3295<=G2660 and G2647;
	G3296<=G3054 and G2650;
	G3298<=G2231 and G2679;
	G3300<=G2232 and G2682;
	G3301<=G218 and G2866;
	G3302<=G212 and G2867;
	G3303<=G2722 and G2890;
	G3304<=G2857 and G1513;
	G3305<=G2960 and G2296;
	G3307<=G2242 and G2692;
	G3309<=G2243 and G2695;
	G3310<=G224 and G2871;
	G3311<=G218 and G2872;
	G3315<=G2701 and G1875;
	G3316<=G2748 and G2894;
	G3317<=G2722 and G2895;
	G3319<=G2688 and G2675;
	G3321<=G2252 and G2713;
	G3323<=G2253 and G2716;
	G3324<=G230 and G2875;
	G3325<=G224 and G2876;
	G3326<=G2734 and G1891;
	G3327<=G2772 and G2906;
	G3328<=G2701 and G1894;
	G3329<=G2748 and G2907;
	G3333<=G2264 and G2728;
	G3334<=G236 and G2883;
	G3335<=G230 and G2884;
	G3336<=G2760 and G1911;
	G3337<=G2796 and G2913;
	G3338<=G3162 and G2914;
	G3339<=G2734 and G1914;
	G3340<=G2772 and G2915;
	G3341<=G2998 and G2709;
	G3344<=G242 and G2885;
	G3345<=G236 and G2886;
	G3349<=G2783 and G1925;
	G3350<=G3150 and G1928;
	G3351<=G2760 and G1931;
	G3352<=G2796 and G2920;
	G3353<=G3162 and G2921;
	G3356<=G248 and G2888;
	G3357<=G242 and G2889;
	G3358<=G2842 and G1369;
	G3359<=G2822 and G2922;
	G3360<=G2783 and G1947;
	G3361<=G3150 and G1950;
	G3362<=G3031 and G2740;
	G3365<=G254 and G2892;
	G3366<=G248 and G2893;
	G3367<=G2809 and G1960;
	G3368<=G2822 and G2923;
	G3371<=G260 and G2904;
	G3372<=G254 and G2905;
	G3373<=G3118 and G2927;
	G3374<=G2809 and G1969;
	G3375<=G260 and G2912;
	G3376<=G3104 and G1979;
	G3377<=G3118 and G2931;
	G3378<=G3136 and G2932;
	G3379<=G3104 and G1988;
	G3381<=G3128 and G1998;
	G3382<=G3136 and G2934;
	G3383<=G3128 and G2004;
	G3421<=G622 and G2846;
	G3425<=G2296 and G3208;
	G3433<=G1359 and G2831 and G905;
	G3434<=G2850 and G857;
	G3437<=G837 and G2853;
	G3449<=G128 and G2946;
	G3454<=G2933 and G1660;
	G3464<=G341 and G2956;
	G3479<=G345 and G2957;
	G3484<=G349 and G2958;
	G3489<=G2607 and G1861;
	G3490<=G353 and G2959;
	G3499<=G357 and G2961;
	G3505<=G2924 and G1749;
	G3512<=G2928 and G1764;
	G3522<=G646 and G2909;
	G3551<=G2937 and G938;
	G3554<=G2941 and G179;
	G3558<=G338 and G3199;
	G3602<=G2688 and G2663;
	G3603<=G2370 and G3019;
	G3608<=G2599 and G2308;
	G3609<=G2706 and G2678;
	G3610<=G2397 and G3034;
	G3611<=G2370 and G3037;
	G3613<=G2604 and G2312;
	G3614<=G2998 and G2691;
	G3615<=G2422 and G3046;
	G3616<=G2397 and G3049;
	G3617<=G2609 and G2317;
	G3618<=G3016 and G2712;
	G3619<=G2449 and G3057;
	G3620<=G2422 and G3060;
	G3625<=G2619 and G2320;
	G3626<=G3031 and G2727;
	G3627<=G2473 and G3067;
	G3628<=G2449 and G3070;
	G3629<=G2809 and G2738;
	G3630<=G3167 and G1756;
	G3631<=G2631 and G2324;
	G3632<=G3043 and G2743;
	G3633<=G2497 and G3076;
	G3634<=G2179 and G2744;
	G3635<=G2473 and G3079;
	G3636<=G2701 and G2327;
	G3637<=G2822 and G2752;
	G3641<=G2644 and G2333;
	G3642<=G3054 and G2754;
	G3643<=G2518 and G3086;
	G3644<=G2197 and G2755;
	G3645<=G2497 and G3090;
	G3646<=G2179 and G2756;
	G3648<=G2722 and G2343;
	G3649<=G3104 and G2764;
	G3650<=G2660 and G2347;
	G3651<=G3064 and G2766;
	G3652<=G2544 and G3096;
	G3653<=G2215 and G2767;
	G3654<=G2518 and G3100;
	G3655<=G2197 and G2768;
	G3657<=G2734 and G2357;
	G3658<=G3118 and G2776;
	G3659<=G2672 and G2361;
	G3660<=G2568 and G3110;
	G3661<=G2234 and G2778;
	G3662<=G2544 and G3114;
	G3663<=G2215 and G2779;
	G3665<=G2748 and G2378;
	G3666<=G3128 and G2787;
	G3667<=G2245 and G2789;
	G3668<=G2568 and G3124;
	G3669<=G2234 and G2790;
	G3670<=G2234 and G2792;
	G3671<=G2760 and G2405;
	G3672<=G3136 and G2800;
	G3678<=G2256 and G2802;
	G3679<=G2245 and G2803;
	G3680<=G2245 and G2805;
	G3681<=G2234 and G2806;
	G3682<=G2772 and G2430;
	G3683<=G3150 and G2813;
	G3684<=G2268 and G2817;
	G3685<=G2256 and G2818;
	G3686<=G2256 and G2819;
	G3687<=G2245 and G2820;
	G3688<=G2783 and G2457;
	G3689<=G3162 and G2826;
	G3690<=G2276 and G2827;
	G3691<=G2268 and G2828;
	G3692<=G2268 and G2829;
	G3693<=G2256 and G2830;
	G3694<=G3147 and G64;
	G3697<=G2796 and G2481;
	G3698<=G2284 and G2835;
	G3699<=G2276 and G2836;
	G3700<=G2276 and G2837;
	G3701<=G2268 and G2838;
	G3702<=G2284 and G2839;
	G3703<=G2284 and G2840;
	G3704<=G2276 and G2841;
	G3709<=G2284 and G2845;
	G3718<=G1743 and G3140 and G1157;
	G3724<=G117 and G3251;
	G3725<=G118 and G3251;
	G3726<=G119 and G3251;
	G3727<=G122 and G3251;
	G3728<=G326 and G3441;
	G3729<=G327 and G3441;
	G3730<=G328 and G3441;
	G3731<=G331 and G3441;
	G3755<=G2604 and G3481;
	G3757<=G2619 and G3487;
	G3758<=G545 and G3461;
	G3759<=G2644 and G3498;
	G3760<=G548 and G3465;
	G3762<=G2672 and G3500;
	G3763<=G3064 and G3501;
	G3764<=G551 and G3480;
	G3765<=G554 and G3485;
	G3767<=G2706 and G3504;
	G3768<=G3448 and G1528;
	G3774<=G3016 and G3510;
	G3780<=G3043 and G3519;
	G3784<=G114 and G3251;
	G3806<=G3384 and G2024;
	G3810<=G625 and G3421;
	G3814<=G913 and G3546;
	G3816<=G3434 and G861;
	G3819<=G964 and G3437;
	G3831<=G2330 and G3425;
	G3843<=G2856 and G945 and G3533;
	G3844<=G3540 and G1665;
	G3887<=G3276 and G1861;
	G3899<=G323 and G3441;
	G3907<=G650 and G3522;
	G3910<=G3546 and G1049;
	G3924<=G3505 and G471;
	G3928<=G3512 and G478;
	G3936<=G3551 and G940;
	G3953<=G3554 and G188;
	G3997<=G1250 and G3425 and G2849;
	G4015<=G445 and G3388;
	G4032<=G441 and G3388;
	G4033<=G426 and G3388;
	G4035<=G437 and G3388;
	G4037<=G2896 and G3388;
	G4038<=G430 and G3388;
	G4039<=G402 and G3388;
	G4041<=G461 and G3388;
	G4042<=G406 and G3388;
	G4043<=G457 and G3388;
	G4044<=G410 and G3388;
	G4045<=G3425 and G123;
	G4046<=I5351 and I5352;
	G4047<=G453 and G3388;
	G4048<=G414 and G3388;
	G4050<=I5359 and I5360;
	G4051<=G449 and G3388;
	G4052<=G418 and G3388;
	G4053<=G3387 and G1415;
	G4054<=G3694 and G69;
	G4057<=G422 and G3388;
	G4058<=G3424 and G1246;
	G4156<=G3926 and G2078;
	G4157<=G3830 and G1533;
	G4159<=G370 and G3890;
	G4160<=G3923 and G1345;
	G4161<=G3931 and G2087;
	G4163<=G374 and G3892;
	G4164<=G3958 and G2091;
	G4165<=G3927 and G1352;
	G4167<=G378 and G3898;
	G4168<=G3925 and G1355;
	G4169<=G3966 and G2099;
	G4170<=G382 and G3900;
	G4171<=G3956 and G2104;
	G4172<=G3930 and G1366;
	G4176<=G386 and G3901;
	G4177<=G3933 and G1372;
	G4178<=G3959 and G2110;
	G4179<=G390 and G3902;
	G4180<=G3929 and G2119;
	G4181<=G3939 and G1381;
	G4182<=G394 and G3904;
	G4183<=G3965 and G1391;
	G4184<=G3934 and G2136;
	G4185<=G398 and G3906;
	G4186<=G3973 and G1395;
	G4199<=G628 and G3810;
	G4209<=G3816 and G865;
	G4214<=G1822 and G4045;
	G4219<=G3911 and G1655;
	G4230<=G3756 and G1861;
	G4236<=G654 and G3907;
	G4244<=G1749 and G4004 and G1609;
	G4247<=G1764 and G4007 and G1628;
	G4253<=G1861 and G3819;
	G4271<=G2121 and G1749 and G4004;
	G4277<=G3936 and G942;
	G4280<=G2138 and G1764 and G4007;
	G4333<=G3964 and G3284;
	G4339<=G3971 and G3289;
	G4340<=G3972 and G3291;
	G4341<=G3977 and G3297;
	G4342<=G3978 and G3299;
	G4344<=G3981 and G3306;
	G4345<=G3982 and G3308;
	G4346<=G157 and G3773;
	G4347<=G3986 and G3320;
	G4348<=G3987 and G3322;
	G4349<=G441 and G3775;
	G4351<=G166 and G3776;
	G4352<=G3988 and G3331;
	G4353<=G3989 and G3332;
	G4354<=G437 and G3777;
	G4355<=G430 and G3778;
	G4356<=G175 and G3779;
	G4357<=G3990 and G3342;
	G4358<=G3991 and G3343;
	G4359<=G434 and G3782;
	G4360<=G184 and G3785;
	G4361<=G3995 and G3354;
	G4362<=G3996 and G3355;
	G4363<=G402 and G3786;
	G4367<=G193 and G3788;
	G4368<=G3998 and G3363;
	G4369<=G3999 and G3364;
	G4371<=G461 and G3789;
	G4372<=G406 and G3790;
	G4373<=G4001 and G3370;
	G4377<=G457 and G3791;
	G4378<=G410 and G3792;
	G4383<=G453 and G3796;
	G4384<=G414 and G3797;
	G4389<=G449 and G3798;
	G4390<=G418 and G3799;
	G4395<=G445 and G3800;
	G4396<=G422 and G3801;
	G4401<=G426 and G3802;
	G4407<=G4054 and G74;
	G4410<=G3903 and G1474;
	G4416<=G3905 and G1481;
	G4429<=G923 and G4253 and G2936;
	G4442<=G4239 and G2882;
	G4445<=G4235 and G1854;
	G4448<=G3815 and G4225;
	G4449<=G4266 and G2887;
	G4452<=G3820 and G4227;
	G4453<=G4238 and G1858;
	G4456<=G3829 and G4229;
	G4457<=G4261 and G2902;
	G4459<=G4245 and G1899;
	G4460<=G4218 and G1539;
	G4461<=G4241 and G2919;
	G4464<=G4272 and G1937;
	G4471<=G4253 and G332;
	G4486<=G716 and G4195;
	G4488<=G1633 and G4202;
	G4489<=G2166 and G4206;
	G4490<=G2941 and G4210;
	G4491<=G3554 and G4215;
	G4495<=G3913 and G4292;
	G4501<=G4250 and G1671;
	G4541<=G631 and G4199;
	G4580<=G706 and G4262;
	G4583<=G1808 and G4267;
	G4588<=G2419 and G4273;
	G4592<=G3147 and G4281;
	G4593<=G4277 and G947;
	G4597<=G3694 and G4286;
	G4598<=G1978 and G4253;
	G4600<=G4054 and G4289;
	G4602<=G4407 and G4293;
	G4611<=G3985 and G119 and G4300;
	G4616<=G4231 and G3761;
	G4621<=G3953 and G4364;
	G4648<=G4407 and G79;
	G4661<=G4637 and G4634;
	G4666<=G4630 and G4627;
	G4667<=G4653 and G4651;
	G4668<=G4642 and G4638;
	G4671<=G4645 and G4641;
	G4672<=G4635 and G4631;
	G4673<=G4656 and G4654;
	G4677<=G4652 and G4646;
	G4683<=G4585 and G2066;
	G4684<=G4584 and G1341;
	G4685<=G4591 and G2079;
	G4686<=G4590 and G1348;
	G4687<=G4493 and G1542;
	G4688<=G1474 and G4568;
	G4691<=G4581 and G2098;
	G4694<=G1481 and G4578;
	G4697<=G4589 and G1363;
	G4698<=G4586 and G2106;
	G4701<=G4596 and G1378;
	G4708<=G578 and G4541;
	G4730<=G1423 and G4565;
	G4735<=G2018 and G4577;
	G4739<=G2850 and G4579;
	G4744<=G3434 and G4582;
	G4756<=G3816 and G4587;
	G4759<=G536 and G4500;
	G4761<=G4567 and G1674;
	G4782<=G1624 and G4623;
	G4785<=G2160 and G4625;
	G4787<=G2937 and G4628;
	G4789<=G3551 and G4632;
	G4791<=G3936 and G4636;
	G4792<=G1417 and G4471;
	G4793<=G4277 and G4639;
	G4794<=G4593 and G949;
	G4797<=G4593 and G4643;
	G4800<=G4648 and G4296;
	G4826<=G4209 and G4463;
	G4827<=G4520 and G4515;
	G4828<=G4510 and G4508;
	G4829<=G4526 and G4522;
	G4830<=G4529 and G4525;
	G4831<=G4528 and G4524;
	G4832<=G4517 and G4512;
	G4833<=G4521 and G4516;
	G4834<=G4534 and G4531;
	G4835<=G4533 and G4530;
	G4836<=G4527 and G4523;
	G4838<=G4648 and G84;
	G4863<=G4777 and G2874;
	G4865<=G4776 and G1849;
	G4867<=G4811 and G3872;
	G4868<=G4774 and G2891;
	G4870<=G4779 and G1884;
	G4872<=G4760 and G1549;
	G4873<=G4838 and G4173;
	G4874<=G582 and G4708;
	G4928<=G148 and G4723;
	G4932<=G157 and G4727;
	G4937<=G166 and G4732;
	G4942<=G175 and G4736;
	G4947<=G184 and G4741;
	G4949<=G193 and G4753;
	G5017<=G4784 and G1679;
	G5023<=G3935 and G4804;
	G5043<=G3941 and G4805;
	G5047<=G3954 and G4806;
	G5050<=G4285 and G4807;
	G5053<=G4599 and G4808;
	G5095<=G4794 and G951;
	G5096<=G4794 and G4647;
	G5098<=G4021 and G4837;
	G5122<=G193 and G4662;
	G5123<=G4670 and G1936;
	G5142<=G148 and G5099;
	G5143<=G157 and G5099;
	G5144<=G166 and G5099;
	G5145<=G175 and G5099;
	G5146<=G184 and G5099;
	G5149<=G4910 and G1480;
	G5152<=G430 and G4950;
	G5153<=G492 and G4904;
	G5154<=G500 and G4993;
	G5156<=G434 and G4877;
	G5157<=G496 and G4904;
	G5158<=G504 and G4993;
	G5159<=G536 and G4967;
	G5161<=G5095 and G4535;
	G5162<=G5088 and G2105;
	G5163<=G402 and G4950;
	G5164<=G437 and G4877;
	G5165<=G508 and G4993;
	G5166<=G541 and G4967;
	G5167<=G5011 and G1556;
	G5169<=G5093 and G1375;
	G5170<=G5091 and G2111;
	G5171<=G406 and G4950;
	G5172<=G441 and G4877;
	G5173<=G512 and G4993;
	G5175<=G5094 and G1384;
	G5176<=G410 and G4950;
	G5177<=G445 and G4877;
	G5178<=G516 and G4993;
	G5180<=G414 and G4950;
	G5181<=G449 and G4877;
	G5182<=G520 and G4993;
	G5183<=G418 and G4950;
	G5184<=G453 and G4877;
	G5185<=G524 and G4993;
	G5186<=G422 and G4950;
	G5187<=G457 and G4877;
	G5188<=G1043 and G4894;
	G5189<=G528 and G4993;
	G5190<=G426 and G4950;
	G5191<=G461 and G4877;
	G5192<=G1046 and G4894;
	G5193<=G532 and G4967;
	G5194<=G586 and G4874;
	G5197<=G465 and G4967;
	G5198<=G558 and G5025;
	G5200<=G559 and G5025;
	G5201<=G4859 and G5084;
	G5209<=G560 and G5025;
	G5211<=G4860 and G5086;
	G5212<=G561 and G5025;
	G5213<=G4862 and G5087;
	G5214<=G562 and G5025;
	G5215<=G4864 and G5090;
	G5216<=G563 and G5025;
	G5217<=G4866 and G5092;
	G5218<=G564 and G5025;
	G5225<=G669 and G5054;
	G5226<=G672 and G5054;
	G5229<=G545 and G4980;
	G5232<=G548 and G4980;
	G5233<=G551 and G4980;
	G5234<=G197 and G4915;
	G5235<=G554 and G4980;
	G5236<=G269 and G4915;
	G5240<=G293 and G4915;
	G5245<=G297 and G4915;
	G5269<=G557 and G5025;
	G5311<=G5013 and G4468;
	G5317<=G148 and G4869;
	G5349<=G5324 and G3451;
	G5350<=G5325 and G3453;
	G5351<=G5326 and G3459;
	G5353<=G5327 and G3463;
	G5354<=G5249 and G2903;
	G5356<=G5265 and G1902;
	G5357<=G398 and G5220;
	G5359<=G4428 and G5155;
	G5360<=G4431 and G5160;
	G5361<=G4435 and G5168;
	G5362<=G4437 and G5174;
	G5363<=G4439 and G5179;
	G5364<=G574 and G5194;
	G5369<=G143 and G5247;
	G5371<=G152 and G5248;
	G5373<=G161 and G5250;
	G5376<=G170 and G5255;
	G5378<=G179 and G5260;
	G5380<=G188 and G5264;
	G5398<=G366 and G5261;
	G5402<=G370 and G5266;
	G5406<=G374 and G5270;
	G5410<=G378 and G5274;
	G5414<=G382 and G5278;
	G5419<=G386 and G5292;
	G5424<=G390 and G5296;
	G5428<=G394 and G5300;
	G5429<=G398 and G5304;
	G5438<=G5224 and G3769;
	G5441<=G4537 and G5251 and G1558;
	G5443<=G4537 and G5251 and G2307;
	G5444<=G4545 and G5256 and G1574;
	G5446<=G4537 and G5241;
	G5447<=G4545 and G5256 and G2311;
	G5449<=G4545 and G5246;
	G5451<=G5251 and G4544;
	G5452<=G5315 and G4612;
	G5454<=G5256 and G4549;
	G5481<=G366 and G5331;
	G5482<=G370 and G5331;
	G5483<=G374 and G5331;
	G5484<=G378 and G5331;
	G5485<=G382 and G5331;
	G5486<=G386 and G5331;
	G5487<=G390 and G5331;
	G5488<=G394 and G5331;
	G5492<=G5441 and G3452;
	G5494<=G5443 and G3455;
	G5495<=G5444 and G3456;
	G5496<=G5446 and G3457;
	G5497<=G5447 and G3458;
	G5498<=G5449 and G3460;
	G5499<=G5451 and G3462;
	G5500<=G5430 and G5074;
	G5501<=G5454 and G3478;
	G5503<=G366 and G5384;
	G5515<=G590 and G5364;
	G5553<=G5012 and G5440;
	G5555<=G5014 and G5442;
	G5556<=G5015 and G5445;
	G5557<=G5016 and G5448;
	G5558<=G5018 and G5450;
	G5559<=G5024 and G5453;
	G5560<=G5044 and G5456;
	G5562<=G5228 and G5457;
	G5569<=G5348 and G3772;
	G5598<=G5046 and G5509;
	G5599<=G5049 and G5512;
	G5600<=G5502 and G4900;
	G5601<=G5052 and G5518;
	G5602<=G594 and G5515;
	G5603<=G5504 and G4911;
	G5604<=G5059 and G5521;
	G5616<=G5505 and G4929;
	G5617<=G5061 and G5524;
	G5618<=G5506 and G4933;
	G5619<=G5064 and G5527;
	G5620<=G5507 and G4938;
	G5621<=G5508 and G4943;
	G5632<=G4494 and G5538;
	G5633<=G4496 and G5539;
	G5635<=G4498 and G5542;
	G5637<=G4499 and G5543;
	G5646<=G4502 and G5544;
	G5648<=G4507 and G5545;
	G5660<=G4509 and G5549;
	G5663<=G4513 and G5550;
	G5665<=G361 and G5570;
	G5668<=G49 and G5571;
	G5671<=G54 and G5572;
	G5673<=G59 and G5573;
	G5675<=G64 and G5574;
	G5677<=G69 and G5575;
	G5679<=G74 and G5576;
	G5681<=G79 and G5577;
	G5682<=G84 and G5578;
	G5701<=G5683 and G3813;
	G5728<=G5623 and G3889;
	G5883<=G5824 and G3752;
	G5898<=G5800 and G5647;
	G5900<=G5804 and G5658;
	G5902<=G5808 and G5661;
	G5904<=G5812 and G5664;
	G5909<=G5787 and G3384;
	G5910<=G5816 and G5667;
	G5911<=G5817 and G5670;
	G5935<=G5112 and G5784;
	G5936<=G5113 and G5788;
	G5937<=G5775 and G5392;
	G5938<=G5114 and G5791;
	G5939<=G5776 and G5395;
	G5940<=G5115 and G5794;
	G5941<=G5777 and G5399;
	G5942<=G5117 and G5797;
	G5944<=G5778 and G5403;
	G5945<=G5118 and G5801;
	G5948<=G5779 and G5407;
	G5949<=G5119 and G5805;
	G5951<=G5780 and G5411;
	G5952<=G5120 and G5809;
	G5953<=G5781 and G5415;
	G5954<=G5121 and G5813;
	G5955<=G5782 and G5420;
	G5956<=G5783 and G5425;
	G6047<=G5824 and G1692;
	G6055<=G5824 and G1696;
	G6056<=G5824 and G1699;
	G6060<=G5824 and G1703;
	G6061<=G5824 and G1711;
	G6066<=G5824 and G1721;
	G6068<=G5824 and G1726;
	G6077<=G5824 and G1735;
	G6079<=G1236 and G5753;
	G6081<=G1177 and G5731;
	G6082<=G1123 and G5742;
	G6084<=G1123 and G5753;
	G6085<=G1161 and G5731;
	G6086<=G1143 and G5742;
	G6088<=G1143 and G5753;
	G6089<=G1143 and G5731;
	G6090<=G1161 and G5742;
	G6091<=G1161 and G5753;
	G6092<=G1123 and G5731;
	G6093<=G1177 and G5742;
	G6094<=G1177 and G5753;
	G6096<=G1193 and G5753;
	G6098<=G1209 and G5753;
	G6099<=G1222 and G5753;
	G6123<=G5702 and G5958;
	G6124<=G5705 and G5958;
	G6125<=G5708 and G5975;
	G6126<=G5711 and G5958;
	G6127<=G5714 and G5975;
	G6128<=G5590 and G5958;
	G6129<=G5717 and G5975;
	G6130<=G5720 and G5958;
	G6131<=G5593 and G5975;
	G6132<=G3752 and G5880;
	G6133<=G5723 and G5975;
	G6135<=G5584 and G5958;
	G6140<=G5587 and G5975;
	G6141<=G3173 and G5997;
	G6144<=G3183 and G5997;
	G6145<=G3187 and G6015;
	G6146<=G3192 and G5997;
	G6148<=G3196 and G6015;
	G6149<=G3200 and G5997;
	G6150<=G3204 and G6015;
	G6151<=G3209 and G5997;
	G6152<=G3212 and G6015;
	G6153<=G3216 and G5997;
	G6154<=G3219 and G6015;
	G6155<=G2588 and G5997;
	G6156<=G2591 and G6015;
	G6157<=G3158 and G5997;
	G6158<=G2594 and G6015;
	G6159<=G3177 and G6015;
	G6238<=G528 and G5886;
	G6240<=G4205 and G5888;
	G6241<=G1325 and G5887;
	G6243<=G500 and G5890;
	G6244<=G4759 and G5891;
	G6245<=G1329 and G5889;
	G6247<=G504 and G5893;
	G6248<=G465 and G5894;
	G6249<=G1332 and G5892;
	G6250<=G1692 and G6036;
	G6253<=G508 and G5896;
	G6254<=G532 and G5897;
	G6255<=G1335 and G5895;
	G6256<=G1696 and G6040;
	G6258<=G512 and G5899;
	G6259<=G1699 and G6044;
	G6260<=G1703 and G6048;
	G6262<=G516 and G5901;
	G6263<=G1711 and G6052;
	G6265<=G520 and G5903;
	G6266<=G1721 and G6057;
	G6269<=G524 and G5908;
	G6270<=G1726 and G6062;
	G6275<=G1735 and G6070;
	G6288<=G5615 and G6160;
	G6291<=G5210 and G6161;
	G6295<=G5379 and G6162;
	G6299<=G5530 and G6163;
	G6302<=G5740 and G6164;
	G6304<=G5915 and G6165;
	G6311<=G3837 and G6194;
	G6313<=G3841 and G6194;
	G6315<=G3849 and G6194;
	G6316<=G3855 and G6194;
	G6317<=G3862 and G6194;
	G6318<=G3865 and G6212;
	G6320<=G3869 and G6194;
	G6321<=G3873 and G6212;
	G6323<=G3877 and G6194;
	G6324<=G3880 and G6212;
	G6326<=G3833 and G6194;
	G6327<=G3884 and G6212;
	G6329<=G3888 and G6212;
	G6331<=G3891 and G6212;
	G6333<=G3896 and G6212;
	G6334<=G3858 and G6212;
	G6336<=G6246 and G6065;
	G6338<=G6251 and G6067;
	G6340<=G6257 and G6069;
	G6341<=G6261 and G6074;
	G6342<=G6264 and G6076;
	G6343<=G6268 and G6078;
	G6344<=G6272 and G6080;
	G6345<=G6273 and G6083;
	G6346<=G6274 and G6087;
	G6348<=G5869 and G6211;
	G6354<=G5866 and G6193;
	G6468<=G2032 and G6394 and G1609;
	G6469<=G2121 and G2032 and G6394;
	G6473<=G2036 and G6397 and G1628;
	G6474<=G2138 and G2036 and G6397;
	G6555<=G1838 and G6469;
	G6557<=G1595 and G6469;
	G6558<=G1842 and G6474;
	G6559<=G1612 and G6474;
	G6603<=G6581 and G6236;
	G6613<=G932 and G6554;
	G6614<=G932 and G6556;
	G6619<=G6515 and G6115;
	G6620<=G6516 and G6117;
	G6625<=G2121 and G1595 and G6538;
	G6628<=G2138 and G1612 and G6540;
	G6631<=G1838 and G6545;
	G6634<=G1595 and G6545;
	G6637<=G1842 and G6549;
	G6640<=G1612 and G6549;
	G6643<=G6574 and G6229;
	G6644<=G6575 and G6230;
	G6645<=G6576 and G6231;
	G6646<=G6577 and G6232;
	G6647<=G6578 and G6233;
	G6648<=G6579 and G6234;
	G6650<=G6580 and G6235;
	G6692<=G6616 and G6615;
	G6693<=G6618 and G6617;
	G6716<=G6682 and G932;
	G6718<=G4511 and G6661;
	G6719<=G4518 and G6665;
	G6731<=G6717 and G4427;
	G6736<=G6712 and G754 and G5237;
	G6737<=G6714 and G760 and G5237;
	G6738<=G6713 and G809 and G5242;
	G6739<=G6715 and G815 and G5242;
	G6748<=G6733 and G6732;
	G6749<=G6735 and G6734;
	G6766<=G6750 and G2986;
	G6767<=G6754 and G2986;
	G6768<=G6750 and G3477;
	G6769<=G6758 and G2986;
	G6770<=G6754 and G3482;
	G6771<=G6758 and G3483;
	G6772<=G6746 and G3312;
	G6773<=G6762 and G2986;
	G6777<=G6762 and G3488;
	G6798<=G4946 and G6781;
	G6799<=G4948 and G6782;
	G6816<=G6784 and G3346;
	G6828<=G6803 and G5958;
	G6829<=G6806 and G5958;
	G6830<=G6809 and G5975;
	G6831<=G6812 and G5975;
	G6848<=G3741 and G328 and G6843;
	G6851<=G6846 and G2293;
	G6852<=G6847 and G2295;
	G6874<=G6873 and G2060;
	G6908<=G6907 and G3886;
	G6909<=G6896 and G6894;
	G6910<=G6892 and G6891;
	G6911<=G6904 and G6902;
	G6912<=G6899 and G6897;
	G6913<=G6900 and G6898;
	G6914<=G6895 and G6893;
	G6915<=G6906 and G6905;
	G6916<=G6903 and G6901;
	G6923<=G6918 and G6917;
	G6924<=G6920 and G6919;
	G6934<=G6932 and G3605;
	G6935<=G6933 and G3622;
	I2566<=G749 and G743 and G736;
	I2574<=G804 and G798 and G791;
	I4040<=G1279 and G2025 and G1267;
	I5351<=G3511 and G3517 and G3520 and G3525;
	I5352<=G3529 and G3531 and G3535 and G3538;
	I5359<=G3518 and G3521 and G3526 and G3530;
	I5360<=G3532 and G3536 and G3539 and G3544;
	G901<= not (G314 and G310);
	G905<= not (G301 and G319);
	G926<= not (I1952 and I1953);
	G928<= not (I1962 and I1963);
	G930<= not (I1970 and I1971);
	G937<= not (I1979 and I1980);
	G939<= not (I1987 and I1988);
	G941<= not (I1995 and I1996);
	G944<= not (I2004 and I2005);
	G948<= not (I2014 and I2015);
	G950<= not (I2022 and I2023);
	G1036<= not (I2061 and I2062);
	G1042<= not (I2073 and I2074);
	G1044<= not (I2081 and I2082);
	G1047<= not (I2090 and I2091);
	G1075<= not (I2109 and I2110);
	G1138<= not (G102 and G98);
	G1157<= not (G89 and G107);
	G1253<= not (I2245 and I2246);
	G1316<= not (I2300 and I2301);
	G1359<= not (G866 and G306);
	G1387<= not (G862 and G314 and G301);
	G1398<= not (G306 and G889);
	G1402<= not (G310 and G866 and G873);
	G1411<= not (G314 and G873);
	G1417<= not (G873 and G889);
	G1534<= not (I2498 and I2499);
	G1540<= not (I2507 and I2508);
	G1558<= not (I2527 and I2528);
	G1573<= not (G729 and G719 and G766);
	G1574<= not (I2543 and I2544);
	G1582<= not (G784 and G774 and G821);
	G1686<= not (I2675 and I2676);
	G1687<= not (I2682 and I2683);
	G1743<= not (G1064 and G94);
	G1749<= not (I2767 and I2768);
	G1764<= not (I2796 and I2797);
	G1777<= not (G1060 and G102 and G89);
	G1793<= not (G94 and G1084);
	G1797<= not (G98 and G1064 and G1070);
	G1815<= not (G102 and G1070);
	G1822<= not (G1070 and G1084);
	G1829<= not (I2898 and I2899);
	G1845<= not (I2934 and I2935);
	G2008<= not (G866 and G873 and G1784);
	G2009<= not (G901 and G1387 and G905);
	G2010<= not (G1473 and G1470 and G1459);
	G2024<= not (I3126 and I3127);
	G2061<= not (I3169 and I3170);
	G2067<= not (I3178 and I3179);
	G2080<= not (I3189 and I3190);
	G2095<= not (G1584 and G749 and G736);
	G2100<= not (G1588 and G804 and G791);
	G2263<= not (I3399 and I3400);
	G2266<= not (I3412 and I3413);
	G2307<= not (I3446 and I3447);
	G2311<= not (I3456 and I3457);
	G2434<= not (G1064 and G1070 and G1620);
	G2435<= not (G1138 and G1777 and G1157);
	G2582<= not (I3698 and I3699);
	G2607<= not (I3740 and I3741);
	G2698<= not (I3847 and I3848);
	G2719<= not (I3875 and I3876);
	G2731<= not (I3894 and I3895);
	G2745<= not (I3915 and I3916);
	G2757<= not (I3934 and I3935);
	G2769<= not (I3953 and I3954);
	G2780<= not (I3971 and I3972);
	G2791<= not (I3989 and I3990);
	G2795<= not (G1997 and G866);
	G2804<= not (I4009 and I4010);
	G2831<= not (G2007 and G862 and G1784);
	G2858<= not (G1815 and G2577);
	G2940<= not (G197 and G2381);
	G2944<= not (G269 and G2381);
	G2947<= not (G1411 and G2026);
	G2951<= not (G2142 and G1797);
	G2960<= not (I4151 and I4152);
	G2966<= not (I4160 and I4161);
	G2995<= not (I4183 and I4184);
	G3012<= not (I4204 and I4205);
	G3013<= not (I4211 and I4212);
	G3028<= not (I4234 and I4235);
	G3109<= not (G2360 and G1064);
	G3140<= not (G2409 and G1060 and G1620);
	G3207<= not (I4445 and I4446);
	G3215<= not (G2340 and G1402);
	G3246<= not (I4527 and I4528);
	G3276<= not (I4546 and I4547);
	G3330<= not (G1815 and G1797 and G3109);
	G3502<= not (G1411 and G1402 and G2795);
	G3511<= not (G3158 and G3002 and G2976 and G2968);
	G3517<= not (G3173 and G3002 and G2976 and G2179);
	G3518<= not (G3177 and G3023 and G3007 and G2981);
	G3520<= not (G3183 and G3002 and G2197 and G2968);
	G3521<= not (G3187 and G3023 and G3007 and G2179);
	G3525<= not (G3192 and G3002 and G2197 and G2179);
	G3526<= not (G3196 and G3023 and G2197 and G2981);
	G3529<= not (G3200 and G2215 and G2976 and G2968);
	G3530<= not (G3204 and G3023 and G2197 and G2179);
	G3531<= not (G3209 and G2215 and G2976 and G2179);
	G3532<= not (G3212 and G2215 and G3007 and G2981);
	G3535<= not (G3216 and G2215 and G2197 and G2968);
	G3536<= not (G3219 and G2215 and G3007 and G2179);
	G3538<= not (G2588 and G2215 and G2197 and G2179);
	G3539<= not (G2591 and G2215 and G2197 and G2981);
	G3544<= not (G2594 and G2215 and G2197 and G2179);
	G3597<= not (I4783 and I4784);
	G3741<= not (G901 and G3433 and G2340);
	G3742<= not (I4920 and I4921);
	G3756<= not (I4940 and I4941);
	G3893<= not (G3664 and G3656 and G3647);
	G3955<= not (I5188 and I5189);
	G3957<= not (I5196 and I5197);
	G3961<= not (I5208 and I5209);
	G3968<= not (I5227 and I5228);
	G3974<= not (I5243 and I5244);
	G3979<= not (I5258 and I5259);
	G3983<= not (I5270 and I5271);
	G3985<= not (G1138 and G3718 and G2142);
	G4002<= not (I5293 and I5294);
	G4004<= not (I5301 and I5302);
	G4007<= not (I5308 and I5309);
	G4017<= not (G107 and G3425);
	G4049<= not (G3677 and G3425);
	G4151<= not (I5536 and I5537);
	G4221<= not (I5648 and I5649);
	G4223<= not (I5658 and I5659);
	G4237<= not (G4049 and G4017);
	G4300<= not (I5760 and I5761);
	G4301<= not (I5767 and I5768);
	G4319<= not (I5783 and I5784);
	G4465<= not (G319 and G4253);
	G4472<= not (G3380 and G4253);
	G4504<= not (I6027 and I6028);
	G4608<= not (I6176 and I6177);
	G4610<= not (I6186 and I6187);
	G4613<= not (I6195 and I6196);
	G4640<= not (G4402 and G1056);
	G4669<= not (G4550 and G1017 and G1680 and G2897);
	G4670<= not (G4611 and G3528);
	G4674<= not (G4550 and G1514 and G2107 and G2897);
	G4678<= not (G2897 and G2101 and G1514 and G4550);
	G4680<= not (G4550 and G1514 and G1006 and G2897);
	G4762<= not (I6391 and I6392);
	G4803<= not (I6474 and I6475);
	G4812<= not (G4550 and G1560 and G1559 and G2073);
	G4813<= not (G4550 and G965 and G1560 and G2073);
	G4814<= not (G4550 and G1575 and G1550 and G2073);
	G4816<= not (G996 and G4550 and G1518 and G2073);
	G4819<= not (I6500 and I6501);
	G4825<= not (G4472 and G4465);
	G4903<= not (G4717 and G858);
	G5019<= not (I6660 and I6661);
	G5111<= not (I6744 and I6745);
	G5308<= not (I6963 and I6964);
	G5318<= not (G676 and G5060);
	G5431<= not (I7098 and I7099);
	G5455<= not (G2330 and G5311);
	G5502<= not (I7209 and I7210);
	G5504<= not (I7217 and I7218);
	G5505<= not (I7224 and I7225);
	G5506<= not (I7231 and I7232);
	G5507<= not (I7238 and I7239);
	G5508<= not (I7245 and I7246);
	G5565<= not (I7312 and I7313);
	G5634<= not (G5563 and G4767);
	G5636<= not (G5564 and G4769);
	G5683<= not (I7433 and I7434);
	G5684<= not (I7440 and I7441);
	G5686<= not (G5546 and G1017 and G1551 and G2916);
	G5688<= not (G5546 and G1585 and G2084 and G2916);
	G5775<= not (I7521 and I7522);
	G5776<= not (I7528 and I7529);
	G5777<= not (I7535 and I7536);
	G5778<= not (I7542 and I7543);
	G5779<= not (I7549 and I7550);
	G5780<= not (I7556 and I7557);
	G5781<= not (I7563 and I7564);
	G5782<= not (I7570 and I7571);
	G5783<= not (I7577 and I7578);
	G5818<= not (G5638 and G2056 and G1666 and G1661);
	G5821<= not (G5638 and G2056 and G1076 and G1666);
	G5852<= not (G5638 and G2053 and G1661);
	G5853<= not (G5638 and G2053 and G1076);
	G5854<= not (G5638 and G1683 and G1552 and G2062);
	G5857<= not (G5638 and G1552 and G1017 and G2062);
	G5862<= not (G5649 and G1529 and G1535 and G2068);
	G5863<= not (G5649 and G1076 and G1535 and G2068);
	G5864<= not (G5649 and G1529 and G1088 and G2068);
	G5865<= not (G5649 and G1088 and G1076 and G2068);
	G5866<= not (G5649 and G1529 and G2081);
	G5869<= not (G5649 and G1076 and G2081);
	G5872<= not (G5649 and G1557 and G1564 and G2113);
	G5873<= not (G5649 and G1017 and G1564 and G2113);
	G5926<= not (G5741 and G639);
	G5943<= not (G5818 and G2940);
	G5947<= not (G5821 and G2944);
	G6095<= not (G2952 and G5854);
	G6097<= not (G2954 and G5857);
	G6394<= not (I8195 and I8196);
	G6397<= not (I8202 and I8203);
	G6717<= not (G6669 and G5065 and G5062);
	G6740<= not (G6703 and G6457 and G4936);
	G6741<= not (G6705 and G6461 and G4941);
	G6742<= not (G6683 and G932 and G6716);
	G6774<= not (G6754 and G6750);
	G6778<= not (G6762 and G6758);
	G6783<= not (G6747 and G5068 and G5066);
	G6843<= not (I9051 and I9052);
	G6873<= not (G6848 and G3621);
	G6928<= not (G4532 and G6926);
	G6929<= not (G4536 and G6927);
	I1951<= not (G524 and G248);
	I1952<= not (G524 and I1951);
	I1953<= not (G248 and I1951);
	I1961<= not (G520 and G242);
	I1962<= not (G520 and I1961);
	I1963<= not (G242 and I1961);
	I1969<= not (G516 and G236);
	I1970<= not (G516 and I1969);
	I1971<= not (G236 and I1969);
	I1978<= not (G512 and G230);
	I1979<= not (G512 and I1978);
	I1980<= not (G230 and I1978);
	I1986<= not (G508 and G224);
	I1987<= not (G508 and I1986);
	I1988<= not (G224 and I1986);
	I1994<= not (G504 and G218);
	I1995<= not (G504 and I1994);
	I1996<= not (G218 and I1994);
	I2003<= not (G500 and G212);
	I2004<= not (G500 and I2003);
	I2005<= not (G212 and I2003);
	I2013<= not (G532 and G260);
	I2014<= not (G532 and I2013);
	I2015<= not (G260 and I2013);
	I2021<= not (G528 and G254);
	I2022<= not (G528 and I2021);
	I2023<= not (G254 and I2021);
	I2060<= not (G7 and G3);
	I2061<= not (G7 and I2060);
	I2062<= not (G3 and I2060);
	I2072<= not (G15 and G11);
	I2073<= not (G15 and I2072);
	I2074<= not (G11 and I2072);
	I2080<= not (G25 and G19);
	I2081<= not (G25 and I2080);
	I2082<= not (G19 and I2080);
	I2089<= not (G33 and G29);
	I2090<= not (G33 and I2089);
	I2091<= not (G29 and I2089);
	I2108<= not (G602 and G610);
	I2109<= not (G602 and I2108);
	I2110<= not (G610 and I2108);
	I2244<= not (G567 and G598);
	I2245<= not (G567 and I2244);
	I2246<= not (G598 and I2244);
	I2299<= not (G830 and G341);
	I2300<= not (G830 and I2299);
	I2301<= not (G341 and I2299);
	I2497<= not (G1042 and G1036);
	I2498<= not (G1042 and I2497);
	I2499<= not (G1036 and I2497);
	I2506<= not (G1047 and G1044);
	I2507<= not (G1047 and I2506);
	I2508<= not (G1044 and I2506);
	I2526<= not (G766 and G719);
	I2527<= not (G766 and I2526);
	I2528<= not (G719 and I2526);
	I2542<= not (G821 and G774);
	I2543<= not (G821 and I2542);
	I2544<= not (G774 and I2542);
	I2674<= not (G710 and G131);
	I2675<= not (G710 and I2674);
	I2676<= not (G131 and I2674);
	I2681<= not (G918 and G613);
	I2682<= not (G918 and I2681);
	I2683<= not (G613 and I2681);
	I2766<= not (G749 and G743);
	I2767<= not (G749 and I2766);
	I2768<= not (G743 and I2766);
	I2795<= not (G804 and G798);
	I2796<= not (G804 and I2795);
	I2797<= not (G798 and I2795);
	I2897<= not (G1027 and G634);
	I2898<= not (G1027 and I2897);
	I2899<= not (G634 and I2897);
	I2933<= not (G1436 and G345);
	I2934<= not (G1436 and I2933);
	I2935<= not (G345 and I2933);
	I3125<= not (G1279 and G1276);
	I3126<= not (G1279 and I3125);
	I3127<= not (G1276 and I3125);
	I3168<= not (G1540 and G1534);
	I3169<= not (G1540 and I3168);
	I3170<= not (G1534 and I3168);
	I3177<= not (G1706 and G736);
	I3178<= not (G1706 and I3177);
	I3179<= not (G736 and I3177);
	I3188<= not (G1716 and G791);
	I3189<= not (G1716 and I3188);
	I3190<= not (G791 and I3188);
	I3398<= not (G1826 and G135);
	I3399<= not (G1826 and I3398);
	I3400<= not (G135 and I3398);
	I3411<= not (G1419 and G616);
	I3412<= not (G1419 and I3411);
	I3413<= not (G616 and I3411);
	I3445<= not (G1689 and G729);
	I3446<= not (G1689 and I3445);
	I3447<= not (G729 and I3445);
	I3455<= not (G1691 and G784);
	I3456<= not (G1691 and I3455);
	I3457<= not (G784 and I3455);
	I3697<= not (G1570 and G642);
	I3698<= not (G1570 and I3697);
	I3699<= not (G642 and I3697);
	I3739<= not (G2021 and G349);
	I3740<= not (G2021 and I3739);
	I3741<= not (G349 and I3739);
	I3846<= not (G284 and G2370);
	I3847<= not (G284 and I3846);
	I3848<= not (G2370 and I3846);
	I3874<= not (G285 and G2397);
	I3875<= not (G285 and I3874);
	I3876<= not (G2397 and I3874);
	I3893<= not (G286 and G2422);
	I3894<= not (G286 and I3893);
	I3895<= not (G2422 and I3893);
	I3914<= not (G287 and G2449);
	I3915<= not (G287 and I3914);
	I3916<= not (G2449 and I3914);
	I3933<= not (G288 and G2473);
	I3934<= not (G288 and I3933);
	I3935<= not (G2473 and I3933);
	I3952<= not (G289 and G2497);
	I3953<= not (G289 and I3952);
	I3954<= not (G2497 and I3952);
	I3970<= not (G290 and G2518);
	I3971<= not (G290 and I3970);
	I3972<= not (G2518 and I3970);
	I3988<= not (G291 and G2544);
	I3989<= not (G291 and I3988);
	I3990<= not (G2544 and I3988);
	I4008<= not (G292 and G2568);
	I4009<= not (G292 and I4008);
	I4010<= not (G2568 and I4008);
	I4150<= not (G2551 and G139);
	I4151<= not (G2551 and I4150);
	I4152<= not (G139 and I4150);
	I4159<= not (G2015 and G619);
	I4160<= not (G2015 and I4159);
	I4161<= not (G619 and I4159);
	I4182<= not (G2292 and G749);
	I4183<= not (G2292 and I4182);
	I4184<= not (G749 and I4182);
	I4203<= not (G2255 and G743);
	I4204<= not (G2255 and I4203);
	I4205<= not (G743 and I4203);
	I4210<= not (G2294 and G804);
	I4211<= not (G2294 and I4210);
	I4212<= not (G804 and I4210);
	I4233<= not (G2267 and G798);
	I4234<= not (G2267 and I4233);
	I4235<= not (G798 and I4233);
	I4444<= not (G2092 and G606);
	I4445<= not (G2092 and I4444);
	I4446<= not (G606 and I4444);
	I4526<= not (G2909 and G646);
	I4527<= not (G2909 and I4526);
	I4528<= not (G646 and I4526);
	I4545<= not (G2853 and G353);
	I4546<= not (G2853 and I4545);
	I4547<= not (G353 and I4545);
	I4782<= not (G2846 and G622);
	I4783<= not (G2846 and I4782);
	I4784<= not (G622 and I4782);
	I4919<= not (G3522 and G650);
	I4920<= not (G3522 and I4919);
	I4921<= not (G650 and I4919);
	I4939<= not (G3437 and G357);
	I4940<= not (G3437 and I4939);
	I4941<= not (G357 and I4939);
	I5187<= not (G3589 and G3593);
	I5188<= not (G3589 and I5187);
	I5189<= not (G3593 and I5187);
	I5195<= not (G3567 and G3571);
	I5196<= not (G3567 and I5195);
	I5197<= not (G3571 and I5195);
	I5207<= not (G3267 and G3271);
	I5208<= not (G3267 and I5207);
	I5209<= not (G3271 and I5207);
	I5226<= not (G3259 and G3263);
	I5227<= not (G3259 and I5226);
	I5228<= not (G3263 and I5226);
	I5242<= not (G3242 and G3247);
	I5243<= not (G3242 and I5242);
	I5244<= not (G3247 and I5242);
	I5257<= not (G3714 and G3719);
	I5258<= not (G3714 and I5257);
	I5259<= not (G3719 and I5257);
	I5269<= not (G3705 and G3710);
	I5270<= not (G3705 and I5269);
	I5271<= not (G3710 and I5269);
	I5292<= not (G3421 and G625);
	I5293<= not (G3421 and I5292);
	I5294<= not (G625 and I5292);
	I5300<= not (G471 and G3505);
	I5301<= not (G471 and I5300);
	I5302<= not (G3505 and I5300);
	I5307<= not (G478 and G3512);
	I5308<= not (G478 and I5307);
	I5309<= not (G3512 and I5307);
	I5535<= not (G3907 and G654);
	I5536<= not (G3907 and I5535);
	I5537<= not (G654 and I5535);
	I5647<= not (G3974 and G3968);
	I5648<= not (G3974 and I5647);
	I5649<= not (G3968 and I5647);
	I5657<= not (G3983 and G3979);
	I5658<= not (G3983 and I5657);
	I5659<= not (G3979 and I5657);
	I5759<= not (G3836 and G3503);
	I5760<= not (G3836 and I5759);
	I5761<= not (G3503 and I5759);
	I5766<= not (G3961 and G3957);
	I5767<= not (G3961 and I5766);
	I5768<= not (G3957 and I5766);
	I5782<= not (G3810 and G628);
	I5783<= not (G3810 and I5782);
	I5784<= not (G628 and I5782);
	I6026<= not (G4223 and G4221);
	I6027<= not (G4223 and I6026);
	I6028<= not (G4221 and I6026);
	I6175<= not (G4236 and G571);
	I6176<= not (G4236 and I6175);
	I6177<= not (G571 and I6175);
	I6185<= not (G4301 and G3955);
	I6186<= not (G4301 and I6185);
	I6187<= not (G3955 and I6185);
	I6194<= not (G4199 and G631);
	I6195<= not (G4199 and I6194);
	I6196<= not (G631 and I6194);
	I6390<= not (G4504 and G4610);
	I6391<= not (G4504 and I6390);
	I6392<= not (G4610 and I6390);
	I6473<= not (G4541 and G578);
	I6474<= not (G4541 and I6473);
	I6475<= not (G578 and I6473);
	I6499<= not (G4504 and G3541);
	I6500<= not (G4504 and I6499);
	I6501<= not (G3541 and I6499);
	I6659<= not (G4762 and G3541);
	I6660<= not (G4762 and I6659);
	I6661<= not (G3541 and I6659);
	I6743<= not (G4708 and G582);
	I6744<= not (G4708 and I6743);
	I6745<= not (G582 and I6743);
	I6962<= not (G4874 and G586);
	I6963<= not (G4874 and I6962);
	I6964<= not (G586 and I6962);
	I7097<= not (G5194 and G574);
	I7098<= not (G5194 and I7097);
	I7099<= not (G574 and I7097);
	I7208<= not (G143 and G5367);
	I7209<= not (G143 and I7208);
	I7210<= not (G5367 and I7208);
	I7216<= not (G152 and G5368);
	I7217<= not (G152 and I7216);
	I7218<= not (G5368 and I7216);
	I7223<= not (G161 and G5370);
	I7224<= not (G161 and I7223);
	I7225<= not (G5370 and I7223);
	I7230<= not (G170 and G5372);
	I7231<= not (G170 and I7230);
	I7232<= not (G5372 and I7230);
	I7237<= not (G179 and G5374);
	I7238<= not (G179 and I7237);
	I7239<= not (G5374 and I7237);
	I7244<= not (G188 and G5377);
	I7245<= not (G188 and I7244);
	I7246<= not (G5377 and I7244);
	I7311<= not (G5364 and G590);
	I7312<= not (G5364 and I7311);
	I7313<= not (G590 and I7311);
	I7432<= not (G111 and G5554);
	I7433<= not (G111 and I7432);
	I7434<= not (G5554 and I7432);
	I7439<= not (G5515 and G594);
	I7440<= not (G5515 and I7439);
	I7441<= not (G594 and I7439);
	I7520<= not (G361 and G5659);
	I7521<= not (G361 and I7520);
	I7522<= not (G5659 and I7520);
	I7527<= not (G49 and G5662);
	I7528<= not (G49 and I7527);
	I7529<= not (G5662 and I7527);
	I7534<= not (G54 and G5666);
	I7535<= not (G54 and I7534);
	I7536<= not (G5666 and I7534);
	I7541<= not (G59 and G5669);
	I7542<= not (G59 and I7541);
	I7543<= not (G5669 and I7541);
	I7548<= not (G64 and G5672);
	I7549<= not (G64 and I7548);
	I7550<= not (G5672 and I7548);
	I7555<= not (G69 and G5674);
	I7556<= not (G69 and I7555);
	I7557<= not (G5674 and I7555);
	I7562<= not (G74 and G5676);
	I7563<= not (G74 and I7562);
	I7564<= not (G5676 and I7562);
	I7569<= not (G79 and G5678);
	I7570<= not (G79 and I7569);
	I7571<= not (G5678 and I7569);
	I7576<= not (G84 and G5680);
	I7577<= not (G84 and I7576);
	I7578<= not (G5680 and I7576);
	I8194<= not (G471 and G6188);
	I8195<= not (G471 and I8194);
	I8196<= not (G6188 and I8194);
	I8201<= not (G478 and G6192);
	I8202<= not (G478 and I8201);
	I8203<= not (G6192 and I8201);
	I9050<= not (G6832 and G3598);
	I9051<= not (G6832 and I9050);
	I9052<= not (G3598 and I9050);
	G1589<=G1059 or G1045;
	G2896<=G2323 or G1763;
	G2924<=G2095 or G1573;
	G2928<=G2100 or G1582;
	G3503<=G3122 or G3132;
	G3533<=G3154 or G3166;
	G3598<=G2808 or G2821;
	G3599<=G2935 or G1637;
	G3732<=G3324 or G2732;
	G3733<=G3325 or G2733;
	G3739<=G3334 or G2746;
	G3740<=G3335 or G2747;
	G3743<=G3344 or G2758;
	G3744<=G3345 or G2759;
	G3745<=G3356 or G2770;
	G3746<=G3357 or G2771;
	G3747<=G3365 or G2781;
	G3748<=G3366 or G2782;
	G3749<=G3371 or G2793;
	G3750<=G3372 or G2794;
	G3751<=G3375 or G2807;
	G3815<=G3282 or G2659;
	G3820<=G3287 or G2671;
	G3821<=G2951 or G3466;
	G3828<=G3304 or G1351;
	G3829<=G3294 or G3305;
	G3833<=G3602 or G3608;
	G3837<=G3609 or G3613;
	G3841<=G3614 or G3617;
	G3842<=G3670 or G3135;
	G3849<=G3618 or G3625;
	G3850<=G3680 or G3145;
	G3851<=G3681 or G3146;
	G3855<=G3626 or G3631;
	G3856<=G3686 or G3157;
	G3857<=G3687 or G3161;
	G3858<=G3629 or G3636;
	G3862<=G3632 or G3641;
	G3863<=G3692 or G3172;
	G3864<=G3693 or G3176;
	G3865<=G3637 or G3648;
	G3869<=G3642 or G3650;
	G3870<=G3700 or G3182;
	G3871<=G3701 or G3186;
	G3873<=G3649 or G3657;
	G3877<=G3651 or G3659;
	G3878<=G3703 or G3191;
	G3879<=G3704 or G3195;
	G3880<=G3658 or G3665;
	G3883<=G3709 or G3203;
	G3884<=G3666 or G3671;
	G3888<=G3672 or G3682;
	G3891<=G3683 or G3688;
	G3896<=G3689 or G3697;
	G3913<=G3449 or G2860;
	G3935<=G3464 or G2868;
	G3941<=G3479 or G2873;
	G3942<=G3215 or G3575;
	G3954<=G3484 or G3489;
	G3964<=G3634 or G3089;
	G3971<=G3644 or G3099;
	G3972<=G3646 or G3103;
	G3977<=G3653 or G3113;
	G3978<=G3655 or G3117;
	G3981<=G3661 or G3123;
	G3982<=G3663 or G3127;
	G3986<=G3667 or G3133;
	G3987<=G3669 or G3134;
	G3988<=G3678 or G3143;
	G3989<=G3679 or G3144;
	G3990<=G3684 or G3155;
	G3991<=G3685 or G3156;
	G3992<=G1555 or G3559;
	G3995<=G3690 or G3170;
	G3996<=G3691 or G3171;
	G3998<=G3698 or G3180;
	G3999<=G3699 or G3181;
	G4001<=G3702 or G3190;
	G4021<=G3558 or G2949;
	G4059<=G3466 or G3425;
	G4068<=G3293 or G2685;
	G4074<=G3301 or G2699;
	G4080<=G3302 or G2700;
	G4086<=G3310 or G2720;
	G4092<=G3311 or G2721;
	G4205<=G3843 or G541;
	G4231<=G3997 or G4000;
	G4233<=G3912 or G471;
	G4234<=G3921 or G478;
	G4243<=G4053 or G4058;
	G4285<=G3490 or G3887;
	G4427<=G4373 or G3668;
	G4430<=G4349 or G4015;
	G4433<=G4354 or G4032;
	G4434<=G4355 or G4033;
	G4436<=G4359 or G4035;
	G4438<=G4363 or G4037;
	G4440<=G4371 or G4038;
	G4441<=G4372 or G4039;
	G4443<=G4377 or G4041;
	G4444<=G4378 or G4042;
	G4446<=G4383 or G4043;
	G4447<=G4384 or G4044;
	G4450<=G4389 or G4047;
	G4451<=G4390 or G4048;
	G4454<=G4395 or G4051;
	G4455<=G4396 or G4052;
	G4458<=G4401 or G4057;
	G4468<=G4214 or G3831;
	G4473<=G3575 or G4253;
	G4497<=G4166 or G3784;
	G4500<=G4243 or G2010;
	G4544<=G4410 or G2995;
	G4549<=G4416 or G3013;
	G4599<=G3499 or G4230;
	G4607<=G4232 or G3899;
	G4627<=G4333 or G3603;
	G4630<=G4339 or G3610;
	G4631<=G4340 or G3611;
	G4634<=G4341 or G3615;
	G4635<=G4342 or G3616;
	G4637<=G4344 or G3619;
	G4638<=G4345 or G3620;
	G4641<=G4347 or G3627;
	G4642<=G4348 or G3628;
	G4645<=G4352 or G3633;
	G4646<=G4353 or G3635;
	G4651<=G4357 or G3643;
	G4652<=G4358 or G3645;
	G4653<=G4361 or G3652;
	G4654<=G4362 or G3654;
	G4655<=G4368 or G3660;
	G4656<=G4369 or G3662;
	G4740<=G4448 or G4154;
	G4745<=G4468 or G4569;
	G4752<=G4452 or G4155;
	G4757<=G4456 or G4158;
	G4773<=G4495 or G4220;
	G4811<=G4429 or G4432;
	G4859<=G4730 or G4486;
	G4860<=G4735 or G4488;
	G4862<=G4739 or G4489;
	G4864<=G4744 or G4490;
	G4866<=G4756 or G4491;
	G4936<=G4827 or G4828;
	G4941<=G4829 or G4832;
	G4946<=G4830 or G4833;
	G4948<=G4834 or G4836;
	G5012<=G4782 or G4580;
	G5013<=G4826 or G4621;
	G5014<=G4785 or G4583;
	G5015<=G4787 or G4588;
	G5016<=G4789 or G4592;
	G5018<=G4791 or G4597;
	G5024<=G4793 or G4600;
	G5044<=G4797 or G4602;
	G5060<=G3491 or G4819;
	G5062<=G4661 or G4666;
	G5065<=G4667 or G4671;
	G5066<=G4668 or G4672;
	G5068<=G4673 or G4677;
	G5069<=G1595 or G4688;
	G5074<=G4792 or G4598;
	G5077<=G1612 or G4694;
	G5083<=G4688 or G4271;
	G5085<=G4694 or G4280;
	G5202<=G4904 or G4914 or G4894;
	G5224<=G5123 or G3630;
	G5228<=G5096 or G4800;
	G5231<=G5048 or G672;
	G5241<=G5069 or G2067;
	G5246<=G5077 or G2080;
	G5277<=G5023 or G4763;
	G5281<=G5074 or G5124;
	G5291<=G5043 or G4764;
	G5295<=G5047 or G4766;
	G5303<=G5053 or G4768;
	G5323<=G5098 or G4802;
	G5326<=G5069 or G4410 or G3012;
	G5327<=G5077 or G4416 or G3028;
	G5348<=G5317 or G5122;
	G5367<=G5199 or G4928;
	G5368<=G5201 or G4932;
	G5370<=G5211 or G4937;
	G5372<=G5213 or G4942;
	G5374<=G5215 or G4947;
	G5377<=G5217 or G4949;
	G5385<=G3992 or G5318;
	G5386<=G5227 or G669;
	G5388<=G5318 or G1589 or G3491;
	G5430<=G5161 or G4873;
	G5458<=G3466 or G5311;
	G5467<=G3868 or G5318 or G3992;
	G5470<=G5359 or G5142;
	G5471<=G5360 or G5143;
	G5472<=G5361 or G5144;
	G5473<=G5362 or G5145;
	G5474<=G5363 or G5146;
	G5531<=G5349 or G3275;
	G5532<=G5350 or G3278;
	G5533<=G5351 or G3290;
	G5535<=G5353 or G3300;
	G5583<=G5569 or G4020;
	G5605<=G3575 or G5500;
	G5622<=G5492 or G3277;
	G5623<=G5503 or G5357;
	G5624<=G5494 or G3280;
	G5625<=G5495 or G3281;
	G5626<=G5496 or G3285;
	G5627<=G5497 or G3286;
	G5628<=G5498 or G3292;
	G5629<=G5499 or G3298;
	G5630<=G5501 or G3309;
	G5659<=G5551 or G5398;
	G5662<=G5553 or G5402;
	G5666<=G5555 or G5406;
	G5669<=G5556 or G5410;
	G5672<=G5557 or G5414;
	G5674<=G5558 or G5419;
	G5676<=G5559 or G5424;
	G5678<=G5560 or G5428;
	G5680<=G5562 or G5429;
	G5693<=G5632 or G5481;
	G5694<=G5633 or G5482;
	G5695<=G5635 or G5483;
	G5696<=G5637 or G5484;
	G5697<=G5646 or G5485;
	G5698<=G5648 or G5486;
	G5699<=G5660 or G5487;
	G5700<=G5663 or G5488;
	G5800<=G5369 or G5600;
	G5804<=G5371 or G5603;
	G5808<=G5373 or G5616;
	G5812<=G5376 or G5618;
	G5816<=G5378 or G5620;
	G5817<=G5380 or G5621;
	G5916<=G5728 or G3781;
	G6108<=G5898 or G5598;
	G6109<=G5900 or G5599;
	G6110<=G5883 or G5996;
	G6113<=G5902 or G5601;
	G6114<=G5904 or G5604;
	G6116<=G5910 or G5617;
	G6118<=G5911 or G5619;
	G6142<=G5909 or G3806;
	G6167<=G6056 or G6039;
	G6170<=G6061 or G6014;
	G6173<=G6066 or G6043;
	G6176<=G6068 or G6033;
	G6179<=G6077 or G6051;
	G6182<=G6047 or G6034;
	G6185<=G6055 or G5995;
	G6189<=G6060 or G6035;
	G6237<=G5912 or G2381;
	G6239<=G2339 or G6073;
	G6242<=G2356 or G6075;
	G6246<=G5665 or G5937;
	G6251<=G5668 or G5939;
	G6252<=G5905 or G2381;
	G6257<=G5671 or G5941;
	G6261<=G5673 or G5944;
	G6264<=G5675 or G5948;
	G6267<=G2953 or G5884;
	G6268<=G5677 or G5951;
	G6271<=G2955 or G5885;
	G6272<=G5679 or G5953;
	G6273<=G5681 or G5955;
	G6274<=G5682 or G5956;
	G6286<=G6238 or G6079;
	G6287<=G6241 or G6082;
	G6289<=G6240 or G6081;
	G6290<=G6245 or G6086;
	G6292<=G6243 or G6084;
	G6293<=G6244 or G6085;
	G6294<=G6249 or G6090;
	G6296<=G6247 or G6088;
	G6297<=G6248 or G6089;
	G6298<=G6255 or G6093;
	G6300<=G6253 or G6091;
	G6301<=G6254 or G6092;
	G6303<=G6258 or G6094;
	G6307<=G6262 or G6096;
	G6309<=G6265 or G6098;
	G6310<=G6269 or G6099;
	G6426<=G6288 or G6119;
	G6437<=G6302 or G6121;
	G6440<=G6336 or G5935;
	G6444<=G6338 or G5936;
	G6447<=G6340 or G5938;
	G6450<=G6341 or G5940;
	G6452<=G6342 or G5942;
	G6453<=G6343 or G5945;
	G6454<=G6344 or G5949;
	G6455<=G6345 or G5952;
	G6456<=G6346 or G5954;
	G6457<=G6352 or G6347;
	G6461<=G6353 or G6351;
	G6479<=I8349 or G6335;
	G6480<=I8360 or G6359;
	G6481<=I8367 or I8368 or I8369 or I8370;
	G6482<=I8376 or I8377 or I8378 or I8379;
	G6483<=I8385 or I8386 or I8387;
	G6485<=I8393 or I8394 or I8395;
	G6545<=G6468 or G4244;
	G6549<=G6473 or G4247;
	G6554<=G6337 or G6466;
	G6556<=G6339 or G6467;
	G6658<=G6132 or G6620;
	G6659<=G6634 or G6631;
	G6660<=G6640 or G6637;
	G6661<=I8773 or I8774;
	G6665<=I8778 or I8779;
	G6669<=G6613 or G4679;
	G6670<=G6557 or G6634 or G4410 or G2948;
	G6673<=G6559 or G6640 or G4416 or G2950;
	G6676<=G6631 or G6555;
	G6679<=G6637 or G6558;
	G6682<=G6478 or G6624 or G6623;
	G6683<=G6465 or G6622 or G6621;
	G6684<=G6250 or G6643;
	G6685<=G6256 or G6644;
	G6686<=G6259 or G6645;
	G6687<=G6260 or G6646;
	G6688<=G6263 or G6647;
	G6689<=G6266 or G6648;
	G6690<=G6270 or G6650;
	G6691<=G6275 or G6603;
	G6702<=G6659 or G496;
	G6703<=G6692 or G4831;
	G6704<=G6660 or G492;
	G6705<=G6693 or G4835;
	G6747<=G6614 or G6731;
	G6750<=G6670 or G6625 or G6736;
	G6754<=G6676 or G6625 or G6737;
	G6758<=G6673 or G6628 or G6738;
	G6762<=G6679 or G6628 or G6739;
	G6781<=G6718 or G6748;
	G6782<=G6719 or G6749;
	G6787<=G3758 or G6766;
	G6788<=G3760 or G6767;
	G6789<=G3764 or G6769;
	G6790<=G3765 or G6773;
	G6791<=G6768 or G3307;
	G6792<=G6770 or G3321;
	G6793<=G6771 or G3323;
	G6794<=G6777 or G3333;
	G6795<=G4867 or G6772;
	G6844<=I9057 or I9058 or I9059;
	G6845<=I9064 or I9065 or I9066;
	G6846<=G5860 or G6834;
	G6847<=G5861 or G6837;
	G6855<=G6851 or G2085;
	G6864<=G6852 or G2089;
	G6907<=G6874 or G3358;
	G6917<=G6909 or G6910;
	G6918<=G6911 or G6913;
	G6919<=G6912 or G6914;
	G6920<=G6915 or G6916;
	G6921<=G6908 or G6816;
	G6926<=G6798 or G6923;
	G6927<=G6799 or G6924;
	G6930<=G6740 or G6928;
	G6931<=G6741 or G6929;
	G6936<=G5438 or G6935;
	G6937<=G4616 or G6934;
	I7969<=G6194 or G5958 or G5975 or G5997;
	I7970<=G6015 or G6212 or G4950 or G4877;
	I7971<=G5202 or G4993 or G4967 or G4980;
	I7972<=G4915 or G5025;
	I7978<=G6194 or G5958 or G5975 or G5997;
	I7979<=G6015 or G6212 or G4950 or G4877;
	I7980<=G5202 or G4993 or G4967 or G4980;
	I7981<=G4915 or G5025;
	I7987<=G6194 or G5958 or G5975 or G5997;
	I7988<=G6015 or G6212 or G4950 or G4877;
	I7989<=G5202 or G4993 or G4967 or G4980;
	I7990<=G4915 or G5025;
	I8079<=G6194 or G5958 or G5975 or G5997;
	I8080<=G6015 or G6212 or G4950 or G4877;
	I8081<=G4894 or G4904 or G4993 or G4967;
	I8082<=G4980 or G4915 or G5025 or G5054;
	I8117<=G6194 or G5958 or G5975 or G5997;
	I8118<=G6015 or G6212 or G4950 or G4877;
	I8119<=G5202 or G4993 or G4967 or G4980;
	I8120<=G4915 or G5025;
	I8126<=G6194 or G5958 or G5975 or G5997;
	I8127<=G6015 or G6212 or G4950 or G4877;
	I8128<=G5202 or G4993 or G4967 or G4980;
	I8129<=G4915 or G5025;
	I8135<=G6194 or G5958 or G5975 or G5997;
	I8136<=G6015 or G6212 or G4950 or G4877;
	I8137<=G4894 or G4904 or G4993 or G4967;
	I8138<=G4980 or G4915 or G5025 or G5054;
	I8208<=G6194 or G5958 or G5975 or G5997;
	I8209<=G6015 or G6212 or G4950 or G4877;
	I8210<=G5202 or G4993 or G4967 or G4980;
	I8211<=G4915 or G5025;
	I8345<=G6326 or G6135 or G6140 or G6157;
	I8346<=G6159 or G6334 or G5163 or G5191;
	I8347<=G5188 or G5157 or G5154 or G5193;
	I8348<=G5229 or G5234 or G5218 or G5225;
	I8349<=I8345 or I8346 or I8347 or I8348;
	I8356<=G6311 or G6123 or G6125 or G6141;
	I8357<=G6145 or G6318 or G5171 or G5187;
	I8358<=G5192 or G5153 or G5158 or G5197;
	I8359<=G5232 or G5236 or G5216 or G5226;
	I8360<=I8356 or I8357 or I8358 or I8359;
	I8367<=G6313 or G6124 or G6127 or G6144;
	I8368<=G6148 or G6321 or G5176 or G5184;
	I8369<=G5165 or G5159 or G5233 or G5240;
	I8370<=G5214 or G6358;
	I8376<=G6315 or G6126 or G6129 or G6146;
	I8377<=G6150 or G6324 or G5180 or G5181;
	I8378<=G5173 or G5166 or G5235 or G5245;
	I8379<=G5212 or G6357;
	I8385<=G6316 or G6128 or G6131 or G6149;
	I8386<=G6152 or G6327 or G5183 or G5177;
	I8387<=G5178 or G5209 or G6281;
	I8393<=G6317 or G6130 or G6133 or G6151;
	I8394<=G6154 or G6329 or G5186 or G5172;
	I8395<=G5182 or G5200 or G6280;
	I8773<=G6610 or G6608 or G6606 or G6604;
	I8774<=G6655 or G6653 or G6651 or G6649;
	I8778<=G6612 or G6611 or G6609 or G6607;
	I8779<=G6605 or G6656 or G6654 or G6652;
	I9057<=G6320 or G6828 or G6830 or G6153;
	I9058<=G6156 or G6331 or G5190 or G5164;
	I9059<=G5185 or G5198 or G6279;
	I9064<=G6323 or G6829 or G6831 or G6155;
	I9065<=G6158 or G6333 or G5152 or G5156;
	I9066<=G5189 or G5269 or G6400;
	G1418<= not (G486 or G943);
	G1422<= not (G1039 or G913);
	G1449<= not (G489 or G1048);
	G1459<= not (G926 or G950 or G948);
	G1470<= not (G937 or G930 or G928);
	G1473<= not (G944 or G941 or G939);
	G1474<= not (G760 or G754);
	G1481<= not (G815 or G809);
	G1518<= not (G980 or G965);
	G1560<= not (G996 or G980);
	G1603<= not (G1039 or G658);
	G1879<= not (G1603 or G1416);
	G2433<= not (G1418 or G1449);
	G2908<= not (G536 or G2010 or G541);
	G3528<= not (G1802 or G3167);
	G3621<= not (G1407 or G2842);
	G3647<= not (G2731 or G2719 or G2698);
	G3656<= not (G2769 or G2757 or G2745);
	G3664<= not (G2804 or G2791 or G2780);
	G3903<= not (G3505 or G471);
	G3905<= not (G3512 or G478);
	G3923<= not (G3378 or G3381);
	G3925<= not (G3303 or G3315);
	G3926<= not (G3338 or G3350);
	G3927<= not (G3382 or G3383);
	G3929<= not (G3373 or G3376);
	G3930<= not (G3317 or G3328);
	G3931<= not (G3353 or G3361);
	G3933<= not (G3327 or G3336);
	G3934<= not (G3377 or G3379);
	G3939<= not (G3340 or G3351);
	G3956<= not (G3337 or G3349);
	G3958<= not (G3316 or G3326);
	G3959<= not (G3352 or G3360);
	G3965<= not (G3359 or G3367);
	G3966<= not (G3329 or G3339);
	G3973<= not (G3368 or G3374);
	G4000<= not (G1250 or G3425);
	G4235<= not (G3780 or G3362);
	G4238<= not (G3755 or G3279);
	G4239<= not (G3763 or G3296);
	G4240<= not (G1589 or G1879 or G3793);
	G4241<= not (G3774 or G3341);
	G4245<= not (G3759 or G3288);
	G4261<= not (G3762 or G3295);
	G4266<= not (G3757 or G3283);
	G4272<= not (G3767 or G3319);
	G4432<= not (G923 or G4253);
	G4568<= not (G4233 or G3924);
	G4578<= not (G4234 or G3928);
	G4581<= not (G4156 or G4160);
	G4584<= not (G4164 or G4168);
	G4585<= not (G4171 or G4177);
	G4586<= not (G4161 or G4165);
	G4589<= not (G4180 or G4183);
	G4590<= not (G4169 or G4172);
	G4591<= not (G4178 or G4181);
	G4596<= not (G4184 or G4186);
	G4774<= not (G4442 or G4445);
	G4776<= not (G4449 or G4453);
	G4777<= not (G4457 or G4459);
	G4779<= not (G4461 or G4464);
	G4877<= not (G952 or G4680);
	G4950<= not (G1472 or G4680);
	G4967<= not (G4674 or G952);
	G4993<= not (G4674 or G1477);
	G5048<= not (G4819 or G3491 or G3559);
	G5088<= not (G4691 or G4697);
	G5091<= not (G4698 or G4701);
	G5093<= not (G4683 or G4684);
	G5094<= not (G4685 or G4686);
	G5227<= not (G5019 or G3559);
	G5249<= not (G4868 or G4870);
	G5265<= not (G4863 or G4865);
	G5324<= not (G5069 or G4410 or G766);
	G5325<= not (G5077 or G4416 or G821);
	G5418<= not (G5162 or G5169);
	G5423<= not (G5170 or G5175);
	G5541<= not (G5388 or G1880);
	G5552<= not (G5354 or G5356);
	G5561<= not (G5391 or G1589 or G3793 or G1880);
	G5731<= not (G952 or G5688);
	G5753<= not (G1477 or G5688);
	G6073<= not (G197 or G5862);
	G6075<= not (G269 or G5863);
	G6279<= not (I7969 or I7970 or I7971 or I7972);
	G6280<= not (I7978 or I7979 or I7980 or I7981);
	G6281<= not (I7987 or I7988 or I7989 or I7990);
	G6335<= not (I8079 or I8080 or I8081 or I8082);
	G6357<= not (I8117 or I8118 or I8119 or I8120);
	G6358<= not (I8126 or I8127 or I8128 or I8129);
	G6359<= not (I8135 or I8136 or I8137 or I8138);
	G6400<= not (I8208 or I8209 or I8210 or I8211);
	G6427<= not (G6376 or G4086 or G4074 or G4068);
	G6429<= not (G6376 or G4086 or G4074 or G4302);
	G6430<= not (G6385 or G3733 or G4092 or G4080);
	G6432<= not (G6376 or G4086 or G4309 or G4068);
	G6433<= not (G6385 or G3733 or G4092 or G4314);
	G6435<= not (G6376 or G4086 or G4309 or G4302);
	G6436<= not (G6385 or G3733 or G4328 or G4080);
	G6438<= not (G6376 or G4323 or G4074 or G4068);
	G6439<= not (G6385 or G3733 or G4328 or G4314);
	G6442<= not (G6376 or G4323 or G4074 or G4302);
	G6443<= not (G6385 or G4334 or G4092 or G4080);
	G6445<= not (G6376 or G4323 or G4309 or G4068);
	G6446<= not (G6385 or G4334 or G4092 or G4314);
	G6448<= not (G6376 or G4323 or G4309 or G4302);
	G6449<= not (G6385 or G4334 or G4328 or G4080);
	G6451<= not (G6385 or G4334 or G4328 or G4314);
	G6492<= not (G6348 or G1734);
	G6494<= not (G952 or G6348);
	G6495<= not (G6354 or G1775);
	G6496<= not (G952 or G6354);
end RTL;
