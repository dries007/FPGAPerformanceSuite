-- File created by Bench2VHDL
-- Name: s1423
-- File: bench/s1423.bench
-- Timestamp: 2019-05-21T22:08:29.256842
--
-- Original File
-- =============
--	# s1423
--	# 17 inputs
--	# 5 outputs
--	# 74 D-type flipflops
--	# 167 inverters
--	# 490 gates (197 ANDs + 64 NANDs + 137 ORs + 92 NORs)
--	
--	INPUT(G0)
--	INPUT(G1)
--	INPUT(G2)
--	INPUT(G3)
--	INPUT(G4)
--	INPUT(G5)
--	INPUT(G6)
--	INPUT(G7)
--	INPUT(G8)
--	INPUT(G9)
--	INPUT(G10)
--	INPUT(G11)
--	INPUT(G12)
--	INPUT(G13)
--	INPUT(G14)
--	INPUT(G15)
--	INPUT(G16)
--	
--	OUTPUT(G726)
--	OUTPUT(G729)
--	OUTPUT(G702)
--	OUTPUT(G727)
--	OUTPUT(G701BF)
--	
--	G22 = DFF(G332BF)
--	G23 = DFF(G328BF)
--	G24 = DFF(G109)
--	G25 = DFF(G113)
--	G26 = DFF(G118)
--	G27 = DFF(G125)
--	G28 = DFF(G129)
--	G29 = DFF(G140)
--	G30 = DFF(G144)
--	G31 = DFF(G149)
--	G32 = DFF(G154)
--	G33 = DFF(G159)
--	G34 = DFF(G166)
--	G35 = DFF(G175)
--	G36 = DFF(G189)
--	G37 = DFF(G193)
--	G38 = DFF(G198)
--	G39 = DFF(G208)
--	G40 = DFF(G214)
--	G41 = DFF(G218)
--	G42 = DFF(G237)
--	G43 = DFF(G242)
--	G44 = DFF(G247)
--	G45 = DFF(G252)
--	G46 = DFF(G260)
--	G47 = DFF(G303)
--	G48 = DFF(G309)
--	G49 = DFF(G315)
--	G50 = DFF(G321)
--	G51 = DFF(G360)
--	G52 = DFF(G365)
--	G53 = DFF(G373)
--	G54 = DFF(G379)
--	G55 = DFF(G384)
--	G56 = DFF(G392)
--	G57 = DFF(G397)
--	G58 = DFF(G405)
--	G59 = DFF(G408)
--	G60 = DFF(G416)
--	G61 = DFF(G424)
--	G62 = DFF(G427)
--	G63 = DFF(G438)
--	G64 = DFF(G441)
--	G65 = DFF(G447)
--	G66 = DFF(G451)
--	G67 = DFF(G459)
--	G68 = DFF(G464)
--	G69 = DFF(G469)
--	G70 = DFF(G477)
--	G71 = DFF(G494)
--	G72 = DFF(G498)
--	G73 = DFF(G503)
--	G74 = DFF(G526)
--	G75 = DFF(G531)
--	G76 = DFF(G536)
--	G77 = DFF(G541)
--	G78 = DFF(G548)
--	G79 = DFF(G565)
--	G80 = DFF(G569)
--	G81 = DFF(G573)
--	G82 = DFF(G577)
--	G83 = DFF(G590)
--	G84 = DFF(G608)
--	G85 = DFF(G613)
--	G86 = DFF(G657)
--	G87 = DFF(G663)
--	G88 = DFF(G669)
--	G89 = DFF(G675)
--	G90 = DFF(G682)
--	G91 = DFF(G687)
--	G92 = DFF(G693)
--	G93 = DFF(G705)
--	G94 = DFF(G707)
--	G95 = DFF(G713)
--	
--	I1 = NOT(G332)
--	G332BF = NOT(I1)
--	I12 = NOT(G328)
--	G328BF = NOT(I12)
--	G108 = NOT(G712)
--	G111 = NOT(G24)
--	G112 = NOT(G712)
--	G117 = NOT(G712)
--	G124 = NOT(G712)
--	G127 = NOT(G27)
--	G128 = NOT(G712)
--	G139 = NOT(G712)
--	G142 = NOT(G29)
--	G143 = NOT(G712)
--	G148 = NOT(G712)
--	G153 = NOT(G712)
--	G158 = NOT(G712)
--	G165 = NOT(G712)
--	G174 = NOT(G712)
--	G176 = NOT(G35)
--	G178 = NOT(G34)
--	G179 = NOT(G180)
--	G180 = NOT(G92)
--	G188 = NOT(G712)
--	G191 = NOT(G36)
--	G192 = NOT(G712)
--	G197 = NOT(G712)
--	G204 = NOT(G38)
--	G207 = NOT(G712)
--	G210 = NOT(G39)
--	G213 = NOT(G712)
--	G216 = NOT(G40)
--	G217 = NOT(G712)
--	G236 = NOT(G259)
--	G241 = NOT(G259)
--	G246 = NOT(G259)
--	G251 = NOT(G259)
--	G258 = NOT(G259)
--	G296 = NOT(G297)
--	G302 = NOT(G712)
--	G305 = NOT(G324)
--	G308 = NOT(G712)
--	G311 = NOT(G324)
--	G314 = NOT(G712)
--	G317 = NOT(G324)
--	G320 = NOT(G712)
--	G323 = NOT(G324)
--	G336 = NOT(G355)
--	G339 = NOT(G355)
--	G343 = NOT(G348)
--	G347 = NOT(G348)
--	G348 = NOT(G91)
--	G351 = NOT(G645)
--	G354 = NOT(G355)
--	G359 = NOT(G372)
--	G364 = NOT(G372)
--	G371 = NOT(G372)
--	G378 = NOT(G391)
--	G383 = NOT(G391)
--	G390 = NOT(G391)
--	G396 = NOT(G404)
--	G403 = NOT(G404)
--	G407 = NOT(G712)
--	G415 = NOT(G423)
--	G422 = NOT(G423)
--	G426 = NOT(G712)
--	G437 = NOT(G712)
--	G440 = NOT(G712)
--	G445 = NOT(G65)
--	G446 = NOT(G712)
--	G449 = NOT(G66)
--	G450 = NOT(G712)
--	G455 = NOT(G456)
--	G458 = NOT(G476)
--	G463 = NOT(G476)
--	G468 = NOT(G476)
--	G475 = NOT(G476)
--	G486 = NOT(G712)
--	G491 = NOT(G500)
--	G495 = NOT(G500)
--	G499 = NOT(G500)
--	G504 = NOT(G511)
--	G507 = NOT(G511)
--	G510 = NOT(G511)
--	G511 = NOT(G63)
--	G525 = NOT(G589)
--	G530 = NOT(G589)
--	G535 = NOT(G589)
--	G540 = NOT(G589)
--	G547 = NOT(G589)
--	G562 = NOT(G610)
--	G566 = NOT(G610)
--	G570 = NOT(G610)
--	G574 = NOT(G610)
--	G588 = NOT(G589)
--	G595 = NOT(G593)
--	G596 = NOT(G597)
--	G600 = NOT(G601)
--	G605 = NOT(G610)
--	G609 = NOT(G610)
--	G614 = NOT(G64)
--	G615 = NOT(G616)
--	G617 = NOT(G645)
--	G620 = NOT(G645)
--	G623 = NOT(G645)
--	G626 = NOT(G645)
--	G629 = NOT(G645)
--	G632 = NOT(G645)
--	G635 = NOT(G645)
--	G638 = NOT(G645)
--	G641 = NOT(G645)
--	G644 = NOT(G645)
--	G645 = NOT(G90)
--	G656 = NOT(G712)
--	G658 = NOT(G659)
--	I1162 = NOT(G13)
--	G659 = NOT(I1162)
--	G661 = NOT(G94)
--	G662 = NOT(G712)
--	G665 = NOT(G678)
--	G668 = NOT(G712)
--	G671 = NOT(G678)
--	G674 = NOT(G712)
--	G677 = NOT(G678)
--	I1183 = NOT(G11)
--	G678 = NOT(I1183)
--	G685 = NOT(G696)
--	G689 = NOT(G696)
--	G695 = NOT(G696)
--	I1203 = NOT(G10)
--	G696 = NOT(I1203)
--	G701 = NOT(G15)
--	I1211 = NOT(G701)
--	G701BF = NOT(I1211)
--	G704 = NOT(G712)
--	G706 = NOT(G712)
--	G711 = NOT(G712)
--	G712 = NOT(G14)
--	G714 = NOT(G701)
--	I1227 = NOT(G6)
--	G715 = NOT(I1227)
--	I1230 = NOT(G7)
--	G716 = NOT(I1230)
--	I1233 = NOT(G8)
--	G717 = NOT(I1233)
--	I1236 = NOT(G9)
--	G718 = NOT(I1236)
--	I1239 = NOT(G12)
--	G719 = NOT(I1239)
--	I1242 = NOT(G0)
--	G720 = NOT(I1242)
--	I1245 = NOT(G1)
--	G721 = NOT(I1245)
--	I1248 = NOT(G2)
--	G722 = NOT(I1248)
--	I1251 = NOT(G3)
--	G723 = NOT(I1251)
--	I1254 = NOT(G4)
--	G724 = NOT(I1254)
--	I1257 = NOT(G5)
--	G725 = NOT(I1257)
--	I1260 = NOT(G93)
--	G726 = NOT(I1260)
--	I1264 = NOT(G16)
--	G728 = NOT(I1264)
--	I1267 = NOT(G95)
--	G729 = NOT(I1267)
--	
--	G101 = AND(G630, G631)
--	G102 = AND(G633, G634)
--	G103 = AND(G636, G637)
--	G104 = AND(G639, G640)
--	G105 = AND(G642, G643)
--	G109 = AND(G106, G108)
--	G113 = AND(G114, G112)
--	G116 = AND(G133, G25)
--	G118 = AND(G119, G117)
--	G121 = AND(G134, G26)
--	G125 = AND(G122, G124)
--	G129 = AND(G130, G128)
--	G132 = AND(G136, G28)
--	G133 = AND(G700, G111)
--	G134 = AND(G133, G25)
--	G135 = AND(G134, G26)
--	G136 = AND(G135, G127)
--	G140 = AND(G137, G139)
--	G144 = AND(G145, G143)
--	G147 = AND(G168, G30)
--	G149 = AND(G150, G148)
--	G152 = AND(G169, G31)
--	G154 = AND(G155, G153)
--	G157 = AND(G170, G32)
--	G159 = AND(G160, G158)
--	G162 = AND(G171, G33)
--	G166 = AND(G163, G165)
--	G168 = AND(G177, G142)
--	G169 = AND(G168, G30)
--	G170 = AND(G169, G31)
--	G171 = AND(G170, G32)
--	G172 = AND(G171, G33)
--	G173 = AND(G172, G34)
--	G175 = AND(G176, G174)
--	G185 = AND(G181, G182)
--	G189 = AND(G186, G188)
--	G193 = AND(G194, G192)
--	G196 = AND(G202, G37)
--	G198 = AND(G199, G197)
--	G201 = AND(G203, G38)
--	G202 = AND(G522, G191)
--	G203 = AND(G202, G37)
--	G208 = AND(G205, G207)
--	G214 = AND(G211, G213)
--	G218 = AND(G219, G217)
--	G221 = AND(G223, G41)
--	G222 = AND(G183, G210)
--	G223 = AND(G222, G216)
--	G224 = AND(G203, G38)
--	G225 = AND(G204, G203)
--	G226 = AND(G136, G28)
--	G227 = AND(G172, G178)
--	G228 = AND(G223, G41)
--	G229 = AND(G432, G62)
--	G237 = AND(G238, G236)
--	G240 = AND(G299, G42)
--	G242 = AND(G243, G241)
--	G245 = AND(G262, G43)
--	G247 = AND(G248, G246)
--	G250 = AND(G263, G44)
--	G252 = AND(G253, G251)
--	G255 = AND(G264, G45)
--	G259 = AND(G624, G625)
--	G260 = AND(G256, G258)
--	G261 = AND(G265, G46)
--	G262 = AND(G299, G42)
--	G263 = AND(G262, G43)
--	G264 = AND(G263, G44)
--	G265 = AND(G264, G45)
--	G271 = AND(G275, G266)
--	G272 = AND(G276, G277)
--	G273 = AND(G278, G279)
--	G274 = AND(G280, G281)
--	G303 = AND(G304, G302)
--	G304 = AND(G306, G307)
--	G309 = AND(G310, G308)
--	G310 = AND(G312, G313)
--	G315 = AND(G316, G314)
--	G316 = AND(G318, G319)
--	G321 = AND(G322, G320)
--	G322 = AND(G325, G326)
--	G329 = AND(G331, G714)
--	G330 = AND(G332, G714)
--	G335 = AND(G337, G338)
--	G342 = AND(G344, G345)
--	G346 = AND(G349, G350)
--	G358 = AND(G523, G53)
--	G360 = AND(G361, G359)
--	G363 = AND(G523, G51)
--	G365 = AND(G366, G364)
--	G368 = AND(G375, G52)
--	G373 = AND(G369, G371)
--	G374 = AND(G376, G53)
--	G375 = AND(G523, G51)
--	G376 = AND(G375, G52)
--	G377 = AND(G183, G54, G56)
--	G379 = AND(G380, G378)
--	G382 = AND(G183, G54)
--	G384 = AND(G385, G383)
--	G387 = AND(G394, G55)
--	G392 = AND(G388, G390)
--	G393 = AND(G395, G56)
--	G394 = AND(G183, G54)
--	G395 = AND(G394, G55)
--	G397 = AND(G398, G396)
--	G400 = AND(G335, G57)
--	G405 = AND(G401, G403)
--	G406 = AND(G412, G58)
--	G408 = AND(G409, G407)
--	G411 = AND(G413, G59)
--	G412 = AND(G335, G57)
--	G413 = AND(G335, G58)
--	G414 = AND(G413, G59)
--	G416 = AND(G417, G415)
--	G419 = AND(G358, G60)
--	G424 = AND(G420, G422)
--	G425 = AND(G431, G61)
--	G427 = AND(G428, G426)
--	G430 = AND(G432, G62)
--	G431 = AND(G358, G60)
--	G432 = AND(G358, G61)
--	G433 = AND(G356, G357)
--	G435 = AND(G340, G341)
--	G436 = AND(G352, G353)
--	G438 = AND(G439, G437)
--	G441 = AND(G442, G440)
--	G443 = AND(G615, G511)
--	G447 = AND(G448, G446)
--	G451 = AND(G452, G450)
--	G453 = AND(G615, G445)
--	G457 = AND(G455, G449, G728)
--	G459 = AND(G460, G458)
--	G462 = AND(G434, G67)
--	G464 = AND(G465, G463)
--	G467 = AND(G479, G68)
--	G469 = AND(G470, G468)
--	G472 = AND(G480, G69)
--	G477 = AND(G473, G475)
--	G478 = AND(G481, G70)
--	G479 = AND(G434, G67)
--	G480 = AND(G479, G68)
--	G481 = AND(G480, G69)
--	G488 = AND(G505, G506)
--	G489 = AND(G508, G509)
--	G490 = AND(G512, G513)
--	G494 = AND(G492, G493)
--	G498 = AND(G496, G497)
--	G503 = AND(G501, G502)
--	G526 = AND(G527, G525)
--	G529 = AND(G604, G74)
--	G531 = AND(G532, G530)
--	G534 = AND(G550, G75)
--	G536 = AND(G537, G535)
--	G539 = AND(G551, G76)
--	G541 = AND(G542, G540)
--	G544 = AND(G552, G77)
--	G548 = AND(G545, G547)
--	G549 = AND(G553, G78)
--	G550 = AND(G604, G74)
--	G551 = AND(G550, G75)
--	G552 = AND(G551, G76)
--	G553 = AND(G552, G77)
--	G565 = AND(G563, G564)
--	G569 = AND(G567, G568)
--	G573 = AND(G571, G572)
--	G577 = AND(G575, G576)
--	G589 = AND(G627, G628)
--	G590 = AND(G591, G588)
--	G592 = AND(G594, G595)
--	G601 = AND(G621, G622)
--	G604 = AND(G433, G524)
--	G608 = AND(G606, G607)
--	G613 = AND(G611, G612)
--	G648 = AND(G646, G647)
--	G649 = AND(G618, G619)
--	G650 = AND(G226, G661)
--	G651 = AND(G227, G87)
--	G652 = AND(G228, G88)
--	G653 = AND(G229, G89)
--	G654 = AND(G90, G476)
--	G655 = AND(G91, G476)
--	G657 = AND(G659, G656)
--	G663 = AND(G664, G662)
--	G664 = AND(G666, G667)
--	G669 = AND(G670, G668)
--	G670 = AND(G672, G673)
--	G675 = AND(G676, G674)
--	G676 = AND(G679, G680)
--	G683 = AND(G684, G685)
--	G688 = AND(G690, G691)
--	G694 = AND(G697, G698)
--	G702 = AND(G703, G645)
--	G705 = AND(G230, G704)
--	G707 = AND(G708, G706)
--	G709 = AND(G678, G89)
--	G713 = AND(G599, G711)
--	G727 = AND(G476, G645)
--	
--	G110 = OR(G700, G111)
--	G126 = OR(G135, G127)
--	G141 = OR(G177, G142)
--	G167 = OR(G172, G178)
--	G177 = OR(G180, G226)
--	G181 = OR(G178, G180)
--	G182 = OR(G35, G179)
--	G183 = OR(G180, G227)
--	G184 = OR(G180, G173)
--	G190 = OR(G522, G191)
--	G209 = OR(G183, G210)
--	G215 = OR(G222, G216)
--	G235 = OR(G649, G233)
--	G275 = OR(G101, G42)
--	G276 = OR(G102, G43)
--	G277 = OR(G267, G271)
--	G278 = OR(G103, G44)
--	G279 = OR(G268, G272)
--	G280 = OR(G104, G45)
--	G281 = OR(G269, G273)
--	G282 = OR(G105, G46)
--	G283 = OR(G270, G274)
--	G291 = OR(G42, G101)
--	G292 = OR(G43, G102)
--	G293 = OR(G44, G103)
--	G294 = OR(G45, G104)
--	G295 = OR(G46, G105)
--	G300 = OR(G50, G49, G48, G47)
--	G306 = OR(G47, G324)
--	G307 = OR(G719, G305)
--	G312 = OR(G48, G324)
--	G313 = OR(G47, G311)
--	G318 = OR(G49, G324)
--	G319 = OR(G48, G317)
--	G324 = OR(G377, G348)
--	G325 = OR(G50, G324)
--	G326 = OR(G49, G323)
--	G333 = OR(G300, G714)
--	G334 = OR(G301, G714)
--	G337 = OR(G224, G355)
--	G338 = OR(G183, G336)
--	G340 = OR(G38, G355)
--	G341 = OR(G185, G339)
--	G344 = OR(G229, G348)
--	G345 = OR(G414, G343)
--	G349 = OR(G62, G348)
--	G350 = OR(G59, G347)
--	G352 = OR(G346, G645)
--	G353 = OR(G35, G351)
--	G355 = OR(G457, G645)
--	G356 = OR(G225, G355)
--	G357 = OR(G184, G354)
--	G372 = OR(G712, G358)
--	G391 = OR(G712, G377)
--	G404 = OR(G712, G413)
--	G423 = OR(G712, G432)
--	G434 = OR(G342, G645)
--	G439 = OR(G435, G63)
--	G448 = OR(G615, G65)
--	G456 = OR(G83, G524)
--	G492 = OR(G71, G500)
--	G493 = OR(G488, G491)
--	G496 = OR(G72, G500)
--	G497 = OR(G489, G495)
--	G500 = OR(G654, G712)
--	G501 = OR(G73, G500)
--	G502 = OR(G490, G499)
--	G505 = OR(G723, G511)
--	G506 = OR(G720, G504)
--	G508 = OR(G724, G511)
--	G509 = OR(G721, G507)
--	G512 = OR(G725, G511)
--	G513 = OR(G722, G510)
--	G518 = OR(G71, G67)
--	G519 = OR(G72, G68)
--	G520 = OR(G73, G69)
--	G521 = OR(G487, G70)
--	G522 = OR(G348, G228)
--	G523 = OR(G348, G414)
--	G524 = OR(G554, G555)
--	G563 = OR(G79, G610)
--	G564 = OR(G715, G562)
--	G567 = OR(G80, G610)
--	G568 = OR(G716, G566)
--	G571 = OR(G81, G610)
--	G572 = OR(G717, G570)
--	G575 = OR(G82, G610)
--	G576 = OR(G718, G574)
--	G583 = OR(G79, G74)
--	G584 = OR(G80, G75)
--	G585 = OR(G81, G76)
--	G586 = OR(G82, G77)
--	G587 = OR(G561, G78)
--	G591 = OR(G592, G604)
--	G594 = OR(G83, G593)
--	G602 = OR(G85, G601)
--	G603 = OR(G600, G84)
--	G606 = OR(G84, G610)
--	G607 = OR(G696, G605)
--	G610 = OR(G655, G712)
--	G611 = OR(G85, G610)
--	G612 = OR(G678, G609)
--	G618 = OR(G457, G645)
--	G619 = OR(G715, G617)
--	G621 = OR(G614, G645)
--	G622 = OR(G717, G620)
--	G624 = OR(G476, G645)
--	G625 = OR(G716, G623)
--	G627 = OR(G476, G645)
--	G628 = OR(G718, G626)
--	G630 = OR(G96, G645)
--	G631 = OR(G720, G629)
--	G633 = OR(G97, G645)
--	G634 = OR(G721, G632)
--	G636 = OR(G98, G645)
--	G637 = OR(G722, G635)
--	G639 = OR(G99, G645)
--	G640 = OR(G723, G638)
--	G642 = OR(G100, G645)
--	G643 = OR(G724, G641)
--	G646 = OR(G456, G645)
--	G647 = OR(G725, G644)
--	G666 = OR(G87, G678)
--	G667 = OR(G661, G665)
--	G672 = OR(G88, G678)
--	G673 = OR(G87, G671)
--	G679 = OR(G89, G678)
--	G680 = OR(G88, G677)
--	G682 = OR(G681, G699)
--	G684 = OR(G645, G696)
--	G687 = OR(G686, G699)
--	G690 = OR(G348, G696)
--	G691 = OR(G645, G689)
--	G693 = OR(G692, G699)
--	G697 = OR(G180, G696)
--	G698 = OR(G348, G695)
--	G699 = OR(G658, G712)
--	
--	G96 = NAND(G74, G596)
--	G97 = NAND(G75, G596)
--	G98 = NAND(G76, G596)
--	G99 = NAND(G77, G596)
--	G100 = NAND(G78, G596)
--	G106 = NAND(G107, G110)
--	G107 = NAND(G700, G111)
--	G122 = NAND(G123, G126)
--	G123 = NAND(G135, G127)
--	G137 = NAND(G138, G141)
--	G138 = NAND(G177, G142)
--	G163 = NAND(G164, G167)
--	G164 = NAND(G172, G178)
--	G186 = NAND(G187, G190)
--	G187 = NAND(G522, G191)
--	G205 = NAND(G206, G209)
--	G206 = NAND(G183, G210)
--	G211 = NAND(G212, G215)
--	G212 = NAND(G222, G216)
--	G230 = NAND(G234, G235)
--	G231 = NAND(G435, G648)
--	G232 = NAND(G296, G298, G435)
--	G233 = NAND(G700, G232, G231)
--	G234 = NAND(G649, G436)
--	G266 = NAND(G286, G291)
--	G267 = NAND(G287, G292)
--	G268 = NAND(G288, G293)
--	G269 = NAND(G284, G294)
--	G270 = NAND(G285, G295)
--	G284 = NAND(G45, G104)
--	G285 = NAND(G46, G105)
--	G286 = NAND(G42, G101)
--	G287 = NAND(G43, G102)
--	G288 = NAND(G44, G103)
--	G297 = NAND(G289, G290)
--	G298 = NAND(G297, G700)
--	G301 = NAND(G50, G49, G48, G47)
--	G331 = NAND(G333, G22)
--	G332 = NAND(G334, G331)
--	G476 = NAND(G486, G616)
--	G482 = NAND(G514, G518)
--	G483 = NAND(G515, G519)
--	G484 = NAND(G516, G520)
--	G485 = NAND(G517, G521)
--	G514 = NAND(G71, G67)
--	G515 = NAND(G72, G68)
--	G516 = NAND(G73, G69)
--	G517 = NAND(G487, G70)
--	G554 = NAND(G556, G557, G558)
--	G555 = NAND(G559, G560)
--	G556 = NAND(G578, G583)
--	G557 = NAND(G579, G584)
--	G558 = NAND(G580, G585)
--	G559 = NAND(G581, G586)
--	G560 = NAND(G582, G587)
--	G578 = NAND(G79, G74)
--	G579 = NAND(G80, G75)
--	G580 = NAND(G81, G76)
--	G581 = NAND(G82, G77)
--	G582 = NAND(G561, G78)
--	G597 = NAND(G602, G603)
--	G598 = NAND(G435, G83)
--	G616 = NAND(G482, G483, G484, G485)
--	G700 = NAND(G282, G283)
--	
--	G114 = NOR(G115, G116)
--	G115 = NOR(G133, G25)
--	G119 = NOR(G120, G121)
--	G120 = NOR(G134, G26)
--	G130 = NOR(G131, G132)
--	G131 = NOR(G136, G28)
--	G145 = NOR(G146, G147)
--	G146 = NOR(G168, G30)
--	G150 = NOR(G151, G152)
--	G151 = NOR(G169, G31)
--	G155 = NOR(G156, G157)
--	G156 = NOR(G170, G32)
--	G160 = NOR(G161, G162)
--	G161 = NOR(G171, G33)
--	G194 = NOR(G195, G196)
--	G195 = NOR(G202, G37)
--	G199 = NOR(G200, G201)
--	G200 = NOR(G203, G38)
--	G219 = NOR(G220, G221)
--	G220 = NOR(G223, G41)
--	G238 = NOR(G239, G240)
--	G239 = NOR(G299, G42)
--	G243 = NOR(G244, G245)
--	G244 = NOR(G262, G43)
--	G248 = NOR(G249, G250)
--	G249 = NOR(G263, G44)
--	G253 = NOR(G254, G255)
--	G254 = NOR(G264, G45)
--	G256 = NOR(G257, G261)
--	G257 = NOR(G265, G46)
--	G289 = NOR(G270, G269, G268)
--	G290 = NOR(G267, G266)
--	G299 = NOR(G301, G328)
--	G327 = NOR(G330, G23)
--	G328 = NOR(G329, G327)
--	G361 = NOR(G362, G363)
--	G362 = NOR(G523, G51)
--	G366 = NOR(G367, G368)
--	G367 = NOR(G375, G52)
--	G369 = NOR(G370, G374)
--	G370 = NOR(G376, G53)
--	G380 = NOR(G381, G382)
--	G381 = NOR(G183, G54)
--	G385 = NOR(G386, G387)
--	G386 = NOR(G394, G55)
--	G388 = NOR(G389, G393)
--	G389 = NOR(G395, G56)
--	G398 = NOR(G399, G400)
--	G399 = NOR(G335, G57)
--	G401 = NOR(G402, G406)
--	G402 = NOR(G412, G58)
--	G409 = NOR(G410, G411)
--	G410 = NOR(G413, G59)
--	G417 = NOR(G418, G419)
--	G418 = NOR(G358, G60)
--	G420 = NOR(G421, G425)
--	G421 = NOR(G431, G61)
--	G428 = NOR(G429, G430)
--	G429 = NOR(G432, G62)
--	G442 = NOR(G443, G444)
--	G444 = NOR(G615, G64)
--	G452 = NOR(G453, G454)
--	G454 = NOR(G615, G66)
--	G460 = NOR(G461, G462)
--	G461 = NOR(G434, G67)
--	G465 = NOR(G466, G467)
--	G466 = NOR(G479, G68)
--	G470 = NOR(G471, G472)
--	G471 = NOR(G480, G69)
--	G473 = NOR(G474, G478)
--	G474 = NOR(G481, G70)
--	G487 = NOR(G71, G72, G73)
--	G527 = NOR(G528, G529)
--	G528 = NOR(G604, G74)
--	G532 = NOR(G533, G534)
--	G533 = NOR(G550, G75)
--	G537 = NOR(G538, G539)
--	G538 = NOR(G551, G76)
--	G542 = NOR(G543, G544)
--	G543 = NOR(G552, G77)
--	G545 = NOR(G546, G549)
--	G546 = NOR(G553, G78)
--	G561 = NOR(G79, G80, G81, G82)
--	G593 = NOR(G435, G524)
--	G599 = NOR(G598, G597)
--	G660 = NOR(G658, G86)
--	G681 = NOR(G683, G660)
--	G686 = NOR(G688, G660)
--	G692 = NOR(G694, G660)
--	G703 = NOR(G650, G651, G652, G653)
--	G708 = NOR(G709, G710)
--	G710 = NOR(G678, G94)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s1423 is
	port (
		CLK: in std_logic;
		G0: in std_logic;
		G1: in std_logic;
		G2: in std_logic;
		G3: in std_logic;
		G4: in std_logic;
		G5: in std_logic;
		G6: in std_logic;
		G7: in std_logic;
		G8: in std_logic;
		G9: in std_logic;
		G10: in std_logic;
		G11: in std_logic;
		G12: in std_logic;
		G13: in std_logic;
		G14: in std_logic;
		G15: in std_logic;
		G16: in std_logic;
		G701BF: out std_logic;
		G702: out std_logic;
		G726: out std_logic;
		G727: out std_logic;
		G729: out std_logic
	);
end entity;

architecture RTL of s1423 is
	attribute dont_touch: boolean;

	signal G22: std_logic; attribute dont_touch of G22: signal is true;
	signal G23: std_logic; attribute dont_touch of G23: signal is true;
	signal G24: std_logic; attribute dont_touch of G24: signal is true;
	signal G25: std_logic; attribute dont_touch of G25: signal is true;
	signal G26: std_logic; attribute dont_touch of G26: signal is true;
	signal G27: std_logic; attribute dont_touch of G27: signal is true;
	signal G28: std_logic; attribute dont_touch of G28: signal is true;
	signal G29: std_logic; attribute dont_touch of G29: signal is true;
	signal G30: std_logic; attribute dont_touch of G30: signal is true;
	signal G31: std_logic; attribute dont_touch of G31: signal is true;
	signal G32: std_logic; attribute dont_touch of G32: signal is true;
	signal G33: std_logic; attribute dont_touch of G33: signal is true;
	signal G34: std_logic; attribute dont_touch of G34: signal is true;
	signal G35: std_logic; attribute dont_touch of G35: signal is true;
	signal G36: std_logic; attribute dont_touch of G36: signal is true;
	signal G37: std_logic; attribute dont_touch of G37: signal is true;
	signal G38: std_logic; attribute dont_touch of G38: signal is true;
	signal G39: std_logic; attribute dont_touch of G39: signal is true;
	signal G40: std_logic; attribute dont_touch of G40: signal is true;
	signal G41: std_logic; attribute dont_touch of G41: signal is true;
	signal G42: std_logic; attribute dont_touch of G42: signal is true;
	signal G43: std_logic; attribute dont_touch of G43: signal is true;
	signal G44: std_logic; attribute dont_touch of G44: signal is true;
	signal G45: std_logic; attribute dont_touch of G45: signal is true;
	signal G46: std_logic; attribute dont_touch of G46: signal is true;
	signal G47: std_logic; attribute dont_touch of G47: signal is true;
	signal G48: std_logic; attribute dont_touch of G48: signal is true;
	signal G49: std_logic; attribute dont_touch of G49: signal is true;
	signal G50: std_logic; attribute dont_touch of G50: signal is true;
	signal G51: std_logic; attribute dont_touch of G51: signal is true;
	signal G52: std_logic; attribute dont_touch of G52: signal is true;
	signal G53: std_logic; attribute dont_touch of G53: signal is true;
	signal G54: std_logic; attribute dont_touch of G54: signal is true;
	signal G55: std_logic; attribute dont_touch of G55: signal is true;
	signal G56: std_logic; attribute dont_touch of G56: signal is true;
	signal G57: std_logic; attribute dont_touch of G57: signal is true;
	signal G58: std_logic; attribute dont_touch of G58: signal is true;
	signal G59: std_logic; attribute dont_touch of G59: signal is true;
	signal G60: std_logic; attribute dont_touch of G60: signal is true;
	signal G61: std_logic; attribute dont_touch of G61: signal is true;
	signal G62: std_logic; attribute dont_touch of G62: signal is true;
	signal G63: std_logic; attribute dont_touch of G63: signal is true;
	signal G64: std_logic; attribute dont_touch of G64: signal is true;
	signal G65: std_logic; attribute dont_touch of G65: signal is true;
	signal G66: std_logic; attribute dont_touch of G66: signal is true;
	signal G67: std_logic; attribute dont_touch of G67: signal is true;
	signal G68: std_logic; attribute dont_touch of G68: signal is true;
	signal G69: std_logic; attribute dont_touch of G69: signal is true;
	signal G70: std_logic; attribute dont_touch of G70: signal is true;
	signal G71: std_logic; attribute dont_touch of G71: signal is true;
	signal G72: std_logic; attribute dont_touch of G72: signal is true;
	signal G73: std_logic; attribute dont_touch of G73: signal is true;
	signal G74: std_logic; attribute dont_touch of G74: signal is true;
	signal G75: std_logic; attribute dont_touch of G75: signal is true;
	signal G76: std_logic; attribute dont_touch of G76: signal is true;
	signal G77: std_logic; attribute dont_touch of G77: signal is true;
	signal G78: std_logic; attribute dont_touch of G78: signal is true;
	signal G79: std_logic; attribute dont_touch of G79: signal is true;
	signal G80: std_logic; attribute dont_touch of G80: signal is true;
	signal G81: std_logic; attribute dont_touch of G81: signal is true;
	signal G82: std_logic; attribute dont_touch of G82: signal is true;
	signal G83: std_logic; attribute dont_touch of G83: signal is true;
	signal G84: std_logic; attribute dont_touch of G84: signal is true;
	signal G85: std_logic; attribute dont_touch of G85: signal is true;
	signal G86: std_logic; attribute dont_touch of G86: signal is true;
	signal G87: std_logic; attribute dont_touch of G87: signal is true;
	signal G88: std_logic; attribute dont_touch of G88: signal is true;
	signal G89: std_logic; attribute dont_touch of G89: signal is true;
	signal G90: std_logic; attribute dont_touch of G90: signal is true;
	signal G91: std_logic; attribute dont_touch of G91: signal is true;
	signal G92: std_logic; attribute dont_touch of G92: signal is true;
	signal G93: std_logic; attribute dont_touch of G93: signal is true;
	signal G94: std_logic; attribute dont_touch of G94: signal is true;
	signal G95: std_logic; attribute dont_touch of G95: signal is true;
	signal G96: std_logic; attribute dont_touch of G96: signal is true;
	signal G97: std_logic; attribute dont_touch of G97: signal is true;
	signal G98: std_logic; attribute dont_touch of G98: signal is true;
	signal G99: std_logic; attribute dont_touch of G99: signal is true;
	signal G100: std_logic; attribute dont_touch of G100: signal is true;
	signal G101: std_logic; attribute dont_touch of G101: signal is true;
	signal G102: std_logic; attribute dont_touch of G102: signal is true;
	signal G103: std_logic; attribute dont_touch of G103: signal is true;
	signal G104: std_logic; attribute dont_touch of G104: signal is true;
	signal G105: std_logic; attribute dont_touch of G105: signal is true;
	signal G106: std_logic; attribute dont_touch of G106: signal is true;
	signal G107: std_logic; attribute dont_touch of G107: signal is true;
	signal G108: std_logic; attribute dont_touch of G108: signal is true;
	signal G109: std_logic; attribute dont_touch of G109: signal is true;
	signal G110: std_logic; attribute dont_touch of G110: signal is true;
	signal G111: std_logic; attribute dont_touch of G111: signal is true;
	signal G112: std_logic; attribute dont_touch of G112: signal is true;
	signal G113: std_logic; attribute dont_touch of G113: signal is true;
	signal G114: std_logic; attribute dont_touch of G114: signal is true;
	signal G115: std_logic; attribute dont_touch of G115: signal is true;
	signal G116: std_logic; attribute dont_touch of G116: signal is true;
	signal G117: std_logic; attribute dont_touch of G117: signal is true;
	signal G118: std_logic; attribute dont_touch of G118: signal is true;
	signal G119: std_logic; attribute dont_touch of G119: signal is true;
	signal G120: std_logic; attribute dont_touch of G120: signal is true;
	signal G121: std_logic; attribute dont_touch of G121: signal is true;
	signal G122: std_logic; attribute dont_touch of G122: signal is true;
	signal G123: std_logic; attribute dont_touch of G123: signal is true;
	signal G124: std_logic; attribute dont_touch of G124: signal is true;
	signal G125: std_logic; attribute dont_touch of G125: signal is true;
	signal G126: std_logic; attribute dont_touch of G126: signal is true;
	signal G127: std_logic; attribute dont_touch of G127: signal is true;
	signal G128: std_logic; attribute dont_touch of G128: signal is true;
	signal G129: std_logic; attribute dont_touch of G129: signal is true;
	signal G130: std_logic; attribute dont_touch of G130: signal is true;
	signal G131: std_logic; attribute dont_touch of G131: signal is true;
	signal G132: std_logic; attribute dont_touch of G132: signal is true;
	signal G133: std_logic; attribute dont_touch of G133: signal is true;
	signal G134: std_logic; attribute dont_touch of G134: signal is true;
	signal G135: std_logic; attribute dont_touch of G135: signal is true;
	signal G136: std_logic; attribute dont_touch of G136: signal is true;
	signal G137: std_logic; attribute dont_touch of G137: signal is true;
	signal G138: std_logic; attribute dont_touch of G138: signal is true;
	signal G139: std_logic; attribute dont_touch of G139: signal is true;
	signal G140: std_logic; attribute dont_touch of G140: signal is true;
	signal G141: std_logic; attribute dont_touch of G141: signal is true;
	signal G142: std_logic; attribute dont_touch of G142: signal is true;
	signal G143: std_logic; attribute dont_touch of G143: signal is true;
	signal G144: std_logic; attribute dont_touch of G144: signal is true;
	signal G145: std_logic; attribute dont_touch of G145: signal is true;
	signal G146: std_logic; attribute dont_touch of G146: signal is true;
	signal G147: std_logic; attribute dont_touch of G147: signal is true;
	signal G148: std_logic; attribute dont_touch of G148: signal is true;
	signal G149: std_logic; attribute dont_touch of G149: signal is true;
	signal G150: std_logic; attribute dont_touch of G150: signal is true;
	signal G151: std_logic; attribute dont_touch of G151: signal is true;
	signal G152: std_logic; attribute dont_touch of G152: signal is true;
	signal G153: std_logic; attribute dont_touch of G153: signal is true;
	signal G154: std_logic; attribute dont_touch of G154: signal is true;
	signal G155: std_logic; attribute dont_touch of G155: signal is true;
	signal G156: std_logic; attribute dont_touch of G156: signal is true;
	signal G157: std_logic; attribute dont_touch of G157: signal is true;
	signal G158: std_logic; attribute dont_touch of G158: signal is true;
	signal G159: std_logic; attribute dont_touch of G159: signal is true;
	signal G160: std_logic; attribute dont_touch of G160: signal is true;
	signal G161: std_logic; attribute dont_touch of G161: signal is true;
	signal G162: std_logic; attribute dont_touch of G162: signal is true;
	signal G163: std_logic; attribute dont_touch of G163: signal is true;
	signal G164: std_logic; attribute dont_touch of G164: signal is true;
	signal G165: std_logic; attribute dont_touch of G165: signal is true;
	signal G166: std_logic; attribute dont_touch of G166: signal is true;
	signal G167: std_logic; attribute dont_touch of G167: signal is true;
	signal G168: std_logic; attribute dont_touch of G168: signal is true;
	signal G169: std_logic; attribute dont_touch of G169: signal is true;
	signal G170: std_logic; attribute dont_touch of G170: signal is true;
	signal G171: std_logic; attribute dont_touch of G171: signal is true;
	signal G172: std_logic; attribute dont_touch of G172: signal is true;
	signal G173: std_logic; attribute dont_touch of G173: signal is true;
	signal G174: std_logic; attribute dont_touch of G174: signal is true;
	signal G175: std_logic; attribute dont_touch of G175: signal is true;
	signal G176: std_logic; attribute dont_touch of G176: signal is true;
	signal G177: std_logic; attribute dont_touch of G177: signal is true;
	signal G178: std_logic; attribute dont_touch of G178: signal is true;
	signal G179: std_logic; attribute dont_touch of G179: signal is true;
	signal G180: std_logic; attribute dont_touch of G180: signal is true;
	signal G181: std_logic; attribute dont_touch of G181: signal is true;
	signal G182: std_logic; attribute dont_touch of G182: signal is true;
	signal G183: std_logic; attribute dont_touch of G183: signal is true;
	signal G184: std_logic; attribute dont_touch of G184: signal is true;
	signal G185: std_logic; attribute dont_touch of G185: signal is true;
	signal G186: std_logic; attribute dont_touch of G186: signal is true;
	signal G187: std_logic; attribute dont_touch of G187: signal is true;
	signal G188: std_logic; attribute dont_touch of G188: signal is true;
	signal G189: std_logic; attribute dont_touch of G189: signal is true;
	signal G190: std_logic; attribute dont_touch of G190: signal is true;
	signal G191: std_logic; attribute dont_touch of G191: signal is true;
	signal G192: std_logic; attribute dont_touch of G192: signal is true;
	signal G193: std_logic; attribute dont_touch of G193: signal is true;
	signal G194: std_logic; attribute dont_touch of G194: signal is true;
	signal G195: std_logic; attribute dont_touch of G195: signal is true;
	signal G196: std_logic; attribute dont_touch of G196: signal is true;
	signal G197: std_logic; attribute dont_touch of G197: signal is true;
	signal G198: std_logic; attribute dont_touch of G198: signal is true;
	signal G199: std_logic; attribute dont_touch of G199: signal is true;
	signal G200: std_logic; attribute dont_touch of G200: signal is true;
	signal G201: std_logic; attribute dont_touch of G201: signal is true;
	signal G202: std_logic; attribute dont_touch of G202: signal is true;
	signal G203: std_logic; attribute dont_touch of G203: signal is true;
	signal G204: std_logic; attribute dont_touch of G204: signal is true;
	signal G205: std_logic; attribute dont_touch of G205: signal is true;
	signal G206: std_logic; attribute dont_touch of G206: signal is true;
	signal G207: std_logic; attribute dont_touch of G207: signal is true;
	signal G208: std_logic; attribute dont_touch of G208: signal is true;
	signal G209: std_logic; attribute dont_touch of G209: signal is true;
	signal G210: std_logic; attribute dont_touch of G210: signal is true;
	signal G211: std_logic; attribute dont_touch of G211: signal is true;
	signal G212: std_logic; attribute dont_touch of G212: signal is true;
	signal G213: std_logic; attribute dont_touch of G213: signal is true;
	signal G214: std_logic; attribute dont_touch of G214: signal is true;
	signal G215: std_logic; attribute dont_touch of G215: signal is true;
	signal G216: std_logic; attribute dont_touch of G216: signal is true;
	signal G217: std_logic; attribute dont_touch of G217: signal is true;
	signal G218: std_logic; attribute dont_touch of G218: signal is true;
	signal G219: std_logic; attribute dont_touch of G219: signal is true;
	signal G220: std_logic; attribute dont_touch of G220: signal is true;
	signal G221: std_logic; attribute dont_touch of G221: signal is true;
	signal G222: std_logic; attribute dont_touch of G222: signal is true;
	signal G223: std_logic; attribute dont_touch of G223: signal is true;
	signal G224: std_logic; attribute dont_touch of G224: signal is true;
	signal G225: std_logic; attribute dont_touch of G225: signal is true;
	signal G226: std_logic; attribute dont_touch of G226: signal is true;
	signal G227: std_logic; attribute dont_touch of G227: signal is true;
	signal G228: std_logic; attribute dont_touch of G228: signal is true;
	signal G229: std_logic; attribute dont_touch of G229: signal is true;
	signal G230: std_logic; attribute dont_touch of G230: signal is true;
	signal G231: std_logic; attribute dont_touch of G231: signal is true;
	signal G232: std_logic; attribute dont_touch of G232: signal is true;
	signal G233: std_logic; attribute dont_touch of G233: signal is true;
	signal G234: std_logic; attribute dont_touch of G234: signal is true;
	signal G235: std_logic; attribute dont_touch of G235: signal is true;
	signal G236: std_logic; attribute dont_touch of G236: signal is true;
	signal G237: std_logic; attribute dont_touch of G237: signal is true;
	signal G238: std_logic; attribute dont_touch of G238: signal is true;
	signal G239: std_logic; attribute dont_touch of G239: signal is true;
	signal G240: std_logic; attribute dont_touch of G240: signal is true;
	signal G241: std_logic; attribute dont_touch of G241: signal is true;
	signal G242: std_logic; attribute dont_touch of G242: signal is true;
	signal G243: std_logic; attribute dont_touch of G243: signal is true;
	signal G244: std_logic; attribute dont_touch of G244: signal is true;
	signal G245: std_logic; attribute dont_touch of G245: signal is true;
	signal G246: std_logic; attribute dont_touch of G246: signal is true;
	signal G247: std_logic; attribute dont_touch of G247: signal is true;
	signal G248: std_logic; attribute dont_touch of G248: signal is true;
	signal G249: std_logic; attribute dont_touch of G249: signal is true;
	signal G250: std_logic; attribute dont_touch of G250: signal is true;
	signal G251: std_logic; attribute dont_touch of G251: signal is true;
	signal G252: std_logic; attribute dont_touch of G252: signal is true;
	signal G253: std_logic; attribute dont_touch of G253: signal is true;
	signal G254: std_logic; attribute dont_touch of G254: signal is true;
	signal G255: std_logic; attribute dont_touch of G255: signal is true;
	signal G256: std_logic; attribute dont_touch of G256: signal is true;
	signal G257: std_logic; attribute dont_touch of G257: signal is true;
	signal G258: std_logic; attribute dont_touch of G258: signal is true;
	signal G259: std_logic; attribute dont_touch of G259: signal is true;
	signal G260: std_logic; attribute dont_touch of G260: signal is true;
	signal G261: std_logic; attribute dont_touch of G261: signal is true;
	signal G262: std_logic; attribute dont_touch of G262: signal is true;
	signal G263: std_logic; attribute dont_touch of G263: signal is true;
	signal G264: std_logic; attribute dont_touch of G264: signal is true;
	signal G265: std_logic; attribute dont_touch of G265: signal is true;
	signal G266: std_logic; attribute dont_touch of G266: signal is true;
	signal G267: std_logic; attribute dont_touch of G267: signal is true;
	signal G268: std_logic; attribute dont_touch of G268: signal is true;
	signal G269: std_logic; attribute dont_touch of G269: signal is true;
	signal G270: std_logic; attribute dont_touch of G270: signal is true;
	signal G271: std_logic; attribute dont_touch of G271: signal is true;
	signal G272: std_logic; attribute dont_touch of G272: signal is true;
	signal G273: std_logic; attribute dont_touch of G273: signal is true;
	signal G274: std_logic; attribute dont_touch of G274: signal is true;
	signal G275: std_logic; attribute dont_touch of G275: signal is true;
	signal G276: std_logic; attribute dont_touch of G276: signal is true;
	signal G277: std_logic; attribute dont_touch of G277: signal is true;
	signal G278: std_logic; attribute dont_touch of G278: signal is true;
	signal G279: std_logic; attribute dont_touch of G279: signal is true;
	signal G280: std_logic; attribute dont_touch of G280: signal is true;
	signal G281: std_logic; attribute dont_touch of G281: signal is true;
	signal G282: std_logic; attribute dont_touch of G282: signal is true;
	signal G283: std_logic; attribute dont_touch of G283: signal is true;
	signal G284: std_logic; attribute dont_touch of G284: signal is true;
	signal G285: std_logic; attribute dont_touch of G285: signal is true;
	signal G286: std_logic; attribute dont_touch of G286: signal is true;
	signal G287: std_logic; attribute dont_touch of G287: signal is true;
	signal G288: std_logic; attribute dont_touch of G288: signal is true;
	signal G289: std_logic; attribute dont_touch of G289: signal is true;
	signal G290: std_logic; attribute dont_touch of G290: signal is true;
	signal G291: std_logic; attribute dont_touch of G291: signal is true;
	signal G292: std_logic; attribute dont_touch of G292: signal is true;
	signal G293: std_logic; attribute dont_touch of G293: signal is true;
	signal G294: std_logic; attribute dont_touch of G294: signal is true;
	signal G295: std_logic; attribute dont_touch of G295: signal is true;
	signal G296: std_logic; attribute dont_touch of G296: signal is true;
	signal G297: std_logic; attribute dont_touch of G297: signal is true;
	signal G298: std_logic; attribute dont_touch of G298: signal is true;
	signal G299: std_logic; attribute dont_touch of G299: signal is true;
	signal G300: std_logic; attribute dont_touch of G300: signal is true;
	signal G301: std_logic; attribute dont_touch of G301: signal is true;
	signal G302: std_logic; attribute dont_touch of G302: signal is true;
	signal G303: std_logic; attribute dont_touch of G303: signal is true;
	signal G304: std_logic; attribute dont_touch of G304: signal is true;
	signal G305: std_logic; attribute dont_touch of G305: signal is true;
	signal G306: std_logic; attribute dont_touch of G306: signal is true;
	signal G307: std_logic; attribute dont_touch of G307: signal is true;
	signal G308: std_logic; attribute dont_touch of G308: signal is true;
	signal G309: std_logic; attribute dont_touch of G309: signal is true;
	signal G310: std_logic; attribute dont_touch of G310: signal is true;
	signal G311: std_logic; attribute dont_touch of G311: signal is true;
	signal G312: std_logic; attribute dont_touch of G312: signal is true;
	signal G313: std_logic; attribute dont_touch of G313: signal is true;
	signal G314: std_logic; attribute dont_touch of G314: signal is true;
	signal G315: std_logic; attribute dont_touch of G315: signal is true;
	signal G316: std_logic; attribute dont_touch of G316: signal is true;
	signal G317: std_logic; attribute dont_touch of G317: signal is true;
	signal G318: std_logic; attribute dont_touch of G318: signal is true;
	signal G319: std_logic; attribute dont_touch of G319: signal is true;
	signal G320: std_logic; attribute dont_touch of G320: signal is true;
	signal G321: std_logic; attribute dont_touch of G321: signal is true;
	signal G322: std_logic; attribute dont_touch of G322: signal is true;
	signal G323: std_logic; attribute dont_touch of G323: signal is true;
	signal G324: std_logic; attribute dont_touch of G324: signal is true;
	signal G325: std_logic; attribute dont_touch of G325: signal is true;
	signal G326: std_logic; attribute dont_touch of G326: signal is true;
	signal G327: std_logic; attribute dont_touch of G327: signal is true;
	signal G328: std_logic; attribute dont_touch of G328: signal is true;
	signal G328BF: std_logic; attribute dont_touch of G328BF: signal is true;
	signal G329: std_logic; attribute dont_touch of G329: signal is true;
	signal G330: std_logic; attribute dont_touch of G330: signal is true;
	signal G331: std_logic; attribute dont_touch of G331: signal is true;
	signal G332: std_logic; attribute dont_touch of G332: signal is true;
	signal G332BF: std_logic; attribute dont_touch of G332BF: signal is true;
	signal G333: std_logic; attribute dont_touch of G333: signal is true;
	signal G334: std_logic; attribute dont_touch of G334: signal is true;
	signal G335: std_logic; attribute dont_touch of G335: signal is true;
	signal G336: std_logic; attribute dont_touch of G336: signal is true;
	signal G337: std_logic; attribute dont_touch of G337: signal is true;
	signal G338: std_logic; attribute dont_touch of G338: signal is true;
	signal G339: std_logic; attribute dont_touch of G339: signal is true;
	signal G340: std_logic; attribute dont_touch of G340: signal is true;
	signal G341: std_logic; attribute dont_touch of G341: signal is true;
	signal G342: std_logic; attribute dont_touch of G342: signal is true;
	signal G343: std_logic; attribute dont_touch of G343: signal is true;
	signal G344: std_logic; attribute dont_touch of G344: signal is true;
	signal G345: std_logic; attribute dont_touch of G345: signal is true;
	signal G346: std_logic; attribute dont_touch of G346: signal is true;
	signal G347: std_logic; attribute dont_touch of G347: signal is true;
	signal G348: std_logic; attribute dont_touch of G348: signal is true;
	signal G349: std_logic; attribute dont_touch of G349: signal is true;
	signal G350: std_logic; attribute dont_touch of G350: signal is true;
	signal G351: std_logic; attribute dont_touch of G351: signal is true;
	signal G352: std_logic; attribute dont_touch of G352: signal is true;
	signal G353: std_logic; attribute dont_touch of G353: signal is true;
	signal G354: std_logic; attribute dont_touch of G354: signal is true;
	signal G355: std_logic; attribute dont_touch of G355: signal is true;
	signal G356: std_logic; attribute dont_touch of G356: signal is true;
	signal G357: std_logic; attribute dont_touch of G357: signal is true;
	signal G358: std_logic; attribute dont_touch of G358: signal is true;
	signal G359: std_logic; attribute dont_touch of G359: signal is true;
	signal G360: std_logic; attribute dont_touch of G360: signal is true;
	signal G361: std_logic; attribute dont_touch of G361: signal is true;
	signal G362: std_logic; attribute dont_touch of G362: signal is true;
	signal G363: std_logic; attribute dont_touch of G363: signal is true;
	signal G364: std_logic; attribute dont_touch of G364: signal is true;
	signal G365: std_logic; attribute dont_touch of G365: signal is true;
	signal G366: std_logic; attribute dont_touch of G366: signal is true;
	signal G367: std_logic; attribute dont_touch of G367: signal is true;
	signal G368: std_logic; attribute dont_touch of G368: signal is true;
	signal G369: std_logic; attribute dont_touch of G369: signal is true;
	signal G370: std_logic; attribute dont_touch of G370: signal is true;
	signal G371: std_logic; attribute dont_touch of G371: signal is true;
	signal G372: std_logic; attribute dont_touch of G372: signal is true;
	signal G373: std_logic; attribute dont_touch of G373: signal is true;
	signal G374: std_logic; attribute dont_touch of G374: signal is true;
	signal G375: std_logic; attribute dont_touch of G375: signal is true;
	signal G376: std_logic; attribute dont_touch of G376: signal is true;
	signal G377: std_logic; attribute dont_touch of G377: signal is true;
	signal G378: std_logic; attribute dont_touch of G378: signal is true;
	signal G379: std_logic; attribute dont_touch of G379: signal is true;
	signal G380: std_logic; attribute dont_touch of G380: signal is true;
	signal G381: std_logic; attribute dont_touch of G381: signal is true;
	signal G382: std_logic; attribute dont_touch of G382: signal is true;
	signal G383: std_logic; attribute dont_touch of G383: signal is true;
	signal G384: std_logic; attribute dont_touch of G384: signal is true;
	signal G385: std_logic; attribute dont_touch of G385: signal is true;
	signal G386: std_logic; attribute dont_touch of G386: signal is true;
	signal G387: std_logic; attribute dont_touch of G387: signal is true;
	signal G388: std_logic; attribute dont_touch of G388: signal is true;
	signal G389: std_logic; attribute dont_touch of G389: signal is true;
	signal G390: std_logic; attribute dont_touch of G390: signal is true;
	signal G391: std_logic; attribute dont_touch of G391: signal is true;
	signal G392: std_logic; attribute dont_touch of G392: signal is true;
	signal G393: std_logic; attribute dont_touch of G393: signal is true;
	signal G394: std_logic; attribute dont_touch of G394: signal is true;
	signal G395: std_logic; attribute dont_touch of G395: signal is true;
	signal G396: std_logic; attribute dont_touch of G396: signal is true;
	signal G397: std_logic; attribute dont_touch of G397: signal is true;
	signal G398: std_logic; attribute dont_touch of G398: signal is true;
	signal G399: std_logic; attribute dont_touch of G399: signal is true;
	signal G400: std_logic; attribute dont_touch of G400: signal is true;
	signal G401: std_logic; attribute dont_touch of G401: signal is true;
	signal G402: std_logic; attribute dont_touch of G402: signal is true;
	signal G403: std_logic; attribute dont_touch of G403: signal is true;
	signal G404: std_logic; attribute dont_touch of G404: signal is true;
	signal G405: std_logic; attribute dont_touch of G405: signal is true;
	signal G406: std_logic; attribute dont_touch of G406: signal is true;
	signal G407: std_logic; attribute dont_touch of G407: signal is true;
	signal G408: std_logic; attribute dont_touch of G408: signal is true;
	signal G409: std_logic; attribute dont_touch of G409: signal is true;
	signal G410: std_logic; attribute dont_touch of G410: signal is true;
	signal G411: std_logic; attribute dont_touch of G411: signal is true;
	signal G412: std_logic; attribute dont_touch of G412: signal is true;
	signal G413: std_logic; attribute dont_touch of G413: signal is true;
	signal G414: std_logic; attribute dont_touch of G414: signal is true;
	signal G415: std_logic; attribute dont_touch of G415: signal is true;
	signal G416: std_logic; attribute dont_touch of G416: signal is true;
	signal G417: std_logic; attribute dont_touch of G417: signal is true;
	signal G418: std_logic; attribute dont_touch of G418: signal is true;
	signal G419: std_logic; attribute dont_touch of G419: signal is true;
	signal G420: std_logic; attribute dont_touch of G420: signal is true;
	signal G421: std_logic; attribute dont_touch of G421: signal is true;
	signal G422: std_logic; attribute dont_touch of G422: signal is true;
	signal G423: std_logic; attribute dont_touch of G423: signal is true;
	signal G424: std_logic; attribute dont_touch of G424: signal is true;
	signal G425: std_logic; attribute dont_touch of G425: signal is true;
	signal G426: std_logic; attribute dont_touch of G426: signal is true;
	signal G427: std_logic; attribute dont_touch of G427: signal is true;
	signal G428: std_logic; attribute dont_touch of G428: signal is true;
	signal G429: std_logic; attribute dont_touch of G429: signal is true;
	signal G430: std_logic; attribute dont_touch of G430: signal is true;
	signal G431: std_logic; attribute dont_touch of G431: signal is true;
	signal G432: std_logic; attribute dont_touch of G432: signal is true;
	signal G433: std_logic; attribute dont_touch of G433: signal is true;
	signal G434: std_logic; attribute dont_touch of G434: signal is true;
	signal G435: std_logic; attribute dont_touch of G435: signal is true;
	signal G436: std_logic; attribute dont_touch of G436: signal is true;
	signal G437: std_logic; attribute dont_touch of G437: signal is true;
	signal G438: std_logic; attribute dont_touch of G438: signal is true;
	signal G439: std_logic; attribute dont_touch of G439: signal is true;
	signal G440: std_logic; attribute dont_touch of G440: signal is true;
	signal G441: std_logic; attribute dont_touch of G441: signal is true;
	signal G442: std_logic; attribute dont_touch of G442: signal is true;
	signal G443: std_logic; attribute dont_touch of G443: signal is true;
	signal G444: std_logic; attribute dont_touch of G444: signal is true;
	signal G445: std_logic; attribute dont_touch of G445: signal is true;
	signal G446: std_logic; attribute dont_touch of G446: signal is true;
	signal G447: std_logic; attribute dont_touch of G447: signal is true;
	signal G448: std_logic; attribute dont_touch of G448: signal is true;
	signal G449: std_logic; attribute dont_touch of G449: signal is true;
	signal G450: std_logic; attribute dont_touch of G450: signal is true;
	signal G451: std_logic; attribute dont_touch of G451: signal is true;
	signal G452: std_logic; attribute dont_touch of G452: signal is true;
	signal G453: std_logic; attribute dont_touch of G453: signal is true;
	signal G454: std_logic; attribute dont_touch of G454: signal is true;
	signal G455: std_logic; attribute dont_touch of G455: signal is true;
	signal G456: std_logic; attribute dont_touch of G456: signal is true;
	signal G457: std_logic; attribute dont_touch of G457: signal is true;
	signal G458: std_logic; attribute dont_touch of G458: signal is true;
	signal G459: std_logic; attribute dont_touch of G459: signal is true;
	signal G460: std_logic; attribute dont_touch of G460: signal is true;
	signal G461: std_logic; attribute dont_touch of G461: signal is true;
	signal G462: std_logic; attribute dont_touch of G462: signal is true;
	signal G463: std_logic; attribute dont_touch of G463: signal is true;
	signal G464: std_logic; attribute dont_touch of G464: signal is true;
	signal G465: std_logic; attribute dont_touch of G465: signal is true;
	signal G466: std_logic; attribute dont_touch of G466: signal is true;
	signal G467: std_logic; attribute dont_touch of G467: signal is true;
	signal G468: std_logic; attribute dont_touch of G468: signal is true;
	signal G469: std_logic; attribute dont_touch of G469: signal is true;
	signal G470: std_logic; attribute dont_touch of G470: signal is true;
	signal G471: std_logic; attribute dont_touch of G471: signal is true;
	signal G472: std_logic; attribute dont_touch of G472: signal is true;
	signal G473: std_logic; attribute dont_touch of G473: signal is true;
	signal G474: std_logic; attribute dont_touch of G474: signal is true;
	signal G475: std_logic; attribute dont_touch of G475: signal is true;
	signal G476: std_logic; attribute dont_touch of G476: signal is true;
	signal G477: std_logic; attribute dont_touch of G477: signal is true;
	signal G478: std_logic; attribute dont_touch of G478: signal is true;
	signal G479: std_logic; attribute dont_touch of G479: signal is true;
	signal G480: std_logic; attribute dont_touch of G480: signal is true;
	signal G481: std_logic; attribute dont_touch of G481: signal is true;
	signal G482: std_logic; attribute dont_touch of G482: signal is true;
	signal G483: std_logic; attribute dont_touch of G483: signal is true;
	signal G484: std_logic; attribute dont_touch of G484: signal is true;
	signal G485: std_logic; attribute dont_touch of G485: signal is true;
	signal G486: std_logic; attribute dont_touch of G486: signal is true;
	signal G487: std_logic; attribute dont_touch of G487: signal is true;
	signal G488: std_logic; attribute dont_touch of G488: signal is true;
	signal G489: std_logic; attribute dont_touch of G489: signal is true;
	signal G490: std_logic; attribute dont_touch of G490: signal is true;
	signal G491: std_logic; attribute dont_touch of G491: signal is true;
	signal G492: std_logic; attribute dont_touch of G492: signal is true;
	signal G493: std_logic; attribute dont_touch of G493: signal is true;
	signal G494: std_logic; attribute dont_touch of G494: signal is true;
	signal G495: std_logic; attribute dont_touch of G495: signal is true;
	signal G496: std_logic; attribute dont_touch of G496: signal is true;
	signal G497: std_logic; attribute dont_touch of G497: signal is true;
	signal G498: std_logic; attribute dont_touch of G498: signal is true;
	signal G499: std_logic; attribute dont_touch of G499: signal is true;
	signal G500: std_logic; attribute dont_touch of G500: signal is true;
	signal G501: std_logic; attribute dont_touch of G501: signal is true;
	signal G502: std_logic; attribute dont_touch of G502: signal is true;
	signal G503: std_logic; attribute dont_touch of G503: signal is true;
	signal G504: std_logic; attribute dont_touch of G504: signal is true;
	signal G505: std_logic; attribute dont_touch of G505: signal is true;
	signal G506: std_logic; attribute dont_touch of G506: signal is true;
	signal G507: std_logic; attribute dont_touch of G507: signal is true;
	signal G508: std_logic; attribute dont_touch of G508: signal is true;
	signal G509: std_logic; attribute dont_touch of G509: signal is true;
	signal G510: std_logic; attribute dont_touch of G510: signal is true;
	signal G511: std_logic; attribute dont_touch of G511: signal is true;
	signal G512: std_logic; attribute dont_touch of G512: signal is true;
	signal G513: std_logic; attribute dont_touch of G513: signal is true;
	signal G514: std_logic; attribute dont_touch of G514: signal is true;
	signal G515: std_logic; attribute dont_touch of G515: signal is true;
	signal G516: std_logic; attribute dont_touch of G516: signal is true;
	signal G517: std_logic; attribute dont_touch of G517: signal is true;
	signal G518: std_logic; attribute dont_touch of G518: signal is true;
	signal G519: std_logic; attribute dont_touch of G519: signal is true;
	signal G520: std_logic; attribute dont_touch of G520: signal is true;
	signal G521: std_logic; attribute dont_touch of G521: signal is true;
	signal G522: std_logic; attribute dont_touch of G522: signal is true;
	signal G523: std_logic; attribute dont_touch of G523: signal is true;
	signal G524: std_logic; attribute dont_touch of G524: signal is true;
	signal G525: std_logic; attribute dont_touch of G525: signal is true;
	signal G526: std_logic; attribute dont_touch of G526: signal is true;
	signal G527: std_logic; attribute dont_touch of G527: signal is true;
	signal G528: std_logic; attribute dont_touch of G528: signal is true;
	signal G529: std_logic; attribute dont_touch of G529: signal is true;
	signal G530: std_logic; attribute dont_touch of G530: signal is true;
	signal G531: std_logic; attribute dont_touch of G531: signal is true;
	signal G532: std_logic; attribute dont_touch of G532: signal is true;
	signal G533: std_logic; attribute dont_touch of G533: signal is true;
	signal G534: std_logic; attribute dont_touch of G534: signal is true;
	signal G535: std_logic; attribute dont_touch of G535: signal is true;
	signal G536: std_logic; attribute dont_touch of G536: signal is true;
	signal G537: std_logic; attribute dont_touch of G537: signal is true;
	signal G538: std_logic; attribute dont_touch of G538: signal is true;
	signal G539: std_logic; attribute dont_touch of G539: signal is true;
	signal G540: std_logic; attribute dont_touch of G540: signal is true;
	signal G541: std_logic; attribute dont_touch of G541: signal is true;
	signal G542: std_logic; attribute dont_touch of G542: signal is true;
	signal G543: std_logic; attribute dont_touch of G543: signal is true;
	signal G544: std_logic; attribute dont_touch of G544: signal is true;
	signal G545: std_logic; attribute dont_touch of G545: signal is true;
	signal G546: std_logic; attribute dont_touch of G546: signal is true;
	signal G547: std_logic; attribute dont_touch of G547: signal is true;
	signal G548: std_logic; attribute dont_touch of G548: signal is true;
	signal G549: std_logic; attribute dont_touch of G549: signal is true;
	signal G550: std_logic; attribute dont_touch of G550: signal is true;
	signal G551: std_logic; attribute dont_touch of G551: signal is true;
	signal G552: std_logic; attribute dont_touch of G552: signal is true;
	signal G553: std_logic; attribute dont_touch of G553: signal is true;
	signal G554: std_logic; attribute dont_touch of G554: signal is true;
	signal G555: std_logic; attribute dont_touch of G555: signal is true;
	signal G556: std_logic; attribute dont_touch of G556: signal is true;
	signal G557: std_logic; attribute dont_touch of G557: signal is true;
	signal G558: std_logic; attribute dont_touch of G558: signal is true;
	signal G559: std_logic; attribute dont_touch of G559: signal is true;
	signal G560: std_logic; attribute dont_touch of G560: signal is true;
	signal G561: std_logic; attribute dont_touch of G561: signal is true;
	signal G562: std_logic; attribute dont_touch of G562: signal is true;
	signal G563: std_logic; attribute dont_touch of G563: signal is true;
	signal G564: std_logic; attribute dont_touch of G564: signal is true;
	signal G565: std_logic; attribute dont_touch of G565: signal is true;
	signal G566: std_logic; attribute dont_touch of G566: signal is true;
	signal G567: std_logic; attribute dont_touch of G567: signal is true;
	signal G568: std_logic; attribute dont_touch of G568: signal is true;
	signal G569: std_logic; attribute dont_touch of G569: signal is true;
	signal G570: std_logic; attribute dont_touch of G570: signal is true;
	signal G571: std_logic; attribute dont_touch of G571: signal is true;
	signal G572: std_logic; attribute dont_touch of G572: signal is true;
	signal G573: std_logic; attribute dont_touch of G573: signal is true;
	signal G574: std_logic; attribute dont_touch of G574: signal is true;
	signal G575: std_logic; attribute dont_touch of G575: signal is true;
	signal G576: std_logic; attribute dont_touch of G576: signal is true;
	signal G577: std_logic; attribute dont_touch of G577: signal is true;
	signal G578: std_logic; attribute dont_touch of G578: signal is true;
	signal G579: std_logic; attribute dont_touch of G579: signal is true;
	signal G580: std_logic; attribute dont_touch of G580: signal is true;
	signal G581: std_logic; attribute dont_touch of G581: signal is true;
	signal G582: std_logic; attribute dont_touch of G582: signal is true;
	signal G583: std_logic; attribute dont_touch of G583: signal is true;
	signal G584: std_logic; attribute dont_touch of G584: signal is true;
	signal G585: std_logic; attribute dont_touch of G585: signal is true;
	signal G586: std_logic; attribute dont_touch of G586: signal is true;
	signal G587: std_logic; attribute dont_touch of G587: signal is true;
	signal G588: std_logic; attribute dont_touch of G588: signal is true;
	signal G589: std_logic; attribute dont_touch of G589: signal is true;
	signal G590: std_logic; attribute dont_touch of G590: signal is true;
	signal G591: std_logic; attribute dont_touch of G591: signal is true;
	signal G592: std_logic; attribute dont_touch of G592: signal is true;
	signal G593: std_logic; attribute dont_touch of G593: signal is true;
	signal G594: std_logic; attribute dont_touch of G594: signal is true;
	signal G595: std_logic; attribute dont_touch of G595: signal is true;
	signal G596: std_logic; attribute dont_touch of G596: signal is true;
	signal G597: std_logic; attribute dont_touch of G597: signal is true;
	signal G598: std_logic; attribute dont_touch of G598: signal is true;
	signal G599: std_logic; attribute dont_touch of G599: signal is true;
	signal G600: std_logic; attribute dont_touch of G600: signal is true;
	signal G601: std_logic; attribute dont_touch of G601: signal is true;
	signal G602: std_logic; attribute dont_touch of G602: signal is true;
	signal G603: std_logic; attribute dont_touch of G603: signal is true;
	signal G604: std_logic; attribute dont_touch of G604: signal is true;
	signal G605: std_logic; attribute dont_touch of G605: signal is true;
	signal G606: std_logic; attribute dont_touch of G606: signal is true;
	signal G607: std_logic; attribute dont_touch of G607: signal is true;
	signal G608: std_logic; attribute dont_touch of G608: signal is true;
	signal G609: std_logic; attribute dont_touch of G609: signal is true;
	signal G610: std_logic; attribute dont_touch of G610: signal is true;
	signal G611: std_logic; attribute dont_touch of G611: signal is true;
	signal G612: std_logic; attribute dont_touch of G612: signal is true;
	signal G613: std_logic; attribute dont_touch of G613: signal is true;
	signal G614: std_logic; attribute dont_touch of G614: signal is true;
	signal G615: std_logic; attribute dont_touch of G615: signal is true;
	signal G616: std_logic; attribute dont_touch of G616: signal is true;
	signal G617: std_logic; attribute dont_touch of G617: signal is true;
	signal G618: std_logic; attribute dont_touch of G618: signal is true;
	signal G619: std_logic; attribute dont_touch of G619: signal is true;
	signal G620: std_logic; attribute dont_touch of G620: signal is true;
	signal G621: std_logic; attribute dont_touch of G621: signal is true;
	signal G622: std_logic; attribute dont_touch of G622: signal is true;
	signal G623: std_logic; attribute dont_touch of G623: signal is true;
	signal G624: std_logic; attribute dont_touch of G624: signal is true;
	signal G625: std_logic; attribute dont_touch of G625: signal is true;
	signal G626: std_logic; attribute dont_touch of G626: signal is true;
	signal G627: std_logic; attribute dont_touch of G627: signal is true;
	signal G628: std_logic; attribute dont_touch of G628: signal is true;
	signal G629: std_logic; attribute dont_touch of G629: signal is true;
	signal G630: std_logic; attribute dont_touch of G630: signal is true;
	signal G631: std_logic; attribute dont_touch of G631: signal is true;
	signal G632: std_logic; attribute dont_touch of G632: signal is true;
	signal G633: std_logic; attribute dont_touch of G633: signal is true;
	signal G634: std_logic; attribute dont_touch of G634: signal is true;
	signal G635: std_logic; attribute dont_touch of G635: signal is true;
	signal G636: std_logic; attribute dont_touch of G636: signal is true;
	signal G637: std_logic; attribute dont_touch of G637: signal is true;
	signal G638: std_logic; attribute dont_touch of G638: signal is true;
	signal G639: std_logic; attribute dont_touch of G639: signal is true;
	signal G640: std_logic; attribute dont_touch of G640: signal is true;
	signal G641: std_logic; attribute dont_touch of G641: signal is true;
	signal G642: std_logic; attribute dont_touch of G642: signal is true;
	signal G643: std_logic; attribute dont_touch of G643: signal is true;
	signal G644: std_logic; attribute dont_touch of G644: signal is true;
	signal G645: std_logic; attribute dont_touch of G645: signal is true;
	signal G646: std_logic; attribute dont_touch of G646: signal is true;
	signal G647: std_logic; attribute dont_touch of G647: signal is true;
	signal G648: std_logic; attribute dont_touch of G648: signal is true;
	signal G649: std_logic; attribute dont_touch of G649: signal is true;
	signal G650: std_logic; attribute dont_touch of G650: signal is true;
	signal G651: std_logic; attribute dont_touch of G651: signal is true;
	signal G652: std_logic; attribute dont_touch of G652: signal is true;
	signal G653: std_logic; attribute dont_touch of G653: signal is true;
	signal G654: std_logic; attribute dont_touch of G654: signal is true;
	signal G655: std_logic; attribute dont_touch of G655: signal is true;
	signal G656: std_logic; attribute dont_touch of G656: signal is true;
	signal G657: std_logic; attribute dont_touch of G657: signal is true;
	signal G658: std_logic; attribute dont_touch of G658: signal is true;
	signal G659: std_logic; attribute dont_touch of G659: signal is true;
	signal G660: std_logic; attribute dont_touch of G660: signal is true;
	signal G661: std_logic; attribute dont_touch of G661: signal is true;
	signal G662: std_logic; attribute dont_touch of G662: signal is true;
	signal G663: std_logic; attribute dont_touch of G663: signal is true;
	signal G664: std_logic; attribute dont_touch of G664: signal is true;
	signal G665: std_logic; attribute dont_touch of G665: signal is true;
	signal G666: std_logic; attribute dont_touch of G666: signal is true;
	signal G667: std_logic; attribute dont_touch of G667: signal is true;
	signal G668: std_logic; attribute dont_touch of G668: signal is true;
	signal G669: std_logic; attribute dont_touch of G669: signal is true;
	signal G670: std_logic; attribute dont_touch of G670: signal is true;
	signal G671: std_logic; attribute dont_touch of G671: signal is true;
	signal G672: std_logic; attribute dont_touch of G672: signal is true;
	signal G673: std_logic; attribute dont_touch of G673: signal is true;
	signal G674: std_logic; attribute dont_touch of G674: signal is true;
	signal G675: std_logic; attribute dont_touch of G675: signal is true;
	signal G676: std_logic; attribute dont_touch of G676: signal is true;
	signal G677: std_logic; attribute dont_touch of G677: signal is true;
	signal G678: std_logic; attribute dont_touch of G678: signal is true;
	signal G679: std_logic; attribute dont_touch of G679: signal is true;
	signal G680: std_logic; attribute dont_touch of G680: signal is true;
	signal G681: std_logic; attribute dont_touch of G681: signal is true;
	signal G682: std_logic; attribute dont_touch of G682: signal is true;
	signal G683: std_logic; attribute dont_touch of G683: signal is true;
	signal G684: std_logic; attribute dont_touch of G684: signal is true;
	signal G685: std_logic; attribute dont_touch of G685: signal is true;
	signal G686: std_logic; attribute dont_touch of G686: signal is true;
	signal G687: std_logic; attribute dont_touch of G687: signal is true;
	signal G688: std_logic; attribute dont_touch of G688: signal is true;
	signal G689: std_logic; attribute dont_touch of G689: signal is true;
	signal G690: std_logic; attribute dont_touch of G690: signal is true;
	signal G691: std_logic; attribute dont_touch of G691: signal is true;
	signal G692: std_logic; attribute dont_touch of G692: signal is true;
	signal G693: std_logic; attribute dont_touch of G693: signal is true;
	signal G694: std_logic; attribute dont_touch of G694: signal is true;
	signal G695: std_logic; attribute dont_touch of G695: signal is true;
	signal G696: std_logic; attribute dont_touch of G696: signal is true;
	signal G697: std_logic; attribute dont_touch of G697: signal is true;
	signal G698: std_logic; attribute dont_touch of G698: signal is true;
	signal G699: std_logic; attribute dont_touch of G699: signal is true;
	signal G700: std_logic; attribute dont_touch of G700: signal is true;
	signal G701: std_logic; attribute dont_touch of G701: signal is true;
	signal G703: std_logic; attribute dont_touch of G703: signal is true;
	signal G704: std_logic; attribute dont_touch of G704: signal is true;
	signal G705: std_logic; attribute dont_touch of G705: signal is true;
	signal G706: std_logic; attribute dont_touch of G706: signal is true;
	signal G707: std_logic; attribute dont_touch of G707: signal is true;
	signal G708: std_logic; attribute dont_touch of G708: signal is true;
	signal G709: std_logic; attribute dont_touch of G709: signal is true;
	signal G710: std_logic; attribute dont_touch of G710: signal is true;
	signal G711: std_logic; attribute dont_touch of G711: signal is true;
	signal G712: std_logic; attribute dont_touch of G712: signal is true;
	signal G713: std_logic; attribute dont_touch of G713: signal is true;
	signal G714: std_logic; attribute dont_touch of G714: signal is true;
	signal G715: std_logic; attribute dont_touch of G715: signal is true;
	signal G716: std_logic; attribute dont_touch of G716: signal is true;
	signal G717: std_logic; attribute dont_touch of G717: signal is true;
	signal G718: std_logic; attribute dont_touch of G718: signal is true;
	signal G719: std_logic; attribute dont_touch of G719: signal is true;
	signal G720: std_logic; attribute dont_touch of G720: signal is true;
	signal G721: std_logic; attribute dont_touch of G721: signal is true;
	signal G722: std_logic; attribute dont_touch of G722: signal is true;
	signal G723: std_logic; attribute dont_touch of G723: signal is true;
	signal G724: std_logic; attribute dont_touch of G724: signal is true;
	signal G725: std_logic; attribute dont_touch of G725: signal is true;
	signal G728: std_logic; attribute dont_touch of G728: signal is true;
	signal I1: std_logic; attribute dont_touch of I1: signal is true;
	signal I12: std_logic; attribute dont_touch of I12: signal is true;
	signal I1162: std_logic; attribute dont_touch of I1162: signal is true;
	signal I1183: std_logic; attribute dont_touch of I1183: signal is true;
	signal I1203: std_logic; attribute dont_touch of I1203: signal is true;
	signal I1211: std_logic; attribute dont_touch of I1211: signal is true;
	signal I1227: std_logic; attribute dont_touch of I1227: signal is true;
	signal I1230: std_logic; attribute dont_touch of I1230: signal is true;
	signal I1233: std_logic; attribute dont_touch of I1233: signal is true;
	signal I1236: std_logic; attribute dont_touch of I1236: signal is true;
	signal I1239: std_logic; attribute dont_touch of I1239: signal is true;
	signal I1242: std_logic; attribute dont_touch of I1242: signal is true;
	signal I1245: std_logic; attribute dont_touch of I1245: signal is true;
	signal I1248: std_logic; attribute dont_touch of I1248: signal is true;
	signal I1251: std_logic; attribute dont_touch of I1251: signal is true;
	signal I1254: std_logic; attribute dont_touch of I1254: signal is true;
	signal I1257: std_logic; attribute dont_touch of I1257: signal is true;
	signal I1260: std_logic; attribute dont_touch of I1260: signal is true;
	signal I1264: std_logic; attribute dont_touch of I1264: signal is true;
	signal I1267: std_logic; attribute dont_touch of I1267: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			G22<=G332BF;
			G23<=G328BF;
			G24<=G109;
			G25<=G113;
			G26<=G118;
			G27<=G125;
			G28<=G129;
			G29<=G140;
			G30<=G144;
			G31<=G149;
			G32<=G154;
			G33<=G159;
			G34<=G166;
			G35<=G175;
			G36<=G189;
			G37<=G193;
			G38<=G198;
			G39<=G208;
			G40<=G214;
			G41<=G218;
			G42<=G237;
			G43<=G242;
			G44<=G247;
			G45<=G252;
			G46<=G260;
			G47<=G303;
			G48<=G309;
			G49<=G315;
			G50<=G321;
			G51<=G360;
			G52<=G365;
			G53<=G373;
			G54<=G379;
			G55<=G384;
			G56<=G392;
			G57<=G397;
			G58<=G405;
			G59<=G408;
			G60<=G416;
			G61<=G424;
			G62<=G427;
			G63<=G438;
			G64<=G441;
			G65<=G447;
			G66<=G451;
			G67<=G459;
			G68<=G464;
			G69<=G469;
			G70<=G477;
			G71<=G494;
			G72<=G498;
			G73<=G503;
			G74<=G526;
			G75<=G531;
			G76<=G536;
			G77<=G541;
			G78<=G548;
			G79<=G565;
			G80<=G569;
			G81<=G573;
			G82<=G577;
			G83<=G590;
			G84<=G608;
			G85<=G613;
			G86<=G657;
			G87<=G663;
			G88<=G669;
			G89<=G675;
			G90<=G682;
			G91<=G687;
			G92<=G693;
			G93<=G705;
			G94<=G707;
			G95<=G713;
		end if;
	end process;
	G108<= not G712;
	G111<= not G24;
	G112<= not G712;
	G117<= not G712;
	G124<= not G712;
	G127<= not G27;
	G128<= not G712;
	G139<= not G712;
	G142<= not G29;
	G143<= not G712;
	G148<= not G712;
	G153<= not G712;
	G158<= not G712;
	G165<= not G712;
	G174<= not G712;
	G176<= not G35;
	G178<= not G34;
	G179<= not G180;
	G180<= not G92;
	G188<= not G712;
	G191<= not G36;
	G192<= not G712;
	G197<= not G712;
	G204<= not G38;
	G207<= not G712;
	G210<= not G39;
	G213<= not G712;
	G216<= not G40;
	G217<= not G712;
	G236<= not G259;
	G241<= not G259;
	G246<= not G259;
	G251<= not G259;
	G258<= not G259;
	G296<= not G297;
	G302<= not G712;
	G305<= not G324;
	G308<= not G712;
	G311<= not G324;
	G314<= not G712;
	G317<= not G324;
	G320<= not G712;
	G323<= not G324;
	G328BF<= not I12;
	G332BF<= not I1;
	G336<= not G355;
	G339<= not G355;
	G343<= not G348;
	G347<= not G348;
	G348<= not G91;
	G351<= not G645;
	G354<= not G355;
	G359<= not G372;
	G364<= not G372;
	G371<= not G372;
	G378<= not G391;
	G383<= not G391;
	G390<= not G391;
	G396<= not G404;
	G403<= not G404;
	G407<= not G712;
	G415<= not G423;
	G422<= not G423;
	G426<= not G712;
	G437<= not G712;
	G440<= not G712;
	G445<= not G65;
	G446<= not G712;
	G449<= not G66;
	G450<= not G712;
	G455<= not G456;
	G458<= not G476;
	G463<= not G476;
	G468<= not G476;
	G475<= not G476;
	G486<= not G712;
	G491<= not G500;
	G495<= not G500;
	G499<= not G500;
	G504<= not G511;
	G507<= not G511;
	G510<= not G511;
	G511<= not G63;
	G525<= not G589;
	G530<= not G589;
	G535<= not G589;
	G540<= not G589;
	G547<= not G589;
	G562<= not G610;
	G566<= not G610;
	G570<= not G610;
	G574<= not G610;
	G588<= not G589;
	G595<= not G593;
	G596<= not G597;
	G600<= not G601;
	G605<= not G610;
	G609<= not G610;
	G614<= not G64;
	G615<= not G616;
	G617<= not G645;
	G620<= not G645;
	G623<= not G645;
	G626<= not G645;
	G629<= not G645;
	G632<= not G645;
	G635<= not G645;
	G638<= not G645;
	G641<= not G645;
	G644<= not G645;
	G645<= not G90;
	G656<= not G712;
	G658<= not G659;
	G659<= not I1162;
	G661<= not G94;
	G662<= not G712;
	G665<= not G678;
	G668<= not G712;
	G671<= not G678;
	G674<= not G712;
	G677<= not G678;
	G678<= not I1183;
	G685<= not G696;
	G689<= not G696;
	G695<= not G696;
	G696<= not I1203;
	G701BF<= not I1211;
	G701<= not G15;
	G704<= not G712;
	G706<= not G712;
	G711<= not G712;
	G712<= not G14;
	G714<= not G701;
	G715<= not I1227;
	G716<= not I1230;
	G717<= not I1233;
	G718<= not I1236;
	G719<= not I1239;
	G720<= not I1242;
	G721<= not I1245;
	G722<= not I1248;
	G723<= not I1251;
	G724<= not I1254;
	G725<= not I1257;
	G726<= not I1260;
	G728<= not I1264;
	G729<= not I1267;
	I1<= not G332;
	I12<= not G328;
	I1162<= not G13;
	I1183<= not G11;
	I1203<= not G10;
	I1211<= not G701;
	I1227<= not G6;
	I1230<= not G7;
	I1233<= not G8;
	I1236<= not G9;
	I1239<= not G12;
	I1242<= not G0;
	I1245<= not G1;
	I1248<= not G2;
	I1251<= not G3;
	I1254<= not G4;
	I1257<= not G5;
	I1260<= not G93;
	I1264<= not G16;
	I1267<= not G95;
	G101<=G630 and G631;
	G102<=G633 and G634;
	G103<=G636 and G637;
	G104<=G639 and G640;
	G105<=G642 and G643;
	G109<=G106 and G108;
	G113<=G114 and G112;
	G116<=G133 and G25;
	G118<=G119 and G117;
	G121<=G134 and G26;
	G125<=G122 and G124;
	G129<=G130 and G128;
	G132<=G136 and G28;
	G133<=G700 and G111;
	G134<=G133 and G25;
	G135<=G134 and G26;
	G136<=G135 and G127;
	G140<=G137 and G139;
	G144<=G145 and G143;
	G147<=G168 and G30;
	G149<=G150 and G148;
	G152<=G169 and G31;
	G154<=G155 and G153;
	G157<=G170 and G32;
	G159<=G160 and G158;
	G162<=G171 and G33;
	G166<=G163 and G165;
	G168<=G177 and G142;
	G169<=G168 and G30;
	G170<=G169 and G31;
	G171<=G170 and G32;
	G172<=G171 and G33;
	G173<=G172 and G34;
	G175<=G176 and G174;
	G185<=G181 and G182;
	G189<=G186 and G188;
	G193<=G194 and G192;
	G196<=G202 and G37;
	G198<=G199 and G197;
	G201<=G203 and G38;
	G202<=G522 and G191;
	G203<=G202 and G37;
	G208<=G205 and G207;
	G214<=G211 and G213;
	G218<=G219 and G217;
	G221<=G223 and G41;
	G222<=G183 and G210;
	G223<=G222 and G216;
	G224<=G203 and G38;
	G225<=G204 and G203;
	G226<=G136 and G28;
	G227<=G172 and G178;
	G228<=G223 and G41;
	G229<=G432 and G62;
	G237<=G238 and G236;
	G240<=G299 and G42;
	G242<=G243 and G241;
	G245<=G262 and G43;
	G247<=G248 and G246;
	G250<=G263 and G44;
	G252<=G253 and G251;
	G255<=G264 and G45;
	G259<=G624 and G625;
	G260<=G256 and G258;
	G261<=G265 and G46;
	G262<=G299 and G42;
	G263<=G262 and G43;
	G264<=G263 and G44;
	G265<=G264 and G45;
	G271<=G275 and G266;
	G272<=G276 and G277;
	G273<=G278 and G279;
	G274<=G280 and G281;
	G303<=G304 and G302;
	G304<=G306 and G307;
	G309<=G310 and G308;
	G310<=G312 and G313;
	G315<=G316 and G314;
	G316<=G318 and G319;
	G321<=G322 and G320;
	G322<=G325 and G326;
	G329<=G331 and G714;
	G330<=G332 and G714;
	G335<=G337 and G338;
	G342<=G344 and G345;
	G346<=G349 and G350;
	G358<=G523 and G53;
	G360<=G361 and G359;
	G363<=G523 and G51;
	G365<=G366 and G364;
	G368<=G375 and G52;
	G373<=G369 and G371;
	G374<=G376 and G53;
	G375<=G523 and G51;
	G376<=G375 and G52;
	G377<=G183 and G54 and G56;
	G379<=G380 and G378;
	G382<=G183 and G54;
	G384<=G385 and G383;
	G387<=G394 and G55;
	G392<=G388 and G390;
	G393<=G395 and G56;
	G394<=G183 and G54;
	G395<=G394 and G55;
	G397<=G398 and G396;
	G400<=G335 and G57;
	G405<=G401 and G403;
	G406<=G412 and G58;
	G408<=G409 and G407;
	G411<=G413 and G59;
	G412<=G335 and G57;
	G413<=G335 and G58;
	G414<=G413 and G59;
	G416<=G417 and G415;
	G419<=G358 and G60;
	G424<=G420 and G422;
	G425<=G431 and G61;
	G427<=G428 and G426;
	G430<=G432 and G62;
	G431<=G358 and G60;
	G432<=G358 and G61;
	G433<=G356 and G357;
	G435<=G340 and G341;
	G436<=G352 and G353;
	G438<=G439 and G437;
	G441<=G442 and G440;
	G443<=G615 and G511;
	G447<=G448 and G446;
	G451<=G452 and G450;
	G453<=G615 and G445;
	G457<=G455 and G449 and G728;
	G459<=G460 and G458;
	G462<=G434 and G67;
	G464<=G465 and G463;
	G467<=G479 and G68;
	G469<=G470 and G468;
	G472<=G480 and G69;
	G477<=G473 and G475;
	G478<=G481 and G70;
	G479<=G434 and G67;
	G480<=G479 and G68;
	G481<=G480 and G69;
	G488<=G505 and G506;
	G489<=G508 and G509;
	G490<=G512 and G513;
	G494<=G492 and G493;
	G498<=G496 and G497;
	G503<=G501 and G502;
	G526<=G527 and G525;
	G529<=G604 and G74;
	G531<=G532 and G530;
	G534<=G550 and G75;
	G536<=G537 and G535;
	G539<=G551 and G76;
	G541<=G542 and G540;
	G544<=G552 and G77;
	G548<=G545 and G547;
	G549<=G553 and G78;
	G550<=G604 and G74;
	G551<=G550 and G75;
	G552<=G551 and G76;
	G553<=G552 and G77;
	G565<=G563 and G564;
	G569<=G567 and G568;
	G573<=G571 and G572;
	G577<=G575 and G576;
	G589<=G627 and G628;
	G590<=G591 and G588;
	G592<=G594 and G595;
	G601<=G621 and G622;
	G604<=G433 and G524;
	G608<=G606 and G607;
	G613<=G611 and G612;
	G648<=G646 and G647;
	G649<=G618 and G619;
	G650<=G226 and G661;
	G651<=G227 and G87;
	G652<=G228 and G88;
	G653<=G229 and G89;
	G654<=G90 and G476;
	G655<=G91 and G476;
	G657<=G659 and G656;
	G663<=G664 and G662;
	G664<=G666 and G667;
	G669<=G670 and G668;
	G670<=G672 and G673;
	G675<=G676 and G674;
	G676<=G679 and G680;
	G683<=G684 and G685;
	G688<=G690 and G691;
	G694<=G697 and G698;
	G702<=G703 and G645;
	G705<=G230 and G704;
	G707<=G708 and G706;
	G709<=G678 and G89;
	G713<=G599 and G711;
	G727<=G476 and G645;
	G96<= not (G74 and G596);
	G97<= not (G75 and G596);
	G98<= not (G76 and G596);
	G99<= not (G77 and G596);
	G100<= not (G78 and G596);
	G106<= not (G107 and G110);
	G107<= not (G700 and G111);
	G122<= not (G123 and G126);
	G123<= not (G135 and G127);
	G137<= not (G138 and G141);
	G138<= not (G177 and G142);
	G163<= not (G164 and G167);
	G164<= not (G172 and G178);
	G186<= not (G187 and G190);
	G187<= not (G522 and G191);
	G205<= not (G206 and G209);
	G206<= not (G183 and G210);
	G211<= not (G212 and G215);
	G212<= not (G222 and G216);
	G230<= not (G234 and G235);
	G231<= not (G435 and G648);
	G232<= not (G296 and G298 and G435);
	G233<= not (G700 and G232 and G231);
	G234<= not (G649 and G436);
	G266<= not (G286 and G291);
	G267<= not (G287 and G292);
	G268<= not (G288 and G293);
	G269<= not (G284 and G294);
	G270<= not (G285 and G295);
	G284<= not (G45 and G104);
	G285<= not (G46 and G105);
	G286<= not (G42 and G101);
	G287<= not (G43 and G102);
	G288<= not (G44 and G103);
	G297<= not (G289 and G290);
	G298<= not (G297 and G700);
	G301<= not (G50 and G49 and G48 and G47);
	G331<= not (G333 and G22);
	G332<= not (G334 and G331);
	G476<= not (G486 and G616);
	G482<= not (G514 and G518);
	G483<= not (G515 and G519);
	G484<= not (G516 and G520);
	G485<= not (G517 and G521);
	G514<= not (G71 and G67);
	G515<= not (G72 and G68);
	G516<= not (G73 and G69);
	G517<= not (G487 and G70);
	G554<= not (G556 and G557 and G558);
	G555<= not (G559 and G560);
	G556<= not (G578 and G583);
	G557<= not (G579 and G584);
	G558<= not (G580 and G585);
	G559<= not (G581 and G586);
	G560<= not (G582 and G587);
	G578<= not (G79 and G74);
	G579<= not (G80 and G75);
	G580<= not (G81 and G76);
	G581<= not (G82 and G77);
	G582<= not (G561 and G78);
	G597<= not (G602 and G603);
	G598<= not (G435 and G83);
	G616<= not (G482 and G483 and G484 and G485);
	G700<= not (G282 and G283);
	G110<=G700 or G111;
	G126<=G135 or G127;
	G141<=G177 or G142;
	G167<=G172 or G178;
	G177<=G180 or G226;
	G181<=G178 or G180;
	G182<=G35 or G179;
	G183<=G180 or G227;
	G184<=G180 or G173;
	G190<=G522 or G191;
	G209<=G183 or G210;
	G215<=G222 or G216;
	G235<=G649 or G233;
	G275<=G101 or G42;
	G276<=G102 or G43;
	G277<=G267 or G271;
	G278<=G103 or G44;
	G279<=G268 or G272;
	G280<=G104 or G45;
	G281<=G269 or G273;
	G282<=G105 or G46;
	G283<=G270 or G274;
	G291<=G42 or G101;
	G292<=G43 or G102;
	G293<=G44 or G103;
	G294<=G45 or G104;
	G295<=G46 or G105;
	G300<=G50 or G49 or G48 or G47;
	G306<=G47 or G324;
	G307<=G719 or G305;
	G312<=G48 or G324;
	G313<=G47 or G311;
	G318<=G49 or G324;
	G319<=G48 or G317;
	G324<=G377 or G348;
	G325<=G50 or G324;
	G326<=G49 or G323;
	G333<=G300 or G714;
	G334<=G301 or G714;
	G337<=G224 or G355;
	G338<=G183 or G336;
	G340<=G38 or G355;
	G341<=G185 or G339;
	G344<=G229 or G348;
	G345<=G414 or G343;
	G349<=G62 or G348;
	G350<=G59 or G347;
	G352<=G346 or G645;
	G353<=G35 or G351;
	G355<=G457 or G645;
	G356<=G225 or G355;
	G357<=G184 or G354;
	G372<=G712 or G358;
	G391<=G712 or G377;
	G404<=G712 or G413;
	G423<=G712 or G432;
	G434<=G342 or G645;
	G439<=G435 or G63;
	G448<=G615 or G65;
	G456<=G83 or G524;
	G492<=G71 or G500;
	G493<=G488 or G491;
	G496<=G72 or G500;
	G497<=G489 or G495;
	G500<=G654 or G712;
	G501<=G73 or G500;
	G502<=G490 or G499;
	G505<=G723 or G511;
	G506<=G720 or G504;
	G508<=G724 or G511;
	G509<=G721 or G507;
	G512<=G725 or G511;
	G513<=G722 or G510;
	G518<=G71 or G67;
	G519<=G72 or G68;
	G520<=G73 or G69;
	G521<=G487 or G70;
	G522<=G348 or G228;
	G523<=G348 or G414;
	G524<=G554 or G555;
	G563<=G79 or G610;
	G564<=G715 or G562;
	G567<=G80 or G610;
	G568<=G716 or G566;
	G571<=G81 or G610;
	G572<=G717 or G570;
	G575<=G82 or G610;
	G576<=G718 or G574;
	G583<=G79 or G74;
	G584<=G80 or G75;
	G585<=G81 or G76;
	G586<=G82 or G77;
	G587<=G561 or G78;
	G591<=G592 or G604;
	G594<=G83 or G593;
	G602<=G85 or G601;
	G603<=G600 or G84;
	G606<=G84 or G610;
	G607<=G696 or G605;
	G610<=G655 or G712;
	G611<=G85 or G610;
	G612<=G678 or G609;
	G618<=G457 or G645;
	G619<=G715 or G617;
	G621<=G614 or G645;
	G622<=G717 or G620;
	G624<=G476 or G645;
	G625<=G716 or G623;
	G627<=G476 or G645;
	G628<=G718 or G626;
	G630<=G96 or G645;
	G631<=G720 or G629;
	G633<=G97 or G645;
	G634<=G721 or G632;
	G636<=G98 or G645;
	G637<=G722 or G635;
	G639<=G99 or G645;
	G640<=G723 or G638;
	G642<=G100 or G645;
	G643<=G724 or G641;
	G646<=G456 or G645;
	G647<=G725 or G644;
	G666<=G87 or G678;
	G667<=G661 or G665;
	G672<=G88 or G678;
	G673<=G87 or G671;
	G679<=G89 or G678;
	G680<=G88 or G677;
	G682<=G681 or G699;
	G684<=G645 or G696;
	G687<=G686 or G699;
	G690<=G348 or G696;
	G691<=G645 or G689;
	G693<=G692 or G699;
	G697<=G180 or G696;
	G698<=G348 or G695;
	G699<=G658 or G712;
	G114<= not (G115 or G116);
	G115<= not (G133 or G25);
	G119<= not (G120 or G121);
	G120<= not (G134 or G26);
	G130<= not (G131 or G132);
	G131<= not (G136 or G28);
	G145<= not (G146 or G147);
	G146<= not (G168 or G30);
	G150<= not (G151 or G152);
	G151<= not (G169 or G31);
	G155<= not (G156 or G157);
	G156<= not (G170 or G32);
	G160<= not (G161 or G162);
	G161<= not (G171 or G33);
	G194<= not (G195 or G196);
	G195<= not (G202 or G37);
	G199<= not (G200 or G201);
	G200<= not (G203 or G38);
	G219<= not (G220 or G221);
	G220<= not (G223 or G41);
	G238<= not (G239 or G240);
	G239<= not (G299 or G42);
	G243<= not (G244 or G245);
	G244<= not (G262 or G43);
	G248<= not (G249 or G250);
	G249<= not (G263 or G44);
	G253<= not (G254 or G255);
	G254<= not (G264 or G45);
	G256<= not (G257 or G261);
	G257<= not (G265 or G46);
	G289<= not (G270 or G269 or G268);
	G290<= not (G267 or G266);
	G299<= not (G301 or G328);
	G327<= not (G330 or G23);
	G328<= not (G329 or G327);
	G361<= not (G362 or G363);
	G362<= not (G523 or G51);
	G366<= not (G367 or G368);
	G367<= not (G375 or G52);
	G369<= not (G370 or G374);
	G370<= not (G376 or G53);
	G380<= not (G381 or G382);
	G381<= not (G183 or G54);
	G385<= not (G386 or G387);
	G386<= not (G394 or G55);
	G388<= not (G389 or G393);
	G389<= not (G395 or G56);
	G398<= not (G399 or G400);
	G399<= not (G335 or G57);
	G401<= not (G402 or G406);
	G402<= not (G412 or G58);
	G409<= not (G410 or G411);
	G410<= not (G413 or G59);
	G417<= not (G418 or G419);
	G418<= not (G358 or G60);
	G420<= not (G421 or G425);
	G421<= not (G431 or G61);
	G428<= not (G429 or G430);
	G429<= not (G432 or G62);
	G442<= not (G443 or G444);
	G444<= not (G615 or G64);
	G452<= not (G453 or G454);
	G454<= not (G615 or G66);
	G460<= not (G461 or G462);
	G461<= not (G434 or G67);
	G465<= not (G466 or G467);
	G466<= not (G479 or G68);
	G470<= not (G471 or G472);
	G471<= not (G480 or G69);
	G473<= not (G474 or G478);
	G474<= not (G481 or G70);
	G487<= not (G71 or G72 or G73);
	G527<= not (G528 or G529);
	G528<= not (G604 or G74);
	G532<= not (G533 or G534);
	G533<= not (G550 or G75);
	G537<= not (G538 or G539);
	G538<= not (G551 or G76);
	G542<= not (G543 or G544);
	G543<= not (G552 or G77);
	G545<= not (G546 or G549);
	G546<= not (G553 or G78);
	G561<= not (G79 or G80 or G81 or G82);
	G593<= not (G435 or G524);
	G599<= not (G598 or G597);
	G660<= not (G658 or G86);
	G681<= not (G683 or G660);
	G686<= not (G688 or G660);
	G692<= not (G694 or G660);
	G703<= not (G650 or G651 or G652 or G653);
	G708<= not (G709 or G710);
	G710<= not (G678 or G94);
end RTL;
